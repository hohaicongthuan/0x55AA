module layer_10_featuremap_367(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17ae45),
	.w1(32'hbc0f4a2c),
	.w2(32'h3be1052b),
	.w3(32'hbb9af17b),
	.w4(32'h3b9f93e6),
	.w5(32'h3c7fc212),
	.w6(32'hbcbc57e3),
	.w7(32'h3c3906dc),
	.w8(32'h3b94b5b1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df618e),
	.w1(32'h3bbad9f6),
	.w2(32'hbc38b268),
	.w3(32'h3a439070),
	.w4(32'h3c031231),
	.w5(32'hba23bd0b),
	.w6(32'hbc4eed74),
	.w7(32'h3b9d17a5),
	.w8(32'hb9c56a6e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d5e34),
	.w1(32'h3b3139d1),
	.w2(32'h39e096f1),
	.w3(32'h3b9bb93d),
	.w4(32'h3c943283),
	.w5(32'h3b467fb8),
	.w6(32'hbd045939),
	.w7(32'hba3abdcd),
	.w8(32'h3b2c4912),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef92f2),
	.w1(32'h3ce37eea),
	.w2(32'hbba7519c),
	.w3(32'h3cd6b0ba),
	.w4(32'hbcacfbd8),
	.w5(32'h3c273fd8),
	.w6(32'hbb19014d),
	.w7(32'h3c3ecbcb),
	.w8(32'h3bc2b28a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeaee7),
	.w1(32'h3b49d121),
	.w2(32'hbb333576),
	.w3(32'h3ac2f6ba),
	.w4(32'h3b3a3e4f),
	.w5(32'h39a5e813),
	.w6(32'h3bcc67f6),
	.w7(32'h3b528866),
	.w8(32'h3dbc69f2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3bdcd),
	.w1(32'hbc86f41c),
	.w2(32'h3ad5ebad),
	.w3(32'h3989ab27),
	.w4(32'hb8884cb6),
	.w5(32'h3c3fc9e5),
	.w6(32'h3ca1a413),
	.w7(32'hbb878985),
	.w8(32'hbb6f4d06),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3615ea),
	.w1(32'hbb94f1c0),
	.w2(32'hbbb4450a),
	.w3(32'hbc70c26a),
	.w4(32'hbd0d62eb),
	.w5(32'hbc0ba074),
	.w6(32'hbb3a4cc4),
	.w7(32'h3bcedc7e),
	.w8(32'h3c0bda3b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6dd6d),
	.w1(32'h3af947a4),
	.w2(32'h3c2ade74),
	.w3(32'hb9ba94c1),
	.w4(32'h3c3e9555),
	.w5(32'h39d1e750),
	.w6(32'h3c08203e),
	.w7(32'h3acc8c9f),
	.w8(32'hbbc0ce7e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae975f),
	.w1(32'hbc15e288),
	.w2(32'hbd06d4e8),
	.w3(32'h3c3180e8),
	.w4(32'hbb114a49),
	.w5(32'hbbfd2862),
	.w6(32'hbba5d711),
	.w7(32'h39dc582c),
	.w8(32'h3acc97a7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8ad8f),
	.w1(32'hbb2fcedd),
	.w2(32'h3c37ce87),
	.w3(32'hbb7c33a1),
	.w4(32'hbb5ff179),
	.w5(32'hbbbfbc3a),
	.w6(32'hbc46e7d0),
	.w7(32'hbba54168),
	.w8(32'h3bacbaa2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2a25c),
	.w1(32'hbc044a00),
	.w2(32'h3b0c03af),
	.w3(32'h3c71fe14),
	.w4(32'hbc350247),
	.w5(32'h3c973a9e),
	.w6(32'h3bb4da6d),
	.w7(32'hbbd43233),
	.w8(32'h3aa1d05b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54f08c),
	.w1(32'hbbface1b),
	.w2(32'h3cdfc0b9),
	.w3(32'hbbff9f71),
	.w4(32'h3c13c821),
	.w5(32'h3b9a353e),
	.w6(32'hbb49775e),
	.w7(32'hb90496d3),
	.w8(32'h3b26ca51),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8911b6),
	.w1(32'h3c484925),
	.w2(32'h3b4cef51),
	.w3(32'h3a21fec5),
	.w4(32'hba6e72ae),
	.w5(32'h3c102246),
	.w6(32'h3c356090),
	.w7(32'h3bb0f642),
	.w8(32'h3a837e98),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4162e),
	.w1(32'h3cacd9ce),
	.w2(32'hbb5848d6),
	.w3(32'hbab89f1a),
	.w4(32'hbcee4ea2),
	.w5(32'hbc4de5f4),
	.w6(32'h3b0829ed),
	.w7(32'hbb2e1fc0),
	.w8(32'h3938d28f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f6a81),
	.w1(32'h3bb2f756),
	.w2(32'h39e2912e),
	.w3(32'h3a6c7bdb),
	.w4(32'hbc1e89c7),
	.w5(32'h3b419fb8),
	.w6(32'hbbee3689),
	.w7(32'hbb0cda71),
	.w8(32'hba22db6f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b725576),
	.w1(32'h3b69a823),
	.w2(32'h3bb847de),
	.w3(32'h3b754c20),
	.w4(32'hbb02c723),
	.w5(32'hba05ad21),
	.w6(32'h3bcd2b87),
	.w7(32'hbc60927f),
	.w8(32'hbc39fbd9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c900c),
	.w1(32'hbc9a1c21),
	.w2(32'h3adb8360),
	.w3(32'hbad59a99),
	.w4(32'h3a722d2c),
	.w5(32'h3b5b87da),
	.w6(32'h3b740306),
	.w7(32'hbac0b297),
	.w8(32'hba92510c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b52b4),
	.w1(32'hbcae791c),
	.w2(32'h3c1f9d20),
	.w3(32'h3b436b06),
	.w4(32'hbb329b78),
	.w5(32'hbb3c1980),
	.w6(32'h3bd6f22f),
	.w7(32'h3d6f8be7),
	.w8(32'h3b7ccb6b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21beb8),
	.w1(32'hbc6c7c35),
	.w2(32'h3a97f49e),
	.w3(32'h3b2783c4),
	.w4(32'h3ae42c83),
	.w5(32'h3c94818d),
	.w6(32'hbc3555f8),
	.w7(32'h3c817614),
	.w8(32'h3b172622),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fe9ee),
	.w1(32'h3c4ffdaf),
	.w2(32'hb95970ac),
	.w3(32'hbbfa90c7),
	.w4(32'hbda21520),
	.w5(32'h3b91bb79),
	.w6(32'h3bf782a3),
	.w7(32'h3b713c84),
	.w8(32'hbb2b618c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b295928),
	.w1(32'hba3a7e15),
	.w2(32'hbd40f008),
	.w3(32'h3b8a8f52),
	.w4(32'hbb8ce7f6),
	.w5(32'hbba927ae),
	.w6(32'h3bb5fe56),
	.w7(32'h3a6386f3),
	.w8(32'h3ae4fd1a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5adbc0),
	.w1(32'hbad3e135),
	.w2(32'h3a1741c2),
	.w3(32'h3be4a1e3),
	.w4(32'h3a897752),
	.w5(32'hbbcde9b4),
	.w6(32'hbc0508ba),
	.w7(32'h3b6ccdf4),
	.w8(32'h3b898300),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2b1d1),
	.w1(32'h3a5e475e),
	.w2(32'h3cb21608),
	.w3(32'hb98f4c03),
	.w4(32'h3a9a119c),
	.w5(32'hbbd34194),
	.w6(32'h3be49a39),
	.w7(32'hbc1093d0),
	.w8(32'hbc2dca4b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc490f32),
	.w1(32'hbaf8a5bc),
	.w2(32'hbaa3c4c2),
	.w3(32'hbb0b33d3),
	.w4(32'hbb587e7b),
	.w5(32'hb82653d1),
	.w6(32'hba0443be),
	.w7(32'hbbd7c010),
	.w8(32'hbbd565ae),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3a627),
	.w1(32'h3c8ac97d),
	.w2(32'h3b9e87dd),
	.w3(32'h3be565ec),
	.w4(32'hbd4f7d06),
	.w5(32'hbb83792d),
	.w6(32'h3b0e2c13),
	.w7(32'hbbad2a95),
	.w8(32'hbcdb053f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b573559),
	.w1(32'hbb9ce8d6),
	.w2(32'hb87197eb),
	.w3(32'hbb55aee7),
	.w4(32'h3a3ec633),
	.w5(32'hbbc42d01),
	.w6(32'hbb043491),
	.w7(32'hba11e5fd),
	.w8(32'h3ae6102f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4a541),
	.w1(32'hbc359ac5),
	.w2(32'h3ba35b0b),
	.w3(32'hb92312d4),
	.w4(32'hb9fcb7da),
	.w5(32'h3b2af346),
	.w6(32'h3c04ea88),
	.w7(32'h3c07506b),
	.w8(32'h3b616e38),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4f388),
	.w1(32'hbbe520ae),
	.w2(32'h3c9b6dab),
	.w3(32'h3bd00290),
	.w4(32'h3c086dea),
	.w5(32'h3bff5935),
	.w6(32'h3adad043),
	.w7(32'hba749ae3),
	.w8(32'hbb68fdab),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e6d49),
	.w1(32'hbb5bd0d6),
	.w2(32'hbc9e7606),
	.w3(32'h3b812d9c),
	.w4(32'hbbe18bb6),
	.w5(32'hba439169),
	.w6(32'h3af11c86),
	.w7(32'h3ab2be40),
	.w8(32'hbb5709f2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd68223),
	.w1(32'h39a1f22a),
	.w2(32'h3b915dcf),
	.w3(32'h3a3e5674),
	.w4(32'h3d2a4e95),
	.w5(32'hbb298274),
	.w6(32'h3ba8a956),
	.w7(32'h3b617e81),
	.w8(32'hbc0e760f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bc38a),
	.w1(32'hbab427e0),
	.w2(32'hbcb49cc0),
	.w3(32'h3b8fad33),
	.w4(32'h3b349c59),
	.w5(32'h39031a4d),
	.w6(32'hbb98a4b9),
	.w7(32'h3b87f652),
	.w8(32'h3c8cdece),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be07ae0),
	.w1(32'h39e5cf57),
	.w2(32'hbbc5e5a1),
	.w3(32'h3b93048a),
	.w4(32'h3b7916cb),
	.w5(32'hbcbdc0ce),
	.w6(32'h3c5047b6),
	.w7(32'hbc87ac3d),
	.w8(32'h3bf46316),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc385c3d),
	.w1(32'h3ad76f73),
	.w2(32'hbc6c77f2),
	.w3(32'hbb31b9bd),
	.w4(32'h3b5e363e),
	.w5(32'hbc7fa9f4),
	.w6(32'h3b85ab0c),
	.w7(32'h3ba44dbe),
	.w8(32'hbb96ba84),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d9599),
	.w1(32'h3d0f859d),
	.w2(32'h3a3fe230),
	.w3(32'hbba8e694),
	.w4(32'hbbbe68ef),
	.w5(32'h3aa53a64),
	.w6(32'hbab2aa2e),
	.w7(32'hbab6ffde),
	.w8(32'hbb66117f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c344482),
	.w1(32'h3b0e62e0),
	.w2(32'hba1c31e5),
	.w3(32'hbac1fcc7),
	.w4(32'hbbf7def5),
	.w5(32'hbba3c036),
	.w6(32'hbb294bd0),
	.w7(32'hbbf8c7c4),
	.w8(32'hbd3d35db),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d37db),
	.w1(32'hbca8399f),
	.w2(32'hbc08d447),
	.w3(32'hbaba1ba2),
	.w4(32'hbc3f3b4e),
	.w5(32'hbab5042d),
	.w6(32'hbbae67ed),
	.w7(32'hbc71da0f),
	.w8(32'h3a67f074),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fb471),
	.w1(32'hbb267326),
	.w2(32'h3aea4d94),
	.w3(32'hbb6dff47),
	.w4(32'hbb6b022e),
	.w5(32'hbc97132a),
	.w6(32'hbbe37e8e),
	.w7(32'h3baa57b0),
	.w8(32'h3bb825e2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec2418),
	.w1(32'hbc5ad307),
	.w2(32'hbbe4d279),
	.w3(32'h3b820db5),
	.w4(32'h3cf8ffcc),
	.w5(32'hb936a15f),
	.w6(32'h3c154b9b),
	.w7(32'h3b94bcc4),
	.w8(32'hba9ee3ff),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6a3ea),
	.w1(32'hbb48ae8f),
	.w2(32'h3b976f1c),
	.w3(32'h3b5453ff),
	.w4(32'h3b815426),
	.w5(32'h3c8361b1),
	.w6(32'hbba9dfee),
	.w7(32'h3b47e34a),
	.w8(32'hbca65d0e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c94568),
	.w1(32'hbbac3c82),
	.w2(32'hbb152f2a),
	.w3(32'hba40c26b),
	.w4(32'h388580c4),
	.w5(32'hba9a84a9),
	.w6(32'h3c1e531c),
	.w7(32'hbb542572),
	.w8(32'h3c33be58),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72c69b6),
	.w1(32'h3bb699cf),
	.w2(32'hbc66641d),
	.w3(32'h3cc5a1a8),
	.w4(32'hbc8c2b7f),
	.w5(32'h3be8c04c),
	.w6(32'hbaf91b38),
	.w7(32'hbadcb28b),
	.w8(32'hbb52a440),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba935854),
	.w1(32'hbacf68d8),
	.w2(32'hbd10455d),
	.w3(32'h3bf36f3f),
	.w4(32'hbd37f217),
	.w5(32'h3b990c03),
	.w6(32'hbabce434),
	.w7(32'hba60ced6),
	.w8(32'hbccdcc0c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcffd310),
	.w1(32'hbb138fa1),
	.w2(32'hbbac5a98),
	.w3(32'hbc0e3ad3),
	.w4(32'hbc1b4705),
	.w5(32'hba9dd93a),
	.w6(32'hbbfbb0da),
	.w7(32'h3acd35ad),
	.w8(32'hbc1f7ba4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea0798),
	.w1(32'h3b5a29a0),
	.w2(32'h3bdcd5c8),
	.w3(32'hba51249f),
	.w4(32'hba8de7e8),
	.w5(32'h3a80200d),
	.w6(32'h3b9eaea6),
	.w7(32'h3c82b65d),
	.w8(32'hba86ba38),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e5ca9),
	.w1(32'hbd04a973),
	.w2(32'h3b776803),
	.w3(32'hb941bb52),
	.w4(32'h3bc8a6d1),
	.w5(32'hbc79d1bd),
	.w6(32'h3bd135e1),
	.w7(32'h3b4b10b3),
	.w8(32'h3a28842d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c498c),
	.w1(32'h3a8ef045),
	.w2(32'hbc215788),
	.w3(32'h3a3e3807),
	.w4(32'h3bf679b5),
	.w5(32'h3cfa2547),
	.w6(32'h3b05fb36),
	.w7(32'hbb90ad2b),
	.w8(32'hbbad2750),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d34229f),
	.w1(32'h3b3f9504),
	.w2(32'hbaeaaf06),
	.w3(32'h3c043eb8),
	.w4(32'h3c0daf4f),
	.w5(32'h3bd1b550),
	.w6(32'h3b85a284),
	.w7(32'hbb60f40c),
	.w8(32'h3b1a8772),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7660cc),
	.w1(32'hb939c5d1),
	.w2(32'hbb5c98db),
	.w3(32'hba26ea6f),
	.w4(32'hbcc2e165),
	.w5(32'hbc2566af),
	.w6(32'h3c2705fc),
	.w7(32'hbbe1afd1),
	.w8(32'hbd0d1e7a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1406c9),
	.w1(32'h39e5d397),
	.w2(32'h3cacd3a7),
	.w3(32'h3b67b875),
	.w4(32'hbb5e187c),
	.w5(32'hbb75fd26),
	.w6(32'h3b42ed2e),
	.w7(32'hbba05c03),
	.w8(32'hbc077bdb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3427e6),
	.w1(32'h3c269a39),
	.w2(32'h3c1523ff),
	.w3(32'hbd196b10),
	.w4(32'hbc3d04d2),
	.w5(32'h3a9584f4),
	.w6(32'h3b69513b),
	.w7(32'h3ba3f675),
	.w8(32'hbb0616a4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d76b5),
	.w1(32'h3bbce448),
	.w2(32'hbad0ed37),
	.w3(32'h38a8f119),
	.w4(32'h3c37ae75),
	.w5(32'h3a0ffeef),
	.w6(32'hbbfdc242),
	.w7(32'h3a370dc5),
	.w8(32'h3b654395),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf5d3d),
	.w1(32'hbcadb4c3),
	.w2(32'hbb01238b),
	.w3(32'hbb642643),
	.w4(32'h3c442512),
	.w5(32'hbc2d086d),
	.w6(32'h3a1df3b4),
	.w7(32'h3b9a2bf7),
	.w8(32'hbb43cefa),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b989b),
	.w1(32'h3bd378be),
	.w2(32'h3c17e53f),
	.w3(32'hb8f86284),
	.w4(32'hb88810c9),
	.w5(32'hbcab2be3),
	.w6(32'hbb116b1f),
	.w7(32'hbc17c0c1),
	.w8(32'h3abf60ad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf7519),
	.w1(32'hbb25b972),
	.w2(32'hbc271f02),
	.w3(32'hbb363d6e),
	.w4(32'h3c38b13e),
	.w5(32'hb964852a),
	.w6(32'h3c03bd7a),
	.w7(32'hbc839f66),
	.w8(32'hbc1491fa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15f04e),
	.w1(32'hba0a89ca),
	.w2(32'h3b25fe13),
	.w3(32'hbb4c9610),
	.w4(32'hbbc7053c),
	.w5(32'hbba2edc5),
	.w6(32'hba94f74b),
	.w7(32'h39d31728),
	.w8(32'h3b9e9c85),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a993794),
	.w1(32'hbbe3d2f6),
	.w2(32'hbb085097),
	.w3(32'hbc369b07),
	.w4(32'hbc84fe06),
	.w5(32'h3c2072bf),
	.w6(32'h3b25d000),
	.w7(32'h3c8a6551),
	.w8(32'h398ddf09),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4afa5),
	.w1(32'hba205d52),
	.w2(32'h3c35223b),
	.w3(32'h3c90c9e0),
	.w4(32'hbad625fb),
	.w5(32'hbb9b0999),
	.w6(32'hbc63d79e),
	.w7(32'h3bc6bf78),
	.w8(32'hbbb3e945),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dcba8d),
	.w1(32'h3b0db321),
	.w2(32'h3ce26894),
	.w3(32'h3cc977d1),
	.w4(32'hb9cf9b30),
	.w5(32'h3b5a86b7),
	.w6(32'h3ac643cc),
	.w7(32'h3be21bf2),
	.w8(32'h3bfe89aa),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb21593),
	.w1(32'hbbb9fb00),
	.w2(32'hbbc592fd),
	.w3(32'hba541184),
	.w4(32'hbb7e0a01),
	.w5(32'h3be3d553),
	.w6(32'hbc7f4308),
	.w7(32'hbbd921a7),
	.w8(32'hbb9af2cb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea8e9a),
	.w1(32'h3c10d501),
	.w2(32'h3aea4521),
	.w3(32'h3ba07f77),
	.w4(32'hbc114062),
	.w5(32'hbc20442f),
	.w6(32'hbba27ce7),
	.w7(32'hbc3e2ef3),
	.w8(32'hbc9b0a98),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a643821),
	.w1(32'hbab47247),
	.w2(32'hbb8868f4),
	.w3(32'hbb5e3c9d),
	.w4(32'hbbe22946),
	.w5(32'hbcb242b3),
	.w6(32'hbc2122d9),
	.w7(32'hbb6c1848),
	.w8(32'hbc8523be),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0c2f),
	.w1(32'hbcd9a430),
	.w2(32'h3ae45e1d),
	.w3(32'hba06e95c),
	.w4(32'hbb17082d),
	.w5(32'hbcdb52ec),
	.w6(32'hba7ffdbf),
	.w7(32'hbaad1507),
	.w8(32'h3b132375),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74df2c),
	.w1(32'hbb6be0a1),
	.w2(32'h3cbe6b13),
	.w3(32'hba011403),
	.w4(32'hb9798bba),
	.w5(32'hbc9b85ee),
	.w6(32'hbc232a17),
	.w7(32'hbbc57a22),
	.w8(32'h3bbba423),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a61b4),
	.w1(32'h3beabc62),
	.w2(32'hbc3c2bff),
	.w3(32'hbbf76515),
	.w4(32'hbaa0ed6f),
	.w5(32'h3a89999a),
	.w6(32'h3c183bfb),
	.w7(32'hbc370378),
	.w8(32'h3c38b58d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0090e),
	.w1(32'h3ca4bd30),
	.w2(32'hbb897ab7),
	.w3(32'h3a5448ca),
	.w4(32'hbb060efa),
	.w5(32'h3c024b50),
	.w6(32'h3b90db5a),
	.w7(32'h3c948eda),
	.w8(32'h3a8c4746),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9782cae),
	.w1(32'hbb5c2f65),
	.w2(32'hbc0606e6),
	.w3(32'hbb855513),
	.w4(32'h3be717ae),
	.w5(32'hbaf431e9),
	.w6(32'h3c48795b),
	.w7(32'hbc1fb128),
	.w8(32'h3b415d6d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9da54),
	.w1(32'h3ab63c7d),
	.w2(32'hbbf93f24),
	.w3(32'h3a15485a),
	.w4(32'hbc3df6a9),
	.w5(32'h3cd4dfa3),
	.w6(32'hbac4d81a),
	.w7(32'h3d0350cc),
	.w8(32'h3bf740a0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c333d61),
	.w1(32'hbaa4a441),
	.w2(32'h3c1d0541),
	.w3(32'hbc75b5f5),
	.w4(32'hbb6c8d34),
	.w5(32'hbd04bedc),
	.w6(32'hbc747281),
	.w7(32'hbc592fbc),
	.w8(32'h3b0c8bd1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d474e8),
	.w1(32'h3bde2f21),
	.w2(32'h3bd3da55),
	.w3(32'hbb264e6b),
	.w4(32'hba24bb74),
	.w5(32'hbc894c3d),
	.w6(32'hbbf551bb),
	.w7(32'h3b0f4371),
	.w8(32'hbd46c156),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9915a),
	.w1(32'hbbcd7974),
	.w2(32'h3caddfb4),
	.w3(32'h3b973155),
	.w4(32'hbc928775),
	.w5(32'hbb372840),
	.w6(32'hb98ba12d),
	.w7(32'hbb0c4f91),
	.w8(32'hbbe4f529),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65149c),
	.w1(32'hbac9a7da),
	.w2(32'hbc7b0600),
	.w3(32'h39f86bf0),
	.w4(32'hbb1a7383),
	.w5(32'hbbbc28d2),
	.w6(32'hbb8f12cb),
	.w7(32'hbc89e2a3),
	.w8(32'hbc877ddc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8c323),
	.w1(32'h3b927dfc),
	.w2(32'hbbc6341d),
	.w3(32'hbc25d332),
	.w4(32'hbc5af68f),
	.w5(32'hbb250e5a),
	.w6(32'h3b75886a),
	.w7(32'h3b57b60e),
	.w8(32'h3c724f88),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d05a0),
	.w1(32'h3a2c545b),
	.w2(32'hba82fc42),
	.w3(32'hbc4b50be),
	.w4(32'hbc2acca9),
	.w5(32'h3bfa542a),
	.w6(32'h3add4e55),
	.w7(32'h3b3d8b1f),
	.w8(32'h3aec4565),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39f877),
	.w1(32'h39fa5751),
	.w2(32'hbc37c9a7),
	.w3(32'hbbb073b8),
	.w4(32'h3bd23362),
	.w5(32'hbc303e0a),
	.w6(32'hbacac88c),
	.w7(32'hbbfa7b52),
	.w8(32'h3cc868a4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e95ea),
	.w1(32'h3c808422),
	.w2(32'hb81a9ff9),
	.w3(32'h3c1f32b2),
	.w4(32'hbc388ee8),
	.w5(32'hbc41a00c),
	.w6(32'hbbb73563),
	.w7(32'hbc9b2d7a),
	.w8(32'h3cc829dd),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4dbbd),
	.w1(32'hbb8b7e64),
	.w2(32'hbbbe5c7a),
	.w3(32'hbc2c0735),
	.w4(32'h3abf6c3c),
	.w5(32'hbb22cb14),
	.w6(32'hbc76817e),
	.w7(32'hbbdc6be5),
	.w8(32'h3a6f1e49),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ce05a),
	.w1(32'h3b1afff1),
	.w2(32'h3b098f09),
	.w3(32'hbc001d4a),
	.w4(32'hbb176243),
	.w5(32'hbbbbc3d9),
	.w6(32'h39d24874),
	.w7(32'h399e85c2),
	.w8(32'hba4d51d2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5501d8),
	.w1(32'h3b86942f),
	.w2(32'h3b7bcc4d),
	.w3(32'h3bac61e5),
	.w4(32'hbc188307),
	.w5(32'h3b0d7048),
	.w6(32'h3afcc3f7),
	.w7(32'hbae76e55),
	.w8(32'hbc53efbf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7602a50),
	.w1(32'hbb12571b),
	.w2(32'hbc52bb3d),
	.w3(32'h3b037fdf),
	.w4(32'h3c11f12e),
	.w5(32'h3bd012cb),
	.w6(32'h3b4f8b53),
	.w7(32'hbac6a779),
	.w8(32'hbb209b7d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f68ae),
	.w1(32'hbb2da5c7),
	.w2(32'h3bc919b2),
	.w3(32'h3b638742),
	.w4(32'hba45b804),
	.w5(32'hbb3f654e),
	.w6(32'h3953dc22),
	.w7(32'h3c427290),
	.w8(32'h3bdae8c2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd0310),
	.w1(32'hbbf1de24),
	.w2(32'hbb31bfa9),
	.w3(32'hbc21c349),
	.w4(32'h3c00b9da),
	.w5(32'h399f85cb),
	.w6(32'h3ca35087),
	.w7(32'hbc06d4b8),
	.w8(32'hba62a36f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d018202),
	.w1(32'hbb92fc18),
	.w2(32'h3c010bb9),
	.w3(32'hbc18e706),
	.w4(32'hbaaf4b75),
	.w5(32'hbb78b3be),
	.w6(32'hbc1347b7),
	.w7(32'h3c98b903),
	.w8(32'h39abface),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8601bb2),
	.w1(32'hbba883c4),
	.w2(32'hba4c3d07),
	.w3(32'hbb49973e),
	.w4(32'h3c93e597),
	.w5(32'hbbb75a64),
	.w6(32'hbc785fb9),
	.w7(32'h3d0af52b),
	.w8(32'h3bfbc988),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa417d),
	.w1(32'hbc5f6188),
	.w2(32'h3b9401b7),
	.w3(32'h3bb457fd),
	.w4(32'h3bbd1784),
	.w5(32'h3c40a6eb),
	.w6(32'hbb6e8780),
	.w7(32'h3c878351),
	.w8(32'hbc4337cc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d860b),
	.w1(32'hbb7e9924),
	.w2(32'hbbdec1c2),
	.w3(32'h3bace56e),
	.w4(32'hbc78a185),
	.w5(32'h3b1887a2),
	.w6(32'h3c4e5497),
	.w7(32'hbc75eeee),
	.w8(32'h3c09dedf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ac712),
	.w1(32'hbb39b5b4),
	.w2(32'hbb2e76de),
	.w3(32'hbc213d10),
	.w4(32'h3b31ce73),
	.w5(32'hbc6e3b03),
	.w6(32'hbb6168f3),
	.w7(32'hbb2c37ea),
	.w8(32'hbb3084b3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974c8ab),
	.w1(32'hba022715),
	.w2(32'hbd13e187),
	.w3(32'h3d0efe71),
	.w4(32'h3c3a9d03),
	.w5(32'h3d03660a),
	.w6(32'hbb3ffe41),
	.w7(32'h3bb6da98),
	.w8(32'h3ba2218a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7ced6),
	.w1(32'h3b88b822),
	.w2(32'h3c240752),
	.w3(32'hb97775ec),
	.w4(32'h3c2b1cf7),
	.w5(32'hbb92b0b0),
	.w6(32'hbc40f05b),
	.w7(32'hbc18646a),
	.w8(32'h3c4d98f8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c0206),
	.w1(32'h3c4363dd),
	.w2(32'h3b541960),
	.w3(32'h3b0ed6f0),
	.w4(32'hbb544a02),
	.w5(32'hbc87e3cc),
	.w6(32'h3b52b328),
	.w7(32'hbbd2026e),
	.w8(32'hbccc6db6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a34ed),
	.w1(32'hbb8ede73),
	.w2(32'h3ca07793),
	.w3(32'hbc2e95f4),
	.w4(32'hbc32aed4),
	.w5(32'h3b6166ef),
	.w6(32'h3cc45a72),
	.w7(32'hbb7979dc),
	.w8(32'h3c52eef3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3be0e),
	.w1(32'h3bfb6a21),
	.w2(32'h3ca227a7),
	.w3(32'h3c018002),
	.w4(32'h3bd7e2e0),
	.w5(32'h3bf0f646),
	.w6(32'hbbee3ed7),
	.w7(32'hbc344cfd),
	.w8(32'h3c8f8f7d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2394d),
	.w1(32'h3c93822a),
	.w2(32'hbc18a6db),
	.w3(32'h3c1bbc02),
	.w4(32'hbbb224dc),
	.w5(32'hbcc0e229),
	.w6(32'hba9824b0),
	.w7(32'h3be55c32),
	.w8(32'hbc19640f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2043f9),
	.w1(32'h3c101848),
	.w2(32'h3cc3fe34),
	.w3(32'h3aec4548),
	.w4(32'h3c74421b),
	.w5(32'hbb1908cc),
	.w6(32'h3c57d9f4),
	.w7(32'h3c15ea7a),
	.w8(32'hbc87a7ae),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd4764c),
	.w1(32'hbbf1b0c0),
	.w2(32'h3d1bd433),
	.w3(32'hbb3bcde8),
	.w4(32'h3c634f3c),
	.w5(32'hbba95dd0),
	.w6(32'h3c84bd18),
	.w7(32'hbcb2351b),
	.w8(32'hbbf4a2b1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47c961),
	.w1(32'h3bf8c56b),
	.w2(32'h3aacd9d9),
	.w3(32'h3c817be9),
	.w4(32'h3b73303a),
	.w5(32'hbbef28e5),
	.w6(32'hb9957ac9),
	.w7(32'hbb63eff7),
	.w8(32'hbc51f711),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf7c3e0),
	.w1(32'hbc7da095),
	.w2(32'h3ba594a1),
	.w3(32'h3b834adc),
	.w4(32'h3c842f97),
	.w5(32'h3c20501f),
	.w6(32'h3cc13d3c),
	.w7(32'hbd249957),
	.w8(32'h3aaec21a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcad923),
	.w1(32'h3c4194d6),
	.w2(32'h3bb3ee91),
	.w3(32'hbc7298ad),
	.w4(32'h3b12e248),
	.w5(32'hbb1adcde),
	.w6(32'hbcd4ab14),
	.w7(32'h3baebe6f),
	.w8(32'hb7cfdbfa),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819d4e),
	.w1(32'hbc85e790),
	.w2(32'hbce625d8),
	.w3(32'hbc31b6eb),
	.w4(32'h3b1fc305),
	.w5(32'hbbad0a42),
	.w6(32'hbc9fe3f9),
	.w7(32'h3bc0c21e),
	.w8(32'hbc7c4457),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97e915),
	.w1(32'h3c69a123),
	.w2(32'hbc7ac2ce),
	.w3(32'h3b887893),
	.w4(32'hbca2594b),
	.w5(32'hbbac69ef),
	.w6(32'h3c8ffd01),
	.w7(32'h3ac6cd69),
	.w8(32'hbcb95192),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c4bd4),
	.w1(32'hbbc38d0a),
	.w2(32'h3c36d136),
	.w3(32'h3c8580a9),
	.w4(32'h3bd4a453),
	.w5(32'hba906e4d),
	.w6(32'h3cfa9b47),
	.w7(32'hbc116f53),
	.w8(32'h3bc2891c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa138f8),
	.w1(32'h3c4ed29a),
	.w2(32'h3a913bba),
	.w3(32'h3b3eb06f),
	.w4(32'h3b7e4de0),
	.w5(32'h3b85bee2),
	.w6(32'h3bf00cef),
	.w7(32'h3c03a8d0),
	.w8(32'h3a50763a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8f983),
	.w1(32'h3a26741d),
	.w2(32'hbbdecec6),
	.w3(32'hbb37f5e4),
	.w4(32'h3b98a0a7),
	.w5(32'h3a5bc233),
	.w6(32'h3bbae5fc),
	.w7(32'h3c3b08b0),
	.w8(32'h3b8f9f36),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e42fe),
	.w1(32'hbc643288),
	.w2(32'hba14fa94),
	.w3(32'hbb9aafcb),
	.w4(32'h3b07b8e7),
	.w5(32'hbbcb94c5),
	.w6(32'hbbd80814),
	.w7(32'hbbac9af4),
	.w8(32'h3b68bcd0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca88035),
	.w1(32'h3cf9a662),
	.w2(32'h3cd5a140),
	.w3(32'h3b998a6b),
	.w4(32'h3b90db2d),
	.w5(32'hbb32a05c),
	.w6(32'hbc2c9bdd),
	.w7(32'hbc5baeaa),
	.w8(32'h3c1532c4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7548ff),
	.w1(32'hbc185460),
	.w2(32'h3c1abee9),
	.w3(32'hbc5a312d),
	.w4(32'hbc0773c2),
	.w5(32'hbc16b572),
	.w6(32'h3a7d7352),
	.w7(32'hba2c573e),
	.w8(32'hbaea59f7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60f24f),
	.w1(32'hbc5fcc0f),
	.w2(32'h3b1e9f0d),
	.w3(32'hbbcfed68),
	.w4(32'hbc034052),
	.w5(32'h3b4b72cf),
	.w6(32'hbb111c77),
	.w7(32'h3c960d13),
	.w8(32'hb9ca32a4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc760d21),
	.w1(32'h3bb0d8c1),
	.w2(32'hba8891b4),
	.w3(32'hbb67ca53),
	.w4(32'h3bb35bec),
	.w5(32'h3b254475),
	.w6(32'h3ba61443),
	.w7(32'h3c3f63a8),
	.w8(32'h3bc9c474),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6445f),
	.w1(32'h3ae8dccb),
	.w2(32'h39321584),
	.w3(32'hbbe87c4d),
	.w4(32'h3aabd114),
	.w5(32'h3a996de0),
	.w6(32'h3c8f09e7),
	.w7(32'hbb30db8c),
	.w8(32'h3bddbb18),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1e528),
	.w1(32'h3bd4d8e1),
	.w2(32'h3d08c6de),
	.w3(32'hbc2d4097),
	.w4(32'h3b76d9fd),
	.w5(32'h3b038b7b),
	.w6(32'hbc7548e8),
	.w7(32'h3c1be872),
	.w8(32'hbbea8362),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021199),
	.w1(32'hbbdc4744),
	.w2(32'hba6ba9f7),
	.w3(32'h3b9727db),
	.w4(32'h3bedad8b),
	.w5(32'hbba57d30),
	.w6(32'hbb9f6cad),
	.w7(32'hbc57ba35),
	.w8(32'h3b932d6f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58ac09),
	.w1(32'hba12e168),
	.w2(32'h3c0c4da4),
	.w3(32'h3c1223a8),
	.w4(32'hbc06f81d),
	.w5(32'h3c4242ae),
	.w6(32'hbbf9db0c),
	.w7(32'hbc556d0e),
	.w8(32'h3c681414),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd5ee1),
	.w1(32'h3d16b0fe),
	.w2(32'h3b051df1),
	.w3(32'hbb16204a),
	.w4(32'h3c2232d7),
	.w5(32'hbb2379fa),
	.w6(32'hbbf883ba),
	.w7(32'h3c99ef6a),
	.w8(32'h3c30142c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36e77f),
	.w1(32'hbc50ba58),
	.w2(32'hbc7ebd91),
	.w3(32'hbbe6ab3c),
	.w4(32'h3bc42acc),
	.w5(32'hbb893695),
	.w6(32'hb8b72720),
	.w7(32'h3bcc8d71),
	.w8(32'hbb4de69e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a1200),
	.w1(32'h3c154607),
	.w2(32'hbc3ac664),
	.w3(32'hbb3463f7),
	.w4(32'h3ba7156d),
	.w5(32'hbc76f18b),
	.w6(32'h3c6f272a),
	.w7(32'hbbc0eea8),
	.w8(32'h39aa3e53),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870010),
	.w1(32'hbc11d36d),
	.w2(32'h3b26b576),
	.w3(32'hbc69000f),
	.w4(32'h3c981b38),
	.w5(32'h3c3fa267),
	.w6(32'hbc0843bc),
	.w7(32'h3c083d08),
	.w8(32'hbb88cf7c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23dc71),
	.w1(32'hbc714536),
	.w2(32'h3b14ec73),
	.w3(32'h3ad4c4d7),
	.w4(32'h3c2f7c4a),
	.w5(32'hbb05bc60),
	.w6(32'hbc0f9e22),
	.w7(32'h39bcec73),
	.w8(32'h3b30de71),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb6b8c),
	.w1(32'hb91d6a7b),
	.w2(32'h3c1afb20),
	.w3(32'hbabfe985),
	.w4(32'hbc4ef159),
	.w5(32'hbcd47736),
	.w6(32'hbb3cc553),
	.w7(32'hbc15c4c8),
	.w8(32'h3b18de8e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f35e4),
	.w1(32'h3c708e44),
	.w2(32'hbad47f1c),
	.w3(32'hbbe0521d),
	.w4(32'h3a3bf382),
	.w5(32'h3c3035a4),
	.w6(32'h3c34dfe8),
	.w7(32'hbbf569c9),
	.w8(32'hbaf42fe3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45f382),
	.w1(32'h3af25606),
	.w2(32'h3a2fab0e),
	.w3(32'hba96c054),
	.w4(32'h3c473353),
	.w5(32'h3c1d51af),
	.w6(32'h3c181787),
	.w7(32'hb96fc913),
	.w8(32'hbaf65524),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0971a5),
	.w1(32'hbc21fd42),
	.w2(32'h3aa3dd07),
	.w3(32'hbbd2963d),
	.w4(32'h3b303376),
	.w5(32'h3bd17948),
	.w6(32'h3a5fc7b4),
	.w7(32'h3d194be9),
	.w8(32'hbc14e27f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a3ce5),
	.w1(32'hbb287776),
	.w2(32'hbacd6b44),
	.w3(32'hbc1ee8ba),
	.w4(32'hbaac45e4),
	.w5(32'h3c7293fb),
	.w6(32'h3aa1a7de),
	.w7(32'hbc59463e),
	.w8(32'h3c8c60fa),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c031b),
	.w1(32'hbba8b939),
	.w2(32'h3c8565a1),
	.w3(32'hbc06c309),
	.w4(32'hbb459b1e),
	.w5(32'h3a8b73bd),
	.w6(32'h3ab89cc5),
	.w7(32'hbac6bf11),
	.w8(32'h3c3af360),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc633073),
	.w1(32'hb943d2e2),
	.w2(32'hbb83fa9c),
	.w3(32'hbb886b13),
	.w4(32'hbc114884),
	.w5(32'hbbf22740),
	.w6(32'hbbfac754),
	.w7(32'hbc7d240a),
	.w8(32'hbbcc67e2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19689f),
	.w1(32'hbb2229f8),
	.w2(32'hbc3654af),
	.w3(32'h3b4dd2c5),
	.w4(32'h3b68587d),
	.w5(32'hbc502302),
	.w6(32'h3c566f97),
	.w7(32'h3b86bbb9),
	.w8(32'h3c13f5b0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d91de),
	.w1(32'h3a990af6),
	.w2(32'hbbb6b050),
	.w3(32'h3c442f3a),
	.w4(32'hbaa08d7e),
	.w5(32'h3b373113),
	.w6(32'hb9dbe450),
	.w7(32'hbc142f84),
	.w8(32'hb9f295d5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18911a),
	.w1(32'h394baf65),
	.w2(32'hbc27839e),
	.w3(32'hbb782da8),
	.w4(32'h3c8f9031),
	.w5(32'hbc185de0),
	.w6(32'h3c0a1a29),
	.w7(32'h3a832dc4),
	.w8(32'h3c4b2697),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56f92a),
	.w1(32'h3bc3debc),
	.w2(32'h3cfa7fc4),
	.w3(32'h3bb78e4f),
	.w4(32'hbbe4a93f),
	.w5(32'hbc6af8b2),
	.w6(32'h3bf553b2),
	.w7(32'hbc0c28a6),
	.w8(32'hbb4ede65),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cd1a7),
	.w1(32'hbbe0bc19),
	.w2(32'h3d087e07),
	.w3(32'hbbfef4cd),
	.w4(32'hbc8c7b52),
	.w5(32'h3a56687f),
	.w6(32'h3b924431),
	.w7(32'hbbaf762d),
	.w8(32'hbab6ecaa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb111d3d),
	.w1(32'hbc2c2f33),
	.w2(32'h3bc44445),
	.w3(32'h3bcb93ee),
	.w4(32'h3b6961e7),
	.w5(32'h3b460246),
	.w6(32'hbba17acf),
	.w7(32'h3b86c775),
	.w8(32'h3b957762),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18fda9),
	.w1(32'hbb92e3d2),
	.w2(32'hbb2832eb),
	.w3(32'h3c03e6ac),
	.w4(32'hbbf69633),
	.w5(32'hbbb13252),
	.w6(32'h3be32833),
	.w7(32'hba41643f),
	.w8(32'hb9a61c0b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7a167),
	.w1(32'h3b4f1538),
	.w2(32'hba9e3554),
	.w3(32'h3b5aec93),
	.w4(32'h3ae52aca),
	.w5(32'h3c865bcf),
	.w6(32'h3a42576c),
	.w7(32'hbaf2d6da),
	.w8(32'hbd21e06c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29b611),
	.w1(32'hbc1dc574),
	.w2(32'hbbd99ba0),
	.w3(32'hbb5a54d6),
	.w4(32'hbc0b5b3e),
	.w5(32'h3c1a8675),
	.w6(32'h3b960dd0),
	.w7(32'h3ba6160f),
	.w8(32'hbc39922a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf9b21),
	.w1(32'h3c956280),
	.w2(32'hbb383539),
	.w3(32'h3bd28c3a),
	.w4(32'h3a832d53),
	.w5(32'hbc3a218f),
	.w6(32'hbbac7d25),
	.w7(32'hbcae74ed),
	.w8(32'hbc312326),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6a938),
	.w1(32'hbba81149),
	.w2(32'h394cf9d8),
	.w3(32'hbc115218),
	.w4(32'hbc077b2a),
	.w5(32'hbd2744c8),
	.w6(32'hbad6420d),
	.w7(32'h3c0091de),
	.w8(32'hbab72975),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcd5e5),
	.w1(32'hbc2ce8a7),
	.w2(32'hba4c3a18),
	.w3(32'hbc257677),
	.w4(32'h3b04475d),
	.w5(32'hbc1e2fcd),
	.w6(32'h392a5e4d),
	.w7(32'hbb6a9c4b),
	.w8(32'hbacbbd22),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab43eb0),
	.w1(32'h3b4f8372),
	.w2(32'h3cf17dfe),
	.w3(32'h3cf48804),
	.w4(32'h3c2a965a),
	.w5(32'h3bef4e4f),
	.w6(32'h3bf3e55a),
	.w7(32'hbc673d2b),
	.w8(32'hbad999ed),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22bf5a),
	.w1(32'h3bb0e31f),
	.w2(32'h3c57ece6),
	.w3(32'h3a3ee0cd),
	.w4(32'h3bec97c3),
	.w5(32'h3c664762),
	.w6(32'h3c1459c2),
	.w7(32'h3b31290b),
	.w8(32'hbbaa55fa),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91c54b),
	.w1(32'h3c5419a4),
	.w2(32'h3c261d98),
	.w3(32'h3add5bca),
	.w4(32'h3b9f75c4),
	.w5(32'hbbd2000c),
	.w6(32'h3b3c15d7),
	.w7(32'h39560bc5),
	.w8(32'hbb0be5b7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2becd2),
	.w1(32'h3c9eefd0),
	.w2(32'hbbca1f08),
	.w3(32'h3b9fe833),
	.w4(32'h3c1dd283),
	.w5(32'h3b089f37),
	.w6(32'hbc8088ce),
	.w7(32'h3ca2137c),
	.w8(32'h3c6c6065),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab08951),
	.w1(32'h3c4ef7cb),
	.w2(32'hbb4e224a),
	.w3(32'h3c5d1927),
	.w4(32'hbb3c1781),
	.w5(32'h3c82d078),
	.w6(32'h3ace3748),
	.w7(32'hbc28d947),
	.w8(32'h3d2629d4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c006339),
	.w1(32'hbbb5e277),
	.w2(32'hbbe8e597),
	.w3(32'hbbf16679),
	.w4(32'hbc2d5849),
	.w5(32'hbacba02a),
	.w6(32'h3ce2a332),
	.w7(32'hbbefc47a),
	.w8(32'hbbd22848),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0532ce),
	.w1(32'hbad56269),
	.w2(32'hbafdec6d),
	.w3(32'hbbe24394),
	.w4(32'hbc7602d5),
	.w5(32'hbb85d0b4),
	.w6(32'h3a875848),
	.w7(32'hbc9652f0),
	.w8(32'hba808b6a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cc202),
	.w1(32'hbaa3d54e),
	.w2(32'h3b179ab0),
	.w3(32'h3bc71129),
	.w4(32'hbc5e771c),
	.w5(32'h3c45b9e9),
	.w6(32'hbc6c9c13),
	.w7(32'h3b3cf73e),
	.w8(32'hba4686ec),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b13e1),
	.w1(32'h3a10c380),
	.w2(32'h3bb9b49a),
	.w3(32'h3b2b7ba5),
	.w4(32'h3942f144),
	.w5(32'h3bb55e55),
	.w6(32'h3d401765),
	.w7(32'hbbaa2633),
	.w8(32'hbce131a9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fc7e4),
	.w1(32'h3a532b36),
	.w2(32'h3c301ae4),
	.w3(32'hba3b834a),
	.w4(32'hbd3badb6),
	.w5(32'h3aef1dd5),
	.w6(32'h3b8552ad),
	.w7(32'hbb55cbf9),
	.w8(32'hbd080bcf),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad9354),
	.w1(32'hbd2a7dae),
	.w2(32'hbc49af9c),
	.w3(32'h3adf46b9),
	.w4(32'h3c7d492c),
	.w5(32'h3b5508f9),
	.w6(32'hbb6f2280),
	.w7(32'h3bb57c27),
	.w8(32'hbb4ab9d0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb235311),
	.w1(32'hbadcca32),
	.w2(32'h3bea2c9a),
	.w3(32'hbb37792f),
	.w4(32'h3bb48623),
	.w5(32'hbb8142e0),
	.w6(32'hbb1740d2),
	.w7(32'hbb825643),
	.w8(32'hba979011),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b7f8d),
	.w1(32'h3afa56c6),
	.w2(32'hbbf763a9),
	.w3(32'hbc12d06d),
	.w4(32'h3ac1f1c1),
	.w5(32'hbb8cd245),
	.w6(32'h3c09fec3),
	.w7(32'h3c060360),
	.w8(32'h3bd3e24e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e6ce),
	.w1(32'h3c07dc09),
	.w2(32'hba0b9a53),
	.w3(32'h3b3d23f5),
	.w4(32'hbbb5ba11),
	.w5(32'hbbcbe837),
	.w6(32'h3bd0df71),
	.w7(32'h3ac7fdf3),
	.w8(32'h3a1d4191),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a266823),
	.w1(32'hbb33c9d2),
	.w2(32'h3b27a506),
	.w3(32'h3b9dfc7d),
	.w4(32'hbb9951fc),
	.w5(32'hbc6ac5a6),
	.w6(32'hbb522134),
	.w7(32'h3b9bff40),
	.w8(32'h3b0954b4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b550c6e),
	.w1(32'h3ae2c3e5),
	.w2(32'h3bba8615),
	.w3(32'h3c58f263),
	.w4(32'hbbea4644),
	.w5(32'h3a770f60),
	.w6(32'h3c6839ca),
	.w7(32'hbcb5c7cd),
	.w8(32'hbba34fee),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7a6fb),
	.w1(32'h3c73784d),
	.w2(32'hbaff7cc2),
	.w3(32'hbbcc30d0),
	.w4(32'hbad4610e),
	.w5(32'h3c540bf9),
	.w6(32'h3cb68c22),
	.w7(32'h3894406e),
	.w8(32'hbbf9255e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2848dd),
	.w1(32'hbb58b26e),
	.w2(32'hbc4aefa2),
	.w3(32'h3c0ee996),
	.w4(32'h3bc0c217),
	.w5(32'hbb256656),
	.w6(32'h3c00b45a),
	.w7(32'h3b606aca),
	.w8(32'h3a9adcfa),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f4f78),
	.w1(32'hbac49bbf),
	.w2(32'hbb752086),
	.w3(32'hbc61f810),
	.w4(32'h3b256612),
	.w5(32'hb9e080e8),
	.w6(32'h3bcacd52),
	.w7(32'h3b025c8d),
	.w8(32'h3ca4fcd1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb908d5d),
	.w1(32'hbb869942),
	.w2(32'h3aaa4888),
	.w3(32'h3b8a5338),
	.w4(32'h3b501855),
	.w5(32'h3a1c9da1),
	.w6(32'h3c16e45c),
	.w7(32'hbb794372),
	.w8(32'hbae120e2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c211090),
	.w1(32'hbc22075b),
	.w2(32'hbd037d17),
	.w3(32'hbc3bcd2d),
	.w4(32'hbd0ad67b),
	.w5(32'hbc4cf51d),
	.w6(32'hbd9c36fe),
	.w7(32'h3b0e6ddc),
	.w8(32'h3ab38e0e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80aea8),
	.w1(32'hbb8d234a),
	.w2(32'hbc0f59cf),
	.w3(32'hbc7e1997),
	.w4(32'hbb1e6639),
	.w5(32'h3b8d8204),
	.w6(32'hbc8d4fd5),
	.w7(32'hbb4145b7),
	.w8(32'hbacdaa69),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48eae2),
	.w1(32'h3c977a89),
	.w2(32'hbaf20ac3),
	.w3(32'hba9c30fd),
	.w4(32'h3b7d317b),
	.w5(32'hb93dab80),
	.w6(32'hbb58621d),
	.w7(32'hb9ff601b),
	.w8(32'h3ac12276),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca33fa),
	.w1(32'h3b943c69),
	.w2(32'h3a21ef6c),
	.w3(32'hbc71d5a6),
	.w4(32'h3b884b32),
	.w5(32'hbb81fcac),
	.w6(32'h3bc4effb),
	.w7(32'hba49b00c),
	.w8(32'hba373284),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2d5d7),
	.w1(32'hbbec25f3),
	.w2(32'h3c459a59),
	.w3(32'hb9c0152d),
	.w4(32'hbb78f15e),
	.w5(32'h3c0ff36c),
	.w6(32'h3b9ce0ed),
	.w7(32'h3ce997d7),
	.w8(32'hba2bba36),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e585),
	.w1(32'hbb1129c5),
	.w2(32'hbb3d4ce4),
	.w3(32'hbb2ee1ab),
	.w4(32'hbbd9928a),
	.w5(32'hbc190a2d),
	.w6(32'h3b08cf9a),
	.w7(32'hbbf6f050),
	.w8(32'hbab527e2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd235a6),
	.w1(32'h3ba04f43),
	.w2(32'h3b877faa),
	.w3(32'hbb1160dd),
	.w4(32'hbc56dc07),
	.w5(32'h3b9abc5d),
	.w6(32'hbd6f3110),
	.w7(32'h3aebb37a),
	.w8(32'hbba8c163),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc07c8),
	.w1(32'h3aa2fb1c),
	.w2(32'h3c6871c2),
	.w3(32'hbb6be0d5),
	.w4(32'h3c2479b0),
	.w5(32'hbc51bba9),
	.w6(32'h3b118a65),
	.w7(32'hbb9c1545),
	.w8(32'hbbe6fc03),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e50df),
	.w1(32'h39708551),
	.w2(32'h3b066845),
	.w3(32'hbc3dc894),
	.w4(32'hbb18eaa6),
	.w5(32'h3b263baf),
	.w6(32'hbc7ddd04),
	.w7(32'hbc797232),
	.w8(32'hb8fa9c59),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55b35f),
	.w1(32'hbb1ab49f),
	.w2(32'h3b827400),
	.w3(32'h39161477),
	.w4(32'hbac36726),
	.w5(32'h3b828046),
	.w6(32'hba96dedd),
	.w7(32'h39e99869),
	.w8(32'h3c7cd4e6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3983c),
	.w1(32'h3bb64680),
	.w2(32'hbab6f3f1),
	.w3(32'hbbf84862),
	.w4(32'h3c38620a),
	.w5(32'hbb28488f),
	.w6(32'hbb1805b8),
	.w7(32'hbba0b214),
	.w8(32'h3b4a0591),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3efcea),
	.w1(32'h3b7bbc0f),
	.w2(32'h3b5d4f45),
	.w3(32'hbb814947),
	.w4(32'h3b5d5694),
	.w5(32'hbb8f4c8d),
	.w6(32'hbbd2a5f7),
	.w7(32'hbb43bda7),
	.w8(32'h3b28674c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b696b),
	.w1(32'hbb99fb05),
	.w2(32'hb962bc93),
	.w3(32'hbbc4cb02),
	.w4(32'hbc261499),
	.w5(32'hbb221c81),
	.w6(32'h3aa32dc1),
	.w7(32'h3b9ce7b4),
	.w8(32'h3bd0c7fb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68538e),
	.w1(32'hbbf8651e),
	.w2(32'hbb572a89),
	.w3(32'hbb9541fa),
	.w4(32'h3b16e15d),
	.w5(32'hbba06db3),
	.w6(32'h3ba319ae),
	.w7(32'h3b92986e),
	.w8(32'hba480a82),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1fed1),
	.w1(32'h3b88b4c1),
	.w2(32'hba8fa703),
	.w3(32'hbaab970b),
	.w4(32'hbb78398d),
	.w5(32'h3b581936),
	.w6(32'hbb3e1ad4),
	.w7(32'h3850240e),
	.w8(32'h3c400868),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93511e),
	.w1(32'h3a445ad8),
	.w2(32'hbbbd6cf4),
	.w3(32'hbb39bf09),
	.w4(32'hbb8c2e6c),
	.w5(32'h3b7a8252),
	.w6(32'hbc3ba508),
	.w7(32'h3c37026a),
	.w8(32'hb8b429cc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85c833),
	.w1(32'h3c048775),
	.w2(32'hbc3975ab),
	.w3(32'hba79dd98),
	.w4(32'h3be30115),
	.w5(32'h3b1a2192),
	.w6(32'hbb2e7a25),
	.w7(32'hbbc4648f),
	.w8(32'h3c1caca8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a2a0b),
	.w1(32'hbb239a33),
	.w2(32'hbc3854e4),
	.w3(32'h3c1102ec),
	.w4(32'hba801dbf),
	.w5(32'hb904f2f0),
	.w6(32'h38843f01),
	.w7(32'h3b3f063b),
	.w8(32'h3c7ecabe),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b032),
	.w1(32'hbc1b5574),
	.w2(32'hbbadde7f),
	.w3(32'h3c81efa6),
	.w4(32'hbba9f857),
	.w5(32'hbba69d85),
	.w6(32'h39b32c44),
	.w7(32'h3b932f9f),
	.w8(32'h3c08f42f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd167a0e),
	.w1(32'h38d681aa),
	.w2(32'h3bb56d93),
	.w3(32'h3adf0faa),
	.w4(32'hbb5bf198),
	.w5(32'h3c45f220),
	.w6(32'h3b0ba0f5),
	.w7(32'h3c031fa9),
	.w8(32'hbc7a60c9),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d3063),
	.w1(32'h38cd33af),
	.w2(32'hbb027574),
	.w3(32'hbbdc78be),
	.w4(32'h39abdfc3),
	.w5(32'hbb8aa48c),
	.w6(32'h3ad857e1),
	.w7(32'h3d82f722),
	.w8(32'hbb989575),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12f639),
	.w1(32'hbba2220d),
	.w2(32'h3c4be8de),
	.w3(32'hbac54910),
	.w4(32'h37e56af7),
	.w5(32'hbc6bd807),
	.w6(32'hbbdee2bb),
	.w7(32'hbc0b6c2f),
	.w8(32'h3bd9e0d6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56a347),
	.w1(32'hbbccff77),
	.w2(32'h3b2ca850),
	.w3(32'hbc80e23d),
	.w4(32'hbc41e3a5),
	.w5(32'h38f8432d),
	.w6(32'h3b998862),
	.w7(32'h3ccc8ece),
	.w8(32'h3c1b3fac),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34315e),
	.w1(32'hba8cfb90),
	.w2(32'h3bd30e3f),
	.w3(32'h3bad3ba4),
	.w4(32'hbb63733d),
	.w5(32'h3b29f2c5),
	.w6(32'hbc3a7dd0),
	.w7(32'hbc0fa896),
	.w8(32'hbb9d5561),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3e0ee),
	.w1(32'h3c1d0343),
	.w2(32'hbce7fad0),
	.w3(32'h3c0530d9),
	.w4(32'h3b5fb1ed),
	.w5(32'h3bc4add0),
	.w6(32'hbb5b27d4),
	.w7(32'hbbcab4ab),
	.w8(32'hbcaccbd0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5aff1),
	.w1(32'hbb35a494),
	.w2(32'hbc8e4188),
	.w3(32'h3bcfd376),
	.w4(32'h389e7daa),
	.w5(32'hbc11c51d),
	.w6(32'hbc7f470c),
	.w7(32'hba28eedd),
	.w8(32'hbaf884ed),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a8937),
	.w1(32'hbb28120e),
	.w2(32'hbbc0f6ed),
	.w3(32'h3be17406),
	.w4(32'hbbf8133c),
	.w5(32'hbadf9ad8),
	.w6(32'h3b833ec6),
	.w7(32'hbad5cfe9),
	.w8(32'hbb3f21f3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ae4d1),
	.w1(32'hbc15ec0d),
	.w2(32'hbc3c9124),
	.w3(32'hbbe7f510),
	.w4(32'hb915a0ae),
	.w5(32'hb977c846),
	.w6(32'hb9524cfe),
	.w7(32'h3c4b8b26),
	.w8(32'hbb96c6a9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5814f),
	.w1(32'h3c141ee9),
	.w2(32'h3c06e0f2),
	.w3(32'hbb9ae3cc),
	.w4(32'h3c39dd80),
	.w5(32'h3bab7a64),
	.w6(32'hbbbe6d96),
	.w7(32'h3bc4eec9),
	.w8(32'hbb95573c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc9f45),
	.w1(32'hbaea8a47),
	.w2(32'hbc9d886d),
	.w3(32'h3d0454c2),
	.w4(32'h3b4b1e6e),
	.w5(32'h3c132c75),
	.w6(32'h3c4f49fa),
	.w7(32'h39ecaa48),
	.w8(32'h3a2bf2ca),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c2ba6),
	.w1(32'h3bbdeb01),
	.w2(32'h3adef10b),
	.w3(32'h3c0bd08a),
	.w4(32'hbb4d50d2),
	.w5(32'hbb7b73fe),
	.w6(32'hbbe3b620),
	.w7(32'h3b2a7ad0),
	.w8(32'hbc862ecb),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44c499),
	.w1(32'h3c3dbff7),
	.w2(32'hbafd4e39),
	.w3(32'hbbd51e4d),
	.w4(32'hb8d6c77b),
	.w5(32'hbc023c5a),
	.w6(32'hba0c1aab),
	.w7(32'hbd231a5e),
	.w8(32'h3bb9ce83),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d98d1),
	.w1(32'hbba142a6),
	.w2(32'hbbf9596f),
	.w3(32'h39374bac),
	.w4(32'hbc04c16e),
	.w5(32'hbbcbebdd),
	.w6(32'h3affb317),
	.w7(32'hbb6ba6b7),
	.w8(32'h3c277f13),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c4486),
	.w1(32'hbbad22d0),
	.w2(32'h3958281e),
	.w3(32'hbc2d5b80),
	.w4(32'hbb82a86c),
	.w5(32'hb9c0602b),
	.w6(32'h3d03f9d7),
	.w7(32'hbb41064d),
	.w8(32'h3b909a0d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb979c0f8),
	.w1(32'hba33f065),
	.w2(32'h3c9bdf65),
	.w3(32'h3c02309c),
	.w4(32'hbc426d24),
	.w5(32'hbc81fc77),
	.w6(32'h3c8a6637),
	.w7(32'hba86e229),
	.w8(32'h3b65445a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62e690),
	.w1(32'hbb85d7bb),
	.w2(32'h3aa23b4c),
	.w3(32'hbcf6acc7),
	.w4(32'hb9f5841a),
	.w5(32'h3b27a661),
	.w6(32'h3c3630c8),
	.w7(32'hb95d1771),
	.w8(32'h3baf390a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e64cd),
	.w1(32'hbcc41c21),
	.w2(32'hbc0fc870),
	.w3(32'h3c594617),
	.w4(32'hbc2998e5),
	.w5(32'hbb67a77b),
	.w6(32'hbc0b803f),
	.w7(32'h3baab8b8),
	.w8(32'h3b680993),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ed2dd),
	.w1(32'h3b7179ab),
	.w2(32'h3a8587b4),
	.w3(32'hbb086bb7),
	.w4(32'h3a657e0f),
	.w5(32'hbb21df1f),
	.w6(32'hb713493e),
	.w7(32'h3c12020c),
	.w8(32'hba86ce4e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376e2946),
	.w1(32'h3c8fb754),
	.w2(32'hbae02360),
	.w3(32'hbbd5a67c),
	.w4(32'hbc20b301),
	.w5(32'h3ac7b31a),
	.w6(32'h3bb7e44e),
	.w7(32'h3ba56153),
	.w8(32'h3b973f84),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb369f49),
	.w1(32'h3c04fa19),
	.w2(32'h3c0946a2),
	.w3(32'h3ca7f93b),
	.w4(32'h3a6755fe),
	.w5(32'h3bc9ef6d),
	.w6(32'hbca44cb8),
	.w7(32'hbb00d221),
	.w8(32'h397ac5b9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21929d),
	.w1(32'hbaafbb48),
	.w2(32'hbc827d12),
	.w3(32'h3c4f259e),
	.w4(32'h3ba9e17d),
	.w5(32'h3c1d6609),
	.w6(32'h3ad050b7),
	.w7(32'hbc78978e),
	.w8(32'h3b16de0e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aa6f0),
	.w1(32'h3c01c8a4),
	.w2(32'h3b29cd65),
	.w3(32'h3c5307ad),
	.w4(32'h3a9f3099),
	.w5(32'h3b89d289),
	.w6(32'hbb245e55),
	.w7(32'hba9fd2b6),
	.w8(32'hbac1eea3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77bd1e),
	.w1(32'hbc47db1b),
	.w2(32'h38c00c45),
	.w3(32'hbb3d70a2),
	.w4(32'hbb8d7d44),
	.w5(32'hbb10f490),
	.w6(32'hba624c40),
	.w7(32'hbbdc24d9),
	.w8(32'hbb4f034a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18f3e0),
	.w1(32'hbbd15173),
	.w2(32'hbb00be3e),
	.w3(32'h3ad9a855),
	.w4(32'hbc62c822),
	.w5(32'h3baf3797),
	.w6(32'h3be4b922),
	.w7(32'hbb97f757),
	.w8(32'hbbcf597f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16f0b6),
	.w1(32'h3c5a5195),
	.w2(32'hbbb5c883),
	.w3(32'h3a727ef4),
	.w4(32'hbb3d7526),
	.w5(32'hbb02d296),
	.w6(32'hbb4b4aef),
	.w7(32'h3b587fe9),
	.w8(32'h3c75012a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25b89e),
	.w1(32'hbb942f71),
	.w2(32'h3b68daa7),
	.w3(32'hbdc52bfc),
	.w4(32'h3c618ccf),
	.w5(32'h3c0b7ce2),
	.w6(32'h3b17f0a6),
	.w7(32'hbb8d09e4),
	.w8(32'hbb37234f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf89891),
	.w1(32'hbcd2cd4d),
	.w2(32'h3b8b3081),
	.w3(32'hbae33538),
	.w4(32'hba4ae03d),
	.w5(32'h3b8e8dd5),
	.w6(32'hbb1fffb0),
	.w7(32'h3b98af02),
	.w8(32'h3ae6c83b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812c0e),
	.w1(32'h3b8aedc6),
	.w2(32'h3bf51742),
	.w3(32'h3ba68ad6),
	.w4(32'h3c2ee7ed),
	.w5(32'hbb997791),
	.w6(32'hbc2fad91),
	.w7(32'h3c930550),
	.w8(32'hbbc63170),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2ce89),
	.w1(32'h3c4dd944),
	.w2(32'hba509a1c),
	.w3(32'h3b5b3bbd),
	.w4(32'h3b55e7f2),
	.w5(32'h3c015aa4),
	.w6(32'h3bb1326c),
	.w7(32'h3c3c00a3),
	.w8(32'h3a6bd7a1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d7af2),
	.w1(32'hbbeceffb),
	.w2(32'h39623225),
	.w3(32'h39819d70),
	.w4(32'hbba1f34c),
	.w5(32'hbb96e254),
	.w6(32'hb9c43a34),
	.w7(32'hbb6b2d22),
	.w8(32'h3c1d1a30),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96620f),
	.w1(32'h3b9c4e70),
	.w2(32'hbbe8c268),
	.w3(32'hbbe5f636),
	.w4(32'h3bb183d1),
	.w5(32'hba6fd5ef),
	.w6(32'hbc4aacc6),
	.w7(32'hbc85d848),
	.w8(32'hbbfe99af),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ec884),
	.w1(32'hbbca96f1),
	.w2(32'h3b56bf94),
	.w3(32'h3b3b3dba),
	.w4(32'hbaf7cab1),
	.w5(32'h3b4cd2b1),
	.w6(32'h3b972fe7),
	.w7(32'h3b1bfc8f),
	.w8(32'h3bbef58e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf703f6),
	.w1(32'hbabe4064),
	.w2(32'h3b8d5b9d),
	.w3(32'hbcd81c95),
	.w4(32'hbc804404),
	.w5(32'hbc35368d),
	.w6(32'hbba68722),
	.w7(32'hbba17c1b),
	.w8(32'hbaabceb7),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c95be),
	.w1(32'h3bd3c453),
	.w2(32'hbcb76372),
	.w3(32'h3cd4ae73),
	.w4(32'hbb848f93),
	.w5(32'h3b6b0bd6),
	.w6(32'hbb8a44fc),
	.w7(32'hbc0eab23),
	.w8(32'h3b6639a5),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bbaa6),
	.w1(32'hbae6c418),
	.w2(32'hbb9238fe),
	.w3(32'h3b779194),
	.w4(32'h3c121af3),
	.w5(32'hbb03cfcb),
	.w6(32'hbbd52991),
	.w7(32'hbb501054),
	.w8(32'h3cda70f2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeaade),
	.w1(32'hbbb9b2d6),
	.w2(32'hba442999),
	.w3(32'hbc2695f7),
	.w4(32'h3b930416),
	.w5(32'h3ccd9cc3),
	.w6(32'hbb5bdb4f),
	.w7(32'h3bdff357),
	.w8(32'hb7da8592),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ec47d),
	.w1(32'h3afdb026),
	.w2(32'hba346019),
	.w3(32'hbb1d1c94),
	.w4(32'h3bfed0ea),
	.w5(32'hbc3723e0),
	.w6(32'hbb2e32a4),
	.w7(32'h3b6e4ff3),
	.w8(32'h3b0b16df),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d6fc9),
	.w1(32'hbc817531),
	.w2(32'h3c4dde80),
	.w3(32'h3da238e7),
	.w4(32'h3cb9c262),
	.w5(32'hbbca930e),
	.w6(32'hba17ce32),
	.w7(32'hbd4e07fc),
	.w8(32'hb99310bf),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a9cd3),
	.w1(32'hbb4cedd8),
	.w2(32'h3b02e243),
	.w3(32'hbc46314e),
	.w4(32'hbad81033),
	.w5(32'hbae353f3),
	.w6(32'hba9da07d),
	.w7(32'hbb086a5e),
	.w8(32'h3bd8901b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ae0c3),
	.w1(32'h3ba01a1d),
	.w2(32'h3bae904c),
	.w3(32'hb9d46e0e),
	.w4(32'hbac3e8ea),
	.w5(32'h3b1d3840),
	.w6(32'h3c4df2f7),
	.w7(32'h3afe4132),
	.w8(32'hbaeef559),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4b517c),
	.w1(32'hbb34360c),
	.w2(32'hba5fa4c3),
	.w3(32'h3ba5c033),
	.w4(32'h3beaf988),
	.w5(32'hbbc410cb),
	.w6(32'h3c9ed40f),
	.w7(32'h3a5bdc70),
	.w8(32'hbd18a001),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bf11c),
	.w1(32'h3b9a33b6),
	.w2(32'h3cd1105f),
	.w3(32'h3bb70947),
	.w4(32'hbd3486f7),
	.w5(32'h3c54fd3d),
	.w6(32'hbba1fceb),
	.w7(32'hbb9318f9),
	.w8(32'hbc1172e8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba457fb4),
	.w1(32'hbad95d1e),
	.w2(32'hbb2a0427),
	.w3(32'h3c50ef92),
	.w4(32'hb9737be6),
	.w5(32'h3b53f470),
	.w6(32'h3c0a211e),
	.w7(32'hbaf2a92e),
	.w8(32'hbc01ec8d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb152d8a),
	.w1(32'h3c2d1499),
	.w2(32'h3b02edf8),
	.w3(32'h3cfaf8fe),
	.w4(32'h3b6d21d3),
	.w5(32'hbae15c91),
	.w6(32'hbc35239d),
	.w7(32'hbc87258a),
	.w8(32'h3bbcc018),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40cd4d),
	.w1(32'h3b6079bd),
	.w2(32'hbc7a262b),
	.w3(32'hbb995bb2),
	.w4(32'h3b85b1b9),
	.w5(32'hbcdf5b06),
	.w6(32'hba6a52ab),
	.w7(32'h3a0ca0dc),
	.w8(32'h3b28e91c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb931752),
	.w1(32'hbb1c7539),
	.w2(32'h3b852ed9),
	.w3(32'hbbc88cc3),
	.w4(32'h3c874598),
	.w5(32'hbb4e89a7),
	.w6(32'hbbdcb936),
	.w7(32'hba2983e1),
	.w8(32'hbbb2cc54),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95b5bd),
	.w1(32'h3b558c41),
	.w2(32'hbc174410),
	.w3(32'hbb6b71c8),
	.w4(32'h39ee6764),
	.w5(32'h3c1f3e68),
	.w6(32'h3bdf0834),
	.w7(32'h3b6dba13),
	.w8(32'hbc5bc73f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99024f),
	.w1(32'hbc43d340),
	.w2(32'h378deff5),
	.w3(32'h3c34df44),
	.w4(32'h3aea402b),
	.w5(32'hb8a35978),
	.w6(32'h3bd4f708),
	.w7(32'hbb371f30),
	.w8(32'h3b672c56),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea6423),
	.w1(32'h3a989bba),
	.w2(32'hbc23187d),
	.w3(32'hbc190db8),
	.w4(32'h3c56d300),
	.w5(32'hbc295e7e),
	.w6(32'hb9d9e410),
	.w7(32'hbccfdfcb),
	.w8(32'h3b50c2c4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2a709),
	.w1(32'hb93f25a7),
	.w2(32'h3c0eeefd),
	.w3(32'h3bba08bb),
	.w4(32'hbc4e131c),
	.w5(32'h3c141c66),
	.w6(32'h3bcf25fb),
	.w7(32'h3a6221c7),
	.w8(32'h3aa266b5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91dbcb),
	.w1(32'h3bddcaea),
	.w2(32'hbaaa2386),
	.w3(32'hbbc89b54),
	.w4(32'hbd653479),
	.w5(32'hbab3ffb2),
	.w6(32'h3b69a247),
	.w7(32'h3a1fbb10),
	.w8(32'hbba40b67),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06fe60),
	.w1(32'hb99c66b1),
	.w2(32'h3c8d3146),
	.w3(32'h3b0b9957),
	.w4(32'h3c4eba9b),
	.w5(32'h3bf578a3),
	.w6(32'hbae4d82e),
	.w7(32'hbbbcdfe4),
	.w8(32'h3da42997),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22aa00),
	.w1(32'h3adac289),
	.w2(32'hbc0c2e18),
	.w3(32'h3b36d50e),
	.w4(32'h3bb10a37),
	.w5(32'hbdbd224e),
	.w6(32'h3c24083b),
	.w7(32'hbb4f6d64),
	.w8(32'h3856de12),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a735d),
	.w1(32'h3becb4eb),
	.w2(32'hbbbca8bc),
	.w3(32'h3b49a0b2),
	.w4(32'hbb65bebc),
	.w5(32'h3b04d09b),
	.w6(32'h3b17090a),
	.w7(32'hbd303d8d),
	.w8(32'hbb93e067),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92b178),
	.w1(32'h3ba2c8c9),
	.w2(32'h3b8b23d4),
	.w3(32'hbb046b1d),
	.w4(32'h38b1e238),
	.w5(32'h3b73f4dd),
	.w6(32'hbc446c71),
	.w7(32'h38d37b3b),
	.w8(32'h3aa9eedb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2213cf),
	.w1(32'h3b31d409),
	.w2(32'h39a560c4),
	.w3(32'hb9a2b919),
	.w4(32'hb99dcb5f),
	.w5(32'h3b7f6e42),
	.w6(32'h3b482a84),
	.w7(32'h3b82cb38),
	.w8(32'hbd0aa3a3),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ae347),
	.w1(32'h3c06a327),
	.w2(32'hbce7f409),
	.w3(32'h3c50e5bc),
	.w4(32'hbb7c8036),
	.w5(32'hbad440b5),
	.w6(32'h3acbe5dd),
	.w7(32'h3addae1c),
	.w8(32'hbc51a014),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84016d),
	.w1(32'h3a918770),
	.w2(32'hbb08f3b5),
	.w3(32'h3b095d8c),
	.w4(32'h3c0fc363),
	.w5(32'hbc01f73e),
	.w6(32'h3b1de295),
	.w7(32'h3919707c),
	.w8(32'h3c7a4524),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9634e),
	.w1(32'hb90477fa),
	.w2(32'h3cb23522),
	.w3(32'hbaae9292),
	.w4(32'h3c268502),
	.w5(32'h3aa97565),
	.w6(32'hbb3ddd60),
	.w7(32'h3b899d6f),
	.w8(32'h3b8fe10c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96311f),
	.w1(32'h3b47e025),
	.w2(32'h3c18b5ae),
	.w3(32'h38e711c6),
	.w4(32'h3d02d677),
	.w5(32'hbbdd3834),
	.w6(32'h3bd07dae),
	.w7(32'h3b057a15),
	.w8(32'h3aeff098),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c503719),
	.w1(32'h3b8a151f),
	.w2(32'h3ade6bec),
	.w3(32'h3b6a027b),
	.w4(32'hbc2ff830),
	.w5(32'hbbeae32b),
	.w6(32'hbaab72ad),
	.w7(32'h3d0abf77),
	.w8(32'hbbf7c222),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b4ea9),
	.w1(32'hbb934048),
	.w2(32'h3bd11f9c),
	.w3(32'h3ba03d3d),
	.w4(32'hbc33088d),
	.w5(32'hbc8be985),
	.w6(32'hbc30e72d),
	.w7(32'hbbce0b01),
	.w8(32'hbb576db9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c1b37),
	.w1(32'h3bd3c934),
	.w2(32'h3c0c82cc),
	.w3(32'h3c0e202f),
	.w4(32'hbc2d69fc),
	.w5(32'hbbacbb0f),
	.w6(32'h3b58a957),
	.w7(32'hbac744e8),
	.w8(32'h3a3bfcdc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda86e0),
	.w1(32'h3b1229ed),
	.w2(32'h3af36c64),
	.w3(32'h3b2a5ba9),
	.w4(32'h3c198514),
	.w5(32'h3ba25799),
	.w6(32'hbb3d888e),
	.w7(32'hbbd66085),
	.w8(32'h3b30032d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0acb9c),
	.w1(32'h3b4a5ed4),
	.w2(32'h3ab05cc8),
	.w3(32'hba83d6b6),
	.w4(32'hbaf01abf),
	.w5(32'h3bbbe510),
	.w6(32'h3b42701f),
	.w7(32'hbaa8b607),
	.w8(32'h3be6f4c9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f4b0f),
	.w1(32'hbbe87760),
	.w2(32'h3b1bae22),
	.w3(32'hbc1f2b06),
	.w4(32'hbbcff46e),
	.w5(32'hbc5241f3),
	.w6(32'hbbfbd7fb),
	.w7(32'h3c459177),
	.w8(32'h3c72eae2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90676d),
	.w1(32'hbb4624bc),
	.w2(32'h39e14e2f),
	.w3(32'h3a62ffa8),
	.w4(32'h3a5cfdef),
	.w5(32'hbc952a84),
	.w6(32'hb9b367b0),
	.w7(32'h3c01877d),
	.w8(32'h3b57300e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1382ec),
	.w1(32'h3b43c805),
	.w2(32'h3c56dcd6),
	.w3(32'hbaff7c80),
	.w4(32'hbc136cbb),
	.w5(32'h3a3f4b31),
	.w6(32'hb8cbf173),
	.w7(32'h3a5e6b1d),
	.w8(32'hba95b922),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3c7b2),
	.w1(32'h3b7aa635),
	.w2(32'h3a503a7a),
	.w3(32'hbc21b072),
	.w4(32'hbdbf1ea8),
	.w5(32'hbbd7a773),
	.w6(32'hbb137d6d),
	.w7(32'h3a32df7b),
	.w8(32'h3c1a25ad),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a696a45),
	.w1(32'hbc0ab39a),
	.w2(32'h3b4c9781),
	.w3(32'h3ae1a3dd),
	.w4(32'h397e0692),
	.w5(32'h3a5c3ad4),
	.w6(32'hbbb7f026),
	.w7(32'h3c44fa5e),
	.w8(32'h3d0d6baa),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c781cf1),
	.w1(32'hbb9d8352),
	.w2(32'h3add47fd),
	.w3(32'h3c806818),
	.w4(32'h3bb9c24b),
	.w5(32'hb9543493),
	.w6(32'hbacd9a18),
	.w7(32'h3ca8a339),
	.w8(32'hbc3dbad7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb44bc),
	.w1(32'hbc8966f6),
	.w2(32'hbb6b1ca3),
	.w3(32'h3c1796f7),
	.w4(32'hbb254161),
	.w5(32'hbae4a506),
	.w6(32'h3a68689f),
	.w7(32'h3c086420),
	.w8(32'hbc2d9cb7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb578c05),
	.w1(32'h3b50826b),
	.w2(32'h3b8d0fcb),
	.w3(32'hbbab2e4f),
	.w4(32'h3bc1490b),
	.w5(32'hbbd1859f),
	.w6(32'hbada0453),
	.w7(32'h3982653d),
	.w8(32'hba42f708),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e5c80),
	.w1(32'h3b74cb89),
	.w2(32'hbb2eb006),
	.w3(32'hbbc229bb),
	.w4(32'hbb19b7f5),
	.w5(32'hbd0343d7),
	.w6(32'h3b11136d),
	.w7(32'hbc35d0f4),
	.w8(32'h3bd06be7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe30ac1),
	.w1(32'h3ab0a97b),
	.w2(32'hbb48cb5e),
	.w3(32'h3b5af75a),
	.w4(32'h3badf1f3),
	.w5(32'h3b78a9ce),
	.w6(32'h3b7e6274),
	.w7(32'hba6fd9c7),
	.w8(32'h3a0af016),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27a5b9),
	.w1(32'hbb467288),
	.w2(32'hbb4de5c7),
	.w3(32'hbc73d27d),
	.w4(32'h39b113e5),
	.w5(32'hbb00eeea),
	.w6(32'hbde1848b),
	.w7(32'hbcc9e061),
	.w8(32'hbb54cba4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8838844),
	.w1(32'h3b637d83),
	.w2(32'h3b6d2471),
	.w3(32'hbc577e4a),
	.w4(32'hbba9e97a),
	.w5(32'hba74c14b),
	.w6(32'h3b8c6bbb),
	.w7(32'hbb21ea77),
	.w8(32'h3bf84e1d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6eea92),
	.w1(32'hbb5a7b98),
	.w2(32'h3bdb26b8),
	.w3(32'h3c3c186f),
	.w4(32'hbd105fd0),
	.w5(32'h3b2b24d2),
	.w6(32'h3c00a39b),
	.w7(32'hb8c01065),
	.w8(32'hbb873bf5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfd0e1),
	.w1(32'h3a8b28ee),
	.w2(32'h3b850d3d),
	.w3(32'h3c7901e9),
	.w4(32'h3b274ae4),
	.w5(32'h3ba01ef8),
	.w6(32'h3b18e1a0),
	.w7(32'hbb8e54c2),
	.w8(32'hbcc9978e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00cd41),
	.w1(32'hbb7c9b7c),
	.w2(32'hbb3148db),
	.w3(32'h3aad5a24),
	.w4(32'h3b0b9c89),
	.w5(32'hbc1c06f3),
	.w6(32'hbb8dfbe4),
	.w7(32'hb9e72c52),
	.w8(32'hbba68d20),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a7310),
	.w1(32'h3c2f362b),
	.w2(32'hbbd771a0),
	.w3(32'hbbecd654),
	.w4(32'h3aee8291),
	.w5(32'h3b1b248f),
	.w6(32'h3b60e20a),
	.w7(32'hbaca0d1e),
	.w8(32'hbb147f80),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule