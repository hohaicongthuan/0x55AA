module layer_8_featuremap_114(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb81e),
	.w1(32'hbb5d4ea7),
	.w2(32'h3c25c632),
	.w3(32'hbba588e7),
	.w4(32'h3c1ceb9e),
	.w5(32'h3bf2bd19),
	.w6(32'hbb710cb1),
	.w7(32'h3a865fe3),
	.w8(32'hbc027b99),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb632cf),
	.w1(32'h3ba3c2f5),
	.w2(32'h3ac3e89e),
	.w3(32'h3c261818),
	.w4(32'hba373b6b),
	.w5(32'hba8b1262),
	.w6(32'hbb349aa8),
	.w7(32'hbb0edcb7),
	.w8(32'hbb71fea2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89c98a),
	.w1(32'hba6a06b0),
	.w2(32'h3a620355),
	.w3(32'h3a87e7e0),
	.w4(32'hb9bd9d96),
	.w5(32'h3af91c61),
	.w6(32'hbb9e11e2),
	.w7(32'hbbea4dfb),
	.w8(32'hba8de695),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba585557),
	.w1(32'hba87c621),
	.w2(32'hbbbec7a2),
	.w3(32'h3822c079),
	.w4(32'hbbd114e6),
	.w5(32'hbb5ae9c9),
	.w6(32'h3b7fec15),
	.w7(32'h3b96c627),
	.w8(32'h3bcd76f1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b2795),
	.w1(32'hbbb80be1),
	.w2(32'h3ac5094a),
	.w3(32'hbc350cb3),
	.w4(32'h3b1ba641),
	.w5(32'hba7ca474),
	.w6(32'h3b6ef647),
	.w7(32'h3c479d06),
	.w8(32'h3aa395a6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4de0b),
	.w1(32'h3bafb519),
	.w2(32'hbb05effc),
	.w3(32'hb9d4b40a),
	.w4(32'hbbb12b7f),
	.w5(32'hbbd338c2),
	.w6(32'h394a1dcc),
	.w7(32'hbb22943d),
	.w8(32'hbbf7128a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac8017),
	.w1(32'hbbe37f46),
	.w2(32'hbbeb79a4),
	.w3(32'hbb8a8cdf),
	.w4(32'hbba90a78),
	.w5(32'hbb9cd6d4),
	.w6(32'hba6995b4),
	.w7(32'h3b84316a),
	.w8(32'h3ab5523f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d50e5),
	.w1(32'hbbc143ef),
	.w2(32'h38bdb24b),
	.w3(32'hbbb19367),
	.w4(32'hbb874f74),
	.w5(32'hbbe6fb36),
	.w6(32'h3baa3d92),
	.w7(32'h3a1c776c),
	.w8(32'h3aad6ad9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2e7f2),
	.w1(32'hbb1c0cab),
	.w2(32'hbb8503d6),
	.w3(32'hbc21aef1),
	.w4(32'hbb9192fc),
	.w5(32'hbad6dde0),
	.w6(32'hbaff2b96),
	.w7(32'hbb870726),
	.w8(32'h38f09368),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab89292),
	.w1(32'hbb0e31d3),
	.w2(32'hb9e82152),
	.w3(32'hba9786ba),
	.w4(32'hbc1ddb72),
	.w5(32'hbba4a032),
	.w6(32'hbabc76d8),
	.w7(32'h3c0cb9f0),
	.w8(32'h3bb3004e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da9a2),
	.w1(32'h3b0d3876),
	.w2(32'h3b5724ab),
	.w3(32'hbb3965ff),
	.w4(32'h3b47c9cb),
	.w5(32'h3c3004a6),
	.w6(32'h3b197f85),
	.w7(32'hbb70f278),
	.w8(32'h3b3943fc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383916d1),
	.w1(32'hba4fcf91),
	.w2(32'h3b6fa4fe),
	.w3(32'h3b88768d),
	.w4(32'hbac6f49b),
	.w5(32'hba6d71a5),
	.w6(32'h3bce09c0),
	.w7(32'hbac0195d),
	.w8(32'hbba3963c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0adca2),
	.w1(32'h3b988517),
	.w2(32'h3beb87ee),
	.w3(32'h3b47cd2f),
	.w4(32'h3aec9678),
	.w5(32'hbae7a8f1),
	.w6(32'h3b611e3c),
	.w7(32'h3c071d05),
	.w8(32'h3c0538be),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a599b78),
	.w1(32'h3b364803),
	.w2(32'h3bcff694),
	.w3(32'h3acbe85e),
	.w4(32'h3b973529),
	.w5(32'h3bb9e80b),
	.w6(32'h3c1c89ec),
	.w7(32'h3c345f0a),
	.w8(32'h3c563b2e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd12773),
	.w1(32'h3b28f690),
	.w2(32'h3b58910f),
	.w3(32'h3b06da93),
	.w4(32'h3acd388f),
	.w5(32'h3bf46115),
	.w6(32'h3be2c9d1),
	.w7(32'h3be80d04),
	.w8(32'h3c6b2d38),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c146c50),
	.w1(32'h3ba7c8e1),
	.w2(32'hbb9195e1),
	.w3(32'h3b8954f1),
	.w4(32'hbb59cff7),
	.w5(32'hbc0e8dff),
	.w6(32'h3c19c36c),
	.w7(32'hbba9a725),
	.w8(32'hbc1e157f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe4d6a),
	.w1(32'hbbeb9193),
	.w2(32'h3b8b252b),
	.w3(32'hbc08bbd3),
	.w4(32'h3c03f0cd),
	.w5(32'h3b9e595e),
	.w6(32'hbc1b0e58),
	.w7(32'h3bc13b55),
	.w8(32'h3bc66608),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a356c),
	.w1(32'h3b22adda),
	.w2(32'hbc4f194b),
	.w3(32'h3b470861),
	.w4(32'hbbf339a0),
	.w5(32'hbc2421ac),
	.w6(32'h3b5d65a0),
	.w7(32'hbc34ed38),
	.w8(32'hbc6970eb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6518d),
	.w1(32'hbca5c35f),
	.w2(32'hbad54e15),
	.w3(32'hbc777534),
	.w4(32'hbbeaa7be),
	.w5(32'hbbae7e6b),
	.w6(32'hbc67f64e),
	.w7(32'h3a1fe2f9),
	.w8(32'hbbf5252b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ab8ed),
	.w1(32'hbc04aa93),
	.w2(32'hbbaf068f),
	.w3(32'hbba1725c),
	.w4(32'hbb6b1c42),
	.w5(32'hbbc2c5f8),
	.w6(32'hbb203a7a),
	.w7(32'hb9ac7eb6),
	.w8(32'hbb39d0e5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d7c1),
	.w1(32'hbbd21459),
	.w2(32'hbb629a51),
	.w3(32'hbb963560),
	.w4(32'hba5214a3),
	.w5(32'hbc3ffe4c),
	.w6(32'hbb8ff691),
	.w7(32'h3ba8b9c0),
	.w8(32'hbc1231e8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29e8f9),
	.w1(32'hbc21d931),
	.w2(32'hbba17522),
	.w3(32'hbc14a7e1),
	.w4(32'hb9d8a9d4),
	.w5(32'hbb8df8dc),
	.w6(32'hbbdc36c6),
	.w7(32'hbb2eaf15),
	.w8(32'hbc04badc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00e319),
	.w1(32'hbc3365d0),
	.w2(32'h3a3e3a96),
	.w3(32'hbbcb30a3),
	.w4(32'hbc08c4d7),
	.w5(32'hbb25ddc6),
	.w6(32'hbb9edbc0),
	.w7(32'h3b054705),
	.w8(32'h3b064927),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39dc70),
	.w1(32'h3a2a5a11),
	.w2(32'hbc3bc13f),
	.w3(32'hbb2a40a4),
	.w4(32'hbc3a4b44),
	.w5(32'hba3a9cfa),
	.w6(32'hbaa0f462),
	.w7(32'hbc44bd54),
	.w8(32'h3a1d5488),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e92be),
	.w1(32'hbb709429),
	.w2(32'h39363025),
	.w3(32'hbb30d1b1),
	.w4(32'hbad649b5),
	.w5(32'hbb145da0),
	.w6(32'hbade9783),
	.w7(32'hba38e79e),
	.w8(32'hbb4a4123),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba100b3c),
	.w1(32'hba9575bb),
	.w2(32'hbc1bcd6f),
	.w3(32'h3b2ab538),
	.w4(32'h38c1779e),
	.w5(32'h3c0223ad),
	.w6(32'h3b70191a),
	.w7(32'h38978c71),
	.w8(32'h3bd1f724),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0867a8),
	.w1(32'hbc12f715),
	.w2(32'hba7a4f24),
	.w3(32'hbb2ccd2c),
	.w4(32'hbbb05ff4),
	.w5(32'hbb7355bd),
	.w6(32'hbb498623),
	.w7(32'hbbec8d00),
	.w8(32'hbbc5c3df),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc444634),
	.w1(32'hbca20d1a),
	.w2(32'hbb673d81),
	.w3(32'hbc61f028),
	.w4(32'hbc2e25f3),
	.w5(32'h3a38dd1f),
	.w6(32'h3ac9d7f3),
	.w7(32'h3c958de0),
	.w8(32'h3d15398c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17db56),
	.w1(32'h3c7c0d94),
	.w2(32'hbb189358),
	.w3(32'h3c02efcc),
	.w4(32'hbbc3d530),
	.w5(32'h38f03394),
	.w6(32'h3c54398e),
	.w7(32'hbb2712d9),
	.w8(32'h3a97b121),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c60cf),
	.w1(32'hbafbfeca),
	.w2(32'hbb098c12),
	.w3(32'hb86af50f),
	.w4(32'h3bd705ab),
	.w5(32'h3c061fe2),
	.w6(32'h3aea67f4),
	.w7(32'h3c297a86),
	.w8(32'h3c9a4708),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa975c),
	.w1(32'hb8b7fde1),
	.w2(32'h3cac2389),
	.w3(32'h3aac0990),
	.w4(32'h3cbda828),
	.w5(32'h3ce8e00c),
	.w6(32'h3bfe587f),
	.w7(32'h3cf94ae4),
	.w8(32'h3d171e2c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce603a3),
	.w1(32'h3cc2d766),
	.w2(32'hbc28c855),
	.w3(32'h3cdb66d8),
	.w4(32'hbbb8d7fd),
	.w5(32'hbc0ee1b4),
	.w6(32'h3d11f9fb),
	.w7(32'hbbb7b605),
	.w8(32'hbba15068),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3149b6),
	.w1(32'hbc2fb207),
	.w2(32'h3b47b0d2),
	.w3(32'hbb4ff284),
	.w4(32'hbba61f03),
	.w5(32'h3a7c2255),
	.w6(32'hbb568dbb),
	.w7(32'hbb1eb4fa),
	.w8(32'h39761af3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b348991),
	.w1(32'h3c16aba9),
	.w2(32'h3c1c8cdc),
	.w3(32'h3bca681a),
	.w4(32'h3c517346),
	.w5(32'h3c59f7ab),
	.w6(32'h3ba43071),
	.w7(32'h3c6a4dfa),
	.w8(32'h3c8256ae),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cda51),
	.w1(32'h3c12207c),
	.w2(32'hbc3d3ad5),
	.w3(32'h3bdae401),
	.w4(32'hbc3e7c11),
	.w5(32'hbb296d42),
	.w6(32'h3c1f0af5),
	.w7(32'hbc17eca7),
	.w8(32'h3aebc2c4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55423e),
	.w1(32'hbc555549),
	.w2(32'hbb98616c),
	.w3(32'hbc37b9fd),
	.w4(32'hbc16d677),
	.w5(32'hbb97593b),
	.w6(32'hbbec4417),
	.w7(32'hbb2a7005),
	.w8(32'hbb2a1b73),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b8c2d),
	.w1(32'h3c1ceae2),
	.w2(32'h3c333a4a),
	.w3(32'h3b1a4dac),
	.w4(32'h3c041572),
	.w5(32'h3bf6c691),
	.w6(32'h3bc7bee7),
	.w7(32'h3bad4c28),
	.w8(32'h3b84efc1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7582c),
	.w1(32'h3bbb6eab),
	.w2(32'h3c7cc239),
	.w3(32'h3c13b3bd),
	.w4(32'h3c979ad6),
	.w5(32'h3c43e16d),
	.w6(32'h3c29d6c1),
	.w7(32'h3cb0061d),
	.w8(32'h3c570e62),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d9270),
	.w1(32'h3a6a2db0),
	.w2(32'hbbc4ff6d),
	.w3(32'h3be84898),
	.w4(32'hbbdede3e),
	.w5(32'hbc3f0f71),
	.w6(32'h3bc522ba),
	.w7(32'hbc0adf2a),
	.w8(32'hbc404e17),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fc0fe),
	.w1(32'hbbc5681d),
	.w2(32'h393ba76f),
	.w3(32'hbbd351c1),
	.w4(32'h3c3e8531),
	.w5(32'h3be9aeac),
	.w6(32'hbbfee1ac),
	.w7(32'h3be4d70e),
	.w8(32'h3ae648ca),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab08180),
	.w1(32'hbb9ab36c),
	.w2(32'hbb82fa5a),
	.w3(32'h3c0321f2),
	.w4(32'hbb460b99),
	.w5(32'hbc34c2d0),
	.w6(32'h3b997802),
	.w7(32'hbae6c064),
	.w8(32'hbc15c8fa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd500c),
	.w1(32'hbb648a87),
	.w2(32'hbc031f9c),
	.w3(32'hbbb71b59),
	.w4(32'h39f82a3c),
	.w5(32'h3c17b326),
	.w6(32'hbb7ea14b),
	.w7(32'h3a3a4076),
	.w8(32'h3c3936f6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b5928),
	.w1(32'h3b8b1c7c),
	.w2(32'h3b4c396b),
	.w3(32'h3be5cfcc),
	.w4(32'hbc3693ce),
	.w5(32'hb884f5dd),
	.w6(32'h3c221278),
	.w7(32'hbc445f83),
	.w8(32'hbb8c08c3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b393a),
	.w1(32'h3b9b90bd),
	.w2(32'h3bbbdf18),
	.w3(32'hbb65ab4b),
	.w4(32'h3abfd45c),
	.w5(32'hbb761825),
	.w6(32'hbb5fec4b),
	.w7(32'h3c534541),
	.w8(32'h3c30c6a0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc38bc),
	.w1(32'h3ac33d5d),
	.w2(32'hbb90318c),
	.w3(32'hbade0a68),
	.w4(32'hbc336b33),
	.w5(32'hbb9641cf),
	.w6(32'h3c5e8806),
	.w7(32'hbbdc2573),
	.w8(32'hbb388bd7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1a4d),
	.w1(32'hbb4900de),
	.w2(32'hbc5a06f3),
	.w3(32'hbba11c85),
	.w4(32'hbc5aebce),
	.w5(32'h3a946be9),
	.w6(32'hbb3d67d7),
	.w7(32'hbbe935e6),
	.w8(32'h3c2015fa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa295e),
	.w1(32'h3a37ef4f),
	.w2(32'hbc08b02e),
	.w3(32'h3babe015),
	.w4(32'hbc678068),
	.w5(32'hbc3b241c),
	.w6(32'h3c4ced7e),
	.w7(32'hbc3e1955),
	.w8(32'hbc0a8910),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1f6ed),
	.w1(32'hbc16ff17),
	.w2(32'hbb48447f),
	.w3(32'hbc2dcfc7),
	.w4(32'hbbc236ec),
	.w5(32'hbba5ce17),
	.w6(32'hbb9904a4),
	.w7(32'hb8e358f3),
	.w8(32'hbb8f3a3d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03a754),
	.w1(32'hbbf178cd),
	.w2(32'hbc50e9c6),
	.w3(32'hbc0a0f09),
	.w4(32'hbc50d505),
	.w5(32'hbc84945f),
	.w6(32'hbc0c417e),
	.w7(32'hbc591dd0),
	.w8(32'hbc8a9c12),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc942f26),
	.w1(32'hbc380ea9),
	.w2(32'hbc224dc6),
	.w3(32'hbc37ddda),
	.w4(32'hbc315d40),
	.w5(32'hbc11cdbc),
	.w6(32'hbc4b0cee),
	.w7(32'hbc2e7223),
	.w8(32'hbc09df15),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a0687),
	.w1(32'hbc3f9ea6),
	.w2(32'hbc905dba),
	.w3(32'hbc4f871f),
	.w4(32'hbbe28c7e),
	.w5(32'h3aba6fce),
	.w6(32'hbc215677),
	.w7(32'hbc3643f3),
	.w8(32'h39994912),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ef1d3),
	.w1(32'hbcb13401),
	.w2(32'hbab8efe1),
	.w3(32'hbc3df41f),
	.w4(32'hbbdbcdac),
	.w5(32'hbbe40d97),
	.w6(32'hbb9bd11f),
	.w7(32'hbb42e748),
	.w8(32'hbad7bc63),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafaed7e),
	.w1(32'h3bbd91a1),
	.w2(32'hbbc8d6a6),
	.w3(32'h3b930343),
	.w4(32'hbc00f5a2),
	.w5(32'hbbdc9d13),
	.w6(32'h3c236a8a),
	.w7(32'hbb8836e8),
	.w8(32'hbb9b033d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc279962),
	.w1(32'hbc5e6f9e),
	.w2(32'h3bd00f30),
	.w3(32'hbc1b5190),
	.w4(32'h3b16c393),
	.w5(32'h36fe60da),
	.w6(32'hbbf1189b),
	.w7(32'h3c48ac82),
	.w8(32'h3c3973a8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b70e1),
	.w1(32'h3bbd3d14),
	.w2(32'hbc140139),
	.w3(32'h3b57f656),
	.w4(32'hbc5ae8ed),
	.w5(32'hbc902f5a),
	.w6(32'h3c452a44),
	.w7(32'hbc860e8a),
	.w8(32'hbcba9ad8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0e1f5),
	.w1(32'hbcbae889),
	.w2(32'hbb91d5cc),
	.w3(32'hbcad7f48),
	.w4(32'hbb5ab1dc),
	.w5(32'hbbd93395),
	.w6(32'hbca33b7b),
	.w7(32'h3a2091a2),
	.w8(32'hbb957893),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03a0df),
	.w1(32'hbc09b9ce),
	.w2(32'h3aa61634),
	.w3(32'hbbf9ac47),
	.w4(32'h3c3393f0),
	.w5(32'h3c5392c8),
	.w6(32'hbbb8e1f0),
	.w7(32'h3b50f026),
	.w8(32'h3c075820),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef4444),
	.w1(32'h3b2eae24),
	.w2(32'hbaff2994),
	.w3(32'h3c11694e),
	.w4(32'hbc0cef3f),
	.w5(32'hbbeb9ffa),
	.w6(32'h3bc39664),
	.w7(32'hbbd58fba),
	.w8(32'hbbb3bbd6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76b689b),
	.w1(32'h3bac738e),
	.w2(32'h3befe770),
	.w3(32'h39c1d783),
	.w4(32'h3ac2ab16),
	.w5(32'hbb0302dd),
	.w6(32'h3b31209e),
	.w7(32'h3c799c94),
	.w8(32'h3c60560d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4971a0),
	.w1(32'h3bc37eb1),
	.w2(32'hbbffc44f),
	.w3(32'h3b03a7b0),
	.w4(32'hbc15b41a),
	.w5(32'hbb628582),
	.w6(32'h3c6150ee),
	.w7(32'hb841000c),
	.w8(32'h3c06b649),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00c6ba),
	.w1(32'hbb9a1b45),
	.w2(32'hba0ac169),
	.w3(32'hbbd3009d),
	.w4(32'h3a48412f),
	.w5(32'h3ba89def),
	.w6(32'h3b509f46),
	.w7(32'h3bc3f4d6),
	.w8(32'h3c18bdc4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38ad19),
	.w1(32'h3b7f6a9e),
	.w2(32'h3bef80ed),
	.w3(32'hbaa8493a),
	.w4(32'h3b50a5bd),
	.w5(32'h3a9fd868),
	.w6(32'h3c06cce1),
	.w7(32'h3b0b3af6),
	.w8(32'h3a6bfc5b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf4b74),
	.w1(32'h3a547d3e),
	.w2(32'hbc28f9c7),
	.w3(32'hbbb92601),
	.w4(32'hbc5b5439),
	.w5(32'hbc8805dc),
	.w6(32'hbb104bd5),
	.w7(32'hbc1b74ae),
	.w8(32'hbc7f7c9e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95d5d4),
	.w1(32'hbc688c14),
	.w2(32'h3b3ce3a5),
	.w3(32'hbc3aed16),
	.w4(32'h39fa1226),
	.w5(32'h3aa1c86a),
	.w6(32'hbc5c3a72),
	.w7(32'h3a3fbed1),
	.w8(32'h3bc9b83c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f3bc4),
	.w1(32'h3b0ead76),
	.w2(32'h3a46e02b),
	.w3(32'h3bd7c6af),
	.w4(32'hbb9a2f2f),
	.w5(32'hbbacfae5),
	.w6(32'h3bde235f),
	.w7(32'hb767a64c),
	.w8(32'hbb30d5b8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8db450),
	.w1(32'hbaa0107b),
	.w2(32'hbc5ad9b3),
	.w3(32'hbb9d6fdf),
	.w4(32'hbc3e383e),
	.w5(32'hbba2ff8c),
	.w6(32'hbb0b9c99),
	.w7(32'hbc685b87),
	.w8(32'hbc2723dd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0daa2e),
	.w1(32'h3b1e8e05),
	.w2(32'hbc3ec143),
	.w3(32'h3b4dbc47),
	.w4(32'hbc6af565),
	.w5(32'hbc3c7b27),
	.w6(32'h3a86ed50),
	.w7(32'hbc70887c),
	.w8(32'hbc3c2c4d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21f0dc),
	.w1(32'hbbf26d0c),
	.w2(32'h3b2e8eaa),
	.w3(32'hbbf16108),
	.w4(32'hbaddd142),
	.w5(32'hbb7c2a70),
	.w6(32'hbbddbefe),
	.w7(32'h3aec1cc2),
	.w8(32'hbb2e1ba6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a29e3),
	.w1(32'h3c20cfec),
	.w2(32'hbbfb52cf),
	.w3(32'h3b1f4996),
	.w4(32'hbc5673c4),
	.w5(32'hbc7dd3ba),
	.w6(32'h3c28c9a1),
	.w7(32'hbc807395),
	.w8(32'hbc8e6054),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd77fac),
	.w1(32'hbc2b95d7),
	.w2(32'hbb9f86ee),
	.w3(32'hbc742f42),
	.w4(32'hbbfd7146),
	.w5(32'hbc00d473),
	.w6(32'hbc4001e8),
	.w7(32'hbb5cff25),
	.w8(32'hbac00cda),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27f9f1),
	.w1(32'hb9909253),
	.w2(32'hbc3fa892),
	.w3(32'hbb7bd9a3),
	.w4(32'hbc19697d),
	.w5(32'hbc34f43c),
	.w6(32'h3a1ec2a4),
	.w7(32'hbc1ee4d5),
	.w8(32'hbc219641),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e28d0),
	.w1(32'hbbf359f4),
	.w2(32'hbc9fd863),
	.w3(32'hbc427c3f),
	.w4(32'hbca53957),
	.w5(32'hbc57044d),
	.w6(32'hbbfaf1b6),
	.w7(32'hbc89d124),
	.w8(32'hbbfe4bf0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d54a9),
	.w1(32'hbc051589),
	.w2(32'h3c22bd51),
	.w3(32'hbc1eaf16),
	.w4(32'h3bf7a0c0),
	.w5(32'h3bcb7600),
	.w6(32'hbbf1b38f),
	.w7(32'h3c10d155),
	.w8(32'h3bda559e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6baba),
	.w1(32'h3bcf2548),
	.w2(32'hbb8d7f1e),
	.w3(32'h3bb7711a),
	.w4(32'hbc4327dd),
	.w5(32'h3aa78887),
	.w6(32'h3bc22288),
	.w7(32'hbba3b856),
	.w8(32'h3bff5e0a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a8e99),
	.w1(32'hbbcfa90e),
	.w2(32'h3a5fe88e),
	.w3(32'hba6a200d),
	.w4(32'hbb8e15fd),
	.w5(32'hbb80601d),
	.w6(32'h3b1116bd),
	.w7(32'h3ab48677),
	.w8(32'h3b8c05c8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39acc2),
	.w1(32'hbb7a0734),
	.w2(32'hbbcc83c3),
	.w3(32'hbb02cbd6),
	.w4(32'hbb04c1b1),
	.w5(32'hbb9bee20),
	.w6(32'h3b130701),
	.w7(32'h3a0ab232),
	.w8(32'hbb1a07db),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92a3d1),
	.w1(32'hbad5a0f8),
	.w2(32'h3b20d71f),
	.w3(32'hbb1765a8),
	.w4(32'hbaaa7382),
	.w5(32'h3991dac3),
	.w6(32'h3a15a85e),
	.w7(32'hb91d26aa),
	.w8(32'hba820e93),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cb215),
	.w1(32'hbbfa3e15),
	.w2(32'hba2eb172),
	.w3(32'hbb4e3803),
	.w4(32'hbad278cc),
	.w5(32'h3a358c7c),
	.w6(32'hbadff784),
	.w7(32'h3aec93c9),
	.w8(32'h3a7813e0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a3294),
	.w1(32'hbb7da917),
	.w2(32'hba56a8c0),
	.w3(32'hbafeda3b),
	.w4(32'h39e83e91),
	.w5(32'hbb166dac),
	.w6(32'hbb58fc1e),
	.w7(32'hba94cf60),
	.w8(32'hbb051e99),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98a1d7),
	.w1(32'hba0b63a5),
	.w2(32'hbae9069f),
	.w3(32'h386fdeb1),
	.w4(32'hbb263acd),
	.w5(32'hbb86f4b5),
	.w6(32'hba3757c9),
	.w7(32'h3b09ae33),
	.w8(32'hbb18b621),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b3ac8),
	.w1(32'hbb8a5560),
	.w2(32'hbb5435c1),
	.w3(32'h3b6298b7),
	.w4(32'h3a2b8b2d),
	.w5(32'hbc012a5f),
	.w6(32'h3a8d6130),
	.w7(32'h3b9d83f0),
	.w8(32'hbc14c720),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c0b1b),
	.w1(32'hb80aa1bb),
	.w2(32'hbbf9e31e),
	.w3(32'hbb947635),
	.w4(32'hbc33b801),
	.w5(32'hba9341e2),
	.w6(32'h3accf1db),
	.w7(32'hbc5b6fbb),
	.w8(32'h3b46e265),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25db2f),
	.w1(32'hbba7e286),
	.w2(32'h3a88e6fb),
	.w3(32'hbbf1bea7),
	.w4(32'h3b43a415),
	.w5(32'h3c389d00),
	.w6(32'hbabecc66),
	.w7(32'h3c2c0154),
	.w8(32'h3c0219de),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e485),
	.w1(32'h3b20701b),
	.w2(32'hbc56cdb8),
	.w3(32'hbab7cf79),
	.w4(32'hbb46dbeb),
	.w5(32'hbb9933bc),
	.w6(32'h3bbb795e),
	.w7(32'h3ac97620),
	.w8(32'hbbb34041),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40fa89),
	.w1(32'hbbfeb74f),
	.w2(32'h3c699bc5),
	.w3(32'hbad977f4),
	.w4(32'h3a86e3d3),
	.w5(32'h3c21c153),
	.w6(32'h3b008ede),
	.w7(32'h3bf2995f),
	.w8(32'hbb64b563),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d01e8a),
	.w1(32'hbbeb4c9f),
	.w2(32'hbba73bcd),
	.w3(32'h3b96ff6d),
	.w4(32'hbc13c868),
	.w5(32'hbc2feee1),
	.w6(32'h3b06bca2),
	.w7(32'hbba4ab5a),
	.w8(32'hbbbd29a8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0293c7),
	.w1(32'h3b4acf1e),
	.w2(32'h39c8d185),
	.w3(32'hbac53c49),
	.w4(32'h3bb7acda),
	.w5(32'h3c460964),
	.w6(32'hbbc49598),
	.w7(32'hbad15995),
	.w8(32'h3bb870f6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52e51a),
	.w1(32'h3b8292b3),
	.w2(32'hbbd2cb59),
	.w3(32'h3b81e659),
	.w4(32'hbbe274b7),
	.w5(32'hbc1929ce),
	.w6(32'h3bc7807d),
	.w7(32'hbc1b5f05),
	.w8(32'hbc41ae6b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e8d49),
	.w1(32'hbb1933af),
	.w2(32'h3c63f258),
	.w3(32'hbb1029ba),
	.w4(32'h3c8cbf94),
	.w5(32'h3d125977),
	.w6(32'hbb04a912),
	.w7(32'h3c895c0a),
	.w8(32'h3d0b5ad5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d4349),
	.w1(32'h3bcd7be8),
	.w2(32'hbb58a4a7),
	.w3(32'h3c9269cc),
	.w4(32'h3c03124a),
	.w5(32'hbb2d2952),
	.w6(32'h3c113c45),
	.w7(32'h38f6c91a),
	.w8(32'hbc1cac99),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43dcc),
	.w1(32'h3c7dd490),
	.w2(32'hbaae8643),
	.w3(32'hbbdcd549),
	.w4(32'h3be5bbba),
	.w5(32'h39fe8012),
	.w6(32'hbc15d75b),
	.w7(32'h3ba55fe3),
	.w8(32'hba3a8240),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47e129),
	.w1(32'hbb895878),
	.w2(32'hbc03f2ed),
	.w3(32'hbac81994),
	.w4(32'h3ae478f9),
	.w5(32'hbc55f64d),
	.w6(32'hbb4569ac),
	.w7(32'hba981349),
	.w8(32'hbba6320c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba457ea),
	.w1(32'hbba61273),
	.w2(32'hba3be645),
	.w3(32'hbc5d8dec),
	.w4(32'hba0ba03a),
	.w5(32'h3a76bed1),
	.w6(32'hbc284aa9),
	.w7(32'hbbadcd9f),
	.w8(32'h3a086cf5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb18bb2),
	.w1(32'h3b11b1de),
	.w2(32'hbaf999c0),
	.w3(32'hbb4f21e2),
	.w4(32'hbc859da0),
	.w5(32'h3aab82ea),
	.w6(32'hbb0d6775),
	.w7(32'hbb8cf4a2),
	.w8(32'h3b7b172d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6f99e),
	.w1(32'hbc9d03f0),
	.w2(32'h3a1bbdbc),
	.w3(32'hbb31e29d),
	.w4(32'h39803c81),
	.w5(32'h3a8c5e91),
	.w6(32'hbbc1358f),
	.w7(32'h39007686),
	.w8(32'h3a8f9d82),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68cdff),
	.w1(32'h3aa6690f),
	.w2(32'h3b834153),
	.w3(32'h3af3e42c),
	.w4(32'hbb553672),
	.w5(32'hbb84ebf6),
	.w6(32'h3b56f680),
	.w7(32'hbb3143a9),
	.w8(32'hb96466cb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b894ded),
	.w1(32'hbc29305d),
	.w2(32'hbbe33778),
	.w3(32'h3b9f85bb),
	.w4(32'hbb689da3),
	.w5(32'h3c9ed59c),
	.w6(32'hbb6555ac),
	.w7(32'hbaef695a),
	.w8(32'h3b9ec852),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec5817),
	.w1(32'hbb9dd715),
	.w2(32'h3c10fae1),
	.w3(32'h39e24fc6),
	.w4(32'h3abb99fe),
	.w5(32'hbbcae2ba),
	.w6(32'hbba4917c),
	.w7(32'h3b9d9a41),
	.w8(32'hbc1a9385),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d2a16),
	.w1(32'hbc299ed1),
	.w2(32'hbaa7e123),
	.w3(32'hbbc07ffb),
	.w4(32'h3b8604f5),
	.w5(32'hba3fc67e),
	.w6(32'hbb04cdac),
	.w7(32'h3b307ab1),
	.w8(32'hbb26d25b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdecb8e),
	.w1(32'h3a8ac3ec),
	.w2(32'h3c09aef7),
	.w3(32'h3b390c0a),
	.w4(32'h3b873063),
	.w5(32'h3cfcaee7),
	.w6(32'h3b2f6e93),
	.w7(32'h3a58b2f8),
	.w8(32'h3d03a031),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4da27),
	.w1(32'h3c6b70b6),
	.w2(32'h3ae72d67),
	.w3(32'h3c54ca17),
	.w4(32'hbb32a05b),
	.w5(32'h3b4062bb),
	.w6(32'h3caeda9b),
	.w7(32'hbadc9f87),
	.w8(32'hba2ffd54),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd501e9),
	.w1(32'hbc15f822),
	.w2(32'hbc0bbef5),
	.w3(32'hba8387ec),
	.w4(32'h3b453ecc),
	.w5(32'h3cd191a9),
	.w6(32'hbb81ec6d),
	.w7(32'hbab53b01),
	.w8(32'h3cd5baaf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd91194),
	.w1(32'h3cce4b36),
	.w2(32'hbbfa4aed),
	.w3(32'h3cb78be2),
	.w4(32'hb75caddd),
	.w5(32'h3bbed011),
	.w6(32'h3cb214fd),
	.w7(32'hbbb19653),
	.w8(32'h3baf9e35),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb654f82),
	.w1(32'h3b9f960a),
	.w2(32'hbb99cf41),
	.w3(32'h3a3436ea),
	.w4(32'h3aabd148),
	.w5(32'hbabd3481),
	.w6(32'h3a884683),
	.w7(32'hba4da195),
	.w8(32'h3c370ef9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f9b12),
	.w1(32'h3c3aacf1),
	.w2(32'hbbc2ff30),
	.w3(32'hbb2675bc),
	.w4(32'hbae7a7ae),
	.w5(32'hbc335445),
	.w6(32'h3bcc1689),
	.w7(32'h3b2d4439),
	.w8(32'hbc1aad11),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034346),
	.w1(32'hbc5f7688),
	.w2(32'hbb53edcf),
	.w3(32'h3b5e3606),
	.w4(32'h3a9fb2c0),
	.w5(32'hbba764c0),
	.w6(32'hbc2be230),
	.w7(32'h3a3ef784),
	.w8(32'hb95f2011),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372b60a3),
	.w1(32'h3b9809a4),
	.w2(32'h3c2f97d0),
	.w3(32'hbb0c00d0),
	.w4(32'hbb1ccbe1),
	.w5(32'h3b98fb2d),
	.w6(32'h3b7376fc),
	.w7(32'hbaf78e5c),
	.w8(32'hb7b54f18),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f2e71),
	.w1(32'hba1c091f),
	.w2(32'h3b1dbed2),
	.w3(32'h3a9c0f6a),
	.w4(32'hbaa36b9d),
	.w5(32'h39a87226),
	.w6(32'h3b74d1ba),
	.w7(32'h3a794116),
	.w8(32'hb9b1048e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a8d48),
	.w1(32'hbbb948b3),
	.w2(32'h3c36a0ab),
	.w3(32'hbb878c3c),
	.w4(32'hbae69618),
	.w5(32'hbb053792),
	.w6(32'hbba4eb65),
	.w7(32'h3a5e1dca),
	.w8(32'hbb93031b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4bda),
	.w1(32'hbb7fa89c),
	.w2(32'hbba63a36),
	.w3(32'hbc1d8fb1),
	.w4(32'hbc75c598),
	.w5(32'hbc5bebbe),
	.w6(32'hbc19015e),
	.w7(32'hbaec1e02),
	.w8(32'h3ac5c0f2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79af08),
	.w1(32'h3c0da284),
	.w2(32'hba099d2b),
	.w3(32'h3c7e8505),
	.w4(32'h3aad01cc),
	.w5(32'h3b73dcaa),
	.w6(32'h3c95704d),
	.w7(32'h3b6421f7),
	.w8(32'h3c291445),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc47d3),
	.w1(32'h3c1e357c),
	.w2(32'h3bf3dc4b),
	.w3(32'hba51256d),
	.w4(32'h3b5e7086),
	.w5(32'h3c3623b8),
	.w6(32'h3ba3953f),
	.w7(32'h3c1e210c),
	.w8(32'h3c2577cd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c038ab5),
	.w1(32'h3be34087),
	.w2(32'h3c036b6d),
	.w3(32'hbbbb9678),
	.w4(32'h3b03c2bb),
	.w5(32'hbac620ec),
	.w6(32'hbb0ee625),
	.w7(32'h3c11bec3),
	.w8(32'hbafd3e03),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e4c77),
	.w1(32'hbc1cbcd7),
	.w2(32'hbb5ef057),
	.w3(32'h3b2600ce),
	.w4(32'h38506b63),
	.w5(32'h3b7568e6),
	.w6(32'hbb5c4dd5),
	.w7(32'hbb029a3b),
	.w8(32'h3c1b9a3e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8681f),
	.w1(32'hbbd7fca6),
	.w2(32'hbc4126f7),
	.w3(32'h3b37e2f9),
	.w4(32'h3bcf2847),
	.w5(32'h3aa8cb15),
	.w6(32'hbb562991),
	.w7(32'h3b7df20f),
	.w8(32'h3a0961e4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90f0fb),
	.w1(32'h3be7e923),
	.w2(32'hbab5ed00),
	.w3(32'h3bf6c6b4),
	.w4(32'h3b6e8f91),
	.w5(32'hbc682959),
	.w6(32'h3bc8fb12),
	.w7(32'h3bd326fe),
	.w8(32'hbc46b18d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaba3d7),
	.w1(32'hbc4cce1c),
	.w2(32'h3b3e3edf),
	.w3(32'hbbb1f9ec),
	.w4(32'h3abb4afe),
	.w5(32'h3b8d6649),
	.w6(32'hbbdbbfd3),
	.w7(32'hb9489100),
	.w8(32'h3c75a8cb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca38f43),
	.w1(32'hbbd1e06d),
	.w2(32'h3b09840e),
	.w3(32'h3c1812ac),
	.w4(32'hba7f87be),
	.w5(32'h3b07c6e9),
	.w6(32'hbaad2e26),
	.w7(32'h3b327b7a),
	.w8(32'h3aee6e62),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3830ea91),
	.w1(32'hbb381511),
	.w2(32'hbb96c0ec),
	.w3(32'hb9eb0d0b),
	.w4(32'h3bce4d68),
	.w5(32'h3a0b894c),
	.w6(32'hbb02d23b),
	.w7(32'hba86d1f0),
	.w8(32'hbb0d3951),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1541),
	.w1(32'h39e2aec4),
	.w2(32'hbaee60cb),
	.w3(32'hbc1ae05d),
	.w4(32'h39edec10),
	.w5(32'hbc35b4cb),
	.w6(32'h3b6f0727),
	.w7(32'h3b46dd8b),
	.w8(32'hbc254bff),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc045f80),
	.w1(32'hbb9f3fdf),
	.w2(32'hbbc1f2c8),
	.w3(32'hbbec10b3),
	.w4(32'hbc0f2ca4),
	.w5(32'hbc0db136),
	.w6(32'hbbaf44b2),
	.w7(32'hbbe05642),
	.w8(32'hbb822b85),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2ee62),
	.w1(32'hbb00e42e),
	.w2(32'hba725931),
	.w3(32'hbba0e209),
	.w4(32'h3abe87ae),
	.w5(32'hbbd3adb5),
	.w6(32'hba2dcb44),
	.w7(32'h3aec9bdb),
	.w8(32'hba7bcbdc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08036a),
	.w1(32'h3c44da24),
	.w2(32'h3a2e02b0),
	.w3(32'h3b5c8cca),
	.w4(32'hb9df1ff6),
	.w5(32'h3a1c0558),
	.w6(32'h3c23af96),
	.w7(32'h3a81e9d0),
	.w8(32'h38994513),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e7037),
	.w1(32'hbb847c24),
	.w2(32'hbc1a92f6),
	.w3(32'hbb0a7b1b),
	.w4(32'h3a29c956),
	.w5(32'hbb97bd1a),
	.w6(32'hbb2ff3a1),
	.w7(32'hbbcdf638),
	.w8(32'hbbb2aad5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2c39d),
	.w1(32'h3c6239da),
	.w2(32'hbb122c6a),
	.w3(32'h3b699556),
	.w4(32'h3b21ab25),
	.w5(32'h3bce5d76),
	.w6(32'h3c790396),
	.w7(32'hbc34f522),
	.w8(32'h3c665f23),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207fe9),
	.w1(32'hbc181c7b),
	.w2(32'hbc3437b1),
	.w3(32'hbadfc950),
	.w4(32'hbc224257),
	.w5(32'hbbfb704c),
	.w6(32'hbbe3169c),
	.w7(32'hbc54a76b),
	.w8(32'hbc075b10),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e0145),
	.w1(32'hbbab5964),
	.w2(32'hbbaaf294),
	.w3(32'hb7fda2b7),
	.w4(32'hbb9c4b8e),
	.w5(32'h3ae7fab2),
	.w6(32'hbb4e19a8),
	.w7(32'hbb9042d4),
	.w8(32'hbbad1bc5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe923e),
	.w1(32'hbb9d11b9),
	.w2(32'h3b1b7c44),
	.w3(32'hbb14bd5f),
	.w4(32'hbb81be90),
	.w5(32'hba5590af),
	.w6(32'hbc29593e),
	.w7(32'hbb07b5c0),
	.w8(32'hbb06e50e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule