module layer_10_featuremap_478(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbd784),
	.w1(32'h3b059054),
	.w2(32'h3b5971f2),
	.w3(32'hbb72a053),
	.w4(32'hbb61be65),
	.w5(32'h3a5c4b11),
	.w6(32'hbbc12a61),
	.w7(32'h3ad6e67d),
	.w8(32'h3b88075f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba890277),
	.w1(32'hbbb663d7),
	.w2(32'h3ba29575),
	.w3(32'hbabd8351),
	.w4(32'hbc49ac91),
	.w5(32'hb9810afe),
	.w6(32'h3c1e519f),
	.w7(32'hbc9477fa),
	.w8(32'hbbe8b6cf),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ae889),
	.w1(32'h3a34e8e3),
	.w2(32'hbc5286ed),
	.w3(32'h3c939b84),
	.w4(32'h3caba1b0),
	.w5(32'h3c4f017e),
	.w6(32'h3bdb995d),
	.w7(32'h3c64d7d5),
	.w8(32'h3cabbed2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a80af),
	.w1(32'hbc98ca70),
	.w2(32'hbc044b30),
	.w3(32'hbb2f98d8),
	.w4(32'hbc7e1819),
	.w5(32'h39e84040),
	.w6(32'hbb786ca9),
	.w7(32'hbc79fa11),
	.w8(32'hbbbb230f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9093ef),
	.w1(32'hba415851),
	.w2(32'hbb892f16),
	.w3(32'h3a8b0b9b),
	.w4(32'h3ba9d400),
	.w5(32'hbac6c366),
	.w6(32'hbbc5e50e),
	.w7(32'h3c051ddd),
	.w8(32'h3b9edda1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6332e),
	.w1(32'h3a37bdcf),
	.w2(32'hb861dc22),
	.w3(32'h3a01c0ae),
	.w4(32'hbbf8d5d2),
	.w5(32'hbc5641b4),
	.w6(32'h3996b850),
	.w7(32'hbaa8e67a),
	.w8(32'hbbde8732),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c7dc9),
	.w1(32'hbc30afcc),
	.w2(32'hbbdb7ad1),
	.w3(32'h3a9749db),
	.w4(32'h3b6d844b),
	.w5(32'hbb233fd1),
	.w6(32'hbb171e87),
	.w7(32'h3ae80a21),
	.w8(32'hbb7d4d9c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6869b8),
	.w1(32'h3c9fe417),
	.w2(32'h3b52086a),
	.w3(32'h3aad3198),
	.w4(32'hbb2dc5a9),
	.w5(32'hbb563ee3),
	.w6(32'hbbdb890a),
	.w7(32'hbb53463d),
	.w8(32'hbc2a407a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e2b77),
	.w1(32'hbc262efb),
	.w2(32'h3ba34d04),
	.w3(32'hbc173d4c),
	.w4(32'hbc5acc7a),
	.w5(32'h3c9ed5d9),
	.w6(32'hbc35d18a),
	.w7(32'hbc389c47),
	.w8(32'h3bb6886d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a661be8),
	.w1(32'hbc2a56d7),
	.w2(32'hbb9ca3e4),
	.w3(32'h3c6da305),
	.w4(32'h3aa4f81d),
	.w5(32'h3a13a7f0),
	.w6(32'hbb3fb133),
	.w7(32'hba8b45b4),
	.w8(32'hbb27c027),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f178e),
	.w1(32'h3961a1ef),
	.w2(32'h3bbc0d04),
	.w3(32'hba3e1473),
	.w4(32'h3b9cf98f),
	.w5(32'h3a271092),
	.w6(32'hb9be0acb),
	.w7(32'hbbd50462),
	.w8(32'h3a42a13e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fe7ab),
	.w1(32'hbb1d7950),
	.w2(32'hbb96404c),
	.w3(32'h3a80d5ee),
	.w4(32'hbb89b7f8),
	.w5(32'hba545713),
	.w6(32'hbb7597bd),
	.w7(32'hbb8189ce),
	.w8(32'h3acf2d8e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47a461),
	.w1(32'hbc701a0e),
	.w2(32'hbbd622c4),
	.w3(32'h3bfcfd1d),
	.w4(32'hbc59bb8c),
	.w5(32'h3c5341e1),
	.w6(32'h3b0a3a5e),
	.w7(32'hbc85938e),
	.w8(32'h3b82e37c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd36da2),
	.w1(32'hbbfb8ec7),
	.w2(32'hbb69af4b),
	.w3(32'h3c8cc513),
	.w4(32'hbc052314),
	.w5(32'hba61cab5),
	.w6(32'h3c2d54d9),
	.w7(32'hbc6a1cc3),
	.w8(32'hbbfa8d63),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1693b7),
	.w1(32'h39c7fba0),
	.w2(32'hbc7eb13b),
	.w3(32'hbbdfd077),
	.w4(32'h3caeaed6),
	.w5(32'hbcc8c594),
	.w6(32'hbc067c6c),
	.w7(32'h3c96d1b3),
	.w8(32'hbc0c8930),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1da974),
	.w1(32'hbb3ab8f4),
	.w2(32'hbb5edb34),
	.w3(32'hbc7ff70c),
	.w4(32'hbba8f2d8),
	.w5(32'hbc1bca02),
	.w6(32'hbc93125e),
	.w7(32'hbbd0f376),
	.w8(32'hbbf01de3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07b86e),
	.w1(32'h3b967cfd),
	.w2(32'h3bc72444),
	.w3(32'hbc4afc93),
	.w4(32'h3c98a6d0),
	.w5(32'h3c949efe),
	.w6(32'hbc10b073),
	.w7(32'h3c825811),
	.w8(32'h3c655cad),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40950d),
	.w1(32'h3bff975c),
	.w2(32'h3c1edd6a),
	.w3(32'h3ca19c5a),
	.w4(32'h3bcf1f99),
	.w5(32'h3c01eab0),
	.w6(32'h3ba90dad),
	.w7(32'h3ae125d3),
	.w8(32'h3a2810cc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00386c),
	.w1(32'hba8bac12),
	.w2(32'h3c319b7b),
	.w3(32'hbb54eec3),
	.w4(32'hbaa89f7a),
	.w5(32'h3b8531ec),
	.w6(32'hbb453509),
	.w7(32'hbbc0be74),
	.w8(32'hb9ba9a33),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7311f6),
	.w1(32'h3b878a44),
	.w2(32'hb922cbd8),
	.w3(32'h3c6746b8),
	.w4(32'h3c912910),
	.w5(32'hbbdad468),
	.w6(32'h3c1743d1),
	.w7(32'h3c5a9a32),
	.w8(32'h3a50780a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44b840),
	.w1(32'h3c8f8f80),
	.w2(32'hbb34e26e),
	.w3(32'hbb8307e4),
	.w4(32'h3c019de0),
	.w5(32'hbc79d94c),
	.w6(32'hbc057550),
	.w7(32'h3b598249),
	.w8(32'hbc0d5fc9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c5645),
	.w1(32'h3bbf8103),
	.w2(32'hba720de7),
	.w3(32'hbc225b68),
	.w4(32'h3c86e833),
	.w5(32'hbc0b3913),
	.w6(32'hbc0d6e2c),
	.w7(32'h3c0c07f6),
	.w8(32'h3a838375),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30c7cf),
	.w1(32'h3a13bf52),
	.w2(32'h3c3faf7c),
	.w3(32'h3bf75f43),
	.w4(32'h3c202257),
	.w5(32'h3b14bd3e),
	.w6(32'hba942813),
	.w7(32'hbb71c995),
	.w8(32'hbaf62941),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34647b),
	.w1(32'hb7fb155c),
	.w2(32'h3c22d295),
	.w3(32'hb9416d12),
	.w4(32'h3c394a77),
	.w5(32'h3ce36fdb),
	.w6(32'h3a4a0a08),
	.w7(32'hbbbcd8af),
	.w8(32'h3b2a0042),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e04fa),
	.w1(32'hba99e029),
	.w2(32'h3b70d7ae),
	.w3(32'h3b78aa94),
	.w4(32'hbaa3f80d),
	.w5(32'h3b7c9ad8),
	.w6(32'hbbdc219a),
	.w7(32'hbc167548),
	.w8(32'hbbfe614f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef1fbc),
	.w1(32'h3c293b5c),
	.w2(32'hbc0f5341),
	.w3(32'h3b1e3fee),
	.w4(32'hbc164d7f),
	.w5(32'hbc91a387),
	.w6(32'h3974e448),
	.w7(32'h3c1af82d),
	.w8(32'hbc282070),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf3d4f),
	.w1(32'h3c085a89),
	.w2(32'hb9f6cdb1),
	.w3(32'h3b29d753),
	.w4(32'hbb2dde02),
	.w5(32'hbc58751f),
	.w6(32'h3c1edbf8),
	.w7(32'hbb61b8ef),
	.w8(32'hbc08a683),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac15a19),
	.w1(32'hbc617ff2),
	.w2(32'h3a47eea1),
	.w3(32'hb9802395),
	.w4(32'hbb936107),
	.w5(32'h3c00920b),
	.w6(32'h3b9627af),
	.w7(32'hba6d83b8),
	.w8(32'h3b685a8d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30f78f),
	.w1(32'hbb2e8542),
	.w2(32'hb9b50b88),
	.w3(32'hba80ba0f),
	.w4(32'hbb6949ce),
	.w5(32'hbb939863),
	.w6(32'h3b850353),
	.w7(32'h3b0d61cd),
	.w8(32'h3c6e075a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc418cd6),
	.w1(32'hbbc43124),
	.w2(32'hbc037f66),
	.w3(32'hbb3a3455),
	.w4(32'hbbad7035),
	.w5(32'hbc10b01e),
	.w6(32'h3c6e232e),
	.w7(32'hb93d310d),
	.w8(32'hbb47f5b0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2e460),
	.w1(32'h3b7493e7),
	.w2(32'h3bd74630),
	.w3(32'hbb96877a),
	.w4(32'hbb85cba9),
	.w5(32'hbbd7d841),
	.w6(32'hbb300b62),
	.w7(32'h3b0e133e),
	.w8(32'h3b3e2e2a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdd92d),
	.w1(32'h3add8981),
	.w2(32'hbbea2673),
	.w3(32'hbad5274e),
	.w4(32'h3c1b2579),
	.w5(32'hbb1b0f48),
	.w6(32'h3b88c96d),
	.w7(32'hbb3d6604),
	.w8(32'hbb5efdf2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9105d),
	.w1(32'h3c674963),
	.w2(32'h3c9f62cb),
	.w3(32'hbaada934),
	.w4(32'hba9878ff),
	.w5(32'hba6e9f21),
	.w6(32'hbbec5796),
	.w7(32'h3973a664),
	.w8(32'hbc0e92c5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68d6e9),
	.w1(32'h3b0e34f0),
	.w2(32'h3c314578),
	.w3(32'hbbd2f8c7),
	.w4(32'h3b61c411),
	.w5(32'h3b67982d),
	.w6(32'hbbafb800),
	.w7(32'h3c60049c),
	.w8(32'h3bc3c20b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83cc1c),
	.w1(32'h3b52e595),
	.w2(32'h3b205868),
	.w3(32'h3af7b313),
	.w4(32'hbbac26ba),
	.w5(32'h392d0d1e),
	.w6(32'h3c00c57b),
	.w7(32'h3ba0bc8f),
	.w8(32'hbbb4ae76),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79172a),
	.w1(32'hbc023183),
	.w2(32'hbbcf4930),
	.w3(32'hbaf5cda3),
	.w4(32'hbb79df30),
	.w5(32'h3c1831a7),
	.w6(32'hbc078bdc),
	.w7(32'hbbe2b050),
	.w8(32'hbb8f5f8e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac6832),
	.w1(32'h3c098ea1),
	.w2(32'h3b206e98),
	.w3(32'hbc0baf7e),
	.w4(32'h3c43765e),
	.w5(32'hbb02278f),
	.w6(32'hbc8ebf6f),
	.w7(32'h3b96b9f0),
	.w8(32'h3c3ca9ee),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0e740),
	.w1(32'hbc04b9de),
	.w2(32'h3b662c07),
	.w3(32'hbb14c450),
	.w4(32'hbc475484),
	.w5(32'h3bb00099),
	.w6(32'h3c067efd),
	.w7(32'hbc5dadaa),
	.w8(32'hbbf9784c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1c7e2),
	.w1(32'hbafa5303),
	.w2(32'h3a952c75),
	.w3(32'h3c342db0),
	.w4(32'h3b28c82b),
	.w5(32'h3bdcac62),
	.w6(32'h3b856868),
	.w7(32'h3a80cbb9),
	.w8(32'h3bd02dc3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199ea6),
	.w1(32'hbc482681),
	.w2(32'hbbd4efae),
	.w3(32'h3b6a577d),
	.w4(32'hbc823ee3),
	.w5(32'h3b2201bb),
	.w6(32'h3bafab1f),
	.w7(32'hbc366ad2),
	.w8(32'hbbffb050),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b445),
	.w1(32'hbc9b96ab),
	.w2(32'hbacc2ff4),
	.w3(32'h3b3d0f04),
	.w4(32'hbb965f8d),
	.w5(32'h3c98bc78),
	.w6(32'h3abb3435),
	.w7(32'hbc86047f),
	.w8(32'hbc82bd53),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc854dd8),
	.w1(32'h3a2f8299),
	.w2(32'hb9926bd5),
	.w3(32'hbc4a8a14),
	.w4(32'h3c0a75f6),
	.w5(32'hbaa30629),
	.w6(32'hbc9f38ef),
	.w7(32'hb7ce4e42),
	.w8(32'hbb87331c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9745e),
	.w1(32'hbb836cfd),
	.w2(32'hba8abfc0),
	.w3(32'hbb7c3f04),
	.w4(32'hbb8686f8),
	.w5(32'h3b30e724),
	.w6(32'hbc22a4e9),
	.w7(32'hbc0eec62),
	.w8(32'hbb6ee673),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e9eb0),
	.w1(32'hbc546d28),
	.w2(32'h3ba41cc1),
	.w3(32'h3c32b19f),
	.w4(32'hbc5dc914),
	.w5(32'h3c068c84),
	.w6(32'h3b80899a),
	.w7(32'hbc10020a),
	.w8(32'hba9baa68),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c030ff8),
	.w1(32'hbb871ce4),
	.w2(32'h3b46692c),
	.w3(32'h3b9b60f8),
	.w4(32'hbb223682),
	.w5(32'hbbacf3e3),
	.w6(32'h3baedadb),
	.w7(32'hbba75c7e),
	.w8(32'hbb9169ee),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fe1f9),
	.w1(32'hbb98b335),
	.w2(32'hbb09d29f),
	.w3(32'hbbcf35db),
	.w4(32'hbbb8018c),
	.w5(32'hbb9a1ec9),
	.w6(32'hbb72529b),
	.w7(32'hbc5b810d),
	.w8(32'hbc85a1bb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5165a),
	.w1(32'h3b904bc3),
	.w2(32'hbc01d741),
	.w3(32'hbc0767b6),
	.w4(32'hba8affee),
	.w5(32'hbb83dae4),
	.w6(32'hbc2209d1),
	.w7(32'hbc6c98b1),
	.w8(32'hbbae38af),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86eee0),
	.w1(32'h39305d50),
	.w2(32'h3b292db4),
	.w3(32'h3bfb6f37),
	.w4(32'hbbb41907),
	.w5(32'h3bb0869b),
	.w6(32'hbae61456),
	.w7(32'hbb0a1849),
	.w8(32'hbb397285),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b642cd0),
	.w1(32'hbbae5f44),
	.w2(32'h3ad4cbfb),
	.w3(32'h3bb5ae6b),
	.w4(32'hbc83f8d5),
	.w5(32'hba6f74f9),
	.w6(32'h3b85875b),
	.w7(32'hbc72bc8f),
	.w8(32'hbc28c1a7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb747ecf),
	.w1(32'h3ba03537),
	.w2(32'hbab59e9a),
	.w3(32'hbbc726aa),
	.w4(32'h3b2f4121),
	.w5(32'hbadc69d3),
	.w6(32'hbc580de9),
	.w7(32'h393a3c20),
	.w8(32'hbb5376a0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb99823),
	.w1(32'hbb121489),
	.w2(32'hba6114ec),
	.w3(32'hbc4a74c7),
	.w4(32'hbbba647b),
	.w5(32'h3b9b7732),
	.w6(32'hbc4411cc),
	.w7(32'hbb816ae8),
	.w8(32'h3bf1d4c6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1ad65),
	.w1(32'h3b09ac76),
	.w2(32'h3b17a1c4),
	.w3(32'h3b20e388),
	.w4(32'hbb179d0c),
	.w5(32'hba89a73d),
	.w6(32'hbb07f1c4),
	.w7(32'hbc5fbc0a),
	.w8(32'hbbf4b1a5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb855ed9),
	.w1(32'h3c13d4c4),
	.w2(32'h3c1cec8b),
	.w3(32'hbb391fc2),
	.w4(32'h3a8d3af2),
	.w5(32'h3b38acf5),
	.w6(32'hbb00facd),
	.w7(32'h3a2bd289),
	.w8(32'hbb57397f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65adf8),
	.w1(32'h3c6c689e),
	.w2(32'h3c23e926),
	.w3(32'h3c4354ff),
	.w4(32'h3a3f341a),
	.w5(32'hba5ef586),
	.w6(32'hb7d7a0b6),
	.w7(32'hbb884d72),
	.w8(32'hbc17627c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ac0ad),
	.w1(32'hbc403d65),
	.w2(32'hbadd7044),
	.w3(32'hbbc66cd8),
	.w4(32'hbc2fea1a),
	.w5(32'h3c03b8f0),
	.w6(32'hbb579d3a),
	.w7(32'hbc92889c),
	.w8(32'hba95a409),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdb67d),
	.w1(32'hbc09ba07),
	.w2(32'h3c404cf3),
	.w3(32'h3c073a60),
	.w4(32'hbc59a928),
	.w5(32'h3c425560),
	.w6(32'h3ba13fd4),
	.w7(32'hbc6798db),
	.w8(32'hbc12146a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd493b9),
	.w1(32'h3b129eed),
	.w2(32'hbb37e6f4),
	.w3(32'h3c7d90d0),
	.w4(32'hbb25e495),
	.w5(32'hbbbfc98d),
	.w6(32'hbb1c07e4),
	.w7(32'h3bacdfae),
	.w8(32'hbaa9a02f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe96cb4),
	.w1(32'h3a5d54d8),
	.w2(32'hbbbbee92),
	.w3(32'hbbe52320),
	.w4(32'h3b9aa421),
	.w5(32'hbbb0124f),
	.w6(32'hbb739da1),
	.w7(32'h3c66ba63),
	.w8(32'hbbac0c93),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13e631),
	.w1(32'hbc77329d),
	.w2(32'hbc2c87a2),
	.w3(32'hbba0ec79),
	.w4(32'hbc01a3c5),
	.w5(32'hb9ad1a0e),
	.w6(32'hbc2a096f),
	.w7(32'hbc4a3df6),
	.w8(32'hbbefeae7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fbe09),
	.w1(32'h39de124e),
	.w2(32'hba0c51a6),
	.w3(32'h3b9f1a38),
	.w4(32'hbc3bb6e1),
	.w5(32'hba349fe8),
	.w6(32'hbc095658),
	.w7(32'hbc876cc9),
	.w8(32'hbc0818f4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b6aba),
	.w1(32'h3c4bc12e),
	.w2(32'h3b866143),
	.w3(32'h3b966944),
	.w4(32'hbbdd0d5e),
	.w5(32'hbc71a348),
	.w6(32'h3a8cd639),
	.w7(32'h394324d1),
	.w8(32'hbc58df22),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c153f35),
	.w1(32'h399ffd60),
	.w2(32'hbac16ce7),
	.w3(32'hbaa5e30b),
	.w4(32'h3c6953c4),
	.w5(32'hbb15691a),
	.w6(32'h3b2213c7),
	.w7(32'h3bb255f8),
	.w8(32'hbabe91b5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a915f2c),
	.w1(32'h3a71a5a9),
	.w2(32'h3c652603),
	.w3(32'hbb2de756),
	.w4(32'h3c77b1c7),
	.w5(32'h3cc930ad),
	.w6(32'hba7031fa),
	.w7(32'hba6f5771),
	.w8(32'h3c184c12),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c49eb),
	.w1(32'hbbabcd80),
	.w2(32'hba4fcbc6),
	.w3(32'h3c2e487a),
	.w4(32'hbbe8720d),
	.w5(32'h3940d61d),
	.w6(32'h3a37101f),
	.w7(32'h3b8104c4),
	.w8(32'h3c1c923e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4f8c),
	.w1(32'h3b07d0ac),
	.w2(32'h3bbc7b8e),
	.w3(32'h3be17cd4),
	.w4(32'hbc35b3d9),
	.w5(32'h3b1e0d71),
	.w6(32'h3c4fb756),
	.w7(32'hbc39a69d),
	.w8(32'hbc023a36),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a67ca),
	.w1(32'hbb4e006b),
	.w2(32'hbaab513c),
	.w3(32'hbafabffa),
	.w4(32'hbb753602),
	.w5(32'hb9947220),
	.w6(32'hbb9323a0),
	.w7(32'hbb521da1),
	.w8(32'hba0ee1ed),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01cc08),
	.w1(32'hbcd0be2c),
	.w2(32'hbce709bb),
	.w3(32'h3c28e232),
	.w4(32'hbca44184),
	.w5(32'hbca704b1),
	.w6(32'h3b675b73),
	.w7(32'hbb82523b),
	.w8(32'hbc45ca1a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7070da),
	.w1(32'hbbe3e89a),
	.w2(32'hbbbc5d59),
	.w3(32'hbbb0b8e3),
	.w4(32'hbbc6eaf9),
	.w5(32'hbc5bd6c4),
	.w6(32'hbc1bd3b8),
	.w7(32'hbc0b5a9a),
	.w8(32'hbc322ce8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2d77a),
	.w1(32'hbb25b711),
	.w2(32'h3ae46457),
	.w3(32'hbb8d1b5c),
	.w4(32'hbc10a3c2),
	.w5(32'hbac7d1c5),
	.w6(32'hbaf7709a),
	.w7(32'hbc5d225c),
	.w8(32'hbbe6086d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a23ea),
	.w1(32'hbb63ca31),
	.w2(32'hb9feb2ed),
	.w3(32'h3c161d86),
	.w4(32'hbc02c8b0),
	.w5(32'hbb3147c8),
	.w6(32'h3c10521a),
	.w7(32'hbbe953ce),
	.w8(32'hbbb13a3c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a288f),
	.w1(32'hba1d8564),
	.w2(32'hba2c6f6c),
	.w3(32'h38bb811f),
	.w4(32'h3a22f554),
	.w5(32'h3a84babf),
	.w6(32'h3a4e5496),
	.w7(32'h392e6987),
	.w8(32'hb9dd9620),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03c100),
	.w1(32'h3a3c7a2d),
	.w2(32'h38394681),
	.w3(32'hba649392),
	.w4(32'h397beb9f),
	.w5(32'hba0c307f),
	.w6(32'hba58586e),
	.w7(32'hbab454f0),
	.w8(32'hba6f5fb3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba33bd),
	.w1(32'hba4cf901),
	.w2(32'hba344341),
	.w3(32'hbacbea7e),
	.w4(32'hb830d2da),
	.w5(32'h3a76a254),
	.w6(32'hbaacbef9),
	.w7(32'hba7ce2e2),
	.w8(32'h3a283b74),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51053b),
	.w1(32'h3a8e9afc),
	.w2(32'h3ab7e88a),
	.w3(32'h3ab0e9b0),
	.w4(32'h3aa725e7),
	.w5(32'h3b0a57c0),
	.w6(32'h3b264eda),
	.w7(32'h3a8c7152),
	.w8(32'hba8cbad8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6adf0b),
	.w1(32'h3a19beb7),
	.w2(32'h3a85e295),
	.w3(32'hb8b86228),
	.w4(32'h39e5daa1),
	.w5(32'h3b204b4c),
	.w6(32'hba837ae4),
	.w7(32'hba6e5f76),
	.w8(32'h3a738e59),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d7810),
	.w1(32'h3b686c86),
	.w2(32'h3b281097),
	.w3(32'h3b892e5f),
	.w4(32'h3b3ba482),
	.w5(32'h3af621bd),
	.w6(32'hbb20c901),
	.w7(32'h3b06554d),
	.w8(32'h3b0796de),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbed9f),
	.w1(32'h3bdfaa5f),
	.w2(32'h3b1b8c0d),
	.w3(32'h3bc934fc),
	.w4(32'h3b934253),
	.w5(32'h3ab90c19),
	.w6(32'hbb8fb9e6),
	.w7(32'h3984f1dc),
	.w8(32'h3a24fbf9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32d32c),
	.w1(32'hbb2a57a9),
	.w2(32'h3a23f140),
	.w3(32'hba51704f),
	.w4(32'hbb950497),
	.w5(32'hbb58397b),
	.w6(32'h3b0fa563),
	.w7(32'hbb78c4f6),
	.w8(32'hbb5c16d6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac9c15),
	.w1(32'h39ec539c),
	.w2(32'hb9887e5c),
	.w3(32'hba45566e),
	.w4(32'h3a0dac6b),
	.w5(32'hb9a59984),
	.w6(32'hbb2142e7),
	.w7(32'h3a314c8e),
	.w8(32'hba629b93),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a903bcb),
	.w1(32'hba0bcc74),
	.w2(32'hbb0f76ca),
	.w3(32'h3b9e1525),
	.w4(32'h3af6b673),
	.w5(32'h3b133019),
	.w6(32'h3b351483),
	.w7(32'hb9b8b4d8),
	.w8(32'hbad6d945),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5823c),
	.w1(32'h3a41f580),
	.w2(32'h3b8a5ca1),
	.w3(32'h3a8a7e79),
	.w4(32'hb79d13d4),
	.w5(32'h3a75d8af),
	.w6(32'h3b0af0e4),
	.w7(32'h3b046bb9),
	.w8(32'h3b00f829),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7a74b),
	.w1(32'h39aa9160),
	.w2(32'h390bb5b9),
	.w3(32'h3bd4719f),
	.w4(32'h3aa99156),
	.w5(32'h3a5230cb),
	.w6(32'h3b7f3c3a),
	.w7(32'h38caee2a),
	.w8(32'hba9bc222),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e98ae),
	.w1(32'h397a50ed),
	.w2(32'h3a5969e5),
	.w3(32'h398362d0),
	.w4(32'hba199cc5),
	.w5(32'hb9cddb51),
	.w6(32'h39d4496d),
	.w7(32'h39705479),
	.w8(32'h37bf0d28),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e53e31),
	.w1(32'hba87a8bb),
	.w2(32'hba959b89),
	.w3(32'h3a5f2d9c),
	.w4(32'hba4bb2b4),
	.w5(32'h3a58eff7),
	.w6(32'h3aaa2ce0),
	.w7(32'h3996318f),
	.w8(32'hbb10deb0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3afc92),
	.w1(32'hbac98514),
	.w2(32'hbae77a1c),
	.w3(32'hbad5518b),
	.w4(32'hb9f57e60),
	.w5(32'hbabf6527),
	.w6(32'hbb489d1d),
	.w7(32'h39fc5b89),
	.w8(32'hba77947b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed7632),
	.w1(32'hbab82542),
	.w2(32'hba2bb24f),
	.w3(32'hba9cde2b),
	.w4(32'h3a11870e),
	.w5(32'h3aab0095),
	.w6(32'h3a1dd517),
	.w7(32'h39b403b2),
	.w8(32'hbaa65062),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c0e55),
	.w1(32'hbb51ec57),
	.w2(32'hbab44f5a),
	.w3(32'hbbdf6437),
	.w4(32'hbba4fd89),
	.w5(32'hbb8d1a99),
	.w6(32'hbb586c31),
	.w7(32'hbb5b8c66),
	.w8(32'hbb27f0fb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d12a1),
	.w1(32'h36bfff46),
	.w2(32'hba4c8e0c),
	.w3(32'hba426ba6),
	.w4(32'hba08f8e6),
	.w5(32'h3ada0da9),
	.w6(32'hbb28ca7f),
	.w7(32'hba91bb59),
	.w8(32'hba8dd6b6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba052199),
	.w1(32'h3b062fbe),
	.w2(32'h3917444c),
	.w3(32'hbbbdb95c),
	.w4(32'hbb4532a5),
	.w5(32'hb9b1519c),
	.w6(32'hbbbc3f0f),
	.w7(32'hbb8ea5d5),
	.w8(32'hbad6c362),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117c97),
	.w1(32'h3b198c0d),
	.w2(32'h3a9a67a9),
	.w3(32'h3ba8280b),
	.w4(32'h38c0d66f),
	.w5(32'h38dcd7c9),
	.w6(32'hbb4b7d90),
	.w7(32'hbb65707c),
	.w8(32'hbb4dc264),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cbbb4),
	.w1(32'hbb0ab811),
	.w2(32'hb87a7985),
	.w3(32'h3a924ca1),
	.w4(32'hba006a51),
	.w5(32'hba035266),
	.w6(32'h3b0e0e3a),
	.w7(32'h3a36e8aa),
	.w8(32'hbab2deaa),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b970299),
	.w1(32'h3ade2b7a),
	.w2(32'hbbb50797),
	.w3(32'h3b48ceb9),
	.w4(32'h3a98724a),
	.w5(32'hb9c718c6),
	.w6(32'hba4a6ca9),
	.w7(32'hbbc94171),
	.w8(32'hbb98ece0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e2ac2),
	.w1(32'h3a2be728),
	.w2(32'h3a285d6a),
	.w3(32'hba72de0c),
	.w4(32'hba761fc2),
	.w5(32'hbb13505f),
	.w6(32'h3a3746da),
	.w7(32'hba7a95c2),
	.w8(32'hbb67c2b6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9558ae),
	.w1(32'h3af48c8a),
	.w2(32'hba67ea57),
	.w3(32'h3a28b19e),
	.w4(32'h3a627216),
	.w5(32'hbb05439d),
	.w6(32'hbba7cad5),
	.w7(32'hbb2f6bbc),
	.w8(32'hbb948612),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab8add),
	.w1(32'hbb22578e),
	.w2(32'hbb404730),
	.w3(32'hba8f03e3),
	.w4(32'h396f4a8c),
	.w5(32'hb8bad5e5),
	.w6(32'h3964c766),
	.w7(32'hbb815f80),
	.w8(32'hbbd105be),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52aed),
	.w1(32'hba9ff9b9),
	.w2(32'h3a0b1ac9),
	.w3(32'h3b5cdd54),
	.w4(32'h3aab018d),
	.w5(32'h3b59dbd5),
	.w6(32'h3acfbc6e),
	.w7(32'hbace562f),
	.w8(32'hbb7ba3af),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93efb69),
	.w1(32'h3a7ebc96),
	.w2(32'hb9d6bdb4),
	.w3(32'hbaffc61d),
	.w4(32'h39b784a2),
	.w5(32'h3adc8c00),
	.w6(32'h391173aa),
	.w7(32'h39801b8b),
	.w8(32'hbb0798a2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba235fc),
	.w1(32'hb9e11928),
	.w2(32'h3aeaa499),
	.w3(32'h3b350b33),
	.w4(32'hb9c1042c),
	.w5(32'h3a408f6b),
	.w6(32'hbb0c6e01),
	.w7(32'hbb80fd14),
	.w8(32'hbb9a70ba),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8edfa2),
	.w1(32'hba0cb5a2),
	.w2(32'hbb81b33a),
	.w3(32'h3b50c8a8),
	.w4(32'hba0a2696),
	.w5(32'hbb8c5562),
	.w6(32'hb9fe75d7),
	.w7(32'hbb97d9e3),
	.w8(32'hbbd5157b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beffa18),
	.w1(32'h3c49867c),
	.w2(32'h3c02b7af),
	.w3(32'hbb48f8de),
	.w4(32'h3b8e3b5f),
	.w5(32'h391ed2f9),
	.w6(32'hbbd7a9bc),
	.w7(32'h37ebf75c),
	.w8(32'hbaa05139),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb454996),
	.w1(32'h3a6b9fed),
	.w2(32'hbb4e67ed),
	.w3(32'hb996c962),
	.w4(32'h3a5721eb),
	.w5(32'hbaf0504c),
	.w6(32'hb8058a5e),
	.w7(32'h3b440d0f),
	.w8(32'h38ca1c5a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803a5a),
	.w1(32'hbaf6cde5),
	.w2(32'hba8adc57),
	.w3(32'hbb9fa0b9),
	.w4(32'hbbb00be2),
	.w5(32'hbb31d5ab),
	.w6(32'hbad6a504),
	.w7(32'hbb897b6a),
	.w8(32'hbbf07265),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc38c7),
	.w1(32'h3b7fa472),
	.w2(32'hbb30b847),
	.w3(32'h3b05222c),
	.w4(32'h3b9a5e79),
	.w5(32'h3afbbf62),
	.w6(32'hbb8fc672),
	.w7(32'hbaaa1d98),
	.w8(32'h3a4679c8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7edb7e),
	.w1(32'hba7feff1),
	.w2(32'h3a2f02ae),
	.w3(32'hbaa35f29),
	.w4(32'hb9b55307),
	.w5(32'hba269506),
	.w6(32'h39a7e636),
	.w7(32'h39ad666a),
	.w8(32'hbae7aa84),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f8ac7),
	.w1(32'h3be32da2),
	.w2(32'h3a9c0446),
	.w3(32'hbaef72a0),
	.w4(32'h3b4fe59c),
	.w5(32'hbbf0c7a2),
	.w6(32'hbc5ee645),
	.w7(32'hbb993f6b),
	.w8(32'h3ba4e9e5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c9e69),
	.w1(32'hbb3cac01),
	.w2(32'hbb4278eb),
	.w3(32'hbada0d25),
	.w4(32'hbb125b76),
	.w5(32'hbb098440),
	.w6(32'h3a9eea05),
	.w7(32'hb91fe105),
	.w8(32'h3b1cba17),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07a43c),
	.w1(32'h3a27fa7c),
	.w2(32'h3aa6955b),
	.w3(32'h3a816087),
	.w4(32'h3abdc0f6),
	.w5(32'h3965690e),
	.w6(32'h3aad45bf),
	.w7(32'h3ab1601f),
	.w8(32'h3a07e98b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a464922),
	.w1(32'h3b0ba25b),
	.w2(32'h3b04c7e1),
	.w3(32'hbb49032b),
	.w4(32'hbae16268),
	.w5(32'hb9943d0d),
	.w6(32'hba1edbd4),
	.w7(32'hbb6ec3a2),
	.w8(32'hbb13d938),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacf3f2),
	.w1(32'hbb11fd38),
	.w2(32'hbb0fdd05),
	.w3(32'h3ad81b7e),
	.w4(32'hbadc3167),
	.w5(32'hbb2cee09),
	.w6(32'h39bbd6cc),
	.w7(32'hbb5374fc),
	.w8(32'hbb4f4141),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafddf68),
	.w1(32'hbb49a4c5),
	.w2(32'h3a85b5e7),
	.w3(32'hbb635e66),
	.w4(32'hbb51a91e),
	.w5(32'hbacf2d7f),
	.w6(32'h39b11ed7),
	.w7(32'hba84d329),
	.w8(32'hbb004cbd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaee8c8),
	.w1(32'hbb43158f),
	.w2(32'h3b01ff90),
	.w3(32'h3aaf1c88),
	.w4(32'h3a4c7d86),
	.w5(32'hbabf4a86),
	.w6(32'h3bc4ec3f),
	.w7(32'hbaf9e11b),
	.w8(32'hbae587fa),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acddd30),
	.w1(32'hba94d260),
	.w2(32'h39e5ffcf),
	.w3(32'hbae59baa),
	.w4(32'hbb13db79),
	.w5(32'hba2bbc2e),
	.w6(32'hba8a2a2e),
	.w7(32'hbaaf8d54),
	.w8(32'hbb64adb6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1feffc),
	.w1(32'h3c0b81c4),
	.w2(32'h3b852465),
	.w3(32'hbb40c731),
	.w4(32'h3b02f2d5),
	.w5(32'h3baae714),
	.w6(32'hbbeaf123),
	.w7(32'hbb4b3afa),
	.w8(32'hbb962812),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34e78d),
	.w1(32'h3b166fa5),
	.w2(32'h3a5cf011),
	.w3(32'h3a88e985),
	.w4(32'h3a1db5d4),
	.w5(32'h3b1bf1fb),
	.w6(32'h3aa1d2b5),
	.w7(32'hb9a4b6ea),
	.w8(32'h3a6e6691),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6dede),
	.w1(32'h39693235),
	.w2(32'h3a3dd96a),
	.w3(32'hbaea072f),
	.w4(32'hbb5b11e2),
	.w5(32'hba8f64c2),
	.w6(32'hbacd8fe2),
	.w7(32'hbb7dac17),
	.w8(32'hbb4cc559),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb8631),
	.w1(32'hb90488d5),
	.w2(32'hbabaf0c2),
	.w3(32'h3a38a366),
	.w4(32'h3a44e29b),
	.w5(32'hba670540),
	.w6(32'h39f2ac08),
	.w7(32'hb855c957),
	.w8(32'hba4f99da),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad7e7e),
	.w1(32'hb9e7bedc),
	.w2(32'hb85cf153),
	.w3(32'h3a9d5804),
	.w4(32'hbaa09a17),
	.w5(32'hbac94ff0),
	.w6(32'h3aa674ff),
	.w7(32'h39c1ed94),
	.w8(32'hbaefb750),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efe020),
	.w1(32'h390cf7c2),
	.w2(32'h3a629825),
	.w3(32'hba3b1f90),
	.w4(32'hb9bca6c6),
	.w5(32'hbac7a455),
	.w6(32'hb89f2276),
	.w7(32'hba986816),
	.w8(32'hb8bd0cc8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30ae90),
	.w1(32'hb9b01fc3),
	.w2(32'h3992238f),
	.w3(32'h3a76b6dd),
	.w4(32'hb9ab0a09),
	.w5(32'h3a621861),
	.w6(32'h3ad72a6a),
	.w7(32'h39c147ec),
	.w8(32'h3a7b753b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f10f6),
	.w1(32'hba8587d7),
	.w2(32'hb9db18d4),
	.w3(32'hbb2c16fe),
	.w4(32'hbb6217b7),
	.w5(32'h3a076332),
	.w6(32'hbafc215a),
	.w7(32'hbbbe8eba),
	.w8(32'hbb9366ca),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f010f7),
	.w1(32'h3b3186d7),
	.w2(32'h3a10b6a8),
	.w3(32'h3ad9d337),
	.w4(32'h3ae2267e),
	.w5(32'h3ab9e0a7),
	.w6(32'h3a105790),
	.w7(32'h3abb3315),
	.w8(32'h3ade6d62),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f2796),
	.w1(32'h3b2d8582),
	.w2(32'hbaafd990),
	.w3(32'h3bf7ce1f),
	.w4(32'h3b59dacc),
	.w5(32'h3ab05c2c),
	.w6(32'h3b5a3fe6),
	.w7(32'hbad72477),
	.w8(32'hbb1746a7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba40cd6),
	.w1(32'hbabbd9c6),
	.w2(32'hba804283),
	.w3(32'hbb8c927b),
	.w4(32'hbadcda86),
	.w5(32'hb9f97f36),
	.w6(32'h3a4e60ee),
	.w7(32'hba8292ac),
	.w8(32'hbb456f0d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f9add),
	.w1(32'hb9b9743b),
	.w2(32'hb9cd4971),
	.w3(32'hba9d5299),
	.w4(32'hb8c2c824),
	.w5(32'hb894e748),
	.w6(32'h3a745eac),
	.w7(32'h3afc6a6b),
	.w8(32'hbb114968),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68cb2c),
	.w1(32'h380a9e67),
	.w2(32'hba6247e5),
	.w3(32'hba607d41),
	.w4(32'hbab67ee8),
	.w5(32'hbabeed54),
	.w6(32'hbaa4a36a),
	.w7(32'hbac8e333),
	.w8(32'hbacadd63),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b97a7f),
	.w1(32'h39967e22),
	.w2(32'h3a77734f),
	.w3(32'hbb21abe1),
	.w4(32'h3a305d34),
	.w5(32'h39ad55e3),
	.w6(32'hbabf5f80),
	.w7(32'hba09ff9b),
	.w8(32'hba743e87),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b38e4b),
	.w1(32'hbafbf501),
	.w2(32'hb9b8a176),
	.w3(32'hbb0b33bd),
	.w4(32'hbab9c20f),
	.w5(32'h3aad9ee8),
	.w6(32'hba3a4fa4),
	.w7(32'hbaa1537b),
	.w8(32'hba30a9cd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b778ac7),
	.w1(32'h3bdf8b61),
	.w2(32'h3bc2332a),
	.w3(32'h3b07ee12),
	.w4(32'h3b815e49),
	.w5(32'h3c2e2e16),
	.w6(32'hbc05146d),
	.w7(32'hbb4b1a33),
	.w8(32'hbade8409),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1313c8),
	.w1(32'hba57291d),
	.w2(32'h39a86a5a),
	.w3(32'h3b24cfcb),
	.w4(32'h3b066dec),
	.w5(32'h3ac72150),
	.w6(32'hba2fda81),
	.w7(32'h39b3444b),
	.w8(32'hb9d0d541),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b196af5),
	.w1(32'hb999d4a3),
	.w2(32'h398fa091),
	.w3(32'h3b02acfa),
	.w4(32'h39175095),
	.w5(32'hb9b2d063),
	.w6(32'h3b1dd28f),
	.w7(32'hba806b74),
	.w8(32'hba4837c0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399984a9),
	.w1(32'hb9909fbb),
	.w2(32'h3a413f6a),
	.w3(32'hbaf0e533),
	.w4(32'hbad4acb1),
	.w5(32'hba578dd2),
	.w6(32'hbb5edd89),
	.w7(32'hb8891740),
	.w8(32'hba692b62),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef62d6),
	.w1(32'h396ac38f),
	.w2(32'hb84a906e),
	.w3(32'h39e37811),
	.w4(32'hb992d88f),
	.w5(32'hbaab66a2),
	.w6(32'hba095004),
	.w7(32'hbb56214d),
	.w8(32'hbb6a0893),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80eff7),
	.w1(32'hba4dbc7e),
	.w2(32'h3ad0db73),
	.w3(32'hba7cd1f8),
	.w4(32'hb99a9eb3),
	.w5(32'hba29cc79),
	.w6(32'hbac9730e),
	.w7(32'hbafc503d),
	.w8(32'hbb31205c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fd017),
	.w1(32'hba2fd205),
	.w2(32'hb8c35e70),
	.w3(32'hbb0d0e0c),
	.w4(32'hbadf927c),
	.w5(32'h39999e7d),
	.w6(32'hb8ce5e76),
	.w7(32'hba9b13ba),
	.w8(32'hbb18b12f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb4293),
	.w1(32'h3bad66f4),
	.w2(32'h3b544247),
	.w3(32'h3be8baab),
	.w4(32'h3b9ac212),
	.w5(32'h3bbc3de0),
	.w6(32'hba6f9efe),
	.w7(32'h3b5b9a37),
	.w8(32'hba45cab8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb4181),
	.w1(32'hbb20caa0),
	.w2(32'hba0315c3),
	.w3(32'hbad5b0fc),
	.w4(32'hba2b4da7),
	.w5(32'hbaa5babb),
	.w6(32'h3a2faca9),
	.w7(32'h3a20beb0),
	.w8(32'hb9eb2438),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cc456),
	.w1(32'h3a244542),
	.w2(32'hb9dd1c09),
	.w3(32'h3af7f0d7),
	.w4(32'h3b1c1297),
	.w5(32'h3a6c7240),
	.w6(32'hbab3ea7e),
	.w7(32'hba7f4193),
	.w8(32'hbb79eea4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0545c2),
	.w1(32'h3ba02b49),
	.w2(32'h3b44beda),
	.w3(32'h3bdaff4c),
	.w4(32'h3b40575f),
	.w5(32'h3acf8086),
	.w6(32'hbb35892c),
	.w7(32'h3a577991),
	.w8(32'hba33917d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92ca4e),
	.w1(32'h3b06bda7),
	.w2(32'h3a8b8bae),
	.w3(32'hbbb2fcc2),
	.w4(32'hba56fc9b),
	.w5(32'hba8377be),
	.w6(32'hbb6ad723),
	.w7(32'hbb57f30a),
	.w8(32'hbb8f299a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a923662),
	.w1(32'hb998e25f),
	.w2(32'hbaf959ca),
	.w3(32'h3a152876),
	.w4(32'hba655155),
	.w5(32'hba4be460),
	.w6(32'hb814f3fb),
	.w7(32'h39d4ffed),
	.w8(32'hba6936b5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f20e8),
	.w1(32'h3a5336bd),
	.w2(32'h3b16c6d5),
	.w3(32'h3b4788cf),
	.w4(32'h3a062be3),
	.w5(32'h3b3da706),
	.w6(32'h3aae4af1),
	.w7(32'hb9ee321e),
	.w8(32'hb9d2f741),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10dc88),
	.w1(32'hbb09266b),
	.w2(32'hbb1e8a42),
	.w3(32'h3b09e0c7),
	.w4(32'hb996c675),
	.w5(32'hb93b7997),
	.w6(32'h3bc95811),
	.w7(32'h3b2ae198),
	.w8(32'h3a066273),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a035a40),
	.w1(32'hba51b830),
	.w2(32'hba997812),
	.w3(32'h3a682be3),
	.w4(32'hbaa60e9f),
	.w5(32'hbb22fb0e),
	.w6(32'h3828dd74),
	.w7(32'hbb127d45),
	.w8(32'hbb9a6599),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae7ccc),
	.w1(32'hba05984e),
	.w2(32'h3a02b6e0),
	.w3(32'hbab12961),
	.w4(32'h3998c3aa),
	.w5(32'hba0c7587),
	.w6(32'hba78173e),
	.w7(32'hb86a2355),
	.w8(32'hb9c3c12b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a800e54),
	.w1(32'hb9aa885d),
	.w2(32'h39153d97),
	.w3(32'h3a3658c2),
	.w4(32'h399744e6),
	.w5(32'hb9f3ea28),
	.w6(32'hb985caaf),
	.w7(32'h3980a840),
	.w8(32'h38af6533),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadd408),
	.w1(32'hb8c65adb),
	.w2(32'h3acefe13),
	.w3(32'hba228909),
	.w4(32'h3a24e11b),
	.w5(32'h3a8d4d8c),
	.w6(32'h3a153435),
	.w7(32'hba76f34c),
	.w8(32'h3abd86e9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf7cb0),
	.w1(32'hba9912d7),
	.w2(32'hbb18f3c1),
	.w3(32'hb96c5e27),
	.w4(32'hbafa5af9),
	.w5(32'hbafc4e3f),
	.w6(32'h3ae1274f),
	.w7(32'hbabb7b68),
	.w8(32'hbb5236a0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04e18d),
	.w1(32'h3ad9573f),
	.w2(32'h3a005882),
	.w3(32'h3abbc8d2),
	.w4(32'h3a2c8155),
	.w5(32'h3a6316f2),
	.w6(32'hbb3beea1),
	.w7(32'hbb17090c),
	.w8(32'hbb6acde5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e468f),
	.w1(32'h3a0c8dbd),
	.w2(32'h3869b7a9),
	.w3(32'hba74f901),
	.w4(32'h3a81f616),
	.w5(32'hb8f147a9),
	.w6(32'hba1a82b7),
	.w7(32'h3a3018d9),
	.w8(32'hba8eb1e5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3128d8),
	.w1(32'hbb8b0bde),
	.w2(32'hbb2ddc39),
	.w3(32'h3b1cc146),
	.w4(32'hbb8439f4),
	.w5(32'hbabd9255),
	.w6(32'h392d5b5d),
	.w7(32'hbba1ceee),
	.w8(32'hbb63f299),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5525ed),
	.w1(32'hb9f06a06),
	.w2(32'hbab0e52a),
	.w3(32'hba717616),
	.w4(32'hbb250a5a),
	.w5(32'hbab5bf50),
	.w6(32'hbae0daf2),
	.w7(32'hbaa29eda),
	.w8(32'hbb5f88f3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b711e),
	.w1(32'h3bc1d084),
	.w2(32'h3a4e03b7),
	.w3(32'h3b890910),
	.w4(32'h3b5d4b51),
	.w5(32'h39ac90d5),
	.w6(32'hbaf802b8),
	.w7(32'hbb62129f),
	.w8(32'hbba3f9dc),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab21e1),
	.w1(32'hbb9d2cb0),
	.w2(32'h3ae3ec82),
	.w3(32'hba4260ce),
	.w4(32'hbbb87acd),
	.w5(32'hbb05af3f),
	.w6(32'h3b32e801),
	.w7(32'hbb4fb5e1),
	.w8(32'hbbaa0c4c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb323b3e),
	.w1(32'h3abdd341),
	.w2(32'h3aa3853a),
	.w3(32'hbb3796bd),
	.w4(32'h3a8d55ac),
	.w5(32'h3a699b29),
	.w6(32'hbb21c5ee),
	.w7(32'h38c06082),
	.w8(32'hba3d4e2b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ceb07a),
	.w1(32'hba7d349f),
	.w2(32'hba036cba),
	.w3(32'hb8e006c8),
	.w4(32'hb93405ad),
	.w5(32'h3b550009),
	.w6(32'hba750298),
	.w7(32'h3a6e4223),
	.w8(32'h3a12efd7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a26ed),
	.w1(32'hb7aa0585),
	.w2(32'hbb280974),
	.w3(32'hbb12e1ef),
	.w4(32'hbab8d62b),
	.w5(32'hbb38574c),
	.w6(32'hbae26306),
	.w7(32'hbb22bf47),
	.w8(32'hbb915aaf),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7be77),
	.w1(32'h38c11a8a),
	.w2(32'hb98b1021),
	.w3(32'hbb37db17),
	.w4(32'hba80e26a),
	.w5(32'hbaf1f844),
	.w6(32'hba6628dd),
	.w7(32'hbaf15dd1),
	.w8(32'hbb6fd547),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e1ee8),
	.w1(32'hbad6b0b2),
	.w2(32'hba19047e),
	.w3(32'hbb6fbbf1),
	.w4(32'hba2d3b46),
	.w5(32'hba97a8e0),
	.w6(32'hbae54401),
	.w7(32'h3a8f5f51),
	.w8(32'hb79c42c4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69cd2d),
	.w1(32'h3a26a177),
	.w2(32'hb9538b19),
	.w3(32'h3b3f42c0),
	.w4(32'hb90f80b4),
	.w5(32'h39e21064),
	.w6(32'hb9ad2444),
	.w7(32'hba59eb21),
	.w8(32'h3abde48d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9228927),
	.w1(32'hbab6e3c4),
	.w2(32'h383f342b),
	.w3(32'hb7ec9263),
	.w4(32'hba687b94),
	.w5(32'hb9ea93cd),
	.w6(32'h398bf3a5),
	.w7(32'hba4655ac),
	.w8(32'hba1cdfb7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d67a),
	.w1(32'h3a4cc56b),
	.w2(32'h39dc6130),
	.w3(32'h3bb94c6b),
	.w4(32'h38fd292d),
	.w5(32'h390ae806),
	.w6(32'hba75f901),
	.w7(32'hb9a272ec),
	.w8(32'hba78d80f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ec117),
	.w1(32'h3961eb5c),
	.w2(32'hba7c6b0e),
	.w3(32'hbaf55c63),
	.w4(32'hb9226677),
	.w5(32'h396af0c1),
	.w6(32'hb9517a46),
	.w7(32'h39d78eb2),
	.w8(32'hbad1970d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58340f),
	.w1(32'hbb024fdd),
	.w2(32'hb98bf945),
	.w3(32'hbaa0e2e7),
	.w4(32'hbb7bf28e),
	.w5(32'hbb11f0de),
	.w6(32'hb962f56f),
	.w7(32'hbb278b2d),
	.w8(32'hba9479aa),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5b461),
	.w1(32'hb8994dfc),
	.w2(32'h383aa65b),
	.w3(32'hb83ba42d),
	.w4(32'h3a9e2b30),
	.w5(32'h39be711e),
	.w6(32'h3ade39aa),
	.w7(32'h3a17be71),
	.w8(32'h3aa19d62),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b3f45),
	.w1(32'hba1be27c),
	.w2(32'hba8466df),
	.w3(32'h3b5d3a3b),
	.w4(32'h3b0f649d),
	.w5(32'h3b6e79c0),
	.w6(32'hba5e11ae),
	.w7(32'h3ac29721),
	.w8(32'hba432b99),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ba6e3),
	.w1(32'hb9b24973),
	.w2(32'h3a1cf13e),
	.w3(32'hbad4d89f),
	.w4(32'hba178ef4),
	.w5(32'h39fc897b),
	.w6(32'h3823c338),
	.w7(32'h3a17cce3),
	.w8(32'h3b0688bb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92696f),
	.w1(32'h3a550b54),
	.w2(32'h3a3bfb1c),
	.w3(32'h3a7c72e4),
	.w4(32'h3a8841ba),
	.w5(32'h3a71da9f),
	.w6(32'h382f9ea8),
	.w7(32'h39fa38ae),
	.w8(32'hb9ddf05a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa96992),
	.w1(32'hbaf5e61f),
	.w2(32'hbadeb2e1),
	.w3(32'h3b172e89),
	.w4(32'hba1e9efd),
	.w5(32'hbb141d31),
	.w6(32'h3b637c34),
	.w7(32'hba5281a3),
	.w8(32'hbb61e5bd),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8524c9),
	.w1(32'h3bcdd649),
	.w2(32'h3b1970f5),
	.w3(32'h3b823645),
	.w4(32'h3b97c3b2),
	.w5(32'h3bc3d4a9),
	.w6(32'hbb99eb6f),
	.w7(32'hbb5e35d4),
	.w8(32'hbb73b289),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98544f6),
	.w1(32'h3a4d6dcc),
	.w2(32'hbaa8ecb3),
	.w3(32'h3aa3d26d),
	.w4(32'hb95625f9),
	.w5(32'h3a1566aa),
	.w6(32'hb820e81b),
	.w7(32'hba732522),
	.w8(32'hbb1586ca),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba141c0c),
	.w1(32'hbb02b256),
	.w2(32'h39645780),
	.w3(32'hba006125),
	.w4(32'hbaff9e7a),
	.w5(32'hb8fd6034),
	.w6(32'h396e6733),
	.w7(32'hbb53141e),
	.w8(32'hbacb6e28),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e5829),
	.w1(32'hba16af35),
	.w2(32'h3acfcbd5),
	.w3(32'hb9b331a5),
	.w4(32'h3a1bd944),
	.w5(32'hb9f68f48),
	.w6(32'h3a7da506),
	.w7(32'h38ffcf20),
	.w8(32'hb9b21418),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cc9e0),
	.w1(32'hba96ee50),
	.w2(32'h3b121822),
	.w3(32'hb8e5830b),
	.w4(32'hbb1c37c9),
	.w5(32'h3b855a29),
	.w6(32'hba198104),
	.w7(32'hb7de7aca),
	.w8(32'hbaefb068),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a8f73),
	.w1(32'h3a9a1c3f),
	.w2(32'hb939d027),
	.w3(32'h3b430d5f),
	.w4(32'h390303e8),
	.w5(32'hba0a8967),
	.w6(32'hbafaeba3),
	.w7(32'hbb667826),
	.w8(32'hbb5ff736),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b291f07),
	.w1(32'h39ec695a),
	.w2(32'h395b3473),
	.w3(32'h3b179338),
	.w4(32'h3ab03a4f),
	.w5(32'h3b06ded1),
	.w6(32'hbb573735),
	.w7(32'hbab944c7),
	.w8(32'hbb4ee144),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ec180),
	.w1(32'hba8f5bc4),
	.w2(32'hb8b62c31),
	.w3(32'hbae54e30),
	.w4(32'h39c3aa3f),
	.w5(32'h3ab2927f),
	.w6(32'h39727934),
	.w7(32'h398837cb),
	.w8(32'h39eabff3),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d75417),
	.w1(32'hb99f673a),
	.w2(32'h3a09e0a4),
	.w3(32'h3b3b2d79),
	.w4(32'hb8b714a1),
	.w5(32'hb935d3d1),
	.w6(32'h3ae1bba9),
	.w7(32'h3aa8845e),
	.w8(32'hba81d369),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68a088),
	.w1(32'h39a1c380),
	.w2(32'hbab8142d),
	.w3(32'h3937099f),
	.w4(32'hb9f3e938),
	.w5(32'hbb0633dd),
	.w6(32'hba9237ab),
	.w7(32'hba339a1d),
	.w8(32'hba9bcb45),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e5f7e),
	.w1(32'h39c7b22d),
	.w2(32'hb9ba8d96),
	.w3(32'h3b5150de),
	.w4(32'h3a149d77),
	.w5(32'hb9ab14e9),
	.w6(32'h3ae4037e),
	.w7(32'hbaf5771a),
	.w8(32'hbb3f9c30),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadca29d),
	.w1(32'hbaf41104),
	.w2(32'hbb082bea),
	.w3(32'hbaa92b8e),
	.w4(32'hbb00f0d5),
	.w5(32'hba1578ba),
	.w6(32'hba0ce938),
	.w7(32'hbac55707),
	.w8(32'hba8beaf2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59c458),
	.w1(32'hba4b0ebd),
	.w2(32'h398710b0),
	.w3(32'hb9a94679),
	.w4(32'hba8d85e1),
	.w5(32'h3a80ab44),
	.w6(32'hbb19450e),
	.w7(32'h3a87ebc8),
	.w8(32'hb9f3cb84),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab590b6),
	.w1(32'hba44bf98),
	.w2(32'h386f42ea),
	.w3(32'h3adae64b),
	.w4(32'h3a05455e),
	.w5(32'hba539ae7),
	.w6(32'hb9bf2502),
	.w7(32'h3acf8c70),
	.w8(32'h3ab1de2f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a291146),
	.w1(32'hba897d02),
	.w2(32'hbaa19a4e),
	.w3(32'hba6d74b6),
	.w4(32'hb9840f92),
	.w5(32'hb9c670d5),
	.w6(32'hb90d8912),
	.w7(32'hb8171e9f),
	.w8(32'h389a78fe),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2813b6),
	.w1(32'hbacbc3e8),
	.w2(32'h38cc6e17),
	.w3(32'hbb21de25),
	.w4(32'hbb29c113),
	.w5(32'hba6f909b),
	.w6(32'h3ab7b4ea),
	.w7(32'hba8ef5e8),
	.w8(32'hb9ade9e8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1f6c2),
	.w1(32'h3bac961e),
	.w2(32'h3a6aa9c4),
	.w3(32'hbab04030),
	.w4(32'h3a9fd597),
	.w5(32'h39e637a6),
	.w6(32'hbbb4a53c),
	.w7(32'hba4bf128),
	.w8(32'hbb976c83),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8206a7),
	.w1(32'h3b5216a5),
	.w2(32'h3a036e87),
	.w3(32'h3adece60),
	.w4(32'h3addcded),
	.w5(32'hba9c23b9),
	.w6(32'hbb69b939),
	.w7(32'hba98b8d1),
	.w8(32'hb8370860),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b28ae3),
	.w1(32'hb90164fa),
	.w2(32'hb9d67207),
	.w3(32'hb9bbb55d),
	.w4(32'hba26d7dc),
	.w5(32'hb90ef880),
	.w6(32'hbaf53ab4),
	.w7(32'hb9ceb119),
	.w8(32'hb9655ffc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a8c7a),
	.w1(32'h3b29cacd),
	.w2(32'h3b5fecbc),
	.w3(32'h3be13231),
	.w4(32'h3b1a3c64),
	.w5(32'h3b877220),
	.w6(32'hbb1f7d53),
	.w7(32'hbb881482),
	.w8(32'hbbbd97e2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba80977),
	.w1(32'hbc2134ca),
	.w2(32'hba13c1fc),
	.w3(32'hbb01ef5f),
	.w4(32'hbbfb35fc),
	.w5(32'hb9bf23e5),
	.w6(32'h3b9b4f8e),
	.w7(32'hbb7768df),
	.w8(32'hbbab3895),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999809d),
	.w1(32'h39c0c30a),
	.w2(32'hba5b9eac),
	.w3(32'h392e9d76),
	.w4(32'hb9b65ed8),
	.w5(32'hbab1c7f3),
	.w6(32'hba794380),
	.w7(32'h3a1cd014),
	.w8(32'hbaa39441),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ce76c),
	.w1(32'h3ab6d662),
	.w2(32'hba0193ca),
	.w3(32'hba310aeb),
	.w4(32'hb9866c1c),
	.w5(32'hb9c11462),
	.w6(32'h3a846c8d),
	.w7(32'hbb354c86),
	.w8(32'hbaee2f9d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1f609),
	.w1(32'hb921e8c2),
	.w2(32'hba4df94d),
	.w3(32'hbaacf6a6),
	.w4(32'h3a9e79bd),
	.w5(32'hb96927f8),
	.w6(32'hbb0dfc25),
	.w7(32'h390b054b),
	.w8(32'h38ae3246),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a50d5c),
	.w1(32'hb93d9200),
	.w2(32'h3ada935d),
	.w3(32'h3a745e57),
	.w4(32'h3a250d56),
	.w5(32'h39f91118),
	.w6(32'h3ad49fce),
	.w7(32'h3aac4450),
	.w8(32'h3afb7692),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dd2d8),
	.w1(32'h3b1481d8),
	.w2(32'h39e1b9c2),
	.w3(32'h3bc7eaaf),
	.w4(32'h3b6ef0e7),
	.w5(32'h3b8b9dbf),
	.w6(32'h3b27bab5),
	.w7(32'h3b58eb28),
	.w8(32'h3af39973),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49ec0e),
	.w1(32'hba90c101),
	.w2(32'hb9f8056d),
	.w3(32'h3b6cd964),
	.w4(32'h38a926ff),
	.w5(32'hba0086a6),
	.w6(32'hba5b56b3),
	.w7(32'hbb17b731),
	.w8(32'hbb3c9f31),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45d571),
	.w1(32'hb9bb716e),
	.w2(32'h3acb9802),
	.w3(32'hbb443c5b),
	.w4(32'hba21b13d),
	.w5(32'hb9e19671),
	.w6(32'hbb266b1f),
	.w7(32'hbadfd03b),
	.w8(32'hbaefae92),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eaa1f),
	.w1(32'hba57f382),
	.w2(32'hb6f45cdd),
	.w3(32'hbb35fbbd),
	.w4(32'hba2674bb),
	.w5(32'h391635ae),
	.w6(32'hbab8727b),
	.w7(32'hb9e075c1),
	.w8(32'hbad1c075),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c9de3),
	.w1(32'h3a858110),
	.w2(32'h37b652c8),
	.w3(32'h3b223f45),
	.w4(32'h3aafd0a1),
	.w5(32'h3a200f17),
	.w6(32'hbb6a33ff),
	.w7(32'hbb0857a8),
	.w8(32'hbb37641d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa379ab),
	.w1(32'h3ae096b6),
	.w2(32'h3a6636a2),
	.w3(32'hb93aea8a),
	.w4(32'hb91f0059),
	.w5(32'hb965c466),
	.w6(32'h38f87a3e),
	.w7(32'hb9746706),
	.w8(32'h3802d206),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bb57b1),
	.w1(32'hb73db7a1),
	.w2(32'h36c2d642),
	.w3(32'hb77c5207),
	.w4(32'hb72083bd),
	.w5(32'h36da3ae0),
	.w6(32'h3751b3ff),
	.w7(32'h377e6045),
	.w8(32'h380bec01),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bffc9),
	.w1(32'h39bc4ed1),
	.w2(32'hbac23317),
	.w3(32'h3a59ee3b),
	.w4(32'h3a389130),
	.w5(32'hbaa96358),
	.w6(32'hbb056ff3),
	.w7(32'hba31c901),
	.w8(32'h3b020a3e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aefa58),
	.w1(32'hb8156a75),
	.w2(32'h37c5a032),
	.w3(32'hb8764fa5),
	.w4(32'hb7ec9666),
	.w5(32'h382a7d04),
	.w6(32'h3837033e),
	.w7(32'h383d70b7),
	.w8(32'h38c7cc83),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b812ad8),
	.w1(32'h39178e92),
	.w2(32'hba507048),
	.w3(32'h3b501545),
	.w4(32'hb90c95bd),
	.w5(32'hba378f9e),
	.w6(32'hb873d062),
	.w7(32'hbb34f110),
	.w8(32'hbb4d0dd4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee2c67),
	.w1(32'h39ac24c1),
	.w2(32'h3ada0cf5),
	.w3(32'hbba4164f),
	.w4(32'hbb25661e),
	.w5(32'hbaef900d),
	.w6(32'h364e536c),
	.w7(32'hbaf7fda2),
	.w8(32'hbb154a5f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391fe5c1),
	.w1(32'h39d96e75),
	.w2(32'h3944b5a6),
	.w3(32'hba4b543b),
	.w4(32'hbaa1ae42),
	.w5(32'hbab795cd),
	.w6(32'hbab0af27),
	.w7(32'hbb304ef1),
	.w8(32'hbb5c1a0b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39921bd2),
	.w1(32'h39855866),
	.w2(32'hb99a6ff2),
	.w3(32'h3972f1e8),
	.w4(32'h396c57f9),
	.w5(32'hb9cb7028),
	.w6(32'h3991e82b),
	.w7(32'h39170917),
	.w8(32'hb9204bf9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99aba7),
	.w1(32'hba8e163a),
	.w2(32'h3ad90549),
	.w3(32'hbb0414f7),
	.w4(32'hbb1be574),
	.w5(32'hbad5bf98),
	.w6(32'hb79b5f40),
	.w7(32'hbb51d2fb),
	.w8(32'hbb678fff),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7f23d),
	.w1(32'h39c94ac7),
	.w2(32'h393dc928),
	.w3(32'h3a9d4fc2),
	.w4(32'hb9c86c02),
	.w5(32'h38d59725),
	.w6(32'hba97321a),
	.w7(32'hba8f7095),
	.w8(32'hbaaee611),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52a41d),
	.w1(32'h3a63ca6c),
	.w2(32'h3ac64fcb),
	.w3(32'h3aa3b48a),
	.w4(32'hb9f61836),
	.w5(32'h3acd7919),
	.w6(32'hbb4627c0),
	.w7(32'hbb715e5a),
	.w8(32'hbb809504),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388be242),
	.w1(32'h374e338a),
	.w2(32'hb89513ba),
	.w3(32'h38c5f1b0),
	.w4(32'h3686f742),
	.w5(32'hb8e2e795),
	.w6(32'hb6e4c0a6),
	.w7(32'hb809ac9e),
	.w8(32'hb8794d8f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81268a2),
	.w1(32'h37563818),
	.w2(32'h37cda96c),
	.w3(32'hb943b0ee),
	.w4(32'hb961d9c9),
	.w5(32'hb9256149),
	.w6(32'hb7afd085),
	.w7(32'hb754f0f9),
	.w8(32'h36af2e0a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba0df0),
	.w1(32'h3bcf0666),
	.w2(32'h3b1b889e),
	.w3(32'hba143ed4),
	.w4(32'h3b54364a),
	.w5(32'h3b0c78f4),
	.w6(32'hbb9f5860),
	.w7(32'hbb9afd3d),
	.w8(32'hbbba8c7e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba05eab),
	.w1(32'h3aefc34f),
	.w2(32'h397c9c54),
	.w3(32'h3b812579),
	.w4(32'h3b567dfc),
	.w5(32'h3b3ab042),
	.w6(32'hbb41d47b),
	.w7(32'hbb5d1553),
	.w8(32'hbb676654),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f630),
	.w1(32'h3affe904),
	.w2(32'h3a11c07e),
	.w3(32'hbb0b915a),
	.w4(32'hbb06ccae),
	.w5(32'hba28cb14),
	.w6(32'hbb4b2e1c),
	.w7(32'hbb966b2d),
	.w8(32'hbba95588),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71384c),
	.w1(32'hbac1fdf5),
	.w2(32'hbbc1c6e4),
	.w3(32'h3afd8caa),
	.w4(32'hba895a91),
	.w5(32'h3b0691c6),
	.w6(32'h3b0fa750),
	.w7(32'h38ceaa86),
	.w8(32'hb9fdd425),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9888dc3),
	.w1(32'hb7afc749),
	.w2(32'hb90f0dba),
	.w3(32'h3641ca16),
	.w4(32'h3a0cf74b),
	.w5(32'h3a0a41d9),
	.w6(32'h3a0272c2),
	.w7(32'h39baa720),
	.w8(32'h398165f4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a746676),
	.w1(32'h39df6711),
	.w2(32'hb99ac3d1),
	.w3(32'h3a305421),
	.w4(32'h3906d6b4),
	.w5(32'h3a2b45ff),
	.w6(32'hb9a36631),
	.w7(32'h367ad89c),
	.w8(32'hba0fb7d7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb7a50),
	.w1(32'h3bf7f6d0),
	.w2(32'hb8cc2132),
	.w3(32'h3a375b08),
	.w4(32'h3bcd1538),
	.w5(32'h3ad48258),
	.w6(32'hbb0b84c6),
	.w7(32'h3be34b73),
	.w8(32'h3ba8c86c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05ccd8),
	.w1(32'h3b89e7af),
	.w2(32'h3b3e64d1),
	.w3(32'h3bb35ed9),
	.w4(32'h3b5b5ac3),
	.w5(32'h3b38a0f2),
	.w6(32'hbb6fad1a),
	.w7(32'hbab9316c),
	.w8(32'hbb7d9fd3),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8a534),
	.w1(32'h3b33afd9),
	.w2(32'h3a234045),
	.w3(32'h3b604add),
	.w4(32'h3b9afd6e),
	.w5(32'h3afab5e4),
	.w6(32'hbb77a243),
	.w7(32'h3a31b37e),
	.w8(32'h3b3cecad),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae83e0a),
	.w1(32'hbad7e6ca),
	.w2(32'hba96be84),
	.w3(32'hbacdddc2),
	.w4(32'hbae519da),
	.w5(32'hbad31486),
	.w6(32'h39d2e4c2),
	.w7(32'hb97f9da7),
	.w8(32'hb9e5d559),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb152478),
	.w1(32'hbab0fdde),
	.w2(32'h3a469eba),
	.w3(32'hbb187b8b),
	.w4(32'hbb1e0d31),
	.w5(32'hbb01e30d),
	.w6(32'h3a5fd7b5),
	.w7(32'hbaa8630d),
	.w8(32'hbb151217),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb736fa04),
	.w1(32'hb68f3081),
	.w2(32'h3655f8d4),
	.w3(32'hb7059044),
	.w4(32'hb6128ac3),
	.w5(32'h367fef4b),
	.w6(32'h35254f4d),
	.w7(32'h35935a34),
	.w8(32'h37163cad),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7125db8),
	.w1(32'hb6e56390),
	.w2(32'h351d9998),
	.w3(32'hb644e717),
	.w4(32'h36b67be6),
	.w5(32'h375d1ec1),
	.w6(32'h37273b65),
	.w7(32'h37b1636c),
	.w8(32'h37fac023),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4cdd2),
	.w1(32'hba8e66de),
	.w2(32'hbacd55bb),
	.w3(32'h3ae20250),
	.w4(32'h3a02b7f0),
	.w5(32'h3a1c669a),
	.w6(32'hba5cb242),
	.w7(32'hba67583c),
	.w8(32'hbaadc6d2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7360c13),
	.w1(32'hb76ccdb4),
	.w2(32'hb65de3f9),
	.w3(32'hb648547a),
	.w4(32'hb6eae2dd),
	.w5(32'h36f4045c),
	.w6(32'h37cf195f),
	.w7(32'h37d08401),
	.w8(32'h381e5c38),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85b434),
	.w1(32'h3ab116d5),
	.w2(32'h3a2c0575),
	.w3(32'h3b1aa6ee),
	.w4(32'h3b6125c0),
	.w5(32'h3b53e1f5),
	.w6(32'hb96b770b),
	.w7(32'h3b0e4f3b),
	.w8(32'h3b1dec53),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82f09b),
	.w1(32'h3addf3f8),
	.w2(32'h39f1ba96),
	.w3(32'h3b16f202),
	.w4(32'h3ac5e104),
	.w5(32'h3ab66702),
	.w6(32'hbb31a6b5),
	.w7(32'hbb449834),
	.w8(32'hbb62fb37),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab010dc),
	.w1(32'h3a437d68),
	.w2(32'hb94f4220),
	.w3(32'h39740415),
	.w4(32'hb92568ed),
	.w5(32'hba75784b),
	.w6(32'hba61d14d),
	.w7(32'hbb01a00a),
	.w8(32'hbb1cbc9f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e6b003),
	.w1(32'hb5bd7efa),
	.w2(32'h373f7d69),
	.w3(32'hb7cad741),
	.w4(32'hb6debb00),
	.w5(32'h36f88617),
	.w6(32'h3605ce18),
	.w7(32'h362e13f3),
	.w8(32'h3756648b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29af14),
	.w1(32'h3bd01f80),
	.w2(32'h3b2e07f7),
	.w3(32'h3c140926),
	.w4(32'h3bf3c26c),
	.w5(32'h3babd048),
	.w6(32'hbb7da5c4),
	.w7(32'h3b1bea26),
	.w8(32'h3b695582),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeee749),
	.w1(32'h39b977e7),
	.w2(32'h3951d5ee),
	.w3(32'h3ae7b445),
	.w4(32'h3a5dff3f),
	.w5(32'h3a7e29ce),
	.w6(32'hbab237aa),
	.w7(32'hba0b0c43),
	.w8(32'hbaae41c8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3876c163),
	.w1(32'hb8300021),
	.w2(32'hb8ab45cf),
	.w3(32'h37c9db11),
	.w4(32'hb845e2f6),
	.w5(32'hb850a713),
	.w6(32'h38e934c4),
	.w7(32'h38c04a8a),
	.w8(32'h37ce8d8a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbfdb0),
	.w1(32'h3b34ce05),
	.w2(32'h3aa3e241),
	.w3(32'h3b8f9e0e),
	.w4(32'h3af8b7ec),
	.w5(32'h3ac44a33),
	.w6(32'hb8af3c32),
	.w7(32'hb98bbd04),
	.w8(32'hb9bb899d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da9bac),
	.w1(32'hb786371a),
	.w2(32'h367484ed),
	.w3(32'hb7b83d77),
	.w4(32'hb7c34cd5),
	.w5(32'h34572f36),
	.w6(32'h37d95930),
	.w7(32'h37270b94),
	.w8(32'h378ba2e9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70c1187),
	.w1(32'hb895b6d1),
	.w2(32'hb93b8d89),
	.w3(32'h39621376),
	.w4(32'h3982f3bc),
	.w5(32'h38c89564),
	.w6(32'h3862899e),
	.w7(32'h372adcf3),
	.w8(32'hb99a144b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b435d0),
	.w1(32'hb7675a70),
	.w2(32'h37a07035),
	.w3(32'hb86148ec),
	.w4(32'hb823f596),
	.w5(32'hb806712c),
	.w6(32'hb8417531),
	.w7(32'hb7c7b2ab),
	.w8(32'h367ff09f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fd007e),
	.w1(32'h37f4e86c),
	.w2(32'h37388832),
	.w3(32'hb7ad1636),
	.w4(32'hb6e1f27c),
	.w5(32'hb7200345),
	.w6(32'hb7ed5016),
	.w7(32'hb5ea10d5),
	.w8(32'h371c7cad),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1184b9),
	.w1(32'h37ba3ecf),
	.w2(32'h3a72f02a),
	.w3(32'hba1fadf7),
	.w4(32'h362bc58d),
	.w5(32'h38c77d73),
	.w6(32'h381ba6f0),
	.w7(32'h3825fe76),
	.w8(32'hb94b7ef8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb3b13),
	.w1(32'hbb366967),
	.w2(32'hb8a50eee),
	.w3(32'hba0347ec),
	.w4(32'hbb5a446e),
	.w5(32'hb9fcec78),
	.w6(32'hb9ee05c7),
	.w7(32'hbab7f625),
	.w8(32'hbac3e6a0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fb7d8),
	.w1(32'h3b32493b),
	.w2(32'h3aa134c1),
	.w3(32'h3b72af51),
	.w4(32'h3ae15a9a),
	.w5(32'h3a9ab388),
	.w6(32'hba77fe9d),
	.w7(32'hba346bb0),
	.w8(32'hbac2cde2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b524c98),
	.w1(32'hb98fee22),
	.w2(32'hb96c4cc6),
	.w3(32'h3b7a00e3),
	.w4(32'h3ac8e55b),
	.w5(32'h3acdf9d4),
	.w6(32'h3992bb3a),
	.w7(32'hb787ab0a),
	.w8(32'hbaa34d5c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36480a97),
	.w1(32'hb7716808),
	.w2(32'h375d5e6d),
	.w3(32'h37a6210c),
	.w4(32'h36708e32),
	.w5(32'hb7178667),
	.w6(32'h389c4e73),
	.w7(32'h379f4979),
	.w8(32'h37997181),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f62131),
	.w1(32'h3950ead1),
	.w2(32'h385f42f9),
	.w3(32'h396c0975),
	.w4(32'h3960f689),
	.w5(32'h3954785f),
	.w6(32'hb9de83e2),
	.w7(32'h390b8e7e),
	.w8(32'h392317f6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb702ca4e),
	.w1(32'hb6f7f547),
	.w2(32'h3491aacf),
	.w3(32'hb71e77c8),
	.w4(32'hb703fe41),
	.w5(32'h358f83b6),
	.w6(32'h36e8133e),
	.w7(32'h36b3f855),
	.w8(32'h376ac39c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c2a7ef),
	.w1(32'h3763a893),
	.w2(32'h36b2f9b9),
	.w3(32'h36222553),
	.w4(32'hb5bdc12e),
	.w5(32'h372153c8),
	.w6(32'h37c04d0f),
	.w7(32'h379c4860),
	.w8(32'h37b24f89),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f2e76),
	.w1(32'h3a9f2bcc),
	.w2(32'h3accef58),
	.w3(32'h3b8b2cc2),
	.w4(32'h3b0d9f75),
	.w5(32'h3b01b1f1),
	.w6(32'hba34d992),
	.w7(32'h37c40cb1),
	.w8(32'hbaa23b34),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b540a0),
	.w1(32'hb6e3fe73),
	.w2(32'hb6f3a426),
	.w3(32'hb4cd9c58),
	.w4(32'h3606b72b),
	.w5(32'h3736beca),
	.w6(32'h37b69116),
	.w7(32'h38046038),
	.w8(32'h38245ee6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c86429),
	.w1(32'h39a139c7),
	.w2(32'hb7660db1),
	.w3(32'h3820e941),
	.w4(32'h3977520b),
	.w5(32'hb915b54f),
	.w6(32'h38eac0de),
	.w7(32'h396f3a50),
	.w8(32'h38954e24),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4332b),
	.w1(32'h39b98cc5),
	.w2(32'h3a659ea1),
	.w3(32'h3a1629ca),
	.w4(32'h39afb26f),
	.w5(32'h397d01a7),
	.w6(32'h39b05a5b),
	.w7(32'h39d46f35),
	.w8(32'h3ab0a237),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70e780e),
	.w1(32'hb7919393),
	.w2(32'hb78981cb),
	.w3(32'h36ca7cb8),
	.w4(32'h363e6445),
	.w5(32'hb7484a86),
	.w6(32'h36ea07d7),
	.w7(32'h3707fa38),
	.w8(32'h3760dc4e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f0b0a),
	.w1(32'h3a83584b),
	.w2(32'h3a566e88),
	.w3(32'h3abdc3aa),
	.w4(32'h3a6394fe),
	.w5(32'h3a792066),
	.w6(32'hb89ad5b0),
	.w7(32'hb8a66053),
	.w8(32'hb9ea9ec0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9f24a),
	.w1(32'hb8f4c884),
	.w2(32'h3900af36),
	.w3(32'hb9c67100),
	.w4(32'h37131092),
	.w5(32'h391d734a),
	.w6(32'h3802cd5c),
	.w7(32'h39fee2ec),
	.w8(32'h39c90ee8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9943769),
	.w1(32'hba367b22),
	.w2(32'h3bb5c5c1),
	.w3(32'h3b3c0edf),
	.w4(32'h3addfcab),
	.w5(32'h3b79f6b3),
	.w6(32'h3ba08585),
	.w7(32'h398f46b1),
	.w8(32'h396485b0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fd2ec4),
	.w1(32'h390328de),
	.w2(32'h3906bcf7),
	.w3(32'h399519d4),
	.w4(32'h3984d6c5),
	.w5(32'h396e77d3),
	.w6(32'hb92b5927),
	.w7(32'hb7d38c18),
	.w8(32'h38bd40b3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38564b),
	.w1(32'h3baa0aa4),
	.w2(32'h3b880908),
	.w3(32'hbb29aff8),
	.w4(32'h392cd414),
	.w5(32'h3ad95975),
	.w6(32'hbb889baf),
	.w7(32'hbb82a879),
	.w8(32'hbb7c79e7),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule