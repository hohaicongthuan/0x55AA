module layer_10_featuremap_406(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94798e),
	.w1(32'h3a801f69),
	.w2(32'h3ab723af),
	.w3(32'h3baa1f11),
	.w4(32'hbbe41d2a),
	.w5(32'h3c7e08f5),
	.w6(32'h3a801bed),
	.w7(32'hbb3a8920),
	.w8(32'h3b75a224),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14ea0c),
	.w1(32'hbbd1b4df),
	.w2(32'hbbb1bc95),
	.w3(32'hbbfd258e),
	.w4(32'hbbceda40),
	.w5(32'h3b560b48),
	.w6(32'hba01930e),
	.w7(32'hbbf46e3a),
	.w8(32'h3ae0031b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a4fd6),
	.w1(32'hbaeee39b),
	.w2(32'hbadd2d9a),
	.w3(32'hbbcb1378),
	.w4(32'h39bc2db6),
	.w5(32'h39123c62),
	.w6(32'hbb9d022c),
	.w7(32'h3b17dc99),
	.w8(32'hbb3d93c5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fe246),
	.w1(32'hbb4ec9f0),
	.w2(32'hbbf99f44),
	.w3(32'hbb110f53),
	.w4(32'hbb4c5b0b),
	.w5(32'h3b621710),
	.w6(32'h3bc5c098),
	.w7(32'h3a4371c4),
	.w8(32'hbc2199c4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bd69c),
	.w1(32'h3b17a410),
	.w2(32'h3b3045c0),
	.w3(32'h3a183c4c),
	.w4(32'h3b03802b),
	.w5(32'hbb0ce5bd),
	.w6(32'hbacda33c),
	.w7(32'h3ba88d27),
	.w8(32'h3b287d77),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be27356),
	.w1(32'hbc0a3c57),
	.w2(32'h39d49bc5),
	.w3(32'h3c1bbcb2),
	.w4(32'h3b29758e),
	.w5(32'hbba72882),
	.w6(32'hba3a5441),
	.w7(32'hbbe1bd7f),
	.w8(32'h3a6041b9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c685),
	.w1(32'h3aa6f926),
	.w2(32'hbad3d9a5),
	.w3(32'hbbaa06f3),
	.w4(32'hb85322ed),
	.w5(32'hbbe9e054),
	.w6(32'hbb1690f0),
	.w7(32'h3b5156a2),
	.w8(32'h3b3c5f89),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bd365),
	.w1(32'h3b3e9e89),
	.w2(32'h3b58b244),
	.w3(32'hbb5ed9ef),
	.w4(32'h3b0f8c14),
	.w5(32'hbb2bb0d8),
	.w6(32'h3b6e0802),
	.w7(32'hbb40859d),
	.w8(32'hbab7003a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b124560),
	.w1(32'hbbb09375),
	.w2(32'h3a9c3b12),
	.w3(32'hbba8bc2a),
	.w4(32'h3b43379a),
	.w5(32'h3b9585c5),
	.w6(32'h3b0d13f0),
	.w7(32'h3b203768),
	.w8(32'h3b4d37b7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3545a),
	.w1(32'hbb5783d9),
	.w2(32'h3b781c39),
	.w3(32'hbb2919ee),
	.w4(32'h3b9ebd65),
	.w5(32'h3bc6837a),
	.w6(32'hbb156a11),
	.w7(32'hba3889ae),
	.w8(32'h39a29f66),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86d6ea),
	.w1(32'hbc1f7422),
	.w2(32'hba1ec591),
	.w3(32'hbbb960e6),
	.w4(32'hbb959f41),
	.w5(32'hbb24566f),
	.w6(32'h3902e492),
	.w7(32'hbbab147c),
	.w8(32'h3980a72d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51c728),
	.w1(32'h3bbba545),
	.w2(32'h3c770ed4),
	.w3(32'hbbb8a6ca),
	.w4(32'h3b266341),
	.w5(32'hbc8c06d7),
	.w6(32'hba0e6f07),
	.w7(32'h3bb42a3d),
	.w8(32'hbb64b7cc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c354d83),
	.w1(32'h3896680a),
	.w2(32'h3c1d93da),
	.w3(32'h3bbbb4d0),
	.w4(32'hbaa69e02),
	.w5(32'hbc3b4290),
	.w6(32'h3a352e95),
	.w7(32'hba51236a),
	.w8(32'hbb206455),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03edbd),
	.w1(32'h3ad6ecb2),
	.w2(32'hba81e123),
	.w3(32'hbae6d2d3),
	.w4(32'h3b2b2bad),
	.w5(32'h3bd1c0b9),
	.w6(32'hbadcda68),
	.w7(32'hbae54d1e),
	.w8(32'hbb44d3d0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90946c),
	.w1(32'h3afcbe8d),
	.w2(32'h3b19be71),
	.w3(32'h39aa6aae),
	.w4(32'h3852e9d7),
	.w5(32'hbb8ad40a),
	.w6(32'h3af031a1),
	.w7(32'hbaf6376b),
	.w8(32'hba01a8dc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c808e),
	.w1(32'h3b898288),
	.w2(32'h3c49e607),
	.w3(32'hbbcd3269),
	.w4(32'h3c167453),
	.w5(32'hbbf9fb8c),
	.w6(32'hbb803b9e),
	.w7(32'h3bd70c39),
	.w8(32'hbb21078b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1508a),
	.w1(32'hbb5b6d50),
	.w2(32'hba7a202e),
	.w3(32'h3c5ac49e),
	.w4(32'hbb37c936),
	.w5(32'hbbb9a4a4),
	.w6(32'h3b7805dc),
	.w7(32'h3c4e0859),
	.w8(32'h3bd329f4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdfc15),
	.w1(32'hbc624e5a),
	.w2(32'hbb5bb8bb),
	.w3(32'hbaecd569),
	.w4(32'hbb2050c9),
	.w5(32'h3cbfca5d),
	.w6(32'hb9e93b1f),
	.w7(32'hbbd99dcf),
	.w8(32'h3c7ea204),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa12d08),
	.w1(32'hbb2d579a),
	.w2(32'h3b6f3365),
	.w3(32'h3a1e0099),
	.w4(32'h3b11226f),
	.w5(32'hbc1e831f),
	.w6(32'h3b08f09c),
	.w7(32'hb8c67af1),
	.w8(32'hbb921973),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804257),
	.w1(32'hbae419c0),
	.w2(32'hbb824ca8),
	.w3(32'hbc064a9b),
	.w4(32'h3b60c08d),
	.w5(32'hbbba6959),
	.w6(32'hbb956b00),
	.w7(32'hbab9b491),
	.w8(32'h3a6feb3f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcac6e5),
	.w1(32'h3af22755),
	.w2(32'h3c0c4d88),
	.w3(32'hbb9c1644),
	.w4(32'hbaa050dd),
	.w5(32'hbb96f1e9),
	.w6(32'hbc04a53d),
	.w7(32'hba283f5e),
	.w8(32'hb98dab7c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b239bd0),
	.w1(32'hbaf41b17),
	.w2(32'h39bd5eb6),
	.w3(32'hbb809a7c),
	.w4(32'hbb978b23),
	.w5(32'hbb646462),
	.w6(32'h3b800d43),
	.w7(32'hbaf2eaec),
	.w8(32'h39d467ae),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9bff5),
	.w1(32'hbb4f931a),
	.w2(32'h3b92a257),
	.w3(32'hbb877e95),
	.w4(32'hbb4367c3),
	.w5(32'hbc13b411),
	.w6(32'hbbdc1a28),
	.w7(32'h3a0920e5),
	.w8(32'hbabf2359),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0b6ac),
	.w1(32'hbbdfaf52),
	.w2(32'h3bf44d87),
	.w3(32'hbc84286e),
	.w4(32'h3b52205c),
	.w5(32'h3c481ac7),
	.w6(32'h3b0f4571),
	.w7(32'h3b1a5313),
	.w8(32'h3c528f81),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb789c03),
	.w1(32'hbc560531),
	.w2(32'hbc528fc5),
	.w3(32'h3bc7befb),
	.w4(32'hbc2c41c6),
	.w5(32'hbb8cff3f),
	.w6(32'h3b816fad),
	.w7(32'hbc69344a),
	.w8(32'hbc588dec),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf05cab),
	.w1(32'hba349518),
	.w2(32'hbb16095e),
	.w3(32'hba7b954c),
	.w4(32'hbb038cdf),
	.w5(32'hbac37126),
	.w6(32'h3b196f18),
	.w7(32'hbb428c3a),
	.w8(32'hbb28bfa6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e6087),
	.w1(32'h3833ef70),
	.w2(32'hba8b60c2),
	.w3(32'hbc02a92f),
	.w4(32'h3b8aafe4),
	.w5(32'h3b95153f),
	.w6(32'hbba9332e),
	.w7(32'h3badb94e),
	.w8(32'h3c13a93c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164680),
	.w1(32'hbb8ffe96),
	.w2(32'hbb9b637d),
	.w3(32'h3b456a7b),
	.w4(32'hbb3bcd93),
	.w5(32'h3bc0d223),
	.w6(32'h3ca7ee98),
	.w7(32'hbad6f56b),
	.w8(32'hbbad7949),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc272bc4),
	.w1(32'h3aa709f7),
	.w2(32'hbbb078aa),
	.w3(32'hbc043c9f),
	.w4(32'hbba87742),
	.w5(32'hbbbbdf23),
	.w6(32'hbb3eb64d),
	.w7(32'h3b324b7c),
	.w8(32'h3c440545),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d2edd),
	.w1(32'h3ae627db),
	.w2(32'h3c804e79),
	.w3(32'h3af95c0c),
	.w4(32'hbc29b4b7),
	.w5(32'hbc128745),
	.w6(32'h3b908d4b),
	.w7(32'hbafb059e),
	.w8(32'h3b720d03),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1189e8),
	.w1(32'hb8bc2b76),
	.w2(32'h3b1e99c9),
	.w3(32'h3a29d870),
	.w4(32'h3b8683b4),
	.w5(32'hbb73be9f),
	.w6(32'h3ae14ac3),
	.w7(32'hbbf02826),
	.w8(32'hbb278887),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae333e6),
	.w1(32'h3a131d75),
	.w2(32'h3ae32260),
	.w3(32'hbbbb361a),
	.w4(32'hbbed6b68),
	.w5(32'h3b99c0fd),
	.w6(32'hbbf6e58a),
	.w7(32'hbb71f5ce),
	.w8(32'h3b2f0b26),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02e673),
	.w1(32'hbacea70d),
	.w2(32'hbb66e47f),
	.w3(32'h3b64669a),
	.w4(32'hbb507a43),
	.w5(32'hbb4cf607),
	.w6(32'h3b924b11),
	.w7(32'h3ad592d1),
	.w8(32'hbbc86751),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcd2f1),
	.w1(32'hbbe5cd38),
	.w2(32'hbbc18448),
	.w3(32'hbb571cc8),
	.w4(32'hbb198b5c),
	.w5(32'h3b87aeeb),
	.w6(32'hbabdb3bf),
	.w7(32'h3ae6a596),
	.w8(32'h3bab19b8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc201af6),
	.w1(32'h3aba28c6),
	.w2(32'h3b4ee448),
	.w3(32'hbbcb6a94),
	.w4(32'h3b843c23),
	.w5(32'h39bbba10),
	.w6(32'h3adf08e2),
	.w7(32'hbb3ea34d),
	.w8(32'hbb9fb83b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba686d9),
	.w1(32'hbb9f847a),
	.w2(32'hbaaa7f7a),
	.w3(32'hba0749e0),
	.w4(32'hbaccd01d),
	.w5(32'h3b1cd838),
	.w6(32'hbb1f7881),
	.w7(32'h3b1b5ec4),
	.w8(32'hbb06058e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb701eb0),
	.w1(32'hbc0a1ef6),
	.w2(32'hbc0cba26),
	.w3(32'h3ba67a82),
	.w4(32'hbc0c12c1),
	.w5(32'hbb8d278e),
	.w6(32'hbb3291cd),
	.w7(32'hbc06205d),
	.w8(32'hbb234f8e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ca7e2),
	.w1(32'h3bc49e2b),
	.w2(32'h3bbb89f8),
	.w3(32'hbbbb8421),
	.w4(32'h3af90922),
	.w5(32'hba11549d),
	.w6(32'h3bba761b),
	.w7(32'hbbca1e37),
	.w8(32'h3b8a86e0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394786f3),
	.w1(32'hbba2b039),
	.w2(32'hbc444c85),
	.w3(32'hbb8f45d5),
	.w4(32'hbc320c23),
	.w5(32'h3b945fa2),
	.w6(32'hbae8525d),
	.w7(32'hbc11567e),
	.w8(32'hbbd62332),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8e33d),
	.w1(32'h3b7dbcd9),
	.w2(32'hbb3086d1),
	.w3(32'hbc104c13),
	.w4(32'h3aadd0dd),
	.w5(32'h3c912f2f),
	.w6(32'hbc29df37),
	.w7(32'hbb102b4a),
	.w8(32'h3b0efcb4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb1b7),
	.w1(32'h3b63c99e),
	.w2(32'h393f35b3),
	.w3(32'hbbe570e2),
	.w4(32'hbc442a82),
	.w5(32'hbb181d9a),
	.w6(32'hba5b45c0),
	.w7(32'h3b9ececc),
	.w8(32'h3b94293a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e4fd),
	.w1(32'hbc1dff36),
	.w2(32'hbb0bd64d),
	.w3(32'hbb4dfec9),
	.w4(32'hbc24ec25),
	.w5(32'hbba0d6e1),
	.w6(32'hbb82b47b),
	.w7(32'hbc001a13),
	.w8(32'hbb209937),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34ad4c),
	.w1(32'hbb47ccff),
	.w2(32'h3adfc81f),
	.w3(32'hbb86735e),
	.w4(32'hbbdb3cbf),
	.w5(32'hbb30d4dd),
	.w6(32'hbb02b67e),
	.w7(32'hba32388d),
	.w8(32'hbb80120a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5af4e),
	.w1(32'hbb9e6d1e),
	.w2(32'hbc37b023),
	.w3(32'h3ae1e3b6),
	.w4(32'hbc250887),
	.w5(32'h3c29bad3),
	.w6(32'h3b15f8c7),
	.w7(32'hbb8b9778),
	.w8(32'hbb819c7b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b57dd),
	.w1(32'hba92665e),
	.w2(32'h3bc642be),
	.w3(32'hbc41420f),
	.w4(32'hbb3eadc8),
	.w5(32'hba12e3f1),
	.w6(32'hbc1b7b1a),
	.w7(32'h3adccbda),
	.w8(32'h3b3a4f60),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad06259),
	.w1(32'hbb3d4213),
	.w2(32'h3b5476e1),
	.w3(32'h3b0d6f30),
	.w4(32'h3a5a65c8),
	.w5(32'hbb9079c4),
	.w6(32'hb968a258),
	.w7(32'h3b991c58),
	.w8(32'hba8aa17d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9899792),
	.w1(32'h3b092955),
	.w2(32'h3bb69aa5),
	.w3(32'hbb94d122),
	.w4(32'h3bdc1122),
	.w5(32'h3a1cd5eb),
	.w6(32'hbaa3558e),
	.w7(32'hbb857fb6),
	.w8(32'hba6bfa7a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903eeb8),
	.w1(32'h3a959b54),
	.w2(32'hbb37a7a1),
	.w3(32'hbbdcc033),
	.w4(32'h3b3f0f01),
	.w5(32'hbb6d3be1),
	.w6(32'hbb88950c),
	.w7(32'h3a82e269),
	.w8(32'hb9e7c85c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6cec4),
	.w1(32'hbbbb136b),
	.w2(32'hbbe768e8),
	.w3(32'hba9bbcad),
	.w4(32'hbb540b23),
	.w5(32'h3aa5d57e),
	.w6(32'hbb2a9430),
	.w7(32'hbb5acdbb),
	.w8(32'hba07d605),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30ccaa),
	.w1(32'hbb906c04),
	.w2(32'hbb9c27b4),
	.w3(32'hbc127de4),
	.w4(32'hbafc828d),
	.w5(32'h3a2fa4d5),
	.w6(32'hbc46c5d5),
	.w7(32'hbb581a66),
	.w8(32'h39896b52),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc003b0e),
	.w1(32'h3b5a520d),
	.w2(32'h3c3049a2),
	.w3(32'hbb0aa6d6),
	.w4(32'h3c055c54),
	.w5(32'h3add71d0),
	.w6(32'hbbafcda7),
	.w7(32'h3bd853bf),
	.w8(32'h3a963a00),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc54db0),
	.w1(32'h3b8d5a37),
	.w2(32'h3b3f03e7),
	.w3(32'h3bd87eeb),
	.w4(32'h3a43ca14),
	.w5(32'hba1db091),
	.w6(32'h3c085cc2),
	.w7(32'h3b230a36),
	.w8(32'hbb4520e4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb435aee),
	.w1(32'hbbfb5835),
	.w2(32'h3a5e3d84),
	.w3(32'h3ba6d3ff),
	.w4(32'hbab1d2fa),
	.w5(32'h3b61f038),
	.w6(32'hba4a7217),
	.w7(32'hbc1f2da7),
	.w8(32'hbab9fc21),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7de2b8),
	.w1(32'hbb0f572f),
	.w2(32'hbab44f65),
	.w3(32'hbb308b1e),
	.w4(32'h3b52463d),
	.w5(32'h3a6fdbba),
	.w6(32'h3a1f0aed),
	.w7(32'hbbbbdc75),
	.w8(32'hbb80883a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bc96b),
	.w1(32'h3bbcefcb),
	.w2(32'h3b36798b),
	.w3(32'hbb01236d),
	.w4(32'h39c1ab40),
	.w5(32'h3b43d838),
	.w6(32'h3b247968),
	.w7(32'h3b1b3f60),
	.w8(32'hbb1df38e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b316a0d),
	.w1(32'h3af4da04),
	.w2(32'h397f4f1d),
	.w3(32'hb9ec093f),
	.w4(32'hba9d721f),
	.w5(32'h3c1ad082),
	.w6(32'hb9b870c5),
	.w7(32'hbb9e9986),
	.w8(32'h3bb57154),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef04d4),
	.w1(32'h3c0a65a3),
	.w2(32'h3c3b7200),
	.w3(32'hba85265e),
	.w4(32'h3c7f7c55),
	.w5(32'hbcf25f1b),
	.w6(32'h3b555e96),
	.w7(32'h3b9d4662),
	.w8(32'hbb84ea32),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5786b2),
	.w1(32'hbbdaddae),
	.w2(32'hbc3aa40f),
	.w3(32'h3c6b1049),
	.w4(32'hb8c94409),
	.w5(32'hbbeec2e9),
	.w6(32'h3c3850b7),
	.w7(32'h3a1d44bb),
	.w8(32'hb9a9b044),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b246ffc),
	.w1(32'hb99fd210),
	.w2(32'hbc010e59),
	.w3(32'h39cf4855),
	.w4(32'hbc00e8d5),
	.w5(32'hbc3812b8),
	.w6(32'hbb450aad),
	.w7(32'hbb55571e),
	.w8(32'hbc2d16b1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb756b0f),
	.w1(32'hbc6a0999),
	.w2(32'hbc5569c9),
	.w3(32'hbad80615),
	.w4(32'hbc0ae2d9),
	.w5(32'hbc2c5412),
	.w6(32'hbbc53859),
	.w7(32'hbbd0cdd9),
	.w8(32'hbb656779),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e1fbd),
	.w1(32'h3be3b631),
	.w2(32'h3aac74f9),
	.w3(32'hbc50426e),
	.w4(32'h3b9ce1a6),
	.w5(32'hbb80bb19),
	.w6(32'hbbfd385d),
	.w7(32'h3b8659a6),
	.w8(32'h3abc9ac6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb270781),
	.w1(32'h3b82eafa),
	.w2(32'h3b6e3fac),
	.w3(32'hbb408be2),
	.w4(32'hbb4d9d10),
	.w5(32'h3c4c1d81),
	.w6(32'h3c22d898),
	.w7(32'h3aefa6fe),
	.w8(32'h3bf6b40d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398d96),
	.w1(32'hbc0cb3c8),
	.w2(32'hbba8c53b),
	.w3(32'hbb5f018f),
	.w4(32'hbb8b7e22),
	.w5(32'h3c5ce27d),
	.w6(32'h3b08c50a),
	.w7(32'hbae27c7c),
	.w8(32'hbb9c16bf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fdc0d),
	.w1(32'h3c0d0af7),
	.w2(32'h3bd37e5b),
	.w3(32'hba551376),
	.w4(32'h3c3847c4),
	.w5(32'hbce50e87),
	.w6(32'h3aae6244),
	.w7(32'hbb4d4e78),
	.w8(32'hbad1fed5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba0cf1),
	.w1(32'h3c075e67),
	.w2(32'h3c110f0b),
	.w3(32'h3abf6d4d),
	.w4(32'h3b661d7b),
	.w5(32'h3a741d7c),
	.w6(32'h3b89808a),
	.w7(32'h3addec78),
	.w8(32'hba269c06),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61dc49),
	.w1(32'hbbe64053),
	.w2(32'hbba0d806),
	.w3(32'hbad8d413),
	.w4(32'hbb9b2c4a),
	.w5(32'h3c125499),
	.w6(32'hbb691749),
	.w7(32'h3aefa51e),
	.w8(32'h3bd4fff0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9d0dd),
	.w1(32'hbb9c893d),
	.w2(32'hba900977),
	.w3(32'h3b84088c),
	.w4(32'h3b04b59d),
	.w5(32'h3b1aab33),
	.w6(32'h3b4e53ca),
	.w7(32'h3b34a7c0),
	.w8(32'hba111897),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10cb28),
	.w1(32'h3bc1cc68),
	.w2(32'h3c024618),
	.w3(32'hbbb2f1fd),
	.w4(32'h3c1c2221),
	.w5(32'h3c42b51e),
	.w6(32'h3abd2259),
	.w7(32'h3c2fdca3),
	.w8(32'h3c5e6fd9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8efef),
	.w1(32'hbae2a27c),
	.w2(32'hbc0bef49),
	.w3(32'hbc0987a1),
	.w4(32'hbc4997b7),
	.w5(32'hbaa6a0d8),
	.w6(32'h3c3b2562),
	.w7(32'hbbe2c3d6),
	.w8(32'hbbc2d02d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293a77),
	.w1(32'hbb97ce6f),
	.w2(32'hbc350095),
	.w3(32'h3b9a7ffd),
	.w4(32'h3b3e9417),
	.w5(32'hbc13b46e),
	.w6(32'hbb6564ce),
	.w7(32'hbaebc6a3),
	.w8(32'hbba9bb1f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf65ab6),
	.w1(32'hbbe41927),
	.w2(32'hbb3e4480),
	.w3(32'hbae872cf),
	.w4(32'hbb4371e0),
	.w5(32'h3b105daa),
	.w6(32'hb9695ad5),
	.w7(32'h3b769885),
	.w8(32'h3b1b1ea4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23dedf),
	.w1(32'h3b25a983),
	.w2(32'hbb387bef),
	.w3(32'hbb4ba731),
	.w4(32'hbba85c73),
	.w5(32'hbc3363ec),
	.w6(32'hbb4c034f),
	.w7(32'hbb414f08),
	.w8(32'hbbde7cb3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3a24b),
	.w1(32'hbba1b1d0),
	.w2(32'hb9f1c716),
	.w3(32'h3ab7f798),
	.w4(32'hbc3b0f40),
	.w5(32'h3c80aa6e),
	.w6(32'h3c147821),
	.w7(32'hbbf12d2e),
	.w8(32'h38b5ccc3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dc376),
	.w1(32'hbb5e95b4),
	.w2(32'h3baaaea1),
	.w3(32'h3b20a6f1),
	.w4(32'hbb4f4862),
	.w5(32'h3b760ab8),
	.w6(32'h3b98abc3),
	.w7(32'hbb6a56fa),
	.w8(32'hb9202e88),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a4ea5),
	.w1(32'hbc2017ca),
	.w2(32'h3b021ad4),
	.w3(32'hbb730329),
	.w4(32'hbbcaeecb),
	.w5(32'h3a2a4f41),
	.w6(32'hbb852292),
	.w7(32'hbc5f9e82),
	.w8(32'h3b601e49),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a69a3),
	.w1(32'hb9a32188),
	.w2(32'hbbb18a3b),
	.w3(32'h3b984578),
	.w4(32'h3ba17717),
	.w5(32'hbc564e37),
	.w6(32'h3b0d7a9d),
	.w7(32'hbb9ae4e8),
	.w8(32'h3a427e00),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7f2be),
	.w1(32'hbba9ac1e),
	.w2(32'h3b50c81c),
	.w3(32'h39fa72d4),
	.w4(32'hbbb13fd7),
	.w5(32'h3cb75e2a),
	.w6(32'h3b75bf09),
	.w7(32'hb998bc5f),
	.w8(32'h3c1052f0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc480091),
	.w1(32'hba1fb73b),
	.w2(32'hbbba1326),
	.w3(32'hbc06d552),
	.w4(32'hbb9d0516),
	.w5(32'h3bc34577),
	.w6(32'hbc649126),
	.w7(32'hbb99425c),
	.w8(32'hbbaff4cf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a2aca),
	.w1(32'hbadf9274),
	.w2(32'h382ddbd8),
	.w3(32'hba3cfa59),
	.w4(32'hbc1b269d),
	.w5(32'h3c26b6fc),
	.w6(32'hbab6fd1e),
	.w7(32'hbb356b25),
	.w8(32'hbaf6cce0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab67a1),
	.w1(32'hbaf17348),
	.w2(32'h39c70829),
	.w3(32'hbc2f110a),
	.w4(32'h3bd2f5f8),
	.w5(32'hbbaf31d4),
	.w6(32'hbb7f047c),
	.w7(32'h3c062b8e),
	.w8(32'h3aaab33e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f662),
	.w1(32'h3b5e7dd1),
	.w2(32'h3b8f93ee),
	.w3(32'h39ac88b6),
	.w4(32'hbbe3ebbe),
	.w5(32'h3acb03fe),
	.w6(32'hbb8d1f33),
	.w7(32'h3aa5bcce),
	.w8(32'h3ba8d55e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77daf5),
	.w1(32'h38f235d5),
	.w2(32'h3ba42c92),
	.w3(32'hbb32eb36),
	.w4(32'hbbf08d45),
	.w5(32'h3ca59e6d),
	.w6(32'h3b52436a),
	.w7(32'hba78dcc5),
	.w8(32'h3bbd586b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc18a84),
	.w1(32'hbb310ce8),
	.w2(32'hb8d88fa3),
	.w3(32'hbc209fec),
	.w4(32'hbbc82d96),
	.w5(32'hb925fb2f),
	.w6(32'hbb012f1a),
	.w7(32'h39bf004a),
	.w8(32'hbb872fda),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f83595),
	.w1(32'hbb8f02ff),
	.w2(32'h3a21772f),
	.w3(32'h3b21fe6b),
	.w4(32'hbcb5730f),
	.w5(32'h3d863d7f),
	.w6(32'h3b0f2943),
	.w7(32'hba116121),
	.w8(32'h3c7c1a5c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7213c4),
	.w1(32'h3b406203),
	.w2(32'h39f24773),
	.w3(32'hb8828035),
	.w4(32'hbc8c3bed),
	.w5(32'h3cc77ed3),
	.w6(32'h3bca120c),
	.w7(32'hbc1a8625),
	.w8(32'h3bcbb720),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5483df),
	.w1(32'hbb73962c),
	.w2(32'h3a179bed),
	.w3(32'hbba93dc3),
	.w4(32'h3b9b0245),
	.w5(32'hbc1263fd),
	.w6(32'h3b32b6fa),
	.w7(32'h3bdedd1a),
	.w8(32'hbc1f67e3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac42000),
	.w1(32'h3bb40c76),
	.w2(32'hbb6538ab),
	.w3(32'h3c458c43),
	.w4(32'h3b9a20f7),
	.w5(32'hbc72a64d),
	.w6(32'h3b37722d),
	.w7(32'h3c23990f),
	.w8(32'h3a813b2e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad64518),
	.w1(32'hba4cbb66),
	.w2(32'h3aa08f4a),
	.w3(32'h3b548cc3),
	.w4(32'hbbe9ba78),
	.w5(32'hbbe25054),
	.w6(32'hbb778375),
	.w7(32'h3bb77a60),
	.w8(32'h3be61dba),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c131744),
	.w1(32'h3b4daa9b),
	.w2(32'h3c2cdd8f),
	.w3(32'h3c0276a4),
	.w4(32'hbc25c29c),
	.w5(32'h3d2adc94),
	.w6(32'h3c474b07),
	.w7(32'h3c212742),
	.w8(32'h3c883a5f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad06a0c),
	.w1(32'h3bbd6cf0),
	.w2(32'hbab1b461),
	.w3(32'hbbf680e3),
	.w4(32'h3c49608d),
	.w5(32'hbc919422),
	.w6(32'hbb82a5dc),
	.w7(32'h3bc9d362),
	.w8(32'hbbfa1d71),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b833248),
	.w1(32'hbc2d639b),
	.w2(32'hbbe2220c),
	.w3(32'hb8b77bed),
	.w4(32'hbc8e9e8e),
	.w5(32'h3be81626),
	.w6(32'hbab00884),
	.w7(32'hbc05717b),
	.w8(32'hba59a5e8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc017ae3),
	.w1(32'hba6a8be2),
	.w2(32'h3c6dbcc5),
	.w3(32'hbc77f36b),
	.w4(32'h3c398ee4),
	.w5(32'hbc209e7c),
	.w6(32'hbb29ee7d),
	.w7(32'h3c2051c3),
	.w8(32'hbb4f03f6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2986fe),
	.w1(32'hbbdbccfa),
	.w2(32'hba0361ad),
	.w3(32'h3be86c1f),
	.w4(32'hbbcaaf29),
	.w5(32'hbb920dc0),
	.w6(32'h3bb875cd),
	.w7(32'hbb96ceff),
	.w8(32'h39da0ac6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d6e65),
	.w1(32'hba9a010b),
	.w2(32'h3c164587),
	.w3(32'h3a78afc3),
	.w4(32'h39cabe6c),
	.w5(32'hbb431cad),
	.w6(32'h3a57777b),
	.w7(32'h3af3f209),
	.w8(32'h3b7799d7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b592898),
	.w1(32'hbb8b47d4),
	.w2(32'h3bca9817),
	.w3(32'h3a344399),
	.w4(32'h3aa002d8),
	.w5(32'h3b43b1d3),
	.w6(32'h3b9c49be),
	.w7(32'h3c64bcc0),
	.w8(32'hbc5ab0b1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fc88b),
	.w1(32'h3ab973ea),
	.w2(32'h3b293bb0),
	.w3(32'h3bfcf961),
	.w4(32'h3bd3a9c8),
	.w5(32'h3bf870fb),
	.w6(32'h3bb8c856),
	.w7(32'h3bb6963c),
	.w8(32'hbb4caf05),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d9a6b),
	.w1(32'h3aeedb35),
	.w2(32'h3bd558ca),
	.w3(32'h3c01cf9d),
	.w4(32'hbb9e65c2),
	.w5(32'h3cb55092),
	.w6(32'hbb59614e),
	.w7(32'h3b766168),
	.w8(32'h3b400bf2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa672ed),
	.w1(32'h3bd9d77b),
	.w2(32'hbb62cfe3),
	.w3(32'hba99c85c),
	.w4(32'h3a8ea6b0),
	.w5(32'hbb66fde2),
	.w6(32'h3ba893ec),
	.w7(32'h3b2210d6),
	.w8(32'h3a89cd9c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfcd2f),
	.w1(32'hbc3a8983),
	.w2(32'hbbed52bf),
	.w3(32'h3b69cacb),
	.w4(32'hbc052ab6),
	.w5(32'hbad20cef),
	.w6(32'hb85e82c0),
	.w7(32'hbb2e8c58),
	.w8(32'hbbcd5371),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06b1a3),
	.w1(32'h3c429299),
	.w2(32'hbbcdd9e3),
	.w3(32'hbc484e27),
	.w4(32'h3c4e3a80),
	.w5(32'hbc044a95),
	.w6(32'hbc107cf0),
	.w7(32'hba25eec5),
	.w8(32'h3c663b87),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35c5d1),
	.w1(32'hbb0dca24),
	.w2(32'h3c196722),
	.w3(32'h3c49e05b),
	.w4(32'hba00bdaf),
	.w5(32'h3c066cc3),
	.w6(32'h3c100495),
	.w7(32'h3ba4075e),
	.w8(32'hbc06fe0e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90fa1a),
	.w1(32'h3bbece13),
	.w2(32'hbbf1d537),
	.w3(32'hbb0ec0f1),
	.w4(32'h3bc04420),
	.w5(32'hb887002a),
	.w6(32'hbb9c9bd3),
	.w7(32'h3aaab89a),
	.w8(32'h3af2dfad),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f8b23),
	.w1(32'hbc16328f),
	.w2(32'h3bbf2751),
	.w3(32'h3b6fc048),
	.w4(32'hbbe0084d),
	.w5(32'hb9e9b8d6),
	.w6(32'hbad1309b),
	.w7(32'h3b8fd211),
	.w8(32'hbb9c6ce2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac56686),
	.w1(32'h3baeb15b),
	.w2(32'hbbf91028),
	.w3(32'hbabb1987),
	.w4(32'h3a14ee4f),
	.w5(32'h3c6553c6),
	.w6(32'h39e1f172),
	.w7(32'h3bbbbcaa),
	.w8(32'hbb7ebf41),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae40bfe),
	.w1(32'h3b431f4b),
	.w2(32'h3c38f188),
	.w3(32'hbb07290f),
	.w4(32'hba7bab36),
	.w5(32'h3c191ac0),
	.w6(32'hbafd9560),
	.w7(32'h3c1840ea),
	.w8(32'h3c2e22a4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2cb96),
	.w1(32'h3bbfdeee),
	.w2(32'h3bc7003d),
	.w3(32'h3b056234),
	.w4(32'hbb8d70e3),
	.w5(32'h3b317891),
	.w6(32'h397f1ee0),
	.w7(32'h39cc3c0b),
	.w8(32'h3a2b7bf6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb00c2),
	.w1(32'h39eeb4fe),
	.w2(32'h3bc4f61c),
	.w3(32'hbb9f02d0),
	.w4(32'h3c46ca92),
	.w5(32'h3c29c936),
	.w6(32'hbb157d05),
	.w7(32'h3bbd8c2c),
	.w8(32'h3bc7f8e9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba887800),
	.w1(32'hbc3f6579),
	.w2(32'hbbc43611),
	.w3(32'hbbcc7521),
	.w4(32'hbc49b1cf),
	.w5(32'hbc0a1262),
	.w6(32'hbb03319c),
	.w7(32'hbc478611),
	.w8(32'hbc44a020),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba9ce4),
	.w1(32'h3b109b0b),
	.w2(32'hbab0d351),
	.w3(32'h3a96d0b5),
	.w4(32'hbaaaed42),
	.w5(32'hbbdfae76),
	.w6(32'hbb4e65f9),
	.w7(32'hbbb2c78b),
	.w8(32'hbc02dfa5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af52c67),
	.w1(32'hbb3e0c11),
	.w2(32'h3bb9a76d),
	.w3(32'h3a4f30b3),
	.w4(32'h3ad8ca89),
	.w5(32'hbaf61fb7),
	.w6(32'h3b232817),
	.w7(32'hbbd2169e),
	.w8(32'h3b389eca),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba93201),
	.w1(32'hbbdc7f33),
	.w2(32'hbb8574f3),
	.w3(32'h3aab6607),
	.w4(32'h3b66b147),
	.w5(32'hbbbddfea),
	.w6(32'hbbb251df),
	.w7(32'h3ac2f340),
	.w8(32'hba433ce7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb9763),
	.w1(32'h3c063604),
	.w2(32'hbb0dfdd5),
	.w3(32'h3ba651ea),
	.w4(32'h3c5f52e5),
	.w5(32'hbc576816),
	.w6(32'h3b950fdd),
	.w7(32'h3c328cb8),
	.w8(32'hbc1bd19e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b798b66),
	.w1(32'hbb62ae74),
	.w2(32'h3b2e67af),
	.w3(32'h3bc5d1fc),
	.w4(32'hbb671d18),
	.w5(32'h3a0acace),
	.w6(32'h3b9fa49c),
	.w7(32'h3b37a9d9),
	.w8(32'h39c61808),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabae7b3),
	.w1(32'hbb89b57e),
	.w2(32'h3b0af64c),
	.w3(32'hb9d2a3e9),
	.w4(32'hbc97afa0),
	.w5(32'h3cd0b304),
	.w6(32'hba4aa8b7),
	.w7(32'hbb805591),
	.w8(32'h3a819d8b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9edffb),
	.w1(32'hbc372923),
	.w2(32'hbb0ac64b),
	.w3(32'hbbc803a2),
	.w4(32'hbc80d9db),
	.w5(32'hbc15aa30),
	.w6(32'hbb34afd7),
	.w7(32'hbc5e5314),
	.w8(32'hbbdbf8b2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0cf6c),
	.w1(32'hbac3d60c),
	.w2(32'hbc8803c3),
	.w3(32'hb9fbdb2e),
	.w4(32'hbc244068),
	.w5(32'hbce67355),
	.w6(32'h3938e366),
	.w7(32'hbc333a3d),
	.w8(32'hbc8426ae),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf96959),
	.w1(32'h3c1137ef),
	.w2(32'hbb2282ef),
	.w3(32'h39f70494),
	.w4(32'h3b9b3376),
	.w5(32'h3a694051),
	.w6(32'hbad20dc0),
	.w7(32'h3b2a8282),
	.w8(32'hbaed62bf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f210a),
	.w1(32'h3a2aadf9),
	.w2(32'h3bf521ef),
	.w3(32'h3b7bf46a),
	.w4(32'hbb2c7dc9),
	.w5(32'hbb2220b0),
	.w6(32'hb967bf99),
	.w7(32'h3a2efc50),
	.w8(32'h3afefc0e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbe5e4),
	.w1(32'hbb61da36),
	.w2(32'hba2b8b2d),
	.w3(32'hbb261a54),
	.w4(32'hbb608e61),
	.w5(32'hbc22b43d),
	.w6(32'h3b08adc5),
	.w7(32'h3b3e4498),
	.w8(32'h3bf8f239),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a6493),
	.w1(32'hbb9a4c9f),
	.w2(32'h3bbc66bf),
	.w3(32'h3a04bb54),
	.w4(32'hbb48c7d3),
	.w5(32'h3c0d3eb8),
	.w6(32'h3a941619),
	.w7(32'hbb1629d2),
	.w8(32'h39d703e5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47eafb),
	.w1(32'h3b000449),
	.w2(32'h3c221922),
	.w3(32'h3bbfbac8),
	.w4(32'hbbd49d61),
	.w5(32'h3d4e2cb2),
	.w6(32'hba95e988),
	.w7(32'h3b826ae4),
	.w8(32'h3c2207f2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91535b),
	.w1(32'hbb1cbb44),
	.w2(32'hbc0dd729),
	.w3(32'hbba11122),
	.w4(32'hbb03d116),
	.w5(32'hbc83507d),
	.w6(32'hba64b3d6),
	.w7(32'hbb8519e6),
	.w8(32'hbbb64229),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad9db1),
	.w1(32'hba735d21),
	.w2(32'h3bfec548),
	.w3(32'hbbdfcd2c),
	.w4(32'h3898f4b6),
	.w5(32'h3b01919d),
	.w6(32'h3bcac951),
	.w7(32'h3c07401c),
	.w8(32'hbc0aba19),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7dd6c),
	.w1(32'hb97128c2),
	.w2(32'hbc2e1bcc),
	.w3(32'hbbb57cbb),
	.w4(32'h3b2f17cf),
	.w5(32'hbcc3a217),
	.w6(32'h3bb42cb3),
	.w7(32'hba676615),
	.w8(32'hbc3db158),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8db0e4),
	.w1(32'h3b356b10),
	.w2(32'hbb5cfbee),
	.w3(32'h3afd84ce),
	.w4(32'hbb4710bb),
	.w5(32'hbc7a4435),
	.w6(32'hba91ef1f),
	.w7(32'h3a43efe7),
	.w8(32'h3b581b6d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49bc15),
	.w1(32'hbaeb187a),
	.w2(32'h3c199728),
	.w3(32'hb9adb4d0),
	.w4(32'hbc161538),
	.w5(32'h3c525a63),
	.w6(32'h3babb882),
	.w7(32'hbb0fcfed),
	.w8(32'hbc37668d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc66c92),
	.w1(32'hbb12af64),
	.w2(32'h3b48578b),
	.w3(32'hbbf703ca),
	.w4(32'hbb4c8abe),
	.w5(32'h3b950fca),
	.w6(32'h3adf93d3),
	.w7(32'hbb3a5780),
	.w8(32'h3c02d501),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bceb841),
	.w1(32'hbb6fe541),
	.w2(32'h3c0044bc),
	.w3(32'h37ce6392),
	.w4(32'hbc1ef158),
	.w5(32'h3b5561d2),
	.w6(32'h3c08b6b8),
	.w7(32'hbb8d9dd0),
	.w8(32'hbaf94e89),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3dfa),
	.w1(32'hbb6bb680),
	.w2(32'h3bd6b5f2),
	.w3(32'h3b1051e0),
	.w4(32'hbc1d2718),
	.w5(32'hba8ba867),
	.w6(32'h3b77f5f1),
	.w7(32'hbbaf9ea6),
	.w8(32'h3b3fba5a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a7435),
	.w1(32'h398f2bae),
	.w2(32'hbbb45fe3),
	.w3(32'h3c46df2a),
	.w4(32'hbb89fd06),
	.w5(32'hbb869b6e),
	.w6(32'h3ad7590a),
	.w7(32'hbb4ffd57),
	.w8(32'hbabd75cc),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91ab3e),
	.w1(32'h3b89af8e),
	.w2(32'hbae0e69f),
	.w3(32'h375da4db),
	.w4(32'h3c09e429),
	.w5(32'hbc4c8836),
	.w6(32'h3b278ea5),
	.w7(32'hbbdca314),
	.w8(32'hbb2574c3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab971a1),
	.w1(32'h3c33e836),
	.w2(32'h3b66fbba),
	.w3(32'h3a8f0205),
	.w4(32'h3b9bcb57),
	.w5(32'h391476ae),
	.w6(32'hb8d9c36c),
	.w7(32'h3ba3d94d),
	.w8(32'hbc01c259),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09246b),
	.w1(32'h3895824b),
	.w2(32'hbc0e54fc),
	.w3(32'hbb21ee4b),
	.w4(32'h3b01620a),
	.w5(32'hbc030629),
	.w6(32'h3b4831f5),
	.w7(32'hbaadc520),
	.w8(32'hbafccfa5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ffda),
	.w1(32'hbabcac66),
	.w2(32'hbc1c42b5),
	.w3(32'h3aecf52d),
	.w4(32'hbbca11ee),
	.w5(32'hbcb1d257),
	.w6(32'hbbb09c49),
	.w7(32'hbabdd684),
	.w8(32'hbc3049e3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b559081),
	.w1(32'h3bec35df),
	.w2(32'hbafcf1b0),
	.w3(32'h3beaa081),
	.w4(32'h3bcae4b3),
	.w5(32'hbb23ab32),
	.w6(32'h3ba7bd51),
	.w7(32'h39ead3a1),
	.w8(32'h3ba5d0a0),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e03993),
	.w1(32'hbb4670c8),
	.w2(32'h3ae95723),
	.w3(32'h3b385d84),
	.w4(32'hbb7be69c),
	.w5(32'h3a810bd9),
	.w6(32'h3b3d25d8),
	.w7(32'h3abc2074),
	.w8(32'hbb13256d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae02f6a),
	.w1(32'hbb26a21d),
	.w2(32'h3b50a093),
	.w3(32'hb832d05f),
	.w4(32'hbc125004),
	.w5(32'h3c910864),
	.w6(32'hb94c766f),
	.w7(32'hbba235f7),
	.w8(32'hbb00e14d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21cab8),
	.w1(32'hbb023e0f),
	.w2(32'h398a5478),
	.w3(32'h3a0f5d09),
	.w4(32'hbc1b10dc),
	.w5(32'hba97ef2d),
	.w6(32'h3ac2d334),
	.w7(32'h3b4d2980),
	.w8(32'h3a8389cc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06d6c6),
	.w1(32'hbaa4eac4),
	.w2(32'h3b1dc9fc),
	.w3(32'hbc226d8d),
	.w4(32'hbbf67d5f),
	.w5(32'hba0c6347),
	.w6(32'h3b29b3a6),
	.w7(32'hbc09aaf6),
	.w8(32'hbaf797c2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a7a17),
	.w1(32'hbafa21c0),
	.w2(32'h3b9113a8),
	.w3(32'hbbe26447),
	.w4(32'hbc379c26),
	.w5(32'h3cbb485a),
	.w6(32'h3980426e),
	.w7(32'hbb8b2684),
	.w8(32'h3c0d4045),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbc64a),
	.w1(32'h39de521b),
	.w2(32'h3ad31a16),
	.w3(32'hbc5a1b84),
	.w4(32'hbc8606c4),
	.w5(32'h3d01309a),
	.w6(32'hbc0c26fe),
	.w7(32'h3b74e63e),
	.w8(32'hba4e6253),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b2666),
	.w1(32'h3bd91407),
	.w2(32'hbb1b3e91),
	.w3(32'hbbd0d002),
	.w4(32'hb846ce4c),
	.w5(32'hbae235cd),
	.w6(32'h3b5de43f),
	.w7(32'h3b8cc08a),
	.w8(32'hbb5f7fd6),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89e62c),
	.w1(32'h3c3bf944),
	.w2(32'h3a4536c9),
	.w3(32'h3c02afb5),
	.w4(32'hbad5a980),
	.w5(32'h3bea9d2b),
	.w6(32'h3b6f0c6f),
	.w7(32'h37296702),
	.w8(32'h3b2911a8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f979),
	.w1(32'hbafb8ee5),
	.w2(32'hbbcb6de5),
	.w3(32'h3b928d7d),
	.w4(32'hbafdad5c),
	.w5(32'h3c07ad03),
	.w6(32'hbb246a02),
	.w7(32'h3adf7263),
	.w8(32'h3a60403f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad61674),
	.w1(32'hbb38fbc7),
	.w2(32'hbb5fde1c),
	.w3(32'h3badd0de),
	.w4(32'hbc0afcba),
	.w5(32'hbb511575),
	.w6(32'h3b8239d3),
	.w7(32'hba97703b),
	.w8(32'hbba4a272),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb236a),
	.w1(32'h3add6270),
	.w2(32'h3c0f1bef),
	.w3(32'hbc1248e9),
	.w4(32'hba51090d),
	.w5(32'h3c8aaa8a),
	.w6(32'hbc17a028),
	.w7(32'h3b990d86),
	.w8(32'h3b934f6b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b692332),
	.w1(32'h3be3de8c),
	.w2(32'h3be7591c),
	.w3(32'h3cc56000),
	.w4(32'hbaae9e7f),
	.w5(32'h3d0bd6d1),
	.w6(32'h3c21e6be),
	.w7(32'h3babd600),
	.w8(32'h3c0b0535),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01ced0),
	.w1(32'h3b549aa9),
	.w2(32'h3c1da773),
	.w3(32'hbc18070d),
	.w4(32'hbd0c8e2d),
	.w5(32'h3d8c4017),
	.w6(32'hbbda0dd0),
	.w7(32'hbb4c1ef3),
	.w8(32'hbb8f2ea8),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac360f8),
	.w1(32'hbc044b14),
	.w2(32'hbb9665e0),
	.w3(32'hbbe26f1c),
	.w4(32'hbc60aa31),
	.w5(32'h3abb933d),
	.w6(32'h3be373be),
	.w7(32'hbbea13e1),
	.w8(32'hbb945485),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6a79),
	.w1(32'h3b87a567),
	.w2(32'h3824b31c),
	.w3(32'hbc06fbc6),
	.w4(32'hbc734059),
	.w5(32'h3cc06775),
	.w6(32'hbb1f883f),
	.w7(32'hbb14d13f),
	.w8(32'h3c8863c1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c079c45),
	.w1(32'h3c25f343),
	.w2(32'hbb2e3378),
	.w3(32'h3c939133),
	.w4(32'h3be366a8),
	.w5(32'hbc929c8e),
	.w6(32'h3c63c9f7),
	.w7(32'h39dcf586),
	.w8(32'h3bd2398a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9696f44),
	.w1(32'hbb2d2976),
	.w2(32'h3b739744),
	.w3(32'h3c4e18d6),
	.w4(32'hbbe5df99),
	.w5(32'hbb4ca41c),
	.w6(32'h3bbcbf0a),
	.w7(32'hbbce0b66),
	.w8(32'hbbeef9ee),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d0477),
	.w1(32'hbac56478),
	.w2(32'hbc4120e7),
	.w3(32'hbbf67e34),
	.w4(32'hbbe6f94a),
	.w5(32'hbc2a2d40),
	.w6(32'hbc1ef052),
	.w7(32'hbb925711),
	.w8(32'hbc3d527e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f203e6),
	.w1(32'hb8e0aa7f),
	.w2(32'hba9b0bfb),
	.w3(32'h3b908251),
	.w4(32'h3c71ee93),
	.w5(32'hbc5fc280),
	.w6(32'h3c0551b8),
	.w7(32'h3ad0c9c0),
	.w8(32'hbb91e22c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf901b1),
	.w1(32'h3a6f90e8),
	.w2(32'h3bfc158c),
	.w3(32'h3c41cf6e),
	.w4(32'hbc02abf3),
	.w5(32'h3b66eb2c),
	.w6(32'h3c1441d3),
	.w7(32'hbb25bf1c),
	.w8(32'hbb5d3ad0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567dad),
	.w1(32'hba769334),
	.w2(32'h3af84ccd),
	.w3(32'hbb5c7b75),
	.w4(32'hba964ae0),
	.w5(32'h3b8ea7b5),
	.w6(32'hbbaf3f06),
	.w7(32'h3a16be34),
	.w8(32'h3b9f2fbc),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fbb6a),
	.w1(32'h3b4dcb41),
	.w2(32'hbb7a06f3),
	.w3(32'h39478b46),
	.w4(32'h3b6939b3),
	.w5(32'hbbd53d59),
	.w6(32'h3c2cb259),
	.w7(32'hbbc270d2),
	.w8(32'hbc1e9dc6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc054d4a),
	.w1(32'hbaf5f13f),
	.w2(32'h3af59cb4),
	.w3(32'h3a920f69),
	.w4(32'hbbae4032),
	.w5(32'h3a40466c),
	.w6(32'hbc27ba80),
	.w7(32'hba9bff08),
	.w8(32'hbb22022b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b89f4),
	.w1(32'h3c0b6aa7),
	.w2(32'hbbdc0f81),
	.w3(32'hbca1d5fa),
	.w4(32'hbb831044),
	.w5(32'h3ca13f34),
	.w6(32'hbc017e43),
	.w7(32'hbb957969),
	.w8(32'h3c09ad49),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b6e06),
	.w1(32'h3a043973),
	.w2(32'h3a9dc433),
	.w3(32'hb9a41fe2),
	.w4(32'hbad4742b),
	.w5(32'h3c5d232b),
	.w6(32'h3bb35214),
	.w7(32'hbbe2a40a),
	.w8(32'h3bd90ef4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a544f),
	.w1(32'hbab13a19),
	.w2(32'hbb458d1b),
	.w3(32'h3ad4aeb8),
	.w4(32'hbbaafac2),
	.w5(32'hbbc39e8f),
	.w6(32'h3a7a1e98),
	.w7(32'hbc4e21d5),
	.w8(32'hbb019566),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6597da),
	.w1(32'hbbbfdea5),
	.w2(32'h3a895930),
	.w3(32'hba3e4861),
	.w4(32'hba0a37c6),
	.w5(32'hbba151d8),
	.w6(32'h3b395a3a),
	.w7(32'hbb858a13),
	.w8(32'hbc03ae84),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0e09),
	.w1(32'h3b0000a1),
	.w2(32'hbb451934),
	.w3(32'h3a5621b7),
	.w4(32'hbbd0d716),
	.w5(32'hbb41f8b8),
	.w6(32'hbac0efd9),
	.w7(32'h3bbfbc9e),
	.w8(32'hbb61504a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26c17a),
	.w1(32'hbbaf3fc6),
	.w2(32'hbc059d7d),
	.w3(32'h3b10bba1),
	.w4(32'hbbfe8b80),
	.w5(32'hbbb8b2dc),
	.w6(32'h3b4b3632),
	.w7(32'hbad4d984),
	.w8(32'hba481efe),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba319faa),
	.w1(32'hbb8fc0a9),
	.w2(32'hbb7c3a0c),
	.w3(32'hbae76494),
	.w4(32'hbc2b0c3a),
	.w5(32'h376663c8),
	.w6(32'hbb6339a7),
	.w7(32'hbc0cd50b),
	.w8(32'hbba6b0ab),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84764b),
	.w1(32'h3ba4b994),
	.w2(32'h3b32d343),
	.w3(32'h3a067392),
	.w4(32'hbc019e44),
	.w5(32'h3d08d012),
	.w6(32'h3a940aa8),
	.w7(32'hbb652021),
	.w8(32'h3c091232),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c3372),
	.w1(32'hbc08db22),
	.w2(32'h3ab3bf3b),
	.w3(32'hbb4730bb),
	.w4(32'hbb06cbac),
	.w5(32'hbb898900),
	.w6(32'h3af41c69),
	.w7(32'h3baee9c8),
	.w8(32'hbac678cc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dcbf1),
	.w1(32'h3ae76890),
	.w2(32'h3c00f126),
	.w3(32'h3b9794b8),
	.w4(32'hbbd9f70d),
	.w5(32'h3c8215f5),
	.w6(32'hbb13a547),
	.w7(32'hbb14840e),
	.w8(32'h3bc11997),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ce513),
	.w1(32'h3b9c7218),
	.w2(32'h3c1c4a49),
	.w3(32'hbbc87454),
	.w4(32'hbb808d12),
	.w5(32'h3cd63214),
	.w6(32'hbb41fbf3),
	.w7(32'h3a619a90),
	.w8(32'h3acc8f2a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1df46e),
	.w1(32'hbb68ef9d),
	.w2(32'h3c195d74),
	.w3(32'hbbb70f89),
	.w4(32'hbc105d22),
	.w5(32'h3cd5b967),
	.w6(32'hbab6a2a5),
	.w7(32'h3ad16d04),
	.w8(32'h3be3b6dc),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6124ca),
	.w1(32'hbb28f14d),
	.w2(32'hbb8a9314),
	.w3(32'hbb046002),
	.w4(32'hbc812aa0),
	.w5(32'h3beff9cd),
	.w6(32'hba8adc50),
	.w7(32'hbbf5d6df),
	.w8(32'hbc2de568),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba024e20),
	.w1(32'hbc33d1ac),
	.w2(32'hbc86b983),
	.w3(32'h3afe1b12),
	.w4(32'hbc5d8a66),
	.w5(32'hb9b133db),
	.w6(32'hbb94b55d),
	.w7(32'hbc25b507),
	.w8(32'hbc354e3c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18fb20),
	.w1(32'hbc15dbbb),
	.w2(32'hbb9963aa),
	.w3(32'hbc780a92),
	.w4(32'hbc5400b3),
	.w5(32'h3aa0aeb2),
	.w6(32'hbc70270d),
	.w7(32'hbbcf2fad),
	.w8(32'hbbe20501),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a70a),
	.w1(32'hbaf4cacd),
	.w2(32'hbb1ef0cd),
	.w3(32'hbb2bbd0e),
	.w4(32'h3acaffc9),
	.w5(32'h3ba02735),
	.w6(32'h3b5ca6d2),
	.w7(32'h3b5adeb7),
	.w8(32'h3b23c6de),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a580c21),
	.w1(32'h3af50d4f),
	.w2(32'h3b930f76),
	.w3(32'h3955e7ae),
	.w4(32'hba92f57d),
	.w5(32'hbc289432),
	.w6(32'h398ba9cf),
	.w7(32'h3b2a0151),
	.w8(32'hbad3f15d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9efd6e),
	.w1(32'hbc16b6e4),
	.w2(32'hbb3634e8),
	.w3(32'hbbc7d751),
	.w4(32'hbb13e700),
	.w5(32'hbb21ae57),
	.w6(32'hbb902e28),
	.w7(32'h38fd65a6),
	.w8(32'hba8a109e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40cce6),
	.w1(32'h3b960bca),
	.w2(32'hbab6738d),
	.w3(32'hbb8c8ccb),
	.w4(32'h3ae69635),
	.w5(32'h3bc85597),
	.w6(32'hbbd8473b),
	.w7(32'h3bd070a6),
	.w8(32'h3bbffe2a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf37a5b),
	.w1(32'hba76227f),
	.w2(32'h3adfcc77),
	.w3(32'hbacc4d17),
	.w4(32'hb9d8b2b6),
	.w5(32'hbbfce434),
	.w6(32'h3b8776cd),
	.w7(32'h3aa727d8),
	.w8(32'h3ba592ec),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b746fb7),
	.w1(32'h3a911190),
	.w2(32'h3a128dee),
	.w3(32'h3b4a6646),
	.w4(32'hbb979789),
	.w5(32'hb9c2f9d7),
	.w6(32'h38ed6a8d),
	.w7(32'hba638db2),
	.w8(32'hbaf85cb8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad123ab),
	.w1(32'h3a8ef829),
	.w2(32'hba60dce1),
	.w3(32'hbb477b8b),
	.w4(32'h3bc9c564),
	.w5(32'hbaebc83b),
	.w6(32'hbb6205d9),
	.w7(32'hb9cdf4cc),
	.w8(32'hbb14ba9b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc373f4c),
	.w1(32'hbba97c84),
	.w2(32'hbb0dbb24),
	.w3(32'hbb0dd903),
	.w4(32'hbaab0dc8),
	.w5(32'hbc1d36e1),
	.w6(32'hbc0bf2b8),
	.w7(32'h37434d56),
	.w8(32'hbb080f10),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b908f),
	.w1(32'h3b51b800),
	.w2(32'hba14530a),
	.w3(32'h39b5a3ab),
	.w4(32'hbbd09dbc),
	.w5(32'hbc02da66),
	.w6(32'hba990147),
	.w7(32'h3b15da23),
	.w8(32'h3bf245fd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96638e),
	.w1(32'hba851bb0),
	.w2(32'hbbfa904d),
	.w3(32'h3b49cb96),
	.w4(32'hbc8fbac9),
	.w5(32'h3cb2f8a6),
	.w6(32'h3ad0aa38),
	.w7(32'hbb9adfe2),
	.w8(32'h3b760369),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5e1af),
	.w1(32'h3bc9588f),
	.w2(32'hbb031e3d),
	.w3(32'hbbe6affb),
	.w4(32'hbc08977e),
	.w5(32'h3cbb3536),
	.w6(32'hbbf6d25d),
	.w7(32'h38991c01),
	.w8(32'h3c05993d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33791b),
	.w1(32'h3a7b914d),
	.w2(32'hbbb1d2de),
	.w3(32'h3b2f7283),
	.w4(32'h3c19d22a),
	.w5(32'hbc9b2c5e),
	.w6(32'hb9d5391e),
	.w7(32'h3c069647),
	.w8(32'hbba8e427),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcc58c),
	.w1(32'h3b06851b),
	.w2(32'hbbcb4046),
	.w3(32'hbb1430c1),
	.w4(32'h3bc5aabc),
	.w5(32'hbbfdd811),
	.w6(32'hbb92d815),
	.w7(32'hbbb103c8),
	.w8(32'hbc078a6d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d718),
	.w1(32'hbbffab22),
	.w2(32'hbc6ebbf9),
	.w3(32'h3baed3d5),
	.w4(32'hbc8c87c5),
	.w5(32'hbc8dcdbc),
	.w6(32'h3b6b6609),
	.w7(32'hbc43bab7),
	.w8(32'hbc7bb155),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcda3d6),
	.w1(32'hbbd94370),
	.w2(32'hbbfb0a8a),
	.w3(32'h3b82d63a),
	.w4(32'hbc3372a8),
	.w5(32'hbcaed545),
	.w6(32'hbbdde6be),
	.w7(32'hbbbae230),
	.w8(32'hbc3bb8a7),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f60f),
	.w1(32'hbc25869f),
	.w2(32'hbb495271),
	.w3(32'h3befac98),
	.w4(32'hbbffb68f),
	.w5(32'hbbe3d0f2),
	.w6(32'hbb5caa47),
	.w7(32'hbaf70fe8),
	.w8(32'hbb005d9b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa342fa),
	.w1(32'h3b8f09e9),
	.w2(32'h3bc5224d),
	.w3(32'hbb32a404),
	.w4(32'hbbb7a699),
	.w5(32'h3ca7ba96),
	.w6(32'hba0a35ca),
	.w7(32'hbb92f34b),
	.w8(32'h3b4e6ede),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1a4f1),
	.w1(32'h3b7b5676),
	.w2(32'h391e203d),
	.w3(32'hbc3070be),
	.w4(32'hbae30b65),
	.w5(32'h3b8f2f45),
	.w6(32'hbc1a3afe),
	.w7(32'h3b64a108),
	.w8(32'hbb047987),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5813b7),
	.w1(32'h3ba27e78),
	.w2(32'hbb110a54),
	.w3(32'h3c84160d),
	.w4(32'hbb468088),
	.w5(32'h3ac05496),
	.w6(32'h3c14b3e0),
	.w7(32'hbb5f4144),
	.w8(32'hbb25f781),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1b87e),
	.w1(32'h3c08a2ef),
	.w2(32'h3b4dfd35),
	.w3(32'hbbbe21f8),
	.w4(32'h3bc58157),
	.w5(32'h3bd51089),
	.w6(32'hbba1eb34),
	.w7(32'h3c64c75c),
	.w8(32'h3bf9f6c7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e117c),
	.w1(32'hbbd80ac9),
	.w2(32'h3ad1d97f),
	.w3(32'hbae3db1b),
	.w4(32'hbae62978),
	.w5(32'hbb168ead),
	.w6(32'h3bacbecc),
	.w7(32'h3a11c483),
	.w8(32'h3c04c86c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b22c5),
	.w1(32'hbba0bca9),
	.w2(32'h3c087e52),
	.w3(32'h3c36147e),
	.w4(32'hbc3dca9f),
	.w5(32'h3be88891),
	.w6(32'h3c26fa73),
	.w7(32'hb98ec92d),
	.w8(32'hbb269701),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b5e1f),
	.w1(32'h3915b7eb),
	.w2(32'h3ac27ac6),
	.w3(32'hbc3e0990),
	.w4(32'h3882f3e1),
	.w5(32'h3afb337d),
	.w6(32'hbafe63f3),
	.w7(32'h3c0931f2),
	.w8(32'hbb681c8a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63090e),
	.w1(32'hbb5df655),
	.w2(32'hbbf16e4a),
	.w3(32'h3b2a58b3),
	.w4(32'hba13b319),
	.w5(32'hba0a04d4),
	.w6(32'h3baa0090),
	.w7(32'h3b980be2),
	.w8(32'hbb0c70a7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe95b6),
	.w1(32'hbb8a6bfd),
	.w2(32'h3bf4c701),
	.w3(32'hbc050859),
	.w4(32'hbbe229c7),
	.w5(32'hbb3d5777),
	.w6(32'hbc0af691),
	.w7(32'hbbde101e),
	.w8(32'hbbfd1d53),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba6ccb),
	.w1(32'hba8d0a1e),
	.w2(32'h3bc0c622),
	.w3(32'h3aa4ac3d),
	.w4(32'hb980fea0),
	.w5(32'h3b31fe27),
	.w6(32'hbb36f656),
	.w7(32'hbb57b624),
	.w8(32'hbbb4fdd2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab67a7b),
	.w1(32'hb962167d),
	.w2(32'hbbd500b1),
	.w3(32'hbb3df09b),
	.w4(32'hbc103b48),
	.w5(32'hbbb3b662),
	.w6(32'hbb81fb1c),
	.w7(32'hba88b23c),
	.w8(32'hbbe16b37),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87036b),
	.w1(32'h3b352416),
	.w2(32'h3a32681b),
	.w3(32'hbb175369),
	.w4(32'h3a3be1e1),
	.w5(32'hbb623e1f),
	.w6(32'hbaaf294a),
	.w7(32'hb918a8f8),
	.w8(32'hbba31eeb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb747c03),
	.w1(32'hbbb330d3),
	.w2(32'hbbb4dbec),
	.w3(32'hb9a3787d),
	.w4(32'hba67862e),
	.w5(32'h3a9a25fa),
	.w6(32'h3c2b55ca),
	.w7(32'hbb9ded29),
	.w8(32'hbab2af61),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2618),
	.w1(32'hbbcfa3c4),
	.w2(32'hbbfdd39b),
	.w3(32'h3b29de4a),
	.w4(32'hbbd54b6e),
	.w5(32'hbc7bd1c5),
	.w6(32'hbb27599c),
	.w7(32'hbb9d32f0),
	.w8(32'hbbf7c312),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eb204),
	.w1(32'h3b65e258),
	.w2(32'hba709bd4),
	.w3(32'hbbd61859),
	.w4(32'h3c28efed),
	.w5(32'h3c0ba3b7),
	.w6(32'hbba6e072),
	.w7(32'h3a999256),
	.w8(32'h3b2072d0),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3616a),
	.w1(32'h3bc6cd5e),
	.w2(32'h3c3704bb),
	.w3(32'h3b212e1e),
	.w4(32'h3ba49dad),
	.w5(32'h3c02f7b9),
	.w6(32'h3bc4a180),
	.w7(32'hbae80623),
	.w8(32'h3af0694d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46c37b),
	.w1(32'hbbcda0f2),
	.w2(32'hbb81101b),
	.w3(32'h3bfc75d3),
	.w4(32'hbc14509c),
	.w5(32'h3c2e0365),
	.w6(32'h3b165ab9),
	.w7(32'hbc20b47b),
	.w8(32'hbc22e733),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8010a3),
	.w1(32'hb7b9d72d),
	.w2(32'hbb7409a2),
	.w3(32'h3aac5fc9),
	.w4(32'h3b203d5d),
	.w5(32'h3b855916),
	.w6(32'hbbfa753f),
	.w7(32'h3aeab54e),
	.w8(32'h3ac59b2d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf15e71),
	.w1(32'hbba38461),
	.w2(32'h3b32840e),
	.w3(32'hbb5217b4),
	.w4(32'hbba04ed8),
	.w5(32'hb9eecea4),
	.w6(32'hbaae1355),
	.w7(32'hbb4f9895),
	.w8(32'hbbb3d963),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62490b),
	.w1(32'hbb5d7c96),
	.w2(32'hbc3e6ecc),
	.w3(32'hbb6ac68b),
	.w4(32'h3b8f0e16),
	.w5(32'hba3d04a9),
	.w6(32'hbb621e97),
	.w7(32'h3c3cd566),
	.w8(32'h3c6e0f61),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4171da),
	.w1(32'h399e4b3a),
	.w2(32'hba547d4f),
	.w3(32'hbbd1e978),
	.w4(32'h3a266700),
	.w5(32'h3afbb32f),
	.w6(32'h3bdce9e8),
	.w7(32'h3af50ffc),
	.w8(32'h3b47f06a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a827d47),
	.w1(32'hbb868123),
	.w2(32'hbb80a136),
	.w3(32'hbaae6d0f),
	.w4(32'hbaae5723),
	.w5(32'hbb9e007e),
	.w6(32'hbb7cce34),
	.w7(32'h3b0fe430),
	.w8(32'hbafed361),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4026e),
	.w1(32'hbb0f896b),
	.w2(32'h398d7d1c),
	.w3(32'hbae39ead),
	.w4(32'hbb013f88),
	.w5(32'hbb4b1323),
	.w6(32'h3a3cc716),
	.w7(32'hbbdb4d4c),
	.w8(32'hbc06b3ef),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80c446),
	.w1(32'h3ac7c3fc),
	.w2(32'hbb2e072c),
	.w3(32'hbb90bc6f),
	.w4(32'hbb11c071),
	.w5(32'hbb08369a),
	.w6(32'hbc4bf526),
	.w7(32'h3a5bad2c),
	.w8(32'h3a519e4a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109e16),
	.w1(32'h3b87104d),
	.w2(32'h3b867a27),
	.w3(32'hbba65608),
	.w4(32'h3b669314),
	.w5(32'h3af57a28),
	.w6(32'hba7af995),
	.w7(32'hbb4a0380),
	.w8(32'hbbbf2453),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e11f9),
	.w1(32'hbaea5d34),
	.w2(32'hbad85a22),
	.w3(32'h3b1d83b6),
	.w4(32'hbb3316b2),
	.w5(32'h3c12d8fd),
	.w6(32'hbc1dc919),
	.w7(32'hbaf46d91),
	.w8(32'hbb922e12),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb738508),
	.w1(32'hbb10dc64),
	.w2(32'hbc17a68d),
	.w3(32'hb9d39260),
	.w4(32'hbb5be9f6),
	.w5(32'h3b90d66c),
	.w6(32'hbb8712a1),
	.w7(32'hbb191511),
	.w8(32'hbb4d0b03),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d813c),
	.w1(32'h3b133d63),
	.w2(32'h3c2502f6),
	.w3(32'hba130688),
	.w4(32'hbb9ff377),
	.w5(32'hb96d6848),
	.w6(32'hbbcd9204),
	.w7(32'hbb1704be),
	.w8(32'hbb89e372),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111536),
	.w1(32'hbb66b3f1),
	.w2(32'hbb35e1b6),
	.w3(32'hbb043531),
	.w4(32'hbb6fe129),
	.w5(32'h3b639acb),
	.w6(32'hbbd8413c),
	.w7(32'hbbb1b78d),
	.w8(32'h38a95206),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0df6dc),
	.w1(32'hbbdb5f84),
	.w2(32'hbae53771),
	.w3(32'hba10aa80),
	.w4(32'hbb34616b),
	.w5(32'hbba5b44d),
	.w6(32'hbb77576f),
	.w7(32'h39a6eb0e),
	.w8(32'hb8a5c457),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3eb99),
	.w1(32'hba941999),
	.w2(32'hbb4447d6),
	.w3(32'hbbae1009),
	.w4(32'h3bad4a76),
	.w5(32'h3c0052d6),
	.w6(32'hbbf3e9e0),
	.w7(32'hbab1ce33),
	.w8(32'h3ba57444),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bfffe),
	.w1(32'hbbb8faef),
	.w2(32'hbc4667fe),
	.w3(32'h3c4c58bf),
	.w4(32'hba81b382),
	.w5(32'hbb8821a7),
	.w6(32'h3b186092),
	.w7(32'h3b351ee7),
	.w8(32'hb92d3c4c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dd90a),
	.w1(32'h3a950611),
	.w2(32'hbb81257e),
	.w3(32'hbc1d835b),
	.w4(32'h3a07ceea),
	.w5(32'h3bad7914),
	.w6(32'hba97a0fb),
	.w7(32'hbb5492fc),
	.w8(32'h39906c61),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66110c),
	.w1(32'h3aec1cad),
	.w2(32'h3a85311e),
	.w3(32'h3b805a9c),
	.w4(32'hbb51e213),
	.w5(32'h3bc79f1f),
	.w6(32'h3bcd1989),
	.w7(32'hbb9b990d),
	.w8(32'hbc0134d4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b981f66),
	.w1(32'hbb46f8ae),
	.w2(32'h3956424e),
	.w3(32'h3ba8d1d4),
	.w4(32'hbbfbe28f),
	.w5(32'hbc139aed),
	.w6(32'h3aeb9e76),
	.w7(32'hbc315e72),
	.w8(32'hbc895728),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adef39d),
	.w1(32'hbb6e21fe),
	.w2(32'hbbbc2364),
	.w3(32'h3b6198be),
	.w4(32'hbbc5e31c),
	.w5(32'hbb5959fa),
	.w6(32'hbc38293b),
	.w7(32'hbac84081),
	.w8(32'hbab3e580),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3722adc1),
	.w1(32'hbb131eda),
	.w2(32'hbb430517),
	.w3(32'h3bc99582),
	.w4(32'h3b7859cf),
	.w5(32'h3c356d8e),
	.w6(32'hbb931c42),
	.w7(32'h3b31310b),
	.w8(32'h3c822511),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d64e3),
	.w1(32'h3bf2c4cf),
	.w2(32'h3bfcb5cb),
	.w3(32'hb9734daa),
	.w4(32'hba60e2b3),
	.w5(32'hbb3f724c),
	.w6(32'hba032fd1),
	.w7(32'h3ba19b68),
	.w8(32'h3bd047ca),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c0824),
	.w1(32'hbbb5e151),
	.w2(32'hbbf62f1c),
	.w3(32'hbb974195),
	.w4(32'hbae9354d),
	.w5(32'h3a4f8418),
	.w6(32'h3bb4d4be),
	.w7(32'hbb1bded3),
	.w8(32'hbb460802),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd933bf),
	.w1(32'hbc063b8a),
	.w2(32'hbc13d1ab),
	.w3(32'h3b976f87),
	.w4(32'h3a3f87c5),
	.w5(32'h3b2bafc9),
	.w6(32'hbb95f8d1),
	.w7(32'hb8e355bb),
	.w8(32'h3b1ded81),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc297),
	.w1(32'h3849a84b),
	.w2(32'h3a464169),
	.w3(32'hbb575e9c),
	.w4(32'hbad02adf),
	.w5(32'h3b514ed6),
	.w6(32'hbb304577),
	.w7(32'hbb692b26),
	.w8(32'hbb7abec1),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2867e),
	.w1(32'hbbca3411),
	.w2(32'hbbd74ad9),
	.w3(32'h3ba14240),
	.w4(32'hbbaeae10),
	.w5(32'hbbc0f278),
	.w6(32'hbb6995cd),
	.w7(32'hbb2bba18),
	.w8(32'hbbc50272),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc145b3c),
	.w1(32'hbbec3f1c),
	.w2(32'hbbc8dbf9),
	.w3(32'hbb40322c),
	.w4(32'hbba4473b),
	.w5(32'hbb8314ea),
	.w6(32'hbbef0b38),
	.w7(32'hbc197e02),
	.w8(32'hbab2b37e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba33fc5),
	.w1(32'hbb12d107),
	.w2(32'h3a6846a7),
	.w3(32'hbb84e586),
	.w4(32'hbba1fd7a),
	.w5(32'hbb466d32),
	.w6(32'hbb4039c0),
	.w7(32'hbb596029),
	.w8(32'hbb884fed),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b792784),
	.w1(32'hbaac96d1),
	.w2(32'hbb041b39),
	.w3(32'hbba103c1),
	.w4(32'hb9f17633),
	.w5(32'hb9cdc35a),
	.w6(32'hbb123952),
	.w7(32'h3b878efc),
	.w8(32'h3b665168),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba471eb8),
	.w1(32'h3a8ef104),
	.w2(32'hbaf33483),
	.w3(32'hba46f0e3),
	.w4(32'h3ab85acd),
	.w5(32'hb982ca2d),
	.w6(32'h3ade6553),
	.w7(32'hbbc4bc35),
	.w8(32'hbb949e0d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb022db),
	.w1(32'hbc13af7a),
	.w2(32'hbbacf2c8),
	.w3(32'hba1a1dcf),
	.w4(32'hbc0162c6),
	.w5(32'hbb8363fe),
	.w6(32'hbb81bc60),
	.w7(32'h3996dcb9),
	.w8(32'h3b825bb6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e2f4),
	.w1(32'hbb34b454),
	.w2(32'hbb64f802),
	.w3(32'hbbac13ee),
	.w4(32'hbaef2cb3),
	.w5(32'hbbb1e294),
	.w6(32'hbb93f855),
	.w7(32'h39193f2e),
	.w8(32'h39c227a3),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6dd8c),
	.w1(32'hbba87c37),
	.w2(32'h3abb9ae1),
	.w3(32'hbbb422ce),
	.w4(32'hbafec00c),
	.w5(32'h3b47f7d6),
	.w6(32'hbb07af67),
	.w7(32'h3a06da04),
	.w8(32'hbbd358b2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc61c8),
	.w1(32'h3bbb65a2),
	.w2(32'hb848ee22),
	.w3(32'hb9fdc09b),
	.w4(32'hb9236d98),
	.w5(32'h3a89c73f),
	.w6(32'hbb1eddf9),
	.w7(32'h3bc185b4),
	.w8(32'h3c457280),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0c4dc),
	.w1(32'hb9e88ba0),
	.w2(32'h39d24b9c),
	.w3(32'hbb15faa7),
	.w4(32'hbac3be15),
	.w5(32'hba760ef4),
	.w6(32'h3a393f55),
	.w7(32'h3b195ee2),
	.w8(32'h3ab66e0d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3585be),
	.w1(32'hbbca9d97),
	.w2(32'hbbe9e1f3),
	.w3(32'hb9cc4cb9),
	.w4(32'hbb1dfa2e),
	.w5(32'hbba58c29),
	.w6(32'h398052f9),
	.w7(32'h3adb9a39),
	.w8(32'h3ac79ae2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16eb32),
	.w1(32'hbbc54148),
	.w2(32'hbc198124),
	.w3(32'hba592c3a),
	.w4(32'hbac45cd6),
	.w5(32'hbb808bde),
	.w6(32'hbb64a884),
	.w7(32'h3a5ac84c),
	.w8(32'h3b735d20),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc555960),
	.w1(32'hba5cc310),
	.w2(32'hbc08b11c),
	.w3(32'hbb67aa7b),
	.w4(32'h3ab08ead),
	.w5(32'hbb989268),
	.w6(32'h3b40c65a),
	.w7(32'h3c08585c),
	.w8(32'h3be49ee7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e3a3d),
	.w1(32'h3b63700f),
	.w2(32'h3c388c21),
	.w3(32'hbb42fade),
	.w4(32'h3b2694b9),
	.w5(32'h3bd1d7e4),
	.w6(32'h3b90e4a0),
	.w7(32'hb98a5679),
	.w8(32'hbbbd2af0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ca0d),
	.w1(32'hbb24e2a3),
	.w2(32'hbbb722d4),
	.w3(32'h3b60afba),
	.w4(32'h3a664f49),
	.w5(32'h3aa2f8b2),
	.w6(32'hbb7f45ae),
	.w7(32'h3bacfa6b),
	.w8(32'h3b402a17),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0e62),
	.w1(32'h3bbd290f),
	.w2(32'hbb5e2e30),
	.w3(32'h3b8733ea),
	.w4(32'h3ac21f85),
	.w5(32'hba5363cf),
	.w6(32'h3b32f5db),
	.w7(32'h3ad8f922),
	.w8(32'h3b8d59f1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e998f),
	.w1(32'h3abe500d),
	.w2(32'h3b1cde7f),
	.w3(32'h3a2bc1e8),
	.w4(32'hbb3f3c48),
	.w5(32'h3c76bc00),
	.w6(32'h3b8652c9),
	.w7(32'hbc004551),
	.w8(32'hbb6e7e57),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb500fb),
	.w1(32'hbc109b7f),
	.w2(32'hbbf9c005),
	.w3(32'h3c1bc40a),
	.w4(32'hbab577d7),
	.w5(32'hba635e91),
	.w6(32'hb7bbad75),
	.w7(32'hba87ab7d),
	.w8(32'hbbdd3897),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc441bd8),
	.w1(32'h3ae7c3af),
	.w2(32'h3beaeef4),
	.w3(32'hbb592756),
	.w4(32'h39e8742b),
	.w5(32'h3a229ecf),
	.w6(32'h38e8b875),
	.w7(32'hbbae00e8),
	.w8(32'hbb47ee14),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b5acf),
	.w1(32'h3a0fceb4),
	.w2(32'hbb0520b4),
	.w3(32'hb8d60d27),
	.w4(32'hbc101eee),
	.w5(32'hbb58ca38),
	.w6(32'hbb7ec452),
	.w7(32'hbba820c1),
	.w8(32'hbbf2870d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45997),
	.w1(32'hbb9f6448),
	.w2(32'h3a531e41),
	.w3(32'hbc1956e8),
	.w4(32'hbb64afe7),
	.w5(32'h3870dfdb),
	.w6(32'hbbae6cd8),
	.w7(32'hbb3fa843),
	.w8(32'hbaf773a7),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cd80e),
	.w1(32'hbafefd47),
	.w2(32'hbbf68501),
	.w3(32'hbac792af),
	.w4(32'h3b39a35a),
	.w5(32'h3b0e711e),
	.w6(32'hbbcfab4a),
	.w7(32'h3bb81006),
	.w8(32'h3c13cd8e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3e3db),
	.w1(32'h3a84ddf2),
	.w2(32'hbb6f848b),
	.w3(32'h3aee5e64),
	.w4(32'hbb7174b0),
	.w5(32'h3b5ce821),
	.w6(32'h3b5bd3f1),
	.w7(32'h3ad16c7d),
	.w8(32'hbb2c0663),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc2a7c),
	.w1(32'hbadce400),
	.w2(32'h398b5f5c),
	.w3(32'hb9d48b82),
	.w4(32'hba799cd0),
	.w5(32'hbb198702),
	.w6(32'h3ab400c1),
	.w7(32'hba866c94),
	.w8(32'hbb951e97),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb123bb9),
	.w1(32'hbb97c5ae),
	.w2(32'hbaaf12d1),
	.w3(32'hba109808),
	.w4(32'hbb51a212),
	.w5(32'hbbef803a),
	.w6(32'hba3071ac),
	.w7(32'hbb92409e),
	.w8(32'hbbc220ff),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25ce17),
	.w1(32'h3bd89b54),
	.w2(32'h3c30d316),
	.w3(32'hbb2350cd),
	.w4(32'h3bd41995),
	.w5(32'h3aad8d97),
	.w6(32'hbbaa8563),
	.w7(32'hbb96a64d),
	.w8(32'hbb824bee),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule