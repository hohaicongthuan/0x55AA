module layer_10_featuremap_361(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb42053),
	.w1(32'hbc0bf14d),
	.w2(32'hbc15bd55),
	.w3(32'hbc19e12e),
	.w4(32'hbc4a1a5b),
	.w5(32'h3b8cda82),
	.w6(32'hbc15d167),
	.w7(32'hbc3b98bb),
	.w8(32'h3bb44947),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c753589),
	.w1(32'h3cc531b2),
	.w2(32'h3c6e879d),
	.w3(32'h3c69417e),
	.w4(32'h3a9ff788),
	.w5(32'hbb5c43ce),
	.w6(32'h3d7bff3c),
	.w7(32'h3c79a2b2),
	.w8(32'h3bb9cb4e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e38cd),
	.w1(32'h3b1bb58f),
	.w2(32'h3b92faa0),
	.w3(32'hba9b5ad5),
	.w4(32'h3be9ecdc),
	.w5(32'h3c69677a),
	.w6(32'hbbfc5379),
	.w7(32'hbb85369f),
	.w8(32'h3c1876b8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11a84b),
	.w1(32'h3c0dee8e),
	.w2(32'h3bd4a9c5),
	.w3(32'h3baff0f7),
	.w4(32'h3c42088d),
	.w5(32'h3c369a42),
	.w6(32'h3bb431a3),
	.w7(32'h3ba0a8c7),
	.w8(32'h3be2cb5d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5610a9),
	.w1(32'hbb7ce442),
	.w2(32'hb93b11e1),
	.w3(32'h3af79c12),
	.w4(32'h3b8bd7b5),
	.w5(32'h3a798305),
	.w6(32'h3b4d65cd),
	.w7(32'h3ae1a772),
	.w8(32'hbb1315e3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11676e),
	.w1(32'hbb6698fb),
	.w2(32'h391e4dab),
	.w3(32'hbb8595ac),
	.w4(32'h3ad52037),
	.w5(32'hb97f4bc8),
	.w6(32'hb81813f3),
	.w7(32'hbb5868c9),
	.w8(32'h387ce91c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd38403),
	.w1(32'h3c8cac90),
	.w2(32'h3c650645),
	.w3(32'hbbc56051),
	.w4(32'h3c3fef00),
	.w5(32'h3b9e60a3),
	.w6(32'h3b0ef273),
	.w7(32'h3b901306),
	.w8(32'h3b62eba8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb16c7b),
	.w1(32'h3c0ea226),
	.w2(32'h37ea99f0),
	.w3(32'h3b2a549b),
	.w4(32'h3bec6c33),
	.w5(32'hbc47b4dc),
	.w6(32'h3b9676e9),
	.w7(32'h3b67de55),
	.w8(32'hbbc5c837),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc164a57),
	.w1(32'hbc190c94),
	.w2(32'hbc01ce15),
	.w3(32'hbc49b002),
	.w4(32'hbc387cf2),
	.w5(32'h3b923b79),
	.w6(32'hbb63f037),
	.w7(32'hbbe83dd4),
	.w8(32'h3b110ef4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b1163),
	.w1(32'h3c34e89f),
	.w2(32'h3c8da42d),
	.w3(32'hbc0d7fe9),
	.w4(32'hb78bc9fc),
	.w5(32'h3adc4864),
	.w6(32'h3bd9de19),
	.w7(32'h3baf107e),
	.w8(32'h3c76567d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f2d5b),
	.w1(32'h3a7cc4ff),
	.w2(32'h3b118f6c),
	.w3(32'hba34876b),
	.w4(32'h3bab87c5),
	.w5(32'hbb9d0b32),
	.w6(32'h3b870b6a),
	.w7(32'hbaf48972),
	.w8(32'hbb946f8a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08fc70),
	.w1(32'h3b51e4c4),
	.w2(32'h3bb9125d),
	.w3(32'hbbdb3887),
	.w4(32'h3a52d940),
	.w5(32'hbac2368e),
	.w6(32'hbc1da78c),
	.w7(32'hbbc6842c),
	.w8(32'hbb5ad281),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d8fc5),
	.w1(32'h3c6923d6),
	.w2(32'h3c459193),
	.w3(32'hbca3c83c),
	.w4(32'hbc5c0d50),
	.w5(32'hbc1f5aa8),
	.w6(32'h3c210224),
	.w7(32'h3c5ce59d),
	.w8(32'h3a7bc08e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd56fc),
	.w1(32'h3c938451),
	.w2(32'h3c547703),
	.w3(32'h3b0418a4),
	.w4(32'h3b9c3b66),
	.w5(32'h3c0fca69),
	.w6(32'h3b7022bc),
	.w7(32'h3a5c253e),
	.w8(32'h3bb90c4e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cd327),
	.w1(32'hbb651115),
	.w2(32'hb929f098),
	.w3(32'h3b7a85f2),
	.w4(32'h3ad7afa1),
	.w5(32'hbbb4dd3c),
	.w6(32'h3b24923f),
	.w7(32'h3a94ac51),
	.w8(32'hbac67588),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10be55),
	.w1(32'h3c742669),
	.w2(32'h3c933d6b),
	.w3(32'h3bc784a7),
	.w4(32'hbb9fd575),
	.w5(32'hbb4ebbd4),
	.w6(32'h3ca9246d),
	.w7(32'h3bb8eca2),
	.w8(32'h3b4b6e92),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc630b),
	.w1(32'hbb3ccdd1),
	.w2(32'hbbc49663),
	.w3(32'hbc3a9c76),
	.w4(32'hbb954d64),
	.w5(32'hbb87f59a),
	.w6(32'h3c1d8255),
	.w7(32'hbbc3a694),
	.w8(32'hbbad0277),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be57d07),
	.w1(32'h3bc7b768),
	.w2(32'h3c78f136),
	.w3(32'hbbc6ba70),
	.w4(32'hbb73f58b),
	.w5(32'hbba9a50e),
	.w6(32'hb95d8697),
	.w7(32'h3b97ed7e),
	.w8(32'hbbc2b916),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a7695),
	.w1(32'hbc2b788b),
	.w2(32'h3b1e1091),
	.w3(32'hbcb87e6a),
	.w4(32'hbc80c38a),
	.w5(32'h3abeb5e7),
	.w6(32'hbc774edb),
	.w7(32'hbc152a13),
	.w8(32'h3bcbd949),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaa454),
	.w1(32'hbaf54bff),
	.w2(32'hba53448c),
	.w3(32'hbad7d3f8),
	.w4(32'hbb37111c),
	.w5(32'hbb0cc3e6),
	.w6(32'hbc7f9e38),
	.w7(32'hbb97fd5d),
	.w8(32'hbc11c9ff),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc116843),
	.w1(32'hb9c4d3ea),
	.w2(32'h3b2ea9a1),
	.w3(32'hbb1d0cf8),
	.w4(32'hbbe43d6d),
	.w5(32'h3a8e19b0),
	.w6(32'h3c8c4d68),
	.w7(32'hbb3ef82b),
	.w8(32'h3ad8ff42),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9908bbc),
	.w1(32'hbb4b0e13),
	.w2(32'h3a94615d),
	.w3(32'hbb4a9de5),
	.w4(32'hba67c400),
	.w5(32'hbb35f5ee),
	.w6(32'hbbb7344e),
	.w7(32'h3ab5bc49),
	.w8(32'h3aecc112),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb46a2c),
	.w1(32'h3ca8c5ce),
	.w2(32'h3cff6270),
	.w3(32'h3bd0617c),
	.w4(32'hbb5f3d28),
	.w5(32'h3c73f039),
	.w6(32'h3cd263d7),
	.w7(32'h3cb0c900),
	.w8(32'h3d242bce),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a46a5),
	.w1(32'h3bcb6cfb),
	.w2(32'h3bf29e10),
	.w3(32'hbb86776e),
	.w4(32'hbb711502),
	.w5(32'hbb6474df),
	.w6(32'h3c2f7301),
	.w7(32'h3bae7072),
	.w8(32'h3c82ab97),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c454a06),
	.w1(32'h3b10d172),
	.w2(32'h3bbc649c),
	.w3(32'h3b3b5eac),
	.w4(32'hbbfc4aab),
	.w5(32'h3a57cfdc),
	.w6(32'h3cb8df03),
	.w7(32'h3c54264d),
	.w8(32'h3b4d7779),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3f947),
	.w1(32'hbbd9da84),
	.w2(32'h3aa82839),
	.w3(32'hbc055146),
	.w4(32'hbb0a9829),
	.w5(32'h3b63abda),
	.w6(32'hbb855177),
	.w7(32'hbb69b9f1),
	.w8(32'h3b30ae91),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972908c),
	.w1(32'hbb04c9c9),
	.w2(32'h3b035f0a),
	.w3(32'hb88ed5c2),
	.w4(32'h3afcbf41),
	.w5(32'hba7489fc),
	.w6(32'h3baafac1),
	.w7(32'h3a393479),
	.w8(32'hbb61b427),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacaf27),
	.w1(32'hbb49c2bc),
	.w2(32'hbb644aaa),
	.w3(32'hbc1021ca),
	.w4(32'hbc0350c5),
	.w5(32'hbb61b791),
	.w6(32'hbc8da778),
	.w7(32'hbc531e58),
	.w8(32'hbbe9b3c6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33fbc2),
	.w1(32'hbb50d375),
	.w2(32'h3a4f77e7),
	.w3(32'hbbcae528),
	.w4(32'hbb872f90),
	.w5(32'h3b061f07),
	.w6(32'hbbfeaf95),
	.w7(32'hbbd04e40),
	.w8(32'hbb4fb781),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc0f17),
	.w1(32'h3b6b6b00),
	.w2(32'hbb52656a),
	.w3(32'h3990140b),
	.w4(32'h3a9a8d00),
	.w5(32'h3bf1210f),
	.w6(32'h3c1db7aa),
	.w7(32'h3bda288d),
	.w8(32'h3c5a22d5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28da99),
	.w1(32'hbc5c3d13),
	.w2(32'hbc091f48),
	.w3(32'h3bc81b3e),
	.w4(32'h3a2bb703),
	.w5(32'hbbd054cd),
	.w6(32'hbc1bc8ac),
	.w7(32'hbbcf594a),
	.w8(32'hbbeb51e0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04a1fa),
	.w1(32'h3c086cd8),
	.w2(32'hbb2f580a),
	.w3(32'hbb842746),
	.w4(32'hbc04f3a4),
	.w5(32'h3ac833bf),
	.w6(32'hbc914dee),
	.w7(32'hbb9eaa25),
	.w8(32'hbb3d9e56),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1799aa),
	.w1(32'h3a360020),
	.w2(32'h3b98094d),
	.w3(32'hbb8ca9d0),
	.w4(32'hbbaf3866),
	.w5(32'h396679e3),
	.w6(32'h3a063899),
	.w7(32'h3b460c1e),
	.w8(32'hbb2ecc78),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0ecf9),
	.w1(32'hbb5caa31),
	.w2(32'h3aeff940),
	.w3(32'h3b646c8c),
	.w4(32'h3c21afa2),
	.w5(32'h3be0b011),
	.w6(32'h3ae995f8),
	.w7(32'h3c1fab98),
	.w8(32'h3c0ccbeb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d2635),
	.w1(32'hbb7c35d2),
	.w2(32'h3b9d7514),
	.w3(32'h3a14a645),
	.w4(32'h3ae52c60),
	.w5(32'hbc0f2fbb),
	.w6(32'hbc867a89),
	.w7(32'h395f3dd0),
	.w8(32'hbbd6821e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7523f8),
	.w1(32'hbbc5f6d7),
	.w2(32'hbb2937d8),
	.w3(32'hbc01ab61),
	.w4(32'hbb0a4c9f),
	.w5(32'h38b5208e),
	.w6(32'h3b4741b0),
	.w7(32'hbbdba64b),
	.w8(32'hbc1818c8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad1906),
	.w1(32'h3c606b63),
	.w2(32'h3c7b3969),
	.w3(32'h3cbc81fb),
	.w4(32'h3b7358eb),
	.w5(32'h3b3e5e24),
	.w6(32'h3c8e3828),
	.w7(32'h3bb2354a),
	.w8(32'h3b356dba),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbccbc9),
	.w1(32'hbcbf00d2),
	.w2(32'h3bfbdbc1),
	.w3(32'hbc04fa43),
	.w4(32'hbc86d293),
	.w5(32'h3bc8aceb),
	.w6(32'h3c8f79f1),
	.w7(32'hbc02abc0),
	.w8(32'h3bbb7c47),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2054e7),
	.w1(32'hbc12a08b),
	.w2(32'h3c5944c7),
	.w3(32'hbac607b4),
	.w4(32'h3b9696f5),
	.w5(32'h3c9ea0ae),
	.w6(32'h3c23f128),
	.w7(32'h3b17b304),
	.w8(32'h3cc83a00),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f00fb),
	.w1(32'hba8edcc1),
	.w2(32'hbb7c7cc9),
	.w3(32'h3c19ee3f),
	.w4(32'hbc61a676),
	.w5(32'hbbedc5cb),
	.w6(32'hbc1ea4dd),
	.w7(32'h3a4fcbf3),
	.w8(32'h39b330c6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ab15f),
	.w1(32'h3bb7cc87),
	.w2(32'hbc2e7c55),
	.w3(32'h3b0cd681),
	.w4(32'h3ac39ecf),
	.w5(32'h3b952ef2),
	.w6(32'h3b491296),
	.w7(32'h39eab12f),
	.w8(32'h3b5cb5a7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae35b57),
	.w1(32'h3adea186),
	.w2(32'h3bbdb0ff),
	.w3(32'hba827554),
	.w4(32'h3baf84f8),
	.w5(32'hba93840d),
	.w6(32'h3c287b75),
	.w7(32'hba15dd13),
	.w8(32'hbbdfab6f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119f1d),
	.w1(32'hbbf65800),
	.w2(32'h3be90718),
	.w3(32'hbba2e25e),
	.w4(32'hbc2671e9),
	.w5(32'h3c04b501),
	.w6(32'h3bbadec2),
	.w7(32'hbbad323b),
	.w8(32'h3c496ee3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca45b6e),
	.w1(32'h3ca4825b),
	.w2(32'h3cad5755),
	.w3(32'h3b3caf54),
	.w4(32'hbb6429ce),
	.w5(32'h3c3c69ff),
	.w6(32'h3d589724),
	.w7(32'h3c04614f),
	.w8(32'h3d11ef9d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc766ac),
	.w1(32'h3ca36d2c),
	.w2(32'h3c86bb61),
	.w3(32'h3c6bcd5c),
	.w4(32'h3c0472fb),
	.w5(32'hbb3a1dde),
	.w6(32'h3bb711cf),
	.w7(32'h3c966ee0),
	.w8(32'h3b579ce3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5b9e8),
	.w1(32'hbb6283b5),
	.w2(32'h3bca6067),
	.w3(32'hbc95a834),
	.w4(32'hbc5f24e0),
	.w5(32'hbc21e606),
	.w6(32'h3c62b3a2),
	.w7(32'h3c3bbbc9),
	.w8(32'h3c34db04),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64b4a5),
	.w1(32'h3b9d840b),
	.w2(32'h3c5fda5f),
	.w3(32'hbb467d9f),
	.w4(32'hbb84a322),
	.w5(32'hbb28867d),
	.w6(32'h3c14b96a),
	.w7(32'h3c3b0fe7),
	.w8(32'h3bf3ef93),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf35d9c),
	.w1(32'h3bd1ae44),
	.w2(32'h3c6bf5da),
	.w3(32'hbc9ff48d),
	.w4(32'hbc0887e1),
	.w5(32'hbb845372),
	.w6(32'h3bbb5561),
	.w7(32'h3b3fc1be),
	.w8(32'h3c5bdf8d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad005d7),
	.w1(32'hbb19fab6),
	.w2(32'hbbbdf3a2),
	.w3(32'hbc1e026f),
	.w4(32'hbbc3b3c9),
	.w5(32'hb996a11a),
	.w6(32'h3b6cfa13),
	.w7(32'hbba4bcb4),
	.w8(32'h3b19b14e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01c908),
	.w1(32'hba66b1de),
	.w2(32'h3b2a3a77),
	.w3(32'hbb4efdc8),
	.w4(32'h3b71efb1),
	.w5(32'h3c03f897),
	.w6(32'hbb10d576),
	.w7(32'h3b765943),
	.w8(32'h3c75e3a4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8d00),
	.w1(32'h3be4296a),
	.w2(32'hbba7b613),
	.w3(32'h3a975ad0),
	.w4(32'hbb215f12),
	.w5(32'h3c6634ff),
	.w6(32'h3aff211a),
	.w7(32'hbb2dad13),
	.w8(32'h3ca0c0e6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce5c27a),
	.w1(32'h3cc577a1),
	.w2(32'h3caa95b9),
	.w3(32'h3cac3cc4),
	.w4(32'h3c5ff467),
	.w5(32'h3c2d1d93),
	.w6(32'h3c30d9a5),
	.w7(32'h3c85a3ae),
	.w8(32'h3c40b9a9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61c301),
	.w1(32'hbb702158),
	.w2(32'h398e2c9e),
	.w3(32'h3bf164b6),
	.w4(32'h3c2a370c),
	.w5(32'hbafec266),
	.w6(32'h3a8e1bf6),
	.w7(32'h3b9b7748),
	.w8(32'h3b1f3afc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcf82c),
	.w1(32'h3bdfcb4b),
	.w2(32'h3c3887de),
	.w3(32'hbb2acda2),
	.w4(32'hbb42203f),
	.w5(32'h3a4ef1cf),
	.w6(32'hba865db7),
	.w7(32'h3c93cbbf),
	.w8(32'h3c8b60e6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b083e26),
	.w1(32'hbab6841d),
	.w2(32'hbb3c04b3),
	.w3(32'hbb2f4f7c),
	.w4(32'hbacacca5),
	.w5(32'h3badb3af),
	.w6(32'hbbf926e8),
	.w7(32'hbb52e082),
	.w8(32'h3b8d8151),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4463b3),
	.w1(32'h3aa3888f),
	.w2(32'hbbe2b690),
	.w3(32'hbbb9ac63),
	.w4(32'h3a855efd),
	.w5(32'h3afc8a02),
	.w6(32'hbaa05014),
	.w7(32'hbc0d1530),
	.w8(32'h3ac5e12d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac14131),
	.w1(32'h3b3a31a3),
	.w2(32'h39acb3c0),
	.w3(32'h39ff02bf),
	.w4(32'hba7f64b8),
	.w5(32'hbc0f32f1),
	.w6(32'hbaf129e3),
	.w7(32'h3b66fb1e),
	.w8(32'hbbb82e74),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1c419),
	.w1(32'h3aff47ff),
	.w2(32'h3b43b0fb),
	.w3(32'h3b8ff6cc),
	.w4(32'h3afb9253),
	.w5(32'hbaef359e),
	.w6(32'h3c1f2927),
	.w7(32'h3c2d61bb),
	.w8(32'hbade9ae5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dbba0),
	.w1(32'hbbd5e7a3),
	.w2(32'h3a1ae9d0),
	.w3(32'hbbdb7043),
	.w4(32'h3a303699),
	.w5(32'h3b8acd91),
	.w6(32'hbc0712db),
	.w7(32'hbb76e034),
	.w8(32'h3bf8c486),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c265e80),
	.w1(32'h3a06856c),
	.w2(32'h3c00d19e),
	.w3(32'h3a217984),
	.w4(32'h3b8fa5ba),
	.w5(32'h3b2ea07a),
	.w6(32'h3c584d48),
	.w7(32'h3c697db7),
	.w8(32'hbb68511c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba197e2),
	.w1(32'hbb02614f),
	.w2(32'h3b95b227),
	.w3(32'hbb1fa3fa),
	.w4(32'hbb71dd1b),
	.w5(32'h3bd11be3),
	.w6(32'h3b89b93d),
	.w7(32'h3b527d55),
	.w8(32'h3b04e1c6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb6a53),
	.w1(32'h3c13335b),
	.w2(32'h3c7f971d),
	.w3(32'hbb642f50),
	.w4(32'hbb01677a),
	.w5(32'h39593b9d),
	.w6(32'h3bea94fe),
	.w7(32'hbb4001c9),
	.w8(32'h3c13f620),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b8f35),
	.w1(32'hbb2cf1ad),
	.w2(32'h3b35c33b),
	.w3(32'hbb61a8a8),
	.w4(32'h3a3f4acb),
	.w5(32'hbb614b70),
	.w6(32'h3bb450c7),
	.w7(32'h3c2412a9),
	.w8(32'hbb1f2d2c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3372a9),
	.w1(32'h3aa76b3a),
	.w2(32'hbb7b5d97),
	.w3(32'h3a56aca6),
	.w4(32'hb8c1642e),
	.w5(32'h3c2c94a4),
	.w6(32'hbbe49072),
	.w7(32'hbb8112f6),
	.w8(32'h382e7f81),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b492e4a),
	.w1(32'h3be7d9db),
	.w2(32'h3b29faea),
	.w3(32'h3aff4344),
	.w4(32'hbb1c9c23),
	.w5(32'hbb8e5410),
	.w6(32'hbbca8888),
	.w7(32'hbbd23860),
	.w8(32'hbb5e3953),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374a62ff),
	.w1(32'hb9401080),
	.w2(32'hbb5879c0),
	.w3(32'hbb02d7ee),
	.w4(32'hbb2e682f),
	.w5(32'hbb748e3e),
	.w6(32'hbb821576),
	.w7(32'h3b14ff50),
	.w8(32'hba7bb0c6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fd294),
	.w1(32'h3c45894c),
	.w2(32'h3c9ae3d9),
	.w3(32'hbbcaa9e9),
	.w4(32'hbb4e7885),
	.w5(32'hbc1b0459),
	.w6(32'hba58e226),
	.w7(32'hbaa8e7a1),
	.w8(32'h3bfa01a6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacd08b),
	.w1(32'h3c116f79),
	.w2(32'h3c9dcef2),
	.w3(32'hbbc3680c),
	.w4(32'h3c077673),
	.w5(32'h3c156b23),
	.w6(32'h3d35894b),
	.w7(32'h3cd779b2),
	.w8(32'h3cdee4cf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63e434),
	.w1(32'h3c6dd39f),
	.w2(32'h3c60e634),
	.w3(32'hbb7e977c),
	.w4(32'hbb789d11),
	.w5(32'h3c74d9c1),
	.w6(32'h3c18d7ef),
	.w7(32'h3c19a3ce),
	.w8(32'h3cc46815),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa33e30),
	.w1(32'h3aad953c),
	.w2(32'h3c233765),
	.w3(32'hbb534e00),
	.w4(32'hbbc83141),
	.w5(32'h3c674956),
	.w6(32'h3d369cfe),
	.w7(32'h3c169fd0),
	.w8(32'h3ccddc83),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc76fbb),
	.w1(32'hba2eb3e5),
	.w2(32'h3a74fe99),
	.w3(32'h3b8a004c),
	.w4(32'h3b9314a0),
	.w5(32'hbc0cf8a6),
	.w6(32'hbbf0ee81),
	.w7(32'hba1ecc41),
	.w8(32'hbbe57708),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1c704),
	.w1(32'hb8db8786),
	.w2(32'hbb3b6ebc),
	.w3(32'hbb34f308),
	.w4(32'hba96a547),
	.w5(32'hbb66b714),
	.w6(32'h3aaf0381),
	.w7(32'hbbb82cfa),
	.w8(32'hbbdcb365),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0985),
	.w1(32'hbaf4a6fd),
	.w2(32'hbaff6c23),
	.w3(32'hbc0fffae),
	.w4(32'h3a9e1503),
	.w5(32'h3afd1aea),
	.w6(32'hbb9f4298),
	.w7(32'hbc02631a),
	.w8(32'hb9bd3415),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b425a0a),
	.w1(32'h3b812a84),
	.w2(32'h3c17efa9),
	.w3(32'h3c92d6cf),
	.w4(32'hbb099a45),
	.w5(32'hbb2efa63),
	.w6(32'h3d2f813e),
	.w7(32'h3ce15662),
	.w8(32'h3b041c7a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3393dd),
	.w1(32'hbbb39b8d),
	.w2(32'hbb6d442b),
	.w3(32'hbbe5d6a8),
	.w4(32'hbb8b4fa2),
	.w5(32'hbb8d72f1),
	.w6(32'h3b8d217e),
	.w7(32'hbc034a46),
	.w8(32'h3b5788ad),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e1df),
	.w1(32'h3c4e6d7b),
	.w2(32'h3bc3f088),
	.w3(32'h3a0d7778),
	.w4(32'hbae47a4f),
	.w5(32'h3a688a2a),
	.w6(32'h3cc4ddbd),
	.w7(32'h3c329766),
	.w8(32'h3c29482d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8dc09),
	.w1(32'h3be42406),
	.w2(32'h3bd0e9e8),
	.w3(32'hba99513d),
	.w4(32'hbb931fa9),
	.w5(32'hbafb1d01),
	.w6(32'h3c6bf2dc),
	.w7(32'h3bedff20),
	.w8(32'h3b095105),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac98cd),
	.w1(32'h3ae9badf),
	.w2(32'h3a131821),
	.w3(32'hbb8c9a1a),
	.w4(32'h3a6e5402),
	.w5(32'h3c32d896),
	.w6(32'hbc8a3e4e),
	.w7(32'h3b5e3fdc),
	.w8(32'h3c5c36de),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a460b),
	.w1(32'h3a294cc9),
	.w2(32'h3cb4812e),
	.w3(32'h3b8b5661),
	.w4(32'h3c5c3202),
	.w5(32'hbb4e0ce3),
	.w6(32'hbc8d3364),
	.w7(32'h3c0009e2),
	.w8(32'h3b65f035),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395375ea),
	.w1(32'h3a5500f5),
	.w2(32'h3bbf6356),
	.w3(32'hbc88676e),
	.w4(32'hbbd4fbc0),
	.w5(32'h3c975be7),
	.w6(32'h3c0e06f1),
	.w7(32'hbb1eea26),
	.w8(32'h3ceba7ce),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89b9f2),
	.w1(32'h3cd56cda),
	.w2(32'h3c89693f),
	.w3(32'h3cbd0bbc),
	.w4(32'h3bdade70),
	.w5(32'h3ae8d902),
	.w6(32'h3c69fc48),
	.w7(32'h3c319747),
	.w8(32'h3c0437cd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58594c),
	.w1(32'h39b65b09),
	.w2(32'h3bb17481),
	.w3(32'hba1ec099),
	.w4(32'hbb1c67b1),
	.w5(32'h3a11d2ed),
	.w6(32'h3bafeb8a),
	.w7(32'h3be45c9f),
	.w8(32'h3c1e5587),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba504976),
	.w1(32'h3b8bd577),
	.w2(32'hbb2b1e56),
	.w3(32'h3b2f880c),
	.w4(32'h3b7760d7),
	.w5(32'h3ba39c59),
	.w6(32'hb769d557),
	.w7(32'h3bc6094b),
	.w8(32'h3bfc748c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa37c6d),
	.w1(32'h3ad3281c),
	.w2(32'h3ba72334),
	.w3(32'h3b05f1b9),
	.w4(32'h3b3f9562),
	.w5(32'hbb58d128),
	.w6(32'h3d0828bd),
	.w7(32'h3aee128e),
	.w8(32'h3a64f946),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cb070),
	.w1(32'h3b9feed9),
	.w2(32'h3a63e9bd),
	.w3(32'hbb1760e3),
	.w4(32'hbbd5994f),
	.w5(32'hbb5b50e1),
	.w6(32'h3bca9482),
	.w7(32'h3bc65316),
	.w8(32'hbbdec57a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02297d),
	.w1(32'h3adf8246),
	.w2(32'h3b65099d),
	.w3(32'hbbc68daf),
	.w4(32'hbaa5937a),
	.w5(32'hb9f325d4),
	.w6(32'h3b37f081),
	.w7(32'h394cb857),
	.w8(32'hbb7ae93a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70aec6),
	.w1(32'hbb8b1f44),
	.w2(32'h3c0af99f),
	.w3(32'h3b54616f),
	.w4(32'hbb511fa9),
	.w5(32'h3b15d818),
	.w6(32'h3bd2e634),
	.w7(32'h3bc8d223),
	.w8(32'h3c174b4d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3d68c),
	.w1(32'hbb9813f3),
	.w2(32'hbb6a05e6),
	.w3(32'hb8d4f42d),
	.w4(32'hbb5a1d6e),
	.w5(32'hbba44868),
	.w6(32'hba9be7cd),
	.w7(32'h3b8ee421),
	.w8(32'hbbb0c044),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb2ddc),
	.w1(32'hbb0b390b),
	.w2(32'hbbb0f95f),
	.w3(32'hbb7f9f48),
	.w4(32'hbbb590fd),
	.w5(32'hbc15640c),
	.w6(32'h3c8803ae),
	.w7(32'h3bc34242),
	.w8(32'h3b7e8ca9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb10f6),
	.w1(32'h3af8f299),
	.w2(32'hbb72fe8d),
	.w3(32'hbc419069),
	.w4(32'hbac48ca3),
	.w5(32'h3bbc2a18),
	.w6(32'h3bc692f7),
	.w7(32'h3911e49e),
	.w8(32'h3cb4948d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a2d86),
	.w1(32'hbc1f96a3),
	.w2(32'hba4a75a6),
	.w3(32'h3ab431b8),
	.w4(32'hb9e80128),
	.w5(32'h3bdfcdae),
	.w6(32'h3a0ae388),
	.w7(32'hbab60957),
	.w8(32'h3c2e85b9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5efe2),
	.w1(32'h3c998429),
	.w2(32'h3cd5a3b2),
	.w3(32'hbc01c26b),
	.w4(32'h3ba405cf),
	.w5(32'hb9da1266),
	.w6(32'h3bb79ac5),
	.w7(32'h3c4d7e8f),
	.w8(32'h3cc611d2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb432e06),
	.w1(32'h3cb1023e),
	.w2(32'h3b6f6be9),
	.w3(32'h3b97a495),
	.w4(32'h3b738f91),
	.w5(32'h3b27f12d),
	.w6(32'h3c26d2eb),
	.w7(32'h3bc02cd8),
	.w8(32'h3c38e209),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc15ec2),
	.w1(32'h3c57f335),
	.w2(32'h3c5faf9c),
	.w3(32'hbb4cfd53),
	.w4(32'hbb292f4c),
	.w5(32'hbc15b88f),
	.w6(32'h3cafd998),
	.w7(32'h3bf2926e),
	.w8(32'h3a431e32),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36d36b),
	.w1(32'hbb225fa8),
	.w2(32'h3bd8178a),
	.w3(32'hbba6c67f),
	.w4(32'hbaecf684),
	.w5(32'h3b4d210f),
	.w6(32'hba08518d),
	.w7(32'h3bd54028),
	.w8(32'h3b72db7d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc107cf6),
	.w1(32'hbc28a090),
	.w2(32'h3ba9ceae),
	.w3(32'hbc15f436),
	.w4(32'hbbf29ada),
	.w5(32'h3cbf2588),
	.w6(32'hbc954447),
	.w7(32'hbc348f76),
	.w8(32'h3cfd6258),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac5f2f),
	.w1(32'h3c1bbdf8),
	.w2(32'h3c57b390),
	.w3(32'h3c91540c),
	.w4(32'h3c4f7539),
	.w5(32'hbb8b0f12),
	.w6(32'hbc06a85f),
	.w7(32'h3c7c8e5c),
	.w8(32'hbb2ea952),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b806903),
	.w1(32'h3c0d9863),
	.w2(32'hb8cb4c3c),
	.w3(32'hbbf5570c),
	.w4(32'hbb524014),
	.w5(32'h3b97c174),
	.w6(32'hbbcf6b14),
	.w7(32'h3ae0a081),
	.w8(32'h3c78f06f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b1164),
	.w1(32'h3c371f06),
	.w2(32'h3c9568a8),
	.w3(32'hbab317b8),
	.w4(32'h3c28bffe),
	.w5(32'h3c432396),
	.w6(32'h3b78e8dd),
	.w7(32'h3c566061),
	.w8(32'h3c92c0de),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c746cf8),
	.w1(32'h3c9b2fbf),
	.w2(32'h3ca0e0f9),
	.w3(32'h3c1db025),
	.w4(32'h3c29792e),
	.w5(32'h3c257cd2),
	.w6(32'h3c86bb98),
	.w7(32'h3bb908ad),
	.w8(32'h3c8b3fee),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84172f),
	.w1(32'hbc3684ce),
	.w2(32'hbb663f65),
	.w3(32'h3c08e213),
	.w4(32'hbc6846a7),
	.w5(32'hbc1d30aa),
	.w6(32'h3c83c89c),
	.w7(32'hbbb4a479),
	.w8(32'hbc0ad5c0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914679),
	.w1(32'h3b81203a),
	.w2(32'h3ba20eaa),
	.w3(32'h3b1525b1),
	.w4(32'hb99bb4f0),
	.w5(32'h39aade39),
	.w6(32'h3c29e94e),
	.w7(32'h3c3cb3fe),
	.w8(32'h3c14c83e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8836ca),
	.w1(32'h3c7d0939),
	.w2(32'h3c9bc1db),
	.w3(32'h3a96c9ec),
	.w4(32'h3b320992),
	.w5(32'h3a29dd19),
	.w6(32'h3c0c8fa8),
	.w7(32'h3bd11e89),
	.w8(32'h3c1271b7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38f789),
	.w1(32'hbb2a10b3),
	.w2(32'hbb9ef731),
	.w3(32'hbac59e6f),
	.w4(32'hbaef68f8),
	.w5(32'hb9837cf8),
	.w6(32'hbb839636),
	.w7(32'hbb9965e4),
	.w8(32'h3a762d37),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf5a8d),
	.w1(32'h3c9f11bc),
	.w2(32'h3caa881d),
	.w3(32'h3c45231d),
	.w4(32'h3b07233c),
	.w5(32'h3ba732f8),
	.w6(32'h3c990f2f),
	.w7(32'h3b752ab4),
	.w8(32'h3c2a70ed),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b5436),
	.w1(32'h39193637),
	.w2(32'h3c754d3b),
	.w3(32'hbbd9374d),
	.w4(32'h3a012c63),
	.w5(32'h3ca3580b),
	.w6(32'hbc01037a),
	.w7(32'h372a6b84),
	.w8(32'h3c1e4bd2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0425c5),
	.w1(32'hbab48be7),
	.w2(32'h3a723bbf),
	.w3(32'h3a0ec21d),
	.w4(32'h3af99a60),
	.w5(32'h3ba93785),
	.w6(32'hbb50a0c0),
	.w7(32'h3a0e197c),
	.w8(32'h3b8bc62d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c003d4f),
	.w1(32'h3c03e85b),
	.w2(32'h3bcf9d68),
	.w3(32'h3bb3a118),
	.w4(32'h3ae8e631),
	.w5(32'h3bf0f804),
	.w6(32'h3c24c083),
	.w7(32'h3bf5d9f9),
	.w8(32'h3be3e5c3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba289c6),
	.w1(32'h3b5226c8),
	.w2(32'h3c4566da),
	.w3(32'hbba1fa70),
	.w4(32'h3afc1d31),
	.w5(32'h3c0778e8),
	.w6(32'hb997614b),
	.w7(32'h3bc4f12c),
	.w8(32'h3c414bf9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c125fe9),
	.w1(32'h3bb0524b),
	.w2(32'h3c15a55a),
	.w3(32'h3b9bb321),
	.w4(32'hb8c36791),
	.w5(32'hb990c667),
	.w6(32'h3c14343d),
	.w7(32'h3bcbe8e8),
	.w8(32'h3bd19615),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dbad0),
	.w1(32'hbb971338),
	.w2(32'hbaf981a6),
	.w3(32'hba581121),
	.w4(32'hbbca993c),
	.w5(32'hba023b24),
	.w6(32'hb8f858b9),
	.w7(32'hbaccca3f),
	.w8(32'h3b9f1aa9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83b37e),
	.w1(32'h3ba03e89),
	.w2(32'h3bb07c27),
	.w3(32'hb5c9d280),
	.w4(32'hbaf7384c),
	.w5(32'h3c012d71),
	.w6(32'h3b52de47),
	.w7(32'h3b974627),
	.w8(32'h3c5fb0fc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ccc56),
	.w1(32'hbc009d16),
	.w2(32'hbb5de10f),
	.w3(32'hbc505df6),
	.w4(32'hbc2f0abb),
	.w5(32'hbb4e6e8b),
	.w6(32'h3bf16fa4),
	.w7(32'h3ac56aa8),
	.w8(32'h3bd0e80b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c754b62),
	.w1(32'h3c8fc326),
	.w2(32'h3c71de5a),
	.w3(32'h3b1ca866),
	.w4(32'h3b993fd0),
	.w5(32'h3a9588e8),
	.w6(32'h3b6bcbd0),
	.w7(32'h3b8ae0ab),
	.w8(32'h3c2ec247),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51e609),
	.w1(32'h3a27c0a7),
	.w2(32'hba5c94e3),
	.w3(32'h3af65177),
	.w4(32'h3b4ff398),
	.w5(32'h3acf1d5d),
	.w6(32'h3b199c4e),
	.w7(32'h3b7bc919),
	.w8(32'h3b9bbfe4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d776a1),
	.w1(32'hba023d31),
	.w2(32'hba08c90d),
	.w3(32'hba6dbca3),
	.w4(32'hbb07855a),
	.w5(32'hb99a061e),
	.w6(32'hbaa83796),
	.w7(32'hbaa803bd),
	.w8(32'h3b2a6816),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74282c),
	.w1(32'h3b652af2),
	.w2(32'h3ae9fe25),
	.w3(32'hba716931),
	.w4(32'hbafd800b),
	.w5(32'hb8e0a27b),
	.w6(32'h3b75db23),
	.w7(32'h3b0a12f9),
	.w8(32'h3ae0cf2e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab24f2b),
	.w1(32'h3a62a249),
	.w2(32'h3aa8f694),
	.w3(32'h39281917),
	.w4(32'h3b58e7ce),
	.w5(32'h3ba55eca),
	.w6(32'h3a6dc07a),
	.w7(32'h3ab0bc7e),
	.w8(32'hbaf701c4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b77fd),
	.w1(32'hb942e2df),
	.w2(32'h3a7dcf33),
	.w3(32'h39bd9654),
	.w4(32'h3b3c68d0),
	.w5(32'h3bc57cb5),
	.w6(32'hbb8c3aba),
	.w7(32'hbb159f6b),
	.w8(32'h3ae7d2cb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc60d93),
	.w1(32'h3b50d887),
	.w2(32'h3b9d3dd7),
	.w3(32'h3b57280d),
	.w4(32'h3b0f4254),
	.w5(32'hbb7524be),
	.w6(32'h3bc8a2a1),
	.w7(32'h3bdc488f),
	.w8(32'h3b896150),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4565a0),
	.w1(32'hb9999fbb),
	.w2(32'hba9c7ba2),
	.w3(32'h3a89cafc),
	.w4(32'hbacccce1),
	.w5(32'h3b39f2ef),
	.w6(32'h3a7c3a54),
	.w7(32'hba2afbbf),
	.w8(32'hba7bceb5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96f6bc),
	.w1(32'hb9db52bf),
	.w2(32'h3b092c38),
	.w3(32'hbb6ceb98),
	.w4(32'hbb29bf93),
	.w5(32'hbb8f79fa),
	.w6(32'hb9c4029b),
	.w7(32'h3b125a3b),
	.w8(32'hbb5deb4c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9cdfb),
	.w1(32'h3a09c846),
	.w2(32'h3bfc9157),
	.w3(32'hbaa57ec6),
	.w4(32'hbb9cf93e),
	.w5(32'h3c9d3009),
	.w6(32'hba717863),
	.w7(32'h3b231194),
	.w8(32'h3cd917e5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b2dd3),
	.w1(32'hbb02306d),
	.w2(32'h3a7b26c7),
	.w3(32'h39810752),
	.w4(32'hbb58edb5),
	.w5(32'hbb687fac),
	.w6(32'h3bb4ae5b),
	.w7(32'h3a61cd64),
	.w8(32'hbb8b58b3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb366e62),
	.w1(32'hbb6b3352),
	.w2(32'hbb220ba0),
	.w3(32'hbb843e8e),
	.w4(32'hbb540b51),
	.w5(32'h3aa9cdc3),
	.w6(32'hbb23e34e),
	.w7(32'hba6f22a0),
	.w8(32'hbb133340),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12e432),
	.w1(32'hbb02236e),
	.w2(32'hbafb0911),
	.w3(32'h3b656970),
	.w4(32'h3b89debc),
	.w5(32'h3b8014a5),
	.w6(32'hb9c85184),
	.w7(32'h398664d4),
	.w8(32'h3b453a1c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76ca26),
	.w1(32'h3ad299d3),
	.w2(32'h3b48aa54),
	.w3(32'hb8b22f9b),
	.w4(32'hb98e2580),
	.w5(32'h3ac511a7),
	.w6(32'h3b489b95),
	.w7(32'h3b18f2c6),
	.w8(32'h3af5783e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba038611),
	.w1(32'h3bd404df),
	.w2(32'h3b928646),
	.w3(32'hbbe9e4cb),
	.w4(32'h3a551a9b),
	.w5(32'h3c1d8423),
	.w6(32'h3c281222),
	.w7(32'h3c41f53b),
	.w8(32'h3c9b6662),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c873ce4),
	.w1(32'h3c4cd966),
	.w2(32'h3c5d78fc),
	.w3(32'hbb5eaefa),
	.w4(32'hb912fee0),
	.w5(32'hbae84597),
	.w6(32'h3bbfeb67),
	.w7(32'h3c0d0e95),
	.w8(32'h3bf4ddb9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75b1d5),
	.w1(32'hbb19ed30),
	.w2(32'h39ab6dac),
	.w3(32'hbb80d5ee),
	.w4(32'hbb7bb3e1),
	.w5(32'h3b2144d9),
	.w6(32'hbacfadf2),
	.w7(32'hba9d770e),
	.w8(32'h3ae71563),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb7b8),
	.w1(32'h3b76dbd5),
	.w2(32'h3aacb5dd),
	.w3(32'hba48fbc7),
	.w4(32'hba66d873),
	.w5(32'h3bb1dd6a),
	.w6(32'h3b80821b),
	.w7(32'h3b16dc54),
	.w8(32'h3bd77f8d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5c9f0),
	.w1(32'h39c6fb5b),
	.w2(32'hb8608b3b),
	.w3(32'h3ac773e3),
	.w4(32'hb9b3ef75),
	.w5(32'h3bcdf2ba),
	.w6(32'h3b999a63),
	.w7(32'h3b76901b),
	.w8(32'hbb2b362f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b253e77),
	.w1(32'h3b8157dd),
	.w2(32'h3ba52b7c),
	.w3(32'h3b8f8ca8),
	.w4(32'h3bb5e21d),
	.w5(32'h3b691fe6),
	.w6(32'hb6cce756),
	.w7(32'hb9daf13e),
	.w8(32'h3b82cec4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c742989),
	.w1(32'h3c6c97fd),
	.w2(32'h3c375d19),
	.w3(32'h3c263835),
	.w4(32'h3bcfa291),
	.w5(32'h3b7f4732),
	.w6(32'h3c354cb7),
	.w7(32'h3c3e0866),
	.w8(32'h3c78690f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c331824),
	.w1(32'h3c4c1d7d),
	.w2(32'h3ca56197),
	.w3(32'hbbd8ffe1),
	.w4(32'hbb60d7fb),
	.w5(32'h3b9963a3),
	.w6(32'h3b8d53c8),
	.w7(32'h3c24866d),
	.w8(32'h3c574132),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fe305),
	.w1(32'hbab91d4b),
	.w2(32'hbad294f6),
	.w3(32'h3a4caa81),
	.w4(32'hbbe109f2),
	.w5(32'h3a19905f),
	.w6(32'h3b303c51),
	.w7(32'hbb1bdd0f),
	.w8(32'h3b8fddf8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c296859),
	.w1(32'h3c156f59),
	.w2(32'h3bf61e6d),
	.w3(32'hbbcabf42),
	.w4(32'hbbbf27c2),
	.w5(32'h3c0f1a4a),
	.w6(32'h3c041c25),
	.w7(32'h3ba18f72),
	.w8(32'h3c8376eb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2178a4),
	.w1(32'h3c4636ea),
	.w2(32'h3c4982d8),
	.w3(32'h3b15d921),
	.w4(32'h3aa87448),
	.w5(32'h3b67dbab),
	.w6(32'h3c596c1d),
	.w7(32'h3c37c028),
	.w8(32'h3c5e65fc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8aa05),
	.w1(32'hbaba1786),
	.w2(32'hbaad11fe),
	.w3(32'h3ae38fe6),
	.w4(32'hbba65aa5),
	.w5(32'hba6d5af5),
	.w6(32'h3c626532),
	.w7(32'h3bbdba1f),
	.w8(32'h3ba37adb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd920e),
	.w1(32'h3ba28fbd),
	.w2(32'h3bcfca07),
	.w3(32'hb818d206),
	.w4(32'hba0bdfde),
	.w5(32'h3b8e509f),
	.w6(32'h3af6d2f7),
	.w7(32'h3b753879),
	.w8(32'h3c1a2067),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7fd7a),
	.w1(32'h3b58601b),
	.w2(32'h3b456439),
	.w3(32'h3ad5c3fb),
	.w4(32'h3ae246a8),
	.w5(32'hbb26ba80),
	.w6(32'h3b8b5865),
	.w7(32'h3b794b42),
	.w8(32'h3aa56f98),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb383e14),
	.w1(32'hba96e37f),
	.w2(32'hbb94eab8),
	.w3(32'hbb4cd3d0),
	.w4(32'h39d32bd4),
	.w5(32'h3be8cd5e),
	.w6(32'h3b21cc6b),
	.w7(32'h3ba6b0a7),
	.w8(32'h3c8865c5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfac32),
	.w1(32'h3b2a53ec),
	.w2(32'h3a5956e6),
	.w3(32'h3b45402d),
	.w4(32'hb904c81b),
	.w5(32'h3ab64487),
	.w6(32'h3c0ddcd8),
	.w7(32'h3b8b6788),
	.w8(32'h3b9f6659),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b096636),
	.w1(32'hbb0182a9),
	.w2(32'hbaa82fbf),
	.w3(32'hbb3801ee),
	.w4(32'hbae90167),
	.w5(32'h3b4dd1e7),
	.w6(32'hbb515642),
	.w7(32'hbabad421),
	.w8(32'h3b0667f6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3103ad),
	.w1(32'h3b5d1e67),
	.w2(32'h3b10a5d0),
	.w3(32'h38a851bd),
	.w4(32'hbacffbb6),
	.w5(32'h3abcd708),
	.w6(32'h3b0eb162),
	.w7(32'h3a26911d),
	.w8(32'h39d4c894),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b50c1),
	.w1(32'hbae8cc05),
	.w2(32'h3aa2f033),
	.w3(32'hb9236973),
	.w4(32'hbb07d4bb),
	.w5(32'hba70dd1c),
	.w6(32'h3b293962),
	.w7(32'h39dd5676),
	.w8(32'h3b8db800),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7599a4),
	.w1(32'hbb9565c1),
	.w2(32'hbb28b900),
	.w3(32'hb9f0788a),
	.w4(32'hbbb728c6),
	.w5(32'hbb5431b9),
	.w6(32'h3ba72cd2),
	.w7(32'h3aae74d4),
	.w8(32'h3b9cbce1),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10778e),
	.w1(32'h3adc6ca1),
	.w2(32'h3b9fdedc),
	.w3(32'hbc0f5b02),
	.w4(32'hbb593657),
	.w5(32'hbb93bb92),
	.w6(32'hbb844f40),
	.w7(32'h3b73c47b),
	.w8(32'h3bfcadf3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6ec74),
	.w1(32'hbae91657),
	.w2(32'hbad25d2f),
	.w3(32'hbb4addc8),
	.w4(32'hba8e9a4f),
	.w5(32'h3b0fef3b),
	.w6(32'hbb45797e),
	.w7(32'hba93f012),
	.w8(32'h3b81f755),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c806b33),
	.w1(32'h3c51bfb1),
	.w2(32'h3c484f53),
	.w3(32'h3a68cc0b),
	.w4(32'hb993854a),
	.w5(32'h394544f6),
	.w6(32'h3bf3925f),
	.w7(32'h3c144c86),
	.w8(32'h3c21b77b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44508a),
	.w1(32'hb9d186c7),
	.w2(32'h3a355daf),
	.w3(32'hbab2cf91),
	.w4(32'h3a457e66),
	.w5(32'hbbb522bb),
	.w6(32'h3a4ded5a),
	.w7(32'h3b7b1bc4),
	.w8(32'h3b5b11fd),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f1f49),
	.w1(32'h3c42920d),
	.w2(32'h3c255614),
	.w3(32'hbbc7e253),
	.w4(32'hba914a3f),
	.w5(32'hbb18eb79),
	.w6(32'hba7e9688),
	.w7(32'h3b7ddff0),
	.w8(32'h3b8050d1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6377f),
	.w1(32'h3be3d846),
	.w2(32'h3bfb7b4a),
	.w3(32'hbabb15e2),
	.w4(32'h3b6b9ac2),
	.w5(32'h3c5cea46),
	.w6(32'hbb476d7d),
	.w7(32'h3c4d27f0),
	.w8(32'h3ce76729),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c032b4d),
	.w1(32'h3bfb27be),
	.w2(32'h3c1185ea),
	.w3(32'h3befe96d),
	.w4(32'h3b04648a),
	.w5(32'h3ac622c8),
	.w6(32'h3c4098a3),
	.w7(32'h3b939e86),
	.w8(32'h3b6c001a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0341c),
	.w1(32'hbab04223),
	.w2(32'h3a59cb31),
	.w3(32'hbac09fe0),
	.w4(32'h3b2c88c0),
	.w5(32'h3bd0f5a8),
	.w6(32'hba36e726),
	.w7(32'h3ac1dddd),
	.w8(32'h3b36f36d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99d2ab),
	.w1(32'hbad225ad),
	.w2(32'h3b20cd94),
	.w3(32'hba9b7955),
	.w4(32'hbc003779),
	.w5(32'hb6171120),
	.w6(32'h3b9b91ef),
	.w7(32'hbabb8523),
	.w8(32'h3b341822),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e6e76),
	.w1(32'hbb207a63),
	.w2(32'h3b7d8703),
	.w3(32'h3c0343ef),
	.w4(32'hbac71503),
	.w5(32'h3bdd8aeb),
	.w6(32'h3c2b77c6),
	.w7(32'hb89625d4),
	.w8(32'h3bc35f65),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33f566),
	.w1(32'hbbec11fe),
	.w2(32'h3b4de448),
	.w3(32'h3a4925d0),
	.w4(32'hbba2ffc2),
	.w5(32'h3a8e3c3a),
	.w6(32'h3b7818bd),
	.w7(32'hb97e064a),
	.w8(32'h3b40a12d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9b4be),
	.w1(32'h3b8928f1),
	.w2(32'h3bb70eda),
	.w3(32'h3914671b),
	.w4(32'h3b49c265),
	.w5(32'h3a736ce2),
	.w6(32'h3b1dcd7d),
	.w7(32'h3b876b5d),
	.w8(32'h3b369b78),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf5a37),
	.w1(32'h3b40ddb2),
	.w2(32'hba6bc74b),
	.w3(32'h39476bf2),
	.w4(32'h3a8be0ec),
	.w5(32'hb9ffb85f),
	.w6(32'hbad40fce),
	.w7(32'h3ab10090),
	.w8(32'h39a6c184),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6fc7c),
	.w1(32'h3bd74ecb),
	.w2(32'h3c36917f),
	.w3(32'hbb27cbf6),
	.w4(32'hba75f48f),
	.w5(32'hb954f9b2),
	.w6(32'h3bb4c84e),
	.w7(32'h3bbf3e7c),
	.w8(32'h3b541692),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad62b94),
	.w1(32'hbb012a5a),
	.w2(32'h3b002fc5),
	.w3(32'hbac318a0),
	.w4(32'hb9f46fec),
	.w5(32'h3b40ec44),
	.w6(32'hbb1ece0c),
	.w7(32'hbaa622e7),
	.w8(32'hb9095f7d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ea574),
	.w1(32'hbb1e64f4),
	.w2(32'hbb0a17a5),
	.w3(32'h3b52d067),
	.w4(32'h3afa5293),
	.w5(32'h3a99fef7),
	.w6(32'h3b88c7f8),
	.w7(32'h3bb007b3),
	.w8(32'h3bbeeadf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e8b7b),
	.w1(32'h3987e767),
	.w2(32'h3a4a122c),
	.w3(32'hbb2062a1),
	.w4(32'hba8bcb86),
	.w5(32'hba152bb2),
	.w6(32'hbae885a4),
	.w7(32'hbafd5862),
	.w8(32'h3ab13fea),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392daa4f),
	.w1(32'h3bde1c6f),
	.w2(32'h3c7eb809),
	.w3(32'hbc339047),
	.w4(32'h3b866a61),
	.w5(32'h3c405e3c),
	.w6(32'hbb220184),
	.w7(32'h3bfb10ac),
	.w8(32'h3c8374e5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6dd90),
	.w1(32'hb788b85d),
	.w2(32'h3ac4f824),
	.w3(32'h3a4682ba),
	.w4(32'h3b0e9283),
	.w5(32'h3a0ca62d),
	.w6(32'h3ad829c3),
	.w7(32'h39fd4464),
	.w8(32'hbb85082e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb42545),
	.w1(32'hbb799ea7),
	.w2(32'h3a6344d0),
	.w3(32'h3a806e8c),
	.w4(32'hba9f9b1b),
	.w5(32'h3b092256),
	.w6(32'h3b39a7ad),
	.w7(32'h3b6f2960),
	.w8(32'h3b85baa5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2810fe),
	.w1(32'hbb8b9e57),
	.w2(32'hbb204f22),
	.w3(32'h3a9b4b4b),
	.w4(32'hbbb2c3ed),
	.w5(32'hbb65d585),
	.w6(32'h3baaa9e3),
	.w7(32'hbad2c7a3),
	.w8(32'hba81a98d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e9ba4),
	.w1(32'h3ae59314),
	.w2(32'h3bc726aa),
	.w3(32'hba54b591),
	.w4(32'hbbd22c3c),
	.w5(32'h3c295edd),
	.w6(32'h3c932fcc),
	.w7(32'h3ba472d4),
	.w8(32'h3ca747f7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41ed4c),
	.w1(32'h3b727898),
	.w2(32'h3bedb96b),
	.w3(32'h3b4e8fce),
	.w4(32'h3943e2fd),
	.w5(32'h3b03f78c),
	.w6(32'h3bd0f0e1),
	.w7(32'h3b559fa0),
	.w8(32'h3b6a0384),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b252154),
	.w1(32'h3aa4fb70),
	.w2(32'h3b952df0),
	.w3(32'h3a485f2d),
	.w4(32'hb9aa67e8),
	.w5(32'h3a182385),
	.w6(32'h3b9a6d60),
	.w7(32'h3b82057f),
	.w8(32'h3b98afb0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad36d4),
	.w1(32'h39399a78),
	.w2(32'h3aef9e53),
	.w3(32'hba107b69),
	.w4(32'h39d4fce5),
	.w5(32'h3addb0d8),
	.w6(32'hbbae055a),
	.w7(32'hb9b3bada),
	.w8(32'h3b12cf28),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3983b5),
	.w1(32'h3c39fc3d),
	.w2(32'h3c8e2fc3),
	.w3(32'h3b1a79eb),
	.w4(32'hbb86534f),
	.w5(32'h3b572054),
	.w6(32'h3bc6288b),
	.w7(32'h3c32b822),
	.w8(32'h3c6b5bd8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c590a1b),
	.w1(32'h3c2dc6af),
	.w2(32'h3c8ad960),
	.w3(32'h3b0bc016),
	.w4(32'h39f025a2),
	.w5(32'h3b89d9fa),
	.w6(32'h3c0a11d2),
	.w7(32'h3bec1f36),
	.w8(32'h3c030317),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17f7d1),
	.w1(32'h3c388e56),
	.w2(32'h3c1aef50),
	.w3(32'h3ad40ea9),
	.w4(32'h3b0f3f96),
	.w5(32'h3a3f4060),
	.w6(32'h3bd2de55),
	.w7(32'h3c2d4ca1),
	.w8(32'h3c65e3b8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad07a41),
	.w1(32'hba232f20),
	.w2(32'hba03a437),
	.w3(32'hbaeec7dc),
	.w4(32'hbb4d2e7a),
	.w5(32'hb9befac1),
	.w6(32'hba07bcf7),
	.w7(32'hbb01f8ec),
	.w8(32'hb846a3a9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf80be2),
	.w1(32'h3be80823),
	.w2(32'h3b80eca3),
	.w3(32'h3b83d5ff),
	.w4(32'h3ae1ca8f),
	.w5(32'h3b22190c),
	.w6(32'h3bf80476),
	.w7(32'h3beabc32),
	.w8(32'h3c2a956c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e1974),
	.w1(32'h3b071bb2),
	.w2(32'h3ac63f2f),
	.w3(32'h39fb52b9),
	.w4(32'h39e84509),
	.w5(32'hba565ccf),
	.w6(32'h3b1a8b38),
	.w7(32'h3ac04e21),
	.w8(32'hbb365845),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d9740),
	.w1(32'hbaf33034),
	.w2(32'h3b003559),
	.w3(32'h3a498e28),
	.w4(32'h3abf3ab0),
	.w5(32'h3b56a87a),
	.w6(32'hbb0580bd),
	.w7(32'h3ac3a21e),
	.w8(32'h3bcc0dfd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bc119),
	.w1(32'h3abde9bd),
	.w2(32'hba3eff73),
	.w3(32'h3b88dd8a),
	.w4(32'h3bb86efd),
	.w5(32'hbb05a76b),
	.w6(32'h3a542cda),
	.w7(32'hb9d18722),
	.w8(32'hbac63728),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49a906),
	.w1(32'h3b961f1b),
	.w2(32'h3bac640b),
	.w3(32'hb9e43375),
	.w4(32'hbb9838d7),
	.w5(32'h3bb2b91d),
	.w6(32'h3ad5714e),
	.w7(32'h389ebc6a),
	.w8(32'h3c36b101),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ad0d2),
	.w1(32'hb9ea3471),
	.w2(32'h3b22cd96),
	.w3(32'h3b0cbdc5),
	.w4(32'h3bb0bc2d),
	.w5(32'hbaa895e0),
	.w6(32'hb756b7dc),
	.w7(32'h3badfd96),
	.w8(32'hbaa28b7a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f7108),
	.w1(32'hbab3be3d),
	.w2(32'hbb8b39b5),
	.w3(32'h385bafc0),
	.w4(32'hb9d7430b),
	.w5(32'hba9fcf9e),
	.w6(32'hba90815e),
	.w7(32'hba79b454),
	.w8(32'hbb3e0bf1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fb393),
	.w1(32'hbb68ed6a),
	.w2(32'hbad8c34c),
	.w3(32'hbb8f6d0c),
	.w4(32'hbbaf1a57),
	.w5(32'hba8f0c48),
	.w6(32'hbaf7500b),
	.w7(32'hbaf9d45f),
	.w8(32'h3b18a2fc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb79337),
	.w1(32'h3c24ce9a),
	.w2(32'h3c1b9aa2),
	.w3(32'hba12634b),
	.w4(32'h3a54c394),
	.w5(32'h3c0a4bd6),
	.w6(32'h3bf3fe1f),
	.w7(32'h3c0dfc8e),
	.w8(32'h3c7c0701),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c593cea),
	.w1(32'h3c2519b9),
	.w2(32'h3be5582d),
	.w3(32'h3c0cb3b9),
	.w4(32'h3bac27d6),
	.w5(32'h3bd2f00a),
	.w6(32'h3be94a54),
	.w7(32'hb9f7a36e),
	.w8(32'h3beab8ba),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5fd7e),
	.w1(32'h3b80778b),
	.w2(32'h3b608034),
	.w3(32'h3ac2b115),
	.w4(32'h3adc7b19),
	.w5(32'hb984add3),
	.w6(32'h3b9ac2d9),
	.w7(32'h3b712000),
	.w8(32'hba8b71a5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c8243),
	.w1(32'h3c9ad13f),
	.w2(32'h3c8c8ba8),
	.w3(32'hbbb930e4),
	.w4(32'h3a8283a7),
	.w5(32'h3bcafb1b),
	.w6(32'h3af10e9c),
	.w7(32'h3c9ac1da),
	.w8(32'h3ca083a7),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25f52a),
	.w1(32'hbbf9aa52),
	.w2(32'h3bdbf6b1),
	.w3(32'h3c0b4ebe),
	.w4(32'hbc0c4416),
	.w5(32'h3ab3f3a5),
	.w6(32'h3bf30ab6),
	.w7(32'h3b1182f6),
	.w8(32'h3c820348),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dfbbd),
	.w1(32'h3b991d85),
	.w2(32'h3bdea2af),
	.w3(32'hbb45b5ac),
	.w4(32'hbaadbbfc),
	.w5(32'h3bc27e6b),
	.w6(32'h3b14acf1),
	.w7(32'h3b2d29f1),
	.w8(32'h3a7026bb),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c336e),
	.w1(32'hbb1ad2e7),
	.w2(32'hbabb2176),
	.w3(32'h3b7188ac),
	.w4(32'h3b4b7db5),
	.w5(32'h3a95ec1a),
	.w6(32'hba442a8a),
	.w7(32'hb9ae981b),
	.w8(32'h3a85bb06),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39660854),
	.w1(32'hba7683f9),
	.w2(32'hba0ad5fd),
	.w3(32'hb937cf5c),
	.w4(32'hbab454cf),
	.w5(32'hb99e61a7),
	.w6(32'h3a2e57d7),
	.w7(32'h39ad8c51),
	.w8(32'hbaafeda2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f1898),
	.w1(32'hbb8dab40),
	.w2(32'hbb07f386),
	.w3(32'h3a697d40),
	.w4(32'h3a017c56),
	.w5(32'hbaa0823a),
	.w6(32'h3565f08d),
	.w7(32'h3b3910f1),
	.w8(32'hbb6bfca8),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f15be),
	.w1(32'h3a551d53),
	.w2(32'h3b515078),
	.w3(32'hbb6f8eb7),
	.w4(32'h3b2b113a),
	.w5(32'h3bc06e23),
	.w6(32'hbba8033b),
	.w7(32'hb7098df4),
	.w8(32'h3ba6c280),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8f964),
	.w1(32'h3922df8f),
	.w2(32'hbaa1b16a),
	.w3(32'hbbb629bd),
	.w4(32'hbbfdc619),
	.w5(32'h3b2309b9),
	.w6(32'h3c0a67b6),
	.w7(32'h3b941e35),
	.w8(32'h3c284f5c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053f13),
	.w1(32'h3b712ceb),
	.w2(32'h3ba6bf1b),
	.w3(32'h3b543eb3),
	.w4(32'hb996aa87),
	.w5(32'hbc0ea024),
	.w6(32'h3baa2298),
	.w7(32'h3bd81d5e),
	.w8(32'h3a435c76),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83faa2),
	.w1(32'hbb170a60),
	.w2(32'h3a351764),
	.w3(32'hba9aca13),
	.w4(32'hbaa311f5),
	.w5(32'hbab9b1b5),
	.w6(32'h3b035928),
	.w7(32'h3b4020e0),
	.w8(32'h3988414e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba00b42),
	.w1(32'h3bcd8d3d),
	.w2(32'h3c518ee4),
	.w3(32'hbc1d74ed),
	.w4(32'hbbcc7bfa),
	.w5(32'hbab8dcc1),
	.w6(32'h3b54325a),
	.w7(32'h3b6bd4e6),
	.w8(32'h3c486426),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81420a),
	.w1(32'h3b88aaf2),
	.w2(32'h3bc7fea1),
	.w3(32'h3a926467),
	.w4(32'h3b3d876c),
	.w5(32'h3ba77693),
	.w6(32'hb844de15),
	.w7(32'h3b53e393),
	.w8(32'h3b9a8677),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba468b82),
	.w1(32'hbb4ea81a),
	.w2(32'hbaa998c6),
	.w3(32'hbb32e150),
	.w4(32'hbae5cd24),
	.w5(32'hba985322),
	.w6(32'hbb50a1c5),
	.w7(32'hbac36861),
	.w8(32'h3a29bd1a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85765b),
	.w1(32'h3bfd3d73),
	.w2(32'h3c03c803),
	.w3(32'hba9b97ff),
	.w4(32'hbacf1672),
	.w5(32'hb9b74151),
	.w6(32'h3bc29bde),
	.w7(32'h3a340164),
	.w8(32'h379adf3e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf2b4b),
	.w1(32'hb886507b),
	.w2(32'hb91b5a5a),
	.w3(32'h3a5985aa),
	.w4(32'h39902806),
	.w5(32'h3ae5c171),
	.w6(32'h3b2fe2df),
	.w7(32'h3a873eab),
	.w8(32'hb9901f91),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b8730),
	.w1(32'h3b174c6b),
	.w2(32'h3c8164d8),
	.w3(32'hbc193b58),
	.w4(32'hbbcd0a2c),
	.w5(32'h3c80f6b5),
	.w6(32'hbb3c06a6),
	.w7(32'h3b2fc500),
	.w8(32'h3cd8a267),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2a487),
	.w1(32'hbb94f0fd),
	.w2(32'h3baa619a),
	.w3(32'h3bb7d72e),
	.w4(32'hbbda6f21),
	.w5(32'h3be71aa8),
	.w6(32'h3c3628bd),
	.w7(32'hb82fe02e),
	.w8(32'h3c38ca8f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51fec5),
	.w1(32'hba930f86),
	.w2(32'h3b2f9e8b),
	.w3(32'h39a504ae),
	.w4(32'hbb6834c9),
	.w5(32'h3aec2e25),
	.w6(32'h3b8d2cb1),
	.w7(32'h3aaf89ef),
	.w8(32'h3bf3eb0d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc476),
	.w1(32'hbb2458a5),
	.w2(32'h39a31766),
	.w3(32'hbadcc20b),
	.w4(32'hbab5e621),
	.w5(32'h3b45ff2d),
	.w6(32'hbb5d154f),
	.w7(32'hbb827bb7),
	.w8(32'h3aa63a3d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a4d3b),
	.w1(32'hbacb7155),
	.w2(32'h3b5c1503),
	.w3(32'hbaecd7d8),
	.w4(32'hbba4d677),
	.w5(32'h3b8b42d1),
	.w6(32'h3adbb1c4),
	.w7(32'hb8c12a11),
	.w8(32'h3c2e464c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02a1ac),
	.w1(32'h3b97b98c),
	.w2(32'h3be8796b),
	.w3(32'hbaca9a81),
	.w4(32'hbb32de26),
	.w5(32'hbba1e76e),
	.w6(32'h3ba9fd86),
	.w7(32'h3b9c036f),
	.w8(32'h3993cc1d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f4c59),
	.w1(32'hbaebf102),
	.w2(32'h3b6ae93b),
	.w3(32'hbc84868d),
	.w4(32'hbc37c0d4),
	.w5(32'hbb9c3271),
	.w6(32'hbbe4ce74),
	.w7(32'h3b6bc5fb),
	.w8(32'h3bf1b151),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7bbfc),
	.w1(32'hb8f3e761),
	.w2(32'h39070230),
	.w3(32'h39b94cec),
	.w4(32'h3a9266d3),
	.w5(32'h393d751d),
	.w6(32'h3b130972),
	.w7(32'h3a925e0e),
	.w8(32'hbaf5e751),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba157f63),
	.w1(32'h3a4b6dbc),
	.w2(32'h3b0c6b13),
	.w3(32'hbab9d619),
	.w4(32'h37992e7b),
	.w5(32'h3b5d7b8a),
	.w6(32'hba542e0d),
	.w7(32'h3a3cfc9b),
	.w8(32'h3b1ba82b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36d4f3),
	.w1(32'h39b3e77e),
	.w2(32'h3c2e725d),
	.w3(32'hbaec361a),
	.w4(32'hbab1ad59),
	.w5(32'h3b9eedcb),
	.w6(32'h3c76374d),
	.w7(32'h3c41d6da),
	.w8(32'h3c5e89c9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd81045),
	.w1(32'h3bb99676),
	.w2(32'h3bf098a6),
	.w3(32'hba7e514e),
	.w4(32'hba2193c8),
	.w5(32'h3c25ae12),
	.w6(32'h3c681e10),
	.w7(32'h3c6dd2f3),
	.w8(32'h3cbeb1e9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c106c39),
	.w1(32'h3ab8c0a3),
	.w2(32'h3b3add76),
	.w3(32'hb991595c),
	.w4(32'hbb851c1e),
	.w5(32'h3b96e79a),
	.w6(32'h3c2cab21),
	.w7(32'h3c164c2e),
	.w8(32'h3c4a44ca),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4227b),
	.w1(32'h3c2c7441),
	.w2(32'h3c1f88c6),
	.w3(32'hbb24f61c),
	.w4(32'h3b8b3a6f),
	.w5(32'h3b0e4003),
	.w6(32'hbb7f1780),
	.w7(32'h3bbe29ee),
	.w8(32'h3b2652e6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa53d0e),
	.w1(32'hba4ea935),
	.w2(32'hba90ce55),
	.w3(32'h3b1538de),
	.w4(32'h3b908614),
	.w5(32'h3a7e404b),
	.w6(32'hba6c9155),
	.w7(32'h39ff039b),
	.w8(32'h3ab4779d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b940750),
	.w1(32'h3b905e1d),
	.w2(32'h3b20c7e3),
	.w3(32'hb9d32468),
	.w4(32'hb9c67d9a),
	.w5(32'h3c15b4bc),
	.w6(32'h3a995ee1),
	.w7(32'hb9432a92),
	.w8(32'h3b8008d9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba524363),
	.w1(32'h3c1d40ef),
	.w2(32'h3c7789e9),
	.w3(32'h3b2c01d5),
	.w4(32'h3bb84bd8),
	.w5(32'h3bcf6fc0),
	.w6(32'h3bdaa91d),
	.w7(32'hbb955385),
	.w8(32'hbb1cf18d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2a7db),
	.w1(32'h3b9d8902),
	.w2(32'h3be6cb9a),
	.w3(32'hbbe86f77),
	.w4(32'hbb8d6af6),
	.w5(32'hb9eae820),
	.w6(32'h3ab58cf4),
	.w7(32'h3be89081),
	.w8(32'h3c52e3c1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddf10c),
	.w1(32'h3b8d4fd4),
	.w2(32'h3c022ab1),
	.w3(32'h3a488b43),
	.w4(32'h3b0ecf5a),
	.w5(32'h3b4ee88c),
	.w6(32'h3b902c61),
	.w7(32'h3ba0ccc7),
	.w8(32'h3c1c3275),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1776ed),
	.w1(32'hbb0b86a0),
	.w2(32'h3966e084),
	.w3(32'h3bb89ac7),
	.w4(32'h39c7ad0d),
	.w5(32'h3b5d4461),
	.w6(32'h3bc460c9),
	.w7(32'h3b848a9f),
	.w8(32'h3bce729f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27e4e0),
	.w1(32'h3bc22f44),
	.w2(32'h3bfbd304),
	.w3(32'h3c3a7383),
	.w4(32'h3adda17c),
	.w5(32'h3c3c06fc),
	.w6(32'h3c5f72ca),
	.w7(32'h3bf9273a),
	.w8(32'h3c924e3b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bfa7e),
	.w1(32'hba047fc6),
	.w2(32'h3b193cfb),
	.w3(32'h39fdba78),
	.w4(32'h3a9f4654),
	.w5(32'hbab63ba2),
	.w6(32'hba83594f),
	.w7(32'h3a93fe6d),
	.w8(32'hba956612),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88e4137),
	.w1(32'h3aacb561),
	.w2(32'h38449c2e),
	.w3(32'h3adf5c59),
	.w4(32'h3b5e1b03),
	.w5(32'hba8a7c29),
	.w6(32'hbb63abd4),
	.w7(32'hba2f3ff9),
	.w8(32'hbad6885d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0943),
	.w1(32'hbb74a22f),
	.w2(32'hbb529233),
	.w3(32'hbbc03447),
	.w4(32'hbb4f0524),
	.w5(32'hbb0b01e2),
	.w6(32'hbb1dba87),
	.w7(32'hbad9070e),
	.w8(32'h3afab309),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed3d02),
	.w1(32'h3b1d8e99),
	.w2(32'hbb0628b4),
	.w3(32'h3ac2bdcf),
	.w4(32'hbb01e1ca),
	.w5(32'hbb7ca240),
	.w6(32'h3a25afcc),
	.w7(32'hbad2515c),
	.w8(32'hbbbd7620),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb045e27),
	.w1(32'h3a96a418),
	.w2(32'h3ba0baa0),
	.w3(32'hbba7dedc),
	.w4(32'hba9fcf1f),
	.w5(32'h3b93f00d),
	.w6(32'hbb955129),
	.w7(32'hbb1c6fe5),
	.w8(32'hb881efdf),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaa03d),
	.w1(32'h3bf03e35),
	.w2(32'h3ba8c225),
	.w3(32'h3a2d74e3),
	.w4(32'hba15655a),
	.w5(32'h3a82ed5a),
	.w6(32'h3c53cdfc),
	.w7(32'h3c1f73b7),
	.w8(32'h3c1c96b8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300b66),
	.w1(32'hbb4cde22),
	.w2(32'h3a3857d6),
	.w3(32'hbb3403ac),
	.w4(32'hbc1a7585),
	.w5(32'h3b1242de),
	.w6(32'h38066233),
	.w7(32'hbb15b618),
	.w8(32'h3b702034),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88dd71),
	.w1(32'hbacccd91),
	.w2(32'hbbb6b650),
	.w3(32'hbab61596),
	.w4(32'hbb608b04),
	.w5(32'hbaf22232),
	.w6(32'hbbf8242f),
	.w7(32'hbc00fb33),
	.w8(32'hbaedbbb4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48e3db),
	.w1(32'h3c784842),
	.w2(32'h3ca86a9d),
	.w3(32'hbbe66d61),
	.w4(32'h38380cd0),
	.w5(32'h3be80094),
	.w6(32'h3b82025c),
	.w7(32'h3bf15eec),
	.w8(32'h3c45d38d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc523),
	.w1(32'h3c27d7fa),
	.w2(32'h3b523e6f),
	.w3(32'h3c4f6097),
	.w4(32'h3b70e205),
	.w5(32'hbabb32f6),
	.w6(32'h3b368e0e),
	.w7(32'h3ab34362),
	.w8(32'h3b6e37ab),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5de8ce),
	.w1(32'h3ae679ac),
	.w2(32'h3b0499a3),
	.w3(32'hbbf8011e),
	.w4(32'hbb48eab2),
	.w5(32'hba5e7326),
	.w6(32'hbae3930c),
	.w7(32'hbbd368f6),
	.w8(32'h39a5d539),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6171d),
	.w1(32'h3a551516),
	.w2(32'h3ba76a82),
	.w3(32'hbb2f119c),
	.w4(32'h3b4f40b8),
	.w5(32'hbbefe111),
	.w6(32'h3a20e88e),
	.w7(32'h3b8de1c0),
	.w8(32'hbb4c4176),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43849b),
	.w1(32'hbac9031a),
	.w2(32'hbbdc1c77),
	.w3(32'hbc03ef56),
	.w4(32'hbbf6c606),
	.w5(32'hba91f493),
	.w6(32'hbbdd46b7),
	.w7(32'hbba49bf5),
	.w8(32'hbb2101f4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8e822),
	.w1(32'h3afc41ed),
	.w2(32'h39f98d7b),
	.w3(32'hb9eff6bc),
	.w4(32'hbadd3ce0),
	.w5(32'h3af4123d),
	.w6(32'h3ac6c6f9),
	.w7(32'h3ac64115),
	.w8(32'hb88fe9d8),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849406),
	.w1(32'h3b68eabb),
	.w2(32'h3a7d5eee),
	.w3(32'h3b28dda1),
	.w4(32'hba0c8415),
	.w5(32'hbb741c32),
	.w6(32'h3aa1cb50),
	.w7(32'hb9c0839e),
	.w8(32'hbba0a417),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4c28f),
	.w1(32'hbb949f2b),
	.w2(32'hbb0323b7),
	.w3(32'hbba93b28),
	.w4(32'hbb5adcd5),
	.w5(32'h3a1d72eb),
	.w6(32'hbb952272),
	.w7(32'hbb7bdd5b),
	.w8(32'hbad9937a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb357c45),
	.w1(32'hbbc56dde),
	.w2(32'hba99db11),
	.w3(32'h3acaad38),
	.w4(32'hba93a89f),
	.w5(32'h3b794f87),
	.w6(32'h3bed409c),
	.w7(32'h3aa6f598),
	.w8(32'h3afcefff),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f2d82),
	.w1(32'h3cb43a39),
	.w2(32'h3ca263d0),
	.w3(32'h3b8e797c),
	.w4(32'h3bef1f1a),
	.w5(32'hbb7afe54),
	.w6(32'h3b191501),
	.w7(32'h3c747994),
	.w8(32'h3c381442),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ab38a),
	.w1(32'hbb52b449),
	.w2(32'h3b84a45d),
	.w3(32'hbc225683),
	.w4(32'hbbc91f39),
	.w5(32'h3a6d75af),
	.w6(32'hbbb81aa9),
	.w7(32'hbabf35f2),
	.w8(32'h3bd8b6bf),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4682ee),
	.w1(32'h3c2343a0),
	.w2(32'h3c214d40),
	.w3(32'hbbb57e21),
	.w4(32'hbb0a72a5),
	.w5(32'hba9c55f0),
	.w6(32'hbbb107ce),
	.w7(32'h3b2fa985),
	.w8(32'h3860272c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0232c),
	.w1(32'h3b9e649d),
	.w2(32'h3b10c345),
	.w3(32'h3bc9bd1c),
	.w4(32'h3b69b191),
	.w5(32'hba0a5fcc),
	.w6(32'h3bf470aa),
	.w7(32'h3c1f09f1),
	.w8(32'hb9d0794b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c904d),
	.w1(32'h3b05c94f),
	.w2(32'hb7dce98e),
	.w3(32'hbad13ad7),
	.w4(32'hba0c10c6),
	.w5(32'hbb1026a2),
	.w6(32'hbc0ee049),
	.w7(32'hba9b4684),
	.w8(32'hbb07eed1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49c054),
	.w1(32'hb99cf70c),
	.w2(32'hbb1b182d),
	.w3(32'hbabb389e),
	.w4(32'hba56563f),
	.w5(32'hbb65aa08),
	.w6(32'hba310a48),
	.w7(32'hbaaa7e21),
	.w8(32'hba12d118),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac95b5e),
	.w1(32'h3a010d83),
	.w2(32'h3a5244c3),
	.w3(32'hbc2dd9e3),
	.w4(32'hbb495b40),
	.w5(32'hbb089cd6),
	.w6(32'hbb2fe666),
	.w7(32'hbc1cfa7f),
	.w8(32'hbb67d250),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21a832),
	.w1(32'h3bc5e149),
	.w2(32'h3c2a7819),
	.w3(32'hbb3d560e),
	.w4(32'hbb0c7aac),
	.w5(32'h3bcaf532),
	.w6(32'h3b5d66af),
	.w7(32'h3ba336cc),
	.w8(32'h3bf40970),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5b513),
	.w1(32'h3aec489a),
	.w2(32'h3a2dacee),
	.w3(32'h3b8ebee0),
	.w4(32'h3a52f799),
	.w5(32'h3b13d637),
	.w6(32'hbb9cf62f),
	.w7(32'hbbac4faf),
	.w8(32'h3b1b909b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd8867),
	.w1(32'h3bb451bf),
	.w2(32'h3b9f173a),
	.w3(32'h3b18d384),
	.w4(32'hb9cd2191),
	.w5(32'h3a955d39),
	.w6(32'hbb944e10),
	.w7(32'hb9dc3dfc),
	.w8(32'hbb08a4aa),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadcd3b),
	.w1(32'h3b02cfac),
	.w2(32'h3ba28b14),
	.w3(32'h3b016b30),
	.w4(32'hbb588606),
	.w5(32'h3baf1819),
	.w6(32'hbb4f2ced),
	.w7(32'h3a42b162),
	.w8(32'h3ae01bd0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cdc90),
	.w1(32'hba9f4353),
	.w2(32'h3ad98b17),
	.w3(32'h39e70335),
	.w4(32'h39a114a9),
	.w5(32'hbb5f66d6),
	.w6(32'h3b1b7300),
	.w7(32'h3b9ac947),
	.w8(32'hbb74f00a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03fabe),
	.w1(32'h3b32685c),
	.w2(32'h3b78c0d6),
	.w3(32'hbbf97b4c),
	.w4(32'hbc36d582),
	.w5(32'hb9c43723),
	.w6(32'hbb120c69),
	.w7(32'hbb472d08),
	.w8(32'h3b4f48ab),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf76547),
	.w1(32'h3b271df8),
	.w2(32'h3b5c68c3),
	.w3(32'hba7c2356),
	.w4(32'h3ace5dbf),
	.w5(32'h3b22c87c),
	.w6(32'h38723872),
	.w7(32'h3ab26c62),
	.w8(32'h3a8b3077),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94f882),
	.w1(32'h3c8e649c),
	.w2(32'h3ca6336a),
	.w3(32'h3c2644cc),
	.w4(32'hb9f3621c),
	.w5(32'hbb833ef0),
	.w6(32'h3bdf9e0e),
	.w7(32'hbac429b5),
	.w8(32'h3bd0aadb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7b68e),
	.w1(32'h3b2ac1ba),
	.w2(32'h3b220cf3),
	.w3(32'hbae08603),
	.w4(32'hba950fc1),
	.w5(32'h3b3500fe),
	.w6(32'h3af45790),
	.w7(32'h39b64d28),
	.w8(32'h3ad40535),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb980283),
	.w1(32'hbc041994),
	.w2(32'hbc08fa10),
	.w3(32'hbb040cd0),
	.w4(32'hbbc1015f),
	.w5(32'hbbd70399),
	.w6(32'h3c5c6799),
	.w7(32'h3c158333),
	.w8(32'h3bb086be),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule