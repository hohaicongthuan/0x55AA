module layer_8_featuremap_227(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad2bd2),
	.w1(32'hba5f7b02),
	.w2(32'h3ccc88c8),
	.w3(32'h3b9aebe8),
	.w4(32'hba311237),
	.w5(32'h3baa7bee),
	.w6(32'h3c88eecd),
	.w7(32'h3cf41849),
	.w8(32'hbc355697),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed4502),
	.w1(32'hbbe7fa72),
	.w2(32'hbbd63c1f),
	.w3(32'h3b9636ff),
	.w4(32'hbb9a4b6c),
	.w5(32'hbbaec679),
	.w6(32'hbb29cc4f),
	.w7(32'hbc11bf26),
	.w8(32'hbbcaad04),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65b11c),
	.w1(32'hbc16123a),
	.w2(32'hbb03370c),
	.w3(32'hbc3d7a0b),
	.w4(32'hbc012306),
	.w5(32'hbb8d4ad8),
	.w6(32'hbc24f9ab),
	.w7(32'hbc07f517),
	.w8(32'hbc588a56),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63f36b),
	.w1(32'h3b840089),
	.w2(32'h3b0ad4b4),
	.w3(32'hbba283b7),
	.w4(32'h3c22ff0a),
	.w5(32'h3c22a13b),
	.w6(32'h3c8e6555),
	.w7(32'h3b655941),
	.w8(32'hba9c9e4c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc575829),
	.w1(32'hbbb1b965),
	.w2(32'hbb564a18),
	.w3(32'hbc949f34),
	.w4(32'hbb2ad14b),
	.w5(32'h3acb33f7),
	.w6(32'hb97a6b26),
	.w7(32'hbb851a43),
	.w8(32'hbc0cf2d1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad57f04),
	.w1(32'h3b8985d3),
	.w2(32'hbaf49819),
	.w3(32'hbc0c74f1),
	.w4(32'hbb97d166),
	.w5(32'hbc078858),
	.w6(32'hbc8008de),
	.w7(32'hbc8a7d9e),
	.w8(32'h39472149),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dc917),
	.w1(32'h3b264809),
	.w2(32'h3b41e379),
	.w3(32'hbc3a15f5),
	.w4(32'h3ade3f85),
	.w5(32'h3b7b512c),
	.w6(32'hba00c0db),
	.w7(32'h3abaf6c2),
	.w8(32'h3a630898),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba9f93),
	.w1(32'hbc0bcb55),
	.w2(32'hbc252c4d),
	.w3(32'hbb747c5c),
	.w4(32'hbbd5b61b),
	.w5(32'hbc9ddcf8),
	.w6(32'hbbc88d98),
	.w7(32'hbceda88f),
	.w8(32'hbc85fa26),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a22fa),
	.w1(32'hba9e3bda),
	.w2(32'hbc286fab),
	.w3(32'h39c166bd),
	.w4(32'hba726328),
	.w5(32'hbbff6075),
	.w6(32'h3b3670a7),
	.w7(32'hbc490d5b),
	.w8(32'hbc2e20ba),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc14e78),
	.w1(32'hba8d8b2c),
	.w2(32'h3b9ae451),
	.w3(32'hb8fb5114),
	.w4(32'hbbf17ae5),
	.w5(32'hba5bc43f),
	.w6(32'h3b907a96),
	.w7(32'h3be234c1),
	.w8(32'hbc8ab85f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0c4dd),
	.w1(32'h3bbc1d40),
	.w2(32'hbbfb4d4e),
	.w3(32'h3b8646cc),
	.w4(32'h3ba1c9c4),
	.w5(32'hbc099370),
	.w6(32'h3c97d175),
	.w7(32'h3bcd5ff4),
	.w8(32'hba1a90d0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c439790),
	.w1(32'hbb2d6e22),
	.w2(32'h3bc88e91),
	.w3(32'h3c832792),
	.w4(32'h3c0f4bfe),
	.w5(32'h3c1102fe),
	.w6(32'h3a36cd83),
	.w7(32'h3b1bf3e4),
	.w8(32'h3cbac33d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac8c27),
	.w1(32'h3aa6edf5),
	.w2(32'h395ffd85),
	.w3(32'h3d015650),
	.w4(32'hbc4b2274),
	.w5(32'hbbe4127c),
	.w6(32'hbb8b903c),
	.w7(32'h3b2d16d0),
	.w8(32'hbbaf19dd),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c071981),
	.w1(32'h3c1b22ed),
	.w2(32'h3c6d7374),
	.w3(32'h3b962d8b),
	.w4(32'h3c34ec46),
	.w5(32'h3ca6d26b),
	.w6(32'h3c74d881),
	.w7(32'h3b973879),
	.w8(32'hbaaf3eb5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34aabd),
	.w1(32'h3bcd3c51),
	.w2(32'hba55b517),
	.w3(32'hbbf668fd),
	.w4(32'h3b8b6685),
	.w5(32'hba38f5e6),
	.w6(32'h3b2d2bf6),
	.w7(32'hbaec690b),
	.w8(32'hbb1ce0f5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12d266),
	.w1(32'h3be05463),
	.w2(32'h3cf439f8),
	.w3(32'hbb335452),
	.w4(32'h3adbf284),
	.w5(32'h3cb1f45b),
	.w6(32'h3c04f411),
	.w7(32'h3cd62c0b),
	.w8(32'hbb07276d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74841b),
	.w1(32'h3bf793fa),
	.w2(32'h3b4e989a),
	.w3(32'h3cfb7f81),
	.w4(32'hb9fc1d12),
	.w5(32'h3b9f480f),
	.w6(32'h3c295ebb),
	.w7(32'h3c19d621),
	.w8(32'hbaa4eb93),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a2352),
	.w1(32'h3a40edf8),
	.w2(32'h3b23e576),
	.w3(32'hbc6ec955),
	.w4(32'hbb077edb),
	.w5(32'hbc262638),
	.w6(32'h3bd7eca4),
	.w7(32'hbb674333),
	.w8(32'h3bcc79bc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a126d),
	.w1(32'hbc218db0),
	.w2(32'hbbb71fcd),
	.w3(32'h3cf6c54b),
	.w4(32'h3a95e2e6),
	.w5(32'hbc0ca7a5),
	.w6(32'h3cddd0d0),
	.w7(32'hba9c2003),
	.w8(32'hbc2cab95),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39e1ea),
	.w1(32'h3c825aa9),
	.w2(32'h3c16c7cd),
	.w3(32'h3bab826c),
	.w4(32'h3bcb1725),
	.w5(32'h3bf9ab9c),
	.w6(32'h3c1b030b),
	.w7(32'h3bbab651),
	.w8(32'h3c452190),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5af4d7),
	.w1(32'hba4d0d6e),
	.w2(32'h3a8d726f),
	.w3(32'h3aa0b8ab),
	.w4(32'hba287e78),
	.w5(32'h3bd17c04),
	.w6(32'h3b3aebe9),
	.w7(32'h3c3cef8c),
	.w8(32'h3bae5103),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc625996),
	.w1(32'h3b08205c),
	.w2(32'h3c2be6b3),
	.w3(32'hbc5840fb),
	.w4(32'h3a6e01e5),
	.w5(32'h3980ed87),
	.w6(32'hbb86f93c),
	.w7(32'hbb6d5662),
	.w8(32'hbd04a2bd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0cbcd),
	.w1(32'h3aaedb2b),
	.w2(32'h3bfcf564),
	.w3(32'hba77e350),
	.w4(32'h3b31be7a),
	.w5(32'hbbb964b1),
	.w6(32'h3d1a6a80),
	.w7(32'h3ca4e3ff),
	.w8(32'hbc572239),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4319ba),
	.w1(32'h3be6f360),
	.w2(32'h3b0735a9),
	.w3(32'hbc7ec0ef),
	.w4(32'hb97994e6),
	.w5(32'hbb2d262b),
	.w6(32'h3ae69518),
	.w7(32'h3ae8377b),
	.w8(32'hbccef680),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd49a4),
	.w1(32'h3bff9fd8),
	.w2(32'hbc00c2e5),
	.w3(32'hbc962de3),
	.w4(32'h3b2deacb),
	.w5(32'hbbd03d20),
	.w6(32'h3b4ba63f),
	.w7(32'hbc0c7ebd),
	.w8(32'hbc80ae61),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d1ddd),
	.w1(32'h3a05d668),
	.w2(32'h3c0652f7),
	.w3(32'hbc615ac9),
	.w4(32'hbb54cb73),
	.w5(32'h3c239770),
	.w6(32'h3c9610a3),
	.w7(32'h3c6bbb23),
	.w8(32'hbcb77e49),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20c860),
	.w1(32'hbb6b6186),
	.w2(32'h3b330610),
	.w3(32'h3ad4f11a),
	.w4(32'h3ad43e81),
	.w5(32'h3ad5a8f1),
	.w6(32'hbb80754a),
	.w7(32'h3b8e9471),
	.w8(32'hbbc42a29),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4cee1c),
	.w1(32'hbd91b15e),
	.w2(32'h3c8921bf),
	.w3(32'h3cf8d841),
	.w4(32'hbcd97caf),
	.w5(32'hbba7cf65),
	.w6(32'h37859134),
	.w7(32'h3d6dab38),
	.w8(32'hbc9e567b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10647d),
	.w1(32'h3c1780a0),
	.w2(32'h39bc4595),
	.w3(32'h3c36d942),
	.w4(32'h3c727fdf),
	.w5(32'hbb8a87b7),
	.w6(32'h3c5ae4d0),
	.w7(32'h3c05ac92),
	.w8(32'hbba246ef),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05d37d),
	.w1(32'hbb18bf6a),
	.w2(32'hbb9bd2d6),
	.w3(32'hbbeada41),
	.w4(32'hbc3418ae),
	.w5(32'hbc76a5b9),
	.w6(32'hbb3c46a1),
	.w7(32'hbbf318e7),
	.w8(32'h3c94fe7b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6bdf2),
	.w1(32'h3c33fc9f),
	.w2(32'hba94b6d6),
	.w3(32'h3ca67fde),
	.w4(32'h3c0fca6a),
	.w5(32'h3852daeb),
	.w6(32'h3c326a85),
	.w7(32'h3ac34bcf),
	.w8(32'hbc043de5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dd661),
	.w1(32'h3c14b2e8),
	.w2(32'hbb821ce7),
	.w3(32'hbc14c38c),
	.w4(32'h3ae7dab9),
	.w5(32'hbab73aa8),
	.w6(32'h3b443b52),
	.w7(32'hbb750c19),
	.w8(32'h3a81451a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2e7f0),
	.w1(32'h3b89f083),
	.w2(32'hbc139513),
	.w3(32'hbb553ac0),
	.w4(32'h3add1ebe),
	.w5(32'h3aaba5e3),
	.w6(32'hbb8ca55d),
	.w7(32'hbab9899e),
	.w8(32'h3b9bb607),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a26be),
	.w1(32'h3b38ab1c),
	.w2(32'hbaa44252),
	.w3(32'h3b3e31a5),
	.w4(32'hb725795c),
	.w5(32'hb917c16a),
	.w6(32'hbb4851c1),
	.w7(32'hba1dbc7b),
	.w8(32'hbaba7baf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2894),
	.w1(32'h3c08bcf8),
	.w2(32'h3b987cee),
	.w3(32'hbc8ace6e),
	.w4(32'hbb5b3457),
	.w5(32'hbbad949a),
	.w6(32'hbb921216),
	.w7(32'hbb2a4adf),
	.w8(32'hbc05224d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbada8f4),
	.w1(32'hbc854c6e),
	.w2(32'hbc2b66f7),
	.w3(32'h3b70847e),
	.w4(32'hbb78b82e),
	.w5(32'hbb3839f9),
	.w6(32'h3bf2b105),
	.w7(32'h3b2a4851),
	.w8(32'hbb6b88d0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99145c7),
	.w1(32'h391befbf),
	.w2(32'h3b8b4461),
	.w3(32'hbb45bd19),
	.w4(32'h3ba9c6c6),
	.w5(32'h3bf6621e),
	.w6(32'h398fe3f9),
	.w7(32'h3bb0d4c8),
	.w8(32'h3b8029e9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c807),
	.w1(32'h3bb51f35),
	.w2(32'hbb93e48e),
	.w3(32'hbb570f35),
	.w4(32'h3b9167a3),
	.w5(32'hbb65d6fc),
	.w6(32'h3bd44e5c),
	.w7(32'hbb06ee55),
	.w8(32'hbbdd14ec),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e864d),
	.w1(32'h3b80d12d),
	.w2(32'hbb39db84),
	.w3(32'hbc2445a5),
	.w4(32'h39327687),
	.w5(32'h38077a83),
	.w6(32'h3b24f310),
	.w7(32'hbc005e6c),
	.w8(32'hbbdc5940),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebb46c),
	.w1(32'hbad43134),
	.w2(32'h3b87e9df),
	.w3(32'h3bc46c5f),
	.w4(32'h3a5fa137),
	.w5(32'h3bb6555d),
	.w6(32'hb9ff5011),
	.w7(32'hb9917121),
	.w8(32'hbc7f1f14),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffe958),
	.w1(32'h3a2bf6b0),
	.w2(32'h3af04b8f),
	.w3(32'h3c0b117d),
	.w4(32'h3a264b9b),
	.w5(32'hbc1bbb33),
	.w6(32'h3c8ccecc),
	.w7(32'h38f0b7a7),
	.w8(32'hbc423140),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c16dc),
	.w1(32'hbbd61f23),
	.w2(32'h3c151448),
	.w3(32'hbc288edf),
	.w4(32'hbbf48c2f),
	.w5(32'h3be66796),
	.w6(32'hbb001d32),
	.w7(32'h399fe602),
	.w8(32'hbacd5fa4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09033b),
	.w1(32'hbb8e2501),
	.w2(32'hbc0d3190),
	.w3(32'h3b079b46),
	.w4(32'hbb5d0d0e),
	.w5(32'hbb8c7664),
	.w6(32'hbbfd034e),
	.w7(32'hbab0fbd8),
	.w8(32'h3c3cad93),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c286879),
	.w1(32'h3b6dc89b),
	.w2(32'h3b70fad3),
	.w3(32'h3bce7332),
	.w4(32'hbbb5c83e),
	.w5(32'hbc3e1a1d),
	.w6(32'h3c76e7f5),
	.w7(32'h3adc52a8),
	.w8(32'h3cad6dc3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce38678),
	.w1(32'hbbe6fbc1),
	.w2(32'h3bb0892d),
	.w3(32'h3ce2ae3d),
	.w4(32'h3990abfb),
	.w5(32'h3c1dc782),
	.w6(32'h3c3528d1),
	.w7(32'h3bf17402),
	.w8(32'hbd34f2ed),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd47adae),
	.w1(32'h3baaf181),
	.w2(32'hbb8cf3f0),
	.w3(32'hbd00cd9e),
	.w4(32'h3b0c8a0a),
	.w5(32'hbbf4bfda),
	.w6(32'h3ae34a0b),
	.w7(32'hbbe5fe4f),
	.w8(32'hbc3ec87e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12f0ed),
	.w1(32'hbbf7a21a),
	.w2(32'h3b5fecdb),
	.w3(32'hbc0fc8d4),
	.w4(32'hbb5e50d6),
	.w5(32'h3b94e1ac),
	.w6(32'hbb984850),
	.w7(32'hbae00de4),
	.w8(32'hbb162fbc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04be4e),
	.w1(32'hbb7a7c36),
	.w2(32'h3c79453f),
	.w3(32'hbaa3c328),
	.w4(32'h3a7e9e31),
	.w5(32'h3c437ea0),
	.w6(32'h3c04705a),
	.w7(32'h3cb8a110),
	.w8(32'hbc24e1da),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80af53),
	.w1(32'h3b39b365),
	.w2(32'h3c8c5c70),
	.w3(32'hbb8f11c4),
	.w4(32'hb9a1e60d),
	.w5(32'h3bb13b63),
	.w6(32'h3b0bb9e6),
	.w7(32'h3c346e9c),
	.w8(32'hbc353a0f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe427f9),
	.w1(32'h3be4728f),
	.w2(32'h3b9a5ea6),
	.w3(32'hb9a0ca0f),
	.w4(32'h3c1b90ad),
	.w5(32'hbbe1bdab),
	.w6(32'h3c850b3c),
	.w7(32'h3bd51329),
	.w8(32'hb98ccace),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f596b),
	.w1(32'hbb19f2ad),
	.w2(32'h3b0b1737),
	.w3(32'h3b8031cb),
	.w4(32'h3a865ba9),
	.w5(32'h3baffd29),
	.w6(32'hbc18238c),
	.w7(32'hbb52c481),
	.w8(32'h3bc628f2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ad73c),
	.w1(32'h3bfe58bd),
	.w2(32'h3c172b12),
	.w3(32'hbacc7f0c),
	.w4(32'hbb70c4e8),
	.w5(32'hbbfaaec4),
	.w6(32'h3c6128f1),
	.w7(32'hbc1f3364),
	.w8(32'hbc375a01),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b670b37),
	.w1(32'h3c49066f),
	.w2(32'h3ba41fda),
	.w3(32'hb9767c3d),
	.w4(32'h3c2a835c),
	.w5(32'h3bda9dab),
	.w6(32'h3c25bf3e),
	.w7(32'h3b378fef),
	.w8(32'hba9d65e1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18b47c),
	.w1(32'hb9e7989b),
	.w2(32'h3c43e48a),
	.w3(32'hb9bfe645),
	.w4(32'hbb0564dc),
	.w5(32'h3a91f872),
	.w6(32'hbb8bd001),
	.w7(32'hb9175d17),
	.w8(32'h3cceff10),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce29f22),
	.w1(32'h3ba27f65),
	.w2(32'hbc02462a),
	.w3(32'h3c800d90),
	.w4(32'hb963f468),
	.w5(32'hbba5cff3),
	.w6(32'h3bc6d05b),
	.w7(32'hbba8c6b3),
	.w8(32'h3b6e23de),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b56b7),
	.w1(32'hbc048962),
	.w2(32'h3bd4f73f),
	.w3(32'h3be7a0a5),
	.w4(32'hba1466b3),
	.w5(32'hbc4a9fe5),
	.w6(32'h3c142eb9),
	.w7(32'h3c8e3667),
	.w8(32'hbbb0cecd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b4166),
	.w1(32'h3c1fc065),
	.w2(32'hbc02aad7),
	.w3(32'hbb21c6f2),
	.w4(32'hbad21304),
	.w5(32'hbb1319ab),
	.w6(32'h3bbc577c),
	.w7(32'hbaed55af),
	.w8(32'h3b50ae7e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42ce2f),
	.w1(32'hbbca1ebc),
	.w2(32'hbc4cea94),
	.w3(32'hbb0984d4),
	.w4(32'hbbec5084),
	.w5(32'hbc838cd8),
	.w6(32'hbabfb79f),
	.w7(32'hbc9d9290),
	.w8(32'hbc5fc5b3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817068),
	.w1(32'hbbe340d1),
	.w2(32'hbb4f00d8),
	.w3(32'hbb2f1f6f),
	.w4(32'hbaf34148),
	.w5(32'hbb1c5705),
	.w6(32'h3a9a2f3c),
	.w7(32'h3b1e4eda),
	.w8(32'hbab65bb6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1320d8),
	.w1(32'h3c8f22cc),
	.w2(32'h3c3c9593),
	.w3(32'h3c2f670a),
	.w4(32'h3c97be7d),
	.w5(32'h3c32313e),
	.w6(32'h3ca2e647),
	.w7(32'h3c49b0bf),
	.w8(32'hbc98c297),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0131df),
	.w1(32'hbbaeb018),
	.w2(32'hbb6d2ac8),
	.w3(32'hbc91a284),
	.w4(32'hbb69d301),
	.w5(32'hbb58c854),
	.w6(32'hbb87f7ba),
	.w7(32'hbbece65b),
	.w8(32'hbc341cff),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7a606),
	.w1(32'h3c208732),
	.w2(32'h3b6a8071),
	.w3(32'h3aecd98c),
	.w4(32'h3c083cb3),
	.w5(32'h3b047fa0),
	.w6(32'h3c09dc72),
	.w7(32'h3b82e497),
	.w8(32'h3917636b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2e246),
	.w1(32'h3ca70a36),
	.w2(32'h3b1d4cff),
	.w3(32'h3c42ccee),
	.w4(32'h3c9d2cac),
	.w5(32'hbc277a85),
	.w6(32'h3cb12f02),
	.w7(32'h3ac57824),
	.w8(32'hb9d879f3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b963b10),
	.w1(32'hbc680e67),
	.w2(32'hbc5d4c69),
	.w3(32'hbbb0ebf6),
	.w4(32'hbc139f6b),
	.w5(32'hbc03496a),
	.w6(32'hbc64fd39),
	.w7(32'hbc717d55),
	.w8(32'h3c4dc998),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c65c3),
	.w1(32'h3bfb92f7),
	.w2(32'hb9a9a6f8),
	.w3(32'h3cccf0f5),
	.w4(32'h3baeaa31),
	.w5(32'h389a4f3d),
	.w6(32'h3bbb5aff),
	.w7(32'hb9bbaef8),
	.w8(32'h3b397516),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb871d0a),
	.w1(32'hbbb15200),
	.w2(32'h39bc6e31),
	.w3(32'hbb25e75c),
	.w4(32'hbb43516d),
	.w5(32'hbb04e5d5),
	.w6(32'h39c73e6c),
	.w7(32'hbaede8bc),
	.w8(32'hbc61eab2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca00dc7),
	.w1(32'h3b195cc1),
	.w2(32'h3c123697),
	.w3(32'hbca82661),
	.w4(32'hb8fbe4e6),
	.w5(32'h3b8fcca2),
	.w6(32'h3b0899db),
	.w7(32'h3a66292c),
	.w8(32'hbbe58069),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc39836),
	.w1(32'h3ad6a2ce),
	.w2(32'h3c9612a9),
	.w3(32'hbc29a471),
	.w4(32'h3bea73ba),
	.w5(32'h3c4c05a3),
	.w6(32'h3acc42bc),
	.w7(32'h3c453bb2),
	.w8(32'hbbb26668),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7856b3),
	.w1(32'h3c463351),
	.w2(32'h3a91b188),
	.w3(32'h3916ce33),
	.w4(32'h3a0f6138),
	.w5(32'h3ba456e4),
	.w6(32'h3b89aef4),
	.w7(32'h3b48d99f),
	.w8(32'hbc090b9a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b2503),
	.w1(32'h3bc4e8db),
	.w2(32'h3cb4fd62),
	.w3(32'hbc84c181),
	.w4(32'h3c292cd2),
	.w5(32'h3cc48a2b),
	.w6(32'h3ce938f2),
	.w7(32'h3d1d87eb),
	.w8(32'hbca25c62),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99ab0f),
	.w1(32'h3c0d3985),
	.w2(32'hbb70bf34),
	.w3(32'hbc3ecf93),
	.w4(32'h3bfbab2a),
	.w5(32'hbba76067),
	.w6(32'h3b97339e),
	.w7(32'hbb8b2da8),
	.w8(32'hbc0b1750),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc679d30),
	.w1(32'hbc5a5003),
	.w2(32'hbb3cd813),
	.w3(32'hbc864673),
	.w4(32'hbb85d126),
	.w5(32'hb9e4842b),
	.w6(32'hb9b13f5c),
	.w7(32'hba5b33fe),
	.w8(32'hbb7fedcf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c538d),
	.w1(32'hbc17e7e0),
	.w2(32'hbc29a357),
	.w3(32'hbb804540),
	.w4(32'hbb273817),
	.w5(32'h3ab62e53),
	.w6(32'h3ae4e93b),
	.w7(32'hbc29524d),
	.w8(32'hbc440537),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc506b31),
	.w1(32'hbbf1ac6e),
	.w2(32'hbbb521ce),
	.w3(32'h3b7a6cbe),
	.w4(32'hbb8bad1c),
	.w5(32'hbbe1cf0c),
	.w6(32'h3b516287),
	.w7(32'hbaf63d6a),
	.w8(32'hbbac9d00),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef823d),
	.w1(32'h3b3d6a23),
	.w2(32'h39859b29),
	.w3(32'hbbacd09e),
	.w4(32'hbb3f4b22),
	.w5(32'hbb731aa8),
	.w6(32'h3a8ad832),
	.w7(32'h3ba01ec8),
	.w8(32'hbb989754),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba06871),
	.w1(32'h3c5478b3),
	.w2(32'hba4bd346),
	.w3(32'hbc0695aa),
	.w4(32'hbb49e6a7),
	.w5(32'hbb8d8c05),
	.w6(32'h3b0b0781),
	.w7(32'hbb4fb765),
	.w8(32'h3b312e2c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2a5f0),
	.w1(32'h3a9b65fd),
	.w2(32'hbbf5e33e),
	.w3(32'h3c40d882),
	.w4(32'h3a9fd44a),
	.w5(32'hbbec92d5),
	.w6(32'hbb4d3226),
	.w7(32'hbbaae042),
	.w8(32'hba177aa6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c506f),
	.w1(32'hbb47bf77),
	.w2(32'h3b805bc0),
	.w3(32'h3c6676b4),
	.w4(32'h3b24a574),
	.w5(32'h3bb60dd8),
	.w6(32'h3c6d592e),
	.w7(32'h3c80d41d),
	.w8(32'h3b390245),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43ce08),
	.w1(32'h3c066328),
	.w2(32'hbac54312),
	.w3(32'h3c1bfddd),
	.w4(32'h3c124a86),
	.w5(32'h3b69cab8),
	.w6(32'h370dbae4),
	.w7(32'hbb60e1b4),
	.w8(32'hbbc9f32b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54be71),
	.w1(32'h3ab45552),
	.w2(32'h3bec0f6b),
	.w3(32'hbc2beab2),
	.w4(32'h3b127f2b),
	.w5(32'h3b046816),
	.w6(32'hbb31eefd),
	.w7(32'h3bc0e49f),
	.w8(32'hbab0efbf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f72df),
	.w1(32'h395db4a7),
	.w2(32'h398766ac),
	.w3(32'h3c546193),
	.w4(32'hbb59c7ab),
	.w5(32'h3b9052b8),
	.w6(32'h3b3580a9),
	.w7(32'h3b5831d3),
	.w8(32'hbc4edfe8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd51c94),
	.w1(32'h3bd9be82),
	.w2(32'h3c4fca27),
	.w3(32'hbc151731),
	.w4(32'hba2bffd4),
	.w5(32'h3c788fea),
	.w6(32'h3bb9a9d2),
	.w7(32'h3bd3dd22),
	.w8(32'h3bcf19f9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f055f),
	.w1(32'h3c3f8665),
	.w2(32'h3bb76348),
	.w3(32'h3b0c4e7e),
	.w4(32'h3ca46e48),
	.w5(32'h3b646bc7),
	.w6(32'h3cf7dd42),
	.w7(32'h3c393718),
	.w8(32'h3c095038),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05f373),
	.w1(32'h3ce3502d),
	.w2(32'h3cb11d44),
	.w3(32'h3d257a60),
	.w4(32'h3cb23833),
	.w5(32'h3c3bb024),
	.w6(32'h3cb61ba3),
	.w7(32'hbb126546),
	.w8(32'h3bff86c3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe283ca),
	.w1(32'h3c8abff8),
	.w2(32'h3c811672),
	.w3(32'h3b2e0ee3),
	.w4(32'h3c76d055),
	.w5(32'h3c752a17),
	.w6(32'h3d07d811),
	.w7(32'h3c225b18),
	.w8(32'hbb209b19),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6a9ac),
	.w1(32'h3c8399b1),
	.w2(32'h3cbb99ad),
	.w3(32'hb98024ff),
	.w4(32'h3bc52446),
	.w5(32'h3c3ddaa9),
	.w6(32'h3c820e32),
	.w7(32'h3cb33f2c),
	.w8(32'hba862468),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b020d),
	.w1(32'h3b8f74a5),
	.w2(32'h3b3e4ec6),
	.w3(32'hb9a1514e),
	.w4(32'h3ae44240),
	.w5(32'h3b9b7a98),
	.w6(32'h3b1bb33a),
	.w7(32'h3af68590),
	.w8(32'hbb824c8e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0d8df),
	.w1(32'h3bb1dbe9),
	.w2(32'hbb3222be),
	.w3(32'hb7a39afe),
	.w4(32'h3c3332e7),
	.w5(32'hba89b9da),
	.w6(32'h3b528d36),
	.w7(32'hbb3cc5c6),
	.w8(32'hbaf6bb17),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a4197),
	.w1(32'hb8a1f826),
	.w2(32'hbaa08ce2),
	.w3(32'hbbfd72ce),
	.w4(32'hba890a6b),
	.w5(32'hbb79c193),
	.w6(32'h3ac6bd6e),
	.w7(32'h3b0274db),
	.w8(32'hbb9e0c42),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafdf33),
	.w1(32'hba90721f),
	.w2(32'h3b909fc8),
	.w3(32'hbb1e5b4b),
	.w4(32'hbacae87d),
	.w5(32'h3beaeaef),
	.w6(32'h3c3b73db),
	.w7(32'h3bef66ea),
	.w8(32'hbc908fa2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cd2ee),
	.w1(32'hbbb8dbc4),
	.w2(32'hbc00c281),
	.w3(32'hbc0829c8),
	.w4(32'hbc06f89d),
	.w5(32'hbb889cc6),
	.w6(32'hbbd459c5),
	.w7(32'hbb0102c0),
	.w8(32'hbc1241fb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcab1c2),
	.w1(32'h3b8f582f),
	.w2(32'h3b743aa3),
	.w3(32'hbb9a577e),
	.w4(32'h3a26083f),
	.w5(32'h3bd47902),
	.w6(32'hb92792bd),
	.w7(32'h3b976b59),
	.w8(32'h3b422fad),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10cebe),
	.w1(32'hb9835227),
	.w2(32'h3b067fbe),
	.w3(32'hbca19abb),
	.w4(32'hbae03c0a),
	.w5(32'h3b55a54c),
	.w6(32'h3a8bf753),
	.w7(32'hb9ea22e3),
	.w8(32'h3b7b27a8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72ae0d),
	.w1(32'hbbc3e313),
	.w2(32'hba84ed06),
	.w3(32'h3b2fbf6f),
	.w4(32'hbb9d2e58),
	.w5(32'hbb86b15a),
	.w6(32'hb8bda1c2),
	.w7(32'hbb57b14b),
	.w8(32'hbb6ce94f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad43b87),
	.w1(32'hbbcd1cdf),
	.w2(32'hbc6d0e52),
	.w3(32'hbb36717d),
	.w4(32'hbb953dae),
	.w5(32'hbc6efd23),
	.w6(32'hbbfe7d7b),
	.w7(32'hbc4a25d1),
	.w8(32'h3bdaccf3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa83f2e),
	.w1(32'h3b838937),
	.w2(32'h3c40f029),
	.w3(32'hbb0cf8b4),
	.w4(32'h3b8a5526),
	.w5(32'h3c0c0a5a),
	.w6(32'h3c0d680d),
	.w7(32'h3c431840),
	.w8(32'hbb48b060),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8026e3),
	.w1(32'h3cdca329),
	.w2(32'h3c9ff3e0),
	.w3(32'hbb02934f),
	.w4(32'h3bd59d75),
	.w5(32'h3c5e42e8),
	.w6(32'h3cbc2566),
	.w7(32'h3c3b20d0),
	.w8(32'h3b96de99),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12e559),
	.w1(32'h3b96ae84),
	.w2(32'hbbff586d),
	.w3(32'hbb816615),
	.w4(32'hbb33169e),
	.w5(32'hbba13a40),
	.w6(32'h3a784419),
	.w7(32'hbc127cef),
	.w8(32'hbb0dd27a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c144804),
	.w1(32'h3b3aa8ce),
	.w2(32'h3a731cdb),
	.w3(32'h3c63c257),
	.w4(32'hbb96b584),
	.w5(32'h3a8737d6),
	.w6(32'hbac7ffd7),
	.w7(32'hbbb38dbf),
	.w8(32'hbbbaccfa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd49e),
	.w1(32'h3b14ce2a),
	.w2(32'hbbe2df55),
	.w3(32'h3c1b00c3),
	.w4(32'h3c5ad0fc),
	.w5(32'hbc86482f),
	.w6(32'h3a487ab7),
	.w7(32'h3a9cacb9),
	.w8(32'h3b104c48),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb26bcc),
	.w1(32'h3c1010d4),
	.w2(32'hbbe6830c),
	.w3(32'hbbfe9b24),
	.w4(32'h3b246f6b),
	.w5(32'hbafd486c),
	.w6(32'h3c14e817),
	.w7(32'hbba330a6),
	.w8(32'h3cbab787),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35b6cb),
	.w1(32'hbc31309b),
	.w2(32'hbcd64de8),
	.w3(32'hbae41a58),
	.w4(32'hbc39b541),
	.w5(32'hbc554321),
	.w6(32'hbc46b907),
	.w7(32'hbc5d1f2d),
	.w8(32'hbc0fa2d6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b4c87),
	.w1(32'h3b069e17),
	.w2(32'h3c1fb174),
	.w3(32'hbc1c69b8),
	.w4(32'h3b1e0bdd),
	.w5(32'h3c98383a),
	.w6(32'hbb194d45),
	.w7(32'h3a32360b),
	.w8(32'h3b128499),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90e2dc),
	.w1(32'h3c8a537d),
	.w2(32'h3b74e237),
	.w3(32'hbc6861db),
	.w4(32'h3bb1e5f8),
	.w5(32'h3c2f20f6),
	.w6(32'h3c6ad46c),
	.w7(32'h397f97ad),
	.w8(32'hbb152ab7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc022ed7),
	.w1(32'hba9e7287),
	.w2(32'hbbd9bd10),
	.w3(32'h3ac8abb2),
	.w4(32'hbc022113),
	.w5(32'h3c319279),
	.w6(32'hbc35da1f),
	.w7(32'hbadba5f2),
	.w8(32'hbb942bc5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43718),
	.w1(32'h3c5bb5af),
	.w2(32'h3c34ec0d),
	.w3(32'h3cab2abb),
	.w4(32'h3c37b6e4),
	.w5(32'h3bc7a48b),
	.w6(32'h3c87c7ed),
	.w7(32'h3c08c797),
	.w8(32'hbb48e397),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf81d8a),
	.w1(32'h3be97dc1),
	.w2(32'h3b496fe6),
	.w3(32'hbb637676),
	.w4(32'h3bc9e848),
	.w5(32'h3b33f991),
	.w6(32'h3bc8689a),
	.w7(32'h3b79d409),
	.w8(32'hbc289117),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc907bb0),
	.w1(32'h3b740cf7),
	.w2(32'h3a6acd36),
	.w3(32'hbc808203),
	.w4(32'h3b3d92a9),
	.w5(32'h3c3f3bb1),
	.w6(32'hbb97cc54),
	.w7(32'h39b2b4ad),
	.w8(32'hba96e534),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41a0cc),
	.w1(32'h3b806330),
	.w2(32'h3b873032),
	.w3(32'hbb91f9c3),
	.w4(32'h3c0467f0),
	.w5(32'h3b7c8a94),
	.w6(32'h3b0b4cae),
	.w7(32'h3c057e24),
	.w8(32'h3bd845c3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12e02a),
	.w1(32'h3abe1a1b),
	.w2(32'hbacc20af),
	.w3(32'h3a81b69f),
	.w4(32'h3ac35330),
	.w5(32'hb8a705e6),
	.w6(32'h3bedb128),
	.w7(32'hbad439a8),
	.w8(32'hbab0327d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35ded7),
	.w1(32'h3c3ce8ec),
	.w2(32'h3c3263a6),
	.w3(32'hb8df70c1),
	.w4(32'h3bbb7c6e),
	.w5(32'h3c59ce83),
	.w6(32'h3b0f3f20),
	.w7(32'h3b00d50a),
	.w8(32'h3b09e476),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4341f),
	.w1(32'h3a92dc05),
	.w2(32'hba79eec6),
	.w3(32'hbb816598),
	.w4(32'hbb12852e),
	.w5(32'hbb9448eb),
	.w6(32'hbabb4096),
	.w7(32'hbbc36062),
	.w8(32'hbb30391c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a757a),
	.w1(32'h3c0172f9),
	.w2(32'hbc60de8e),
	.w3(32'hbbfe67b1),
	.w4(32'h3a1d9afb),
	.w5(32'hbc0def28),
	.w6(32'h39d505b0),
	.w7(32'hbc4e379c),
	.w8(32'hbac82a0d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a211cf7),
	.w1(32'h3c6bde6a),
	.w2(32'h3c5b631e),
	.w3(32'hbb3c3c0a),
	.w4(32'h3c249f89),
	.w5(32'h3b641733),
	.w6(32'h3c2e199b),
	.w7(32'h3c8fa724),
	.w8(32'hbb31b84f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2be860),
	.w1(32'h3aced5a7),
	.w2(32'hba641218),
	.w3(32'hbc1086a4),
	.w4(32'h3bdb80a9),
	.w5(32'h3bd2b252),
	.w6(32'h3b380c12),
	.w7(32'h3bb444a6),
	.w8(32'h3ac72ad1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8fb38),
	.w1(32'h3bb7355b),
	.w2(32'h3a1075be),
	.w3(32'h3b8b8aa9),
	.w4(32'h3bbbe56e),
	.w5(32'h3acf5641),
	.w6(32'h3bd32c06),
	.w7(32'h3b34bbea),
	.w8(32'h3b09e655),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b287302),
	.w1(32'h3b9795c2),
	.w2(32'h3c06c102),
	.w3(32'h3a2f244e),
	.w4(32'h378af55a),
	.w5(32'h3afd4cfc),
	.w6(32'h3a8b0573),
	.w7(32'h3aa60dde),
	.w8(32'h3c0fd93c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08276e),
	.w1(32'hbb5b9867),
	.w2(32'h3aff05fd),
	.w3(32'h3c21413c),
	.w4(32'h3a6cd8ee),
	.w5(32'hbb4b9e2c),
	.w6(32'h3bff5b15),
	.w7(32'h3a896c9e),
	.w8(32'h3b83b643),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9669c),
	.w1(32'hbb3bb18d),
	.w2(32'h3c0be5d5),
	.w3(32'hbb4a9ffc),
	.w4(32'h3b159596),
	.w5(32'h3b864438),
	.w6(32'h3bd9bea5),
	.w7(32'h3b621dfd),
	.w8(32'h3abf9794),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66eb09),
	.w1(32'h3a626479),
	.w2(32'h3b5e3c66),
	.w3(32'hbc40527a),
	.w4(32'hbb3bb4f2),
	.w5(32'hbb267901),
	.w6(32'hba5952ba),
	.w7(32'h3b45f813),
	.w8(32'h3b9bbd1c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28e3f8),
	.w1(32'h3c361acd),
	.w2(32'h3bf9b556),
	.w3(32'hba5e2a5b),
	.w4(32'h3b4b4bf2),
	.w5(32'hbacfa9e5),
	.w6(32'h3c40d2d5),
	.w7(32'h3baef7fe),
	.w8(32'h3b63cc82),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cd426),
	.w1(32'hbbe1a560),
	.w2(32'h3adcc542),
	.w3(32'hbcc7bc3f),
	.w4(32'hbbc07282),
	.w5(32'h3a4df3b1),
	.w6(32'hba90e538),
	.w7(32'hbbc5edf8),
	.w8(32'hbbbc2017),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53ce46),
	.w1(32'hbb0e2992),
	.w2(32'hbb616a36),
	.w3(32'hbb84e43f),
	.w4(32'h3af2a4fe),
	.w5(32'hbb2d5cf1),
	.w6(32'h3a2b9723),
	.w7(32'hbb8ab0fd),
	.w8(32'hbb02aee0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bd176),
	.w1(32'h3c016c04),
	.w2(32'h3a057db2),
	.w3(32'h3ac51e62),
	.w4(32'h3c32b69f),
	.w5(32'hbbca7e91),
	.w6(32'h3bc1be72),
	.w7(32'hbb6dfa1d),
	.w8(32'hbb4538a5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ffc56),
	.w1(32'h3bcfd489),
	.w2(32'h3c2b3dbb),
	.w3(32'hbbad5beb),
	.w4(32'h3bc64bde),
	.w5(32'h3c51ad9b),
	.w6(32'h3bc0c143),
	.w7(32'hbaed8611),
	.w8(32'hbc63ec78),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84fd8c),
	.w1(32'hbb9c6173),
	.w2(32'h3c888c14),
	.w3(32'hbc23a08c),
	.w4(32'h3be74896),
	.w5(32'h3c817aea),
	.w6(32'h3b88af84),
	.w7(32'h3c8ca706),
	.w8(32'hbb51368a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e1774),
	.w1(32'hba7d4aab),
	.w2(32'hbb4e5ea3),
	.w3(32'hbb139b2e),
	.w4(32'hbab470f5),
	.w5(32'hbb47a598),
	.w6(32'h3a8a43f2),
	.w7(32'hbb742d84),
	.w8(32'hba0be06b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafda213),
	.w1(32'h3b1233c1),
	.w2(32'hbacb2a0a),
	.w3(32'h39b1f3f3),
	.w4(32'h3b5377ff),
	.w5(32'h3ae07250),
	.w6(32'h3c7168d7),
	.w7(32'h3c536ae0),
	.w8(32'hbc1514c5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule