module layer_10_featuremap_255(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a01a),
	.w1(32'hbb9c5185),
	.w2(32'hbac8d33d),
	.w3(32'hbb6974ce),
	.w4(32'h3af54798),
	.w5(32'hbaaa6fa8),
	.w6(32'hbbfbca3b),
	.w7(32'hbb9798a9),
	.w8(32'hbacf3927),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a532ff7),
	.w1(32'h3936183c),
	.w2(32'h3ac0f670),
	.w3(32'h3a03c71c),
	.w4(32'h3b89c5e0),
	.w5(32'h3bd38920),
	.w6(32'hba891c69),
	.w7(32'h3ba3c691),
	.w8(32'h39dfecfa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9674a0),
	.w1(32'hbbf4c9fb),
	.w2(32'h38dc8b49),
	.w3(32'hba8aba19),
	.w4(32'hbb9f43c0),
	.w5(32'h3b3a5f45),
	.w6(32'hbc45dae3),
	.w7(32'hbbd0ce70),
	.w8(32'h3b4c6ab7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba380),
	.w1(32'h3b3482a9),
	.w2(32'h3b90723a),
	.w3(32'h3b96d82e),
	.w4(32'h3b581a1b),
	.w5(32'h3a073508),
	.w6(32'hb88d6bce),
	.w7(32'h3b63fba3),
	.w8(32'hbc614862),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77c0072),
	.w1(32'hbbef24ae),
	.w2(32'hbb126c9f),
	.w3(32'hbbb798bb),
	.w4(32'h3a6f85f2),
	.w5(32'h3a91d19b),
	.w6(32'hbc96f522),
	.w7(32'hbc13007d),
	.w8(32'hbbb7be76),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa89bbb),
	.w1(32'hbc172a41),
	.w2(32'hbb1f0248),
	.w3(32'hbbaca119),
	.w4(32'hbb80c77e),
	.w5(32'h3c18bae6),
	.w6(32'hbca075a3),
	.w7(32'hbc20ca5c),
	.w8(32'h3c0bdc32),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ac78),
	.w1(32'h3bbeeea1),
	.w2(32'h3bb770c5),
	.w3(32'h3c0cbfda),
	.w4(32'h3bd95eec),
	.w5(32'hbb6c5ae7),
	.w6(32'hbb8fba77),
	.w7(32'h3b999cda),
	.w8(32'hbbba6466),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3f9ac),
	.w1(32'hbc422282),
	.w2(32'hbc57ed2f),
	.w3(32'hbbe338b3),
	.w4(32'hbb699f7c),
	.w5(32'h3b874c57),
	.w6(32'hbc436244),
	.w7(32'hbc6c3be0),
	.w8(32'h3a5eaaf0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b86dd5),
	.w1(32'hbb8b0305),
	.w2(32'hbad38d70),
	.w3(32'h393c5edd),
	.w4(32'h3a8f7b2b),
	.w5(32'hbb5d6975),
	.w6(32'hb97f9a77),
	.w7(32'hba4d4f80),
	.w8(32'hbc1fdcbf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5915),
	.w1(32'hbc76a862),
	.w2(32'hbc0953d3),
	.w3(32'hbc2f443e),
	.w4(32'hbc030d0d),
	.w5(32'hba08b3ed),
	.w6(32'hbcd55f95),
	.w7(32'hbc5418cf),
	.w8(32'hbc0fa671),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb809f82),
	.w1(32'hbc090248),
	.w2(32'hba6611c5),
	.w3(32'hbc1b1e2e),
	.w4(32'hbc13675d),
	.w5(32'h3bd59223),
	.w6(32'hbcbca301),
	.w7(32'hbbf07532),
	.w8(32'h3b9eb303),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e50b7),
	.w1(32'hba1ef22d),
	.w2(32'hbae20cc7),
	.w3(32'h3c822c69),
	.w4(32'h3b6bba9b),
	.w5(32'hb977c445),
	.w6(32'h3bac69d2),
	.w7(32'h3b5978e2),
	.w8(32'hbbb8cbf9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78b9dc),
	.w1(32'hbc8ef34d),
	.w2(32'hbbc3ce1a),
	.w3(32'hbbb877e4),
	.w4(32'h3b6bafd9),
	.w5(32'hbbe2d9fd),
	.w6(32'hbc1cf13a),
	.w7(32'hbb8d8824),
	.w8(32'hbb5d97d0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a561cc0),
	.w1(32'hbbe173d5),
	.w2(32'hbb560eec),
	.w3(32'hbc0b83f5),
	.w4(32'hbb0c6271),
	.w5(32'h3bad0d2e),
	.w6(32'hbb9b7e52),
	.w7(32'h3b8b4b2d),
	.w8(32'h3b698b64),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98b08f),
	.w1(32'h3aae7289),
	.w2(32'h3bcf32b4),
	.w3(32'h39d71401),
	.w4(32'h3b686c78),
	.w5(32'h3a87e55d),
	.w6(32'hbbf6fea2),
	.w7(32'h3b4de191),
	.w8(32'h3a9b430b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0d49a),
	.w1(32'h3ade78ae),
	.w2(32'h3bd5fe16),
	.w3(32'hbbd2c2b1),
	.w4(32'h3b8ac05f),
	.w5(32'h3b88143a),
	.w6(32'hbc56420a),
	.w7(32'h3bba6191),
	.w8(32'hbae1dedb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc148d5),
	.w1(32'h3bf769a7),
	.w2(32'h3c144f51),
	.w3(32'hba719375),
	.w4(32'h3bedeec5),
	.w5(32'hb9b1aae6),
	.w6(32'hbc475589),
	.w7(32'h3b170d6e),
	.w8(32'hbaafba3e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a6e95),
	.w1(32'hbbe1e1cb),
	.w2(32'hbb5537ed),
	.w3(32'hbb55a895),
	.w4(32'hbb881c0a),
	.w5(32'hbb8563e5),
	.w6(32'hbb9861f0),
	.w7(32'hbba6aac2),
	.w8(32'hbc2e4650),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaf471),
	.w1(32'hbb5a6c51),
	.w2(32'h3a9aee85),
	.w3(32'hbba8e741),
	.w4(32'hbb8209c2),
	.w5(32'hbb5b14dc),
	.w6(32'hbc353f3c),
	.w7(32'hbb7e56f1),
	.w8(32'h3b50a94e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfb9dd),
	.w1(32'hbb3a1850),
	.w2(32'hbbc2810c),
	.w3(32'hbba92118),
	.w4(32'hbb5ece0c),
	.w5(32'hbbb8f528),
	.w6(32'hbb8438e4),
	.w7(32'h3a2cbaef),
	.w8(32'hbb10ce73),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09f5a7),
	.w1(32'hbbb0fd35),
	.w2(32'hbba156bf),
	.w3(32'hbc2ae383),
	.w4(32'hbb796005),
	.w5(32'h3b980a40),
	.w6(32'hbc185084),
	.w7(32'hbb4e5015),
	.w8(32'h3c287c3f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95dfec),
	.w1(32'h3c2010b2),
	.w2(32'h39e2ca8a),
	.w3(32'h3c57be13),
	.w4(32'h3b743632),
	.w5(32'h3c18c627),
	.w6(32'h3cacdf65),
	.w7(32'h3c070284),
	.w8(32'h3b0e9645),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b713269),
	.w1(32'h3bb1cb6f),
	.w2(32'h395ce2d9),
	.w3(32'h3bd629a7),
	.w4(32'hba30e042),
	.w5(32'hbb9cd276),
	.w6(32'h3af1cb50),
	.w7(32'hbaf5899e),
	.w8(32'hbc564e2f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbced841),
	.w1(32'hbc74f0a9),
	.w2(32'hbb2e36bb),
	.w3(32'hbc57963f),
	.w4(32'hbbd27e68),
	.w5(32'h3b42bc04),
	.w6(32'hbc8b9b5f),
	.w7(32'h3af5868f),
	.w8(32'h3b86bd8d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96ea35),
	.w1(32'h3baf0189),
	.w2(32'h3bae9dbe),
	.w3(32'h3b8b0ad1),
	.w4(32'h3aa8f14f),
	.w5(32'h3ab74073),
	.w6(32'h3bdf5e0b),
	.w7(32'h3b3e9fe4),
	.w8(32'hba5663a8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15ac1e),
	.w1(32'hbb7ad521),
	.w2(32'h3b4a27ea),
	.w3(32'hbb8e93b2),
	.w4(32'hb8effb6a),
	.w5(32'h3b22bd2e),
	.w6(32'hbca918c4),
	.w7(32'hbb91323d),
	.w8(32'h3b68e59b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2081e3),
	.w1(32'h3b9abfc8),
	.w2(32'h3b9ccf46),
	.w3(32'h3b17d8d9),
	.w4(32'h3b2cb296),
	.w5(32'h3ae9d561),
	.w6(32'hbb7783c1),
	.w7(32'h3b938a6f),
	.w8(32'hbaaa19fc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b4bbc),
	.w1(32'hbb89d986),
	.w2(32'hba9f1131),
	.w3(32'h3aa312f5),
	.w4(32'h3b11ba24),
	.w5(32'hba197800),
	.w6(32'h3a3ce5bd),
	.w7(32'hbb8d362c),
	.w8(32'h3bcea0e9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad506a),
	.w1(32'h3b156738),
	.w2(32'hbbc1bc55),
	.w3(32'h3b76118b),
	.w4(32'h3c01eea3),
	.w5(32'h3b5a8774),
	.w6(32'h3b7999c8),
	.w7(32'h3ba940ae),
	.w8(32'h3b8ef84a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d71d7),
	.w1(32'hbad6b1ef),
	.w2(32'hbbcb46fa),
	.w3(32'hbc031fe7),
	.w4(32'hbbc3adb3),
	.w5(32'hbb4f26ea),
	.w6(32'hbc0679ab),
	.w7(32'hbbd4930a),
	.w8(32'h3c3d2a50),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cb6d1),
	.w1(32'h3b4ac9eb),
	.w2(32'h3c4bba77),
	.w3(32'hbc001c39),
	.w4(32'h3b28b2c8),
	.w5(32'h3b978535),
	.w6(32'hbac1373f),
	.w7(32'h3c458e40),
	.w8(32'h3ab0e807),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11dc33),
	.w1(32'h3afc92d6),
	.w2(32'h3b408016),
	.w3(32'h3bd483a9),
	.w4(32'h3bc6ba1b),
	.w5(32'hbb93e837),
	.w6(32'hbb22c01e),
	.w7(32'h3bb58ec0),
	.w8(32'hbb2a7a12),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909ca1a),
	.w1(32'h3b791dc6),
	.w2(32'h3a1c7696),
	.w3(32'hbb6a2d5d),
	.w4(32'h399db60a),
	.w5(32'hbb443bdf),
	.w6(32'hbbfb1db9),
	.w7(32'h381d0582),
	.w8(32'hbbd1001e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cad45),
	.w1(32'hbbb5f9cd),
	.w2(32'hbb702ac1),
	.w3(32'hbb8f20a4),
	.w4(32'hbb9ff10a),
	.w5(32'hbb4d390b),
	.w6(32'hbbde19e7),
	.w7(32'hbbf0f97c),
	.w8(32'hba9fd539),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fddcb),
	.w1(32'h3b319284),
	.w2(32'h3af9cc75),
	.w3(32'h3b7bceeb),
	.w4(32'h3b9861b3),
	.w5(32'hbb808c83),
	.w6(32'h3bcd9a82),
	.w7(32'h3bb8b38c),
	.w8(32'hbc1228d4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07d4be),
	.w1(32'hbb387e56),
	.w2(32'h3c3ce226),
	.w3(32'hbb808b3d),
	.w4(32'hba8afa1c),
	.w5(32'hbb147205),
	.w6(32'hbc14a34d),
	.w7(32'h3a52a8cf),
	.w8(32'h3ad764ad),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b102dc7),
	.w1(32'h3abdda6e),
	.w2(32'h3990f7a0),
	.w3(32'hbbbbaee1),
	.w4(32'hbab2255c),
	.w5(32'h3ad864cc),
	.w6(32'h3a813aef),
	.w7(32'h3b5a1985),
	.w8(32'hbc35a64d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2b68d),
	.w1(32'hbb94dbe9),
	.w2(32'hbaf36064),
	.w3(32'hbbaa806f),
	.w4(32'h3b2d16ce),
	.w5(32'h3b2b847f),
	.w6(32'hbcce0806),
	.w7(32'hbb89723b),
	.w8(32'hba90b401),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec5dc4),
	.w1(32'h3a330306),
	.w2(32'h3a819309),
	.w3(32'h3b5d7fb0),
	.w4(32'h3a4ab5b9),
	.w5(32'h3bcef71f),
	.w6(32'hba87b6f8),
	.w7(32'hbac084d1),
	.w8(32'h3b786c3d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb86618),
	.w1(32'h3c1b8769),
	.w2(32'h3c0bf924),
	.w3(32'h3c4cd834),
	.w4(32'h3b62bc4b),
	.w5(32'hbaa19723),
	.w6(32'h3c06b541),
	.w7(32'h3bf65c8a),
	.w8(32'h3aba19fd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab82500),
	.w1(32'hbb054ccf),
	.w2(32'hbbf70d6a),
	.w3(32'h3b15d5ac),
	.w4(32'hbc23226c),
	.w5(32'h3a32868f),
	.w6(32'h3c35d077),
	.w7(32'hbbda3efd),
	.w8(32'hbae383d2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9aacc),
	.w1(32'hbb0905f3),
	.w2(32'h39b5855c),
	.w3(32'hbb8c4e4b),
	.w4(32'h38f7c82e),
	.w5(32'h3b1be111),
	.w6(32'hbcc4d5cf),
	.w7(32'hbb921136),
	.w8(32'hbb9733cf),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4c9b7),
	.w1(32'h3aa679f0),
	.w2(32'hba1a39b7),
	.w3(32'hbb17a0a4),
	.w4(32'hbb2b8e1f),
	.w5(32'hbad38391),
	.w6(32'hbc0ba3f0),
	.w7(32'hbbbb98b9),
	.w8(32'hbbea30b1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de93c3),
	.w1(32'hbc297717),
	.w2(32'h3c8c355f),
	.w3(32'hbc724762),
	.w4(32'h3bcf2ecf),
	.w5(32'h3c55365e),
	.w6(32'hbcd9f673),
	.w7(32'h3b3cfb72),
	.w8(32'h3c2228f6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5901e6),
	.w1(32'h3c00498f),
	.w2(32'h3c0a5be1),
	.w3(32'h3c41d3af),
	.w4(32'h3c0bd5bd),
	.w5(32'h3b626173),
	.w6(32'hbb87b34d),
	.w7(32'h3b2739e6),
	.w8(32'h3b30215f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f53c1),
	.w1(32'h3b1fe23a),
	.w2(32'h3bc9eb30),
	.w3(32'hbb539d78),
	.w4(32'h3b970a02),
	.w5(32'hbb06b125),
	.w6(32'hbb871066),
	.w7(32'h3ac20ee5),
	.w8(32'hbac1e97a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae440a7),
	.w1(32'hbaedbf0c),
	.w2(32'h3b35c21b),
	.w3(32'hbb3055d1),
	.w4(32'h3b3677f7),
	.w5(32'h3b7f12b1),
	.w6(32'hbc0c1b13),
	.w7(32'h3ab3c1a3),
	.w8(32'h3bb77600),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d9e87),
	.w1(32'h3b26c0c0),
	.w2(32'hbbb1c2ff),
	.w3(32'h3c2c967f),
	.w4(32'h3ac4beb2),
	.w5(32'h3acf4184),
	.w6(32'h3c9c4d8e),
	.w7(32'h3b79344a),
	.w8(32'hbb96d4dc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1b7fe),
	.w1(32'hbb7b6ee3),
	.w2(32'h3b7210be),
	.w3(32'h3ad9ed21),
	.w4(32'h3ba25cdc),
	.w5(32'h3aa9a772),
	.w6(32'hbb44fdd1),
	.w7(32'hbad359de),
	.w8(32'h3b446291),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0782aa),
	.w1(32'h3be46bae),
	.w2(32'h3a7379c5),
	.w3(32'h3be94727),
	.w4(32'h3b8fbe0b),
	.w5(32'h3af9477e),
	.w6(32'h3baf90fd),
	.w7(32'h3baf7e0c),
	.w8(32'hbaf3c2be),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8514d7),
	.w1(32'hbc04ed21),
	.w2(32'h3b2cd233),
	.w3(32'hbbe5cb13),
	.w4(32'hbba6a0aa),
	.w5(32'h3a28e2da),
	.w6(32'hbbf8734b),
	.w7(32'hbb97f366),
	.w8(32'h3a0cb95c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e9c4d),
	.w1(32'hbb87813a),
	.w2(32'hbba744cf),
	.w3(32'h3842bf33),
	.w4(32'h3b2a79e9),
	.w5(32'h3c5591fb),
	.w6(32'hbc140040),
	.w7(32'hbb44a299),
	.w8(32'h3b844681),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba21483),
	.w1(32'h3bb803c9),
	.w2(32'h3c28b034),
	.w3(32'h3b42c646),
	.w4(32'hbbe03241),
	.w5(32'h3c3c896b),
	.w6(32'h3a3ec016),
	.w7(32'h3b27b1e3),
	.w8(32'h3c611554),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d6c91),
	.w1(32'h3c39611c),
	.w2(32'hbb5e3449),
	.w3(32'h3bcbe1bd),
	.w4(32'hbb883092),
	.w5(32'hbb44ff86),
	.w6(32'h3a342b6b),
	.w7(32'hbbae0e5e),
	.w8(32'h3a9cf1bc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaa140),
	.w1(32'hbbadebc1),
	.w2(32'hbbab064b),
	.w3(32'hbbca6ddb),
	.w4(32'hbb3f96a2),
	.w5(32'hba9136d6),
	.w6(32'hbbcb4a51),
	.w7(32'hba2650fc),
	.w8(32'hbbda6c28),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb196f8),
	.w1(32'hbbb53be9),
	.w2(32'hb97079aa),
	.w3(32'h3b8cc348),
	.w4(32'h3b99dcea),
	.w5(32'h39b67e47),
	.w6(32'hbbb95527),
	.w7(32'h3bf15a14),
	.w8(32'h3b7a59e0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9da71),
	.w1(32'hb95dcc36),
	.w2(32'hbbee2536),
	.w3(32'h3b6fcec0),
	.w4(32'hbba8d45f),
	.w5(32'h3a9d32b8),
	.w6(32'h3c494319),
	.w7(32'hbb3f8c4a),
	.w8(32'h3b5c44cf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be42e2c),
	.w1(32'h3a73b82b),
	.w2(32'hba89be38),
	.w3(32'hbb8215b6),
	.w4(32'hba85d2be),
	.w5(32'h3b34bf9f),
	.w6(32'hbc1ed795),
	.w7(32'hbae2df7d),
	.w8(32'h3b767bd1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa5ac4),
	.w1(32'h3bc752e5),
	.w2(32'h3a954bc1),
	.w3(32'h3b8819a5),
	.w4(32'h3b98b3f0),
	.w5(32'h3b27dbfd),
	.w6(32'hba580187),
	.w7(32'h3b7a5be7),
	.w8(32'hbb055caa),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50193c),
	.w1(32'hbb4d8e0c),
	.w2(32'hbc10f3a6),
	.w3(32'h3c15e7d6),
	.w4(32'h3c2fc1ed),
	.w5(32'hbb715bea),
	.w6(32'h3b20b4d6),
	.w7(32'h3ab885ac),
	.w8(32'hbb92e282),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1701f),
	.w1(32'hbb19e7a2),
	.w2(32'hbaedf747),
	.w3(32'hbb85f6d9),
	.w4(32'hbba3fa06),
	.w5(32'hb90d62f6),
	.w6(32'hbbe034e8),
	.w7(32'hbb126a90),
	.w8(32'hbab1ec2f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b60da1),
	.w1(32'h3ab7d688),
	.w2(32'h3c158776),
	.w3(32'hbbd09e5e),
	.w4(32'h3b7e8c9e),
	.w5(32'hbb99c22a),
	.w6(32'hbc88089b),
	.w7(32'h3b2bccde),
	.w8(32'hbc491758),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b529ba6),
	.w1(32'h3b696ee1),
	.w2(32'h3bba2d43),
	.w3(32'h3ab2c0fb),
	.w4(32'h3a9718df),
	.w5(32'h3802859d),
	.w6(32'hbc182be1),
	.w7(32'hbbe71775),
	.w8(32'h3896b3ff),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7595d65),
	.w1(32'hbb7f75ae),
	.w2(32'hbb087eea),
	.w3(32'hbb47d9ea),
	.w4(32'hbb39d91b),
	.w5(32'hbb80de0c),
	.w6(32'h3aaafe96),
	.w7(32'hbac7a151),
	.w8(32'hbaae545a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9c3d0),
	.w1(32'hbc1f2357),
	.w2(32'hbbbdb8be),
	.w3(32'hbb6838e0),
	.w4(32'h3babc05e),
	.w5(32'h3b9f7e40),
	.w6(32'hbc15d9a5),
	.w7(32'h39af4268),
	.w8(32'h3b560408),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf11d48),
	.w1(32'h3b92c1d7),
	.w2(32'h3b461197),
	.w3(32'h3b29ce19),
	.w4(32'hbb440963),
	.w5(32'h37df2724),
	.w6(32'hb8d92611),
	.w7(32'hbae269c6),
	.w8(32'hbb921b73),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a9f45),
	.w1(32'hb9d72848),
	.w2(32'h3c142165),
	.w3(32'hbb45dd8a),
	.w4(32'h3b754e0e),
	.w5(32'h3b839fd6),
	.w6(32'hbc17ba5d),
	.w7(32'h3b6ceff0),
	.w8(32'h3b9dc3e7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97059c),
	.w1(32'hbc1004b1),
	.w2(32'h3b262f9e),
	.w3(32'hbaef27ee),
	.w4(32'h3a8fe048),
	.w5(32'hbb219d6a),
	.w6(32'hbbb5d14e),
	.w7(32'h3a20060c),
	.w8(32'hbbc0420f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d9c4c),
	.w1(32'hbc2a11dc),
	.w2(32'hbb44413f),
	.w3(32'hbc39dcf8),
	.w4(32'h3a30c278),
	.w5(32'hbad08452),
	.w6(32'hbc7e61f6),
	.w7(32'hbb8ee3b7),
	.w8(32'hbbf5de4f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeba104),
	.w1(32'hbba75574),
	.w2(32'h39be5337),
	.w3(32'hbb236716),
	.w4(32'h3933b9ea),
	.w5(32'h3b236dcc),
	.w6(32'hbc863065),
	.w7(32'hbb885b04),
	.w8(32'h3b487ded),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9024cb),
	.w1(32'h3b95a342),
	.w2(32'h3b8a94a4),
	.w3(32'h3b52a85d),
	.w4(32'h3b34f04c),
	.w5(32'h3a80ea24),
	.w6(32'h3a06d34a),
	.w7(32'h3b1fd44a),
	.w8(32'h3be77a36),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee5b4),
	.w1(32'hbbb9d372),
	.w2(32'hbb9461b0),
	.w3(32'h38c99f37),
	.w4(32'h3ad6fea6),
	.w5(32'h3c0bf5da),
	.w6(32'hbb11c060),
	.w7(32'hbb86875c),
	.w8(32'h3adcfb46),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80be33),
	.w1(32'hbbca8a56),
	.w2(32'hbb119b16),
	.w3(32'h3c3d13cd),
	.w4(32'h3bf50c16),
	.w5(32'h3a677e15),
	.w6(32'h3a9716fd),
	.w7(32'h3b15e778),
	.w8(32'hba6780a9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0e9b4),
	.w1(32'h3b43e91e),
	.w2(32'hbb67073b),
	.w3(32'hbada35db),
	.w4(32'hbbc939eb),
	.w5(32'h3af6579e),
	.w6(32'hbb84c2cb),
	.w7(32'hbbe39ff6),
	.w8(32'hbbfb8429),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4d5ca),
	.w1(32'h3ba79cfb),
	.w2(32'h3c11833c),
	.w3(32'hbaff68f4),
	.w4(32'h3b365b94),
	.w5(32'h3bb22786),
	.w6(32'hbbf6ff7f),
	.w7(32'h3ba86ca4),
	.w8(32'h3ae9073b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ba298),
	.w1(32'hbc0e5781),
	.w2(32'hbc02e8f4),
	.w3(32'h3b70cc44),
	.w4(32'h39830ede),
	.w5(32'h3acf4e2b),
	.w6(32'h3b0e2165),
	.w7(32'hbbc2faeb),
	.w8(32'hbb15c4ba),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e1ae0),
	.w1(32'h3a878e5b),
	.w2(32'h3956614a),
	.w3(32'hba645c5b),
	.w4(32'hbbcea403),
	.w5(32'hbbef2d68),
	.w6(32'h3b33c7d4),
	.w7(32'hbaf2e4cb),
	.w8(32'hbc0b9a70),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31adc4),
	.w1(32'hbbbaddb3),
	.w2(32'hba096ff2),
	.w3(32'hbb97d1ef),
	.w4(32'hba940862),
	.w5(32'h3ab3746c),
	.w6(32'hbc696a77),
	.w7(32'hbaca2940),
	.w8(32'hb9544b82),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44cd0f),
	.w1(32'hbc1a081e),
	.w2(32'hbbff666b),
	.w3(32'hba852af4),
	.w4(32'hba16e16d),
	.w5(32'h3baf2e95),
	.w6(32'hbbaeb31b),
	.w7(32'hbc1ba537),
	.w8(32'h3b058388),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfed8b6),
	.w1(32'hbaed817d),
	.w2(32'h3c1bc4e8),
	.w3(32'h3b364a7f),
	.w4(32'h3bccb4ea),
	.w5(32'hb9a67868),
	.w6(32'hbb9042bb),
	.w7(32'h3aeedccc),
	.w8(32'h3b97f7b8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae05c39),
	.w1(32'hbb2a2a9b),
	.w2(32'hbc4126d7),
	.w3(32'h3b5e91d3),
	.w4(32'h3b85e59a),
	.w5(32'hbb474bd1),
	.w6(32'h3c63bf59),
	.w7(32'h3998ea5a),
	.w8(32'hbb68d7ed),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27d10a),
	.w1(32'hbaa32fad),
	.w2(32'hbb0889a8),
	.w3(32'hba7552c9),
	.w4(32'hbb27431c),
	.w5(32'h3a386430),
	.w6(32'hbba48ed4),
	.w7(32'hbbaf493b),
	.w8(32'hbb8ebfb7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84505c),
	.w1(32'hbb738e60),
	.w2(32'h3bf39cfd),
	.w3(32'hbc202640),
	.w4(32'hbb609239),
	.w5(32'h3ae42b72),
	.w6(32'hbc11a449),
	.w7(32'h3aca5d43),
	.w8(32'h3ac14a30),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c4c4f),
	.w1(32'hbbc5f4e4),
	.w2(32'hbb68a8a0),
	.w3(32'hbbe0185a),
	.w4(32'hbbab47c6),
	.w5(32'h3b0850a8),
	.w6(32'hbc555ddc),
	.w7(32'hbba5d2b2),
	.w8(32'hbae10fa8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d399a),
	.w1(32'hba568522),
	.w2(32'h3bd14e53),
	.w3(32'hbb0485af),
	.w4(32'hbb16b556),
	.w5(32'h3ab940f0),
	.w6(32'hbb65c9ee),
	.w7(32'hba9096b0),
	.w8(32'hbb62dce5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e41377),
	.w1(32'hbafc491b),
	.w2(32'hbb06cf50),
	.w3(32'hbb84d4f8),
	.w4(32'hbbb4e5de),
	.w5(32'hbaa677de),
	.w6(32'hbc690484),
	.w7(32'hbc34822d),
	.w8(32'hb769aba6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06b8e5),
	.w1(32'hbb9dffc1),
	.w2(32'hbb998689),
	.w3(32'hbb316d13),
	.w4(32'hbb255c5f),
	.w5(32'h3b1bbb13),
	.w6(32'hbc85bc9a),
	.w7(32'hbb87db25),
	.w8(32'hbb513b43),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba14424),
	.w1(32'h3bb6d9b2),
	.w2(32'h3af8bfb4),
	.w3(32'h3b14d367),
	.w4(32'h3a4f1375),
	.w5(32'h3bb91882),
	.w6(32'hbb35ecf4),
	.w7(32'hbb1fafae),
	.w8(32'h3b5cf078),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9b830),
	.w1(32'h3bdef4a6),
	.w2(32'h3c0cb5d8),
	.w3(32'h3af989b0),
	.w4(32'h3c0a7cda),
	.w5(32'hbc4093a4),
	.w6(32'hbbab73b4),
	.w7(32'h3bfdbddd),
	.w8(32'hbc35ecf0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc483d1b),
	.w1(32'hbbf2304e),
	.w2(32'hbb59f423),
	.w3(32'hbc13e450),
	.w4(32'hbbde601e),
	.w5(32'hbb63eb62),
	.w6(32'hbc1b2e87),
	.w7(32'hbc431933),
	.w8(32'hbc0638c9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf436a0),
	.w1(32'hbc0ead83),
	.w2(32'h3a8cf384),
	.w3(32'hbb380420),
	.w4(32'hbb86ca64),
	.w5(32'hbad8fe7b),
	.w6(32'h3ab828cd),
	.w7(32'h3b7114b4),
	.w8(32'hbb8b6779),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ccdc1),
	.w1(32'hbbcf7fb1),
	.w2(32'hb9086e0e),
	.w3(32'hbb9d0465),
	.w4(32'h3ab45c20),
	.w5(32'hbbad90c2),
	.w6(32'hbc039ec5),
	.w7(32'hbb7d902c),
	.w8(32'hbbe9f86f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf9982),
	.w1(32'hbb811d87),
	.w2(32'h3c487992),
	.w3(32'h3a379437),
	.w4(32'h3bdfdd03),
	.w5(32'hbb03fd14),
	.w6(32'hbc9a4411),
	.w7(32'h3c667abb),
	.w8(32'hbbe1db18),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c1703),
	.w1(32'hbb9deb6e),
	.w2(32'h3c31e95e),
	.w3(32'hbc468ede),
	.w4(32'h3ad1e7a5),
	.w5(32'hbabb15ae),
	.w6(32'hbc325d22),
	.w7(32'hba5a97fb),
	.w8(32'hbbc1c1fc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f9b50),
	.w1(32'hbc1b1a56),
	.w2(32'hb8356acd),
	.w3(32'hbb44573f),
	.w4(32'h3b58c72f),
	.w5(32'h3be57e00),
	.w6(32'hbc51d3ad),
	.w7(32'hbb06103e),
	.w8(32'hbb7e7ebc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e446b),
	.w1(32'hbb56048a),
	.w2(32'h3b357dc6),
	.w3(32'h3b96c392),
	.w4(32'h3c121ee9),
	.w5(32'h3b5a1e80),
	.w6(32'hbc568361),
	.w7(32'h3b3d9d0a),
	.w8(32'hbaa441db),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc04b56),
	.w1(32'hbbd1eb66),
	.w2(32'hbc43efc0),
	.w3(32'h3bb596c3),
	.w4(32'hbb5669a6),
	.w5(32'hb8cb0f1e),
	.w6(32'h3bf7362d),
	.w7(32'hbc00588c),
	.w8(32'h3b832b38),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6876ae),
	.w1(32'h3b13d427),
	.w2(32'h3c5b8216),
	.w3(32'h3b8ce591),
	.w4(32'hbac915e3),
	.w5(32'hbb317501),
	.w6(32'h3bab777f),
	.w7(32'h3aa55a43),
	.w8(32'hbb50203b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae94331),
	.w1(32'hb9a32bbb),
	.w2(32'hba25c9dd),
	.w3(32'h3ae5118e),
	.w4(32'h3b204d4a),
	.w5(32'h3631b7e8),
	.w6(32'h3b0075bd),
	.w7(32'hba4e80f8),
	.w8(32'hbb4e56ac),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d0db4),
	.w1(32'h39b629f4),
	.w2(32'hba9c50c5),
	.w3(32'hbb0b7259),
	.w4(32'hbafca594),
	.w5(32'hbaba8798),
	.w6(32'h3b92fdc5),
	.w7(32'hba622684),
	.w8(32'hbad3c6ea),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98b84e),
	.w1(32'hbb8e5c20),
	.w2(32'hbab62f82),
	.w3(32'hbb28a7e2),
	.w4(32'h3b4f2243),
	.w5(32'h3a7f8a72),
	.w6(32'hbb19d513),
	.w7(32'h3b6f4dea),
	.w8(32'h3b156496),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5e183),
	.w1(32'hbadadeb8),
	.w2(32'hbb33545c),
	.w3(32'hbac2f2ee),
	.w4(32'hbab74803),
	.w5(32'hbb53907b),
	.w6(32'hbb2d736e),
	.w7(32'hbb039008),
	.w8(32'hbab6fc92),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dbd6fe),
	.w1(32'hba22c2f9),
	.w2(32'h3a9311b7),
	.w3(32'h3a546698),
	.w4(32'h3b3973ac),
	.w5(32'h3ab2dcbc),
	.w6(32'h3af9c92b),
	.w7(32'h3a96621a),
	.w8(32'hba0ff7af),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a217e12),
	.w1(32'h3b1b91b6),
	.w2(32'h3b529e39),
	.w3(32'h3a19c867),
	.w4(32'hb9a22416),
	.w5(32'h3ac745e0),
	.w6(32'hba6f72f6),
	.w7(32'h3b3ae1a6),
	.w8(32'h3b1a2cc7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb905afd),
	.w1(32'hbbd0dcea),
	.w2(32'hbbca1ef7),
	.w3(32'hbbb484b8),
	.w4(32'hbb87be98),
	.w5(32'h382dc7e0),
	.w6(32'hba585fa7),
	.w7(32'h38482308),
	.w8(32'hbae45b7c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb872cac0),
	.w1(32'h39fa0a3d),
	.w2(32'hbb09b843),
	.w3(32'h3a64ea69),
	.w4(32'h39d0779b),
	.w5(32'hbb55909f),
	.w6(32'h3ab822d3),
	.w7(32'h3a6510c8),
	.w8(32'hbb15d0ba),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1477a3),
	.w1(32'hba809f79),
	.w2(32'hbb2f0443),
	.w3(32'hbaddf3f8),
	.w4(32'hbb4f907f),
	.w5(32'hba4ad795),
	.w6(32'hbab03236),
	.w7(32'hbb64802b),
	.w8(32'hb9cea816),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7459c4),
	.w1(32'h3a83b759),
	.w2(32'hbaa7e581),
	.w3(32'h399f99c3),
	.w4(32'h3a5841f8),
	.w5(32'hbad9fc04),
	.w6(32'h3ac62f29),
	.w7(32'h378832d8),
	.w8(32'hb860ce07),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cf5b9),
	.w1(32'h3b2ad843),
	.w2(32'hb9641203),
	.w3(32'h3b0e08f6),
	.w4(32'h3aa0b15f),
	.w5(32'hbb2838b0),
	.w6(32'h3b1ac47d),
	.w7(32'h39dde453),
	.w8(32'hbb130938),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a534d75),
	.w1(32'h3a37f262),
	.w2(32'hbb46552c),
	.w3(32'h3a5c7f0c),
	.w4(32'h3a9ea213),
	.w5(32'hba7ba78d),
	.w6(32'h3aadd22c),
	.w7(32'h3a4bf5d1),
	.w8(32'h39f0fce0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e8f95),
	.w1(32'hbae55560),
	.w2(32'hbb5538a2),
	.w3(32'hbac0043c),
	.w4(32'hbb2037b6),
	.w5(32'hba4d38f2),
	.w6(32'h3b06259e),
	.w7(32'hbac04c4d),
	.w8(32'hba745cbb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d981a),
	.w1(32'hbae6d6a7),
	.w2(32'hb9791e4b),
	.w3(32'hbb128b6c),
	.w4(32'hba011c20),
	.w5(32'h39bbdc6f),
	.w6(32'hbaed99f2),
	.w7(32'hb6902c6c),
	.w8(32'hbabe4fac),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9043d86),
	.w1(32'h3a128f96),
	.w2(32'h39e32155),
	.w3(32'h3a84e8c0),
	.w4(32'h3a933c01),
	.w5(32'h3ae723a3),
	.w6(32'h3a343ce5),
	.w7(32'h3b00f20b),
	.w8(32'h3b7a38ef),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940ad72),
	.w1(32'h3a4c5486),
	.w2(32'hba470a33),
	.w3(32'hba744b6c),
	.w4(32'hb71159d2),
	.w5(32'h3b824922),
	.w6(32'hb9a3f892),
	.w7(32'hb908219d),
	.w8(32'h3af69379),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b048ca9),
	.w1(32'h3b298db9),
	.w2(32'h3b5a6f97),
	.w3(32'h3aba9206),
	.w4(32'h3ababd5d),
	.w5(32'hbaea9263),
	.w6(32'h3b5b7dfa),
	.w7(32'h3b01d48a),
	.w8(32'hbb214b8e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eff6c),
	.w1(32'hba4f1021),
	.w2(32'hba0437fd),
	.w3(32'hbb23ba07),
	.w4(32'hba722891),
	.w5(32'hbab8f013),
	.w6(32'hbb402a93),
	.w7(32'hb9b6270c),
	.w8(32'hbb0b6dfc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafd843),
	.w1(32'hba0d9a15),
	.w2(32'h3a17f2f5),
	.w3(32'hba283cbe),
	.w4(32'hb9427946),
	.w5(32'hb84fb66c),
	.w6(32'hbaaddbdb),
	.w7(32'hb9948978),
	.w8(32'h3a3141e0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a21b6),
	.w1(32'h39e1cb9a),
	.w2(32'hba5d399e),
	.w3(32'hba61246b),
	.w4(32'hb98ae5b4),
	.w5(32'h3956594b),
	.w6(32'h3ad190c4),
	.w7(32'hba14d714),
	.w8(32'h3abca0df),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f32f0),
	.w1(32'h3a536024),
	.w2(32'h3aa68d28),
	.w3(32'h3737d0cf),
	.w4(32'h3a732bac),
	.w5(32'hbb0b77cc),
	.w6(32'h39f8dc5c),
	.w7(32'h3ae3e4fa),
	.w8(32'hb9871826),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1214c2),
	.w1(32'h3a0595c4),
	.w2(32'h39b06813),
	.w3(32'hbb1a9d58),
	.w4(32'hb9cab1c7),
	.w5(32'hba9a8e07),
	.w6(32'hbb59c2ad),
	.w7(32'h3a561b35),
	.w8(32'hba92c9bc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1efe5),
	.w1(32'hbaf35a9a),
	.w2(32'hbabd1c15),
	.w3(32'hbaae223c),
	.w4(32'hbadf7e3e),
	.w5(32'hb94b605b),
	.w6(32'hbb4de7fa),
	.w7(32'h3914302a),
	.w8(32'hba2a2c95),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe5f44),
	.w1(32'hbad5b814),
	.w2(32'hba93b03c),
	.w3(32'hb9452231),
	.w4(32'hba82b27d),
	.w5(32'h3a233557),
	.w6(32'h3a869be4),
	.w7(32'hba75d65b),
	.w8(32'hbaa381f9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99d4a2),
	.w1(32'hba16a2cd),
	.w2(32'hbac2256f),
	.w3(32'h3a07ef9d),
	.w4(32'hba881436),
	.w5(32'hb92b7e91),
	.w6(32'hba80898a),
	.w7(32'hba69cd96),
	.w8(32'h3a0c385f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba287a9d),
	.w1(32'hba34ef90),
	.w2(32'hba19d618),
	.w3(32'hba52cd38),
	.w4(32'h3a042c24),
	.w5(32'h3a82a05b),
	.w6(32'hb9ba192c),
	.w7(32'hba9e2e92),
	.w8(32'h3a2cfb76),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bdddb),
	.w1(32'h388f5576),
	.w2(32'hb9bcfd49),
	.w3(32'hb6fbfd7b),
	.w4(32'hba1a7d7a),
	.w5(32'hb836129c),
	.w6(32'h3a02c1e1),
	.w7(32'hba033c75),
	.w8(32'h3aa2f1c8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb877c),
	.w1(32'h3a3ee038),
	.w2(32'h3a7cd0b8),
	.w3(32'hb919e4ac),
	.w4(32'hba63fea9),
	.w5(32'hb9b8fc4c),
	.w6(32'h3b678827),
	.w7(32'h3a02e60c),
	.w8(32'hba998125),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95e59b),
	.w1(32'hb9b0e496),
	.w2(32'h3666fd82),
	.w3(32'h39d67379),
	.w4(32'h398d9db3),
	.w5(32'hb9853398),
	.w6(32'h39e256ed),
	.w7(32'hb898c644),
	.w8(32'h3a0f36f2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42f04c),
	.w1(32'h3a32ddc8),
	.w2(32'hbb10ad19),
	.w3(32'h3b7989ff),
	.w4(32'hba1cec51),
	.w5(32'hbb40c585),
	.w6(32'h3b00da97),
	.w7(32'h3a6d8a04),
	.w8(32'hb9912632),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b089b82),
	.w1(32'hb8e29177),
	.w2(32'hbb2349dc),
	.w3(32'h381b0740),
	.w4(32'h389ef541),
	.w5(32'h3aa3b62f),
	.w6(32'h39fa2999),
	.w7(32'h39aef33f),
	.w8(32'hbb2f6057),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5864a),
	.w1(32'hbb0f5964),
	.w2(32'h3a2effde),
	.w3(32'hb8bad00c),
	.w4(32'h3a4ed632),
	.w5(32'h38931bc7),
	.w6(32'hbae56dc8),
	.w7(32'hbadf8bc2),
	.w8(32'hba633e13),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ae05b),
	.w1(32'hbada0ec0),
	.w2(32'hba44d369),
	.w3(32'hbad8a963),
	.w4(32'hba9fd9cc),
	.w5(32'hb980dafc),
	.w6(32'hbac1cfe8),
	.w7(32'hb923c0a3),
	.w8(32'hba615a3c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1afbe),
	.w1(32'h3991e90f),
	.w2(32'h3a358b5d),
	.w3(32'h39b55a07),
	.w4(32'h3a2c840d),
	.w5(32'h38a41930),
	.w6(32'h3ab6a8d0),
	.w7(32'h3a844335),
	.w8(32'hba752c3b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90d3cf),
	.w1(32'h3b0fbf2c),
	.w2(32'h39a44e6e),
	.w3(32'h3ae34d73),
	.w4(32'hba25c78e),
	.w5(32'hbb2793b3),
	.w6(32'h39c56e99),
	.w7(32'h3ae33830),
	.w8(32'hbaf2948b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb380673),
	.w1(32'hba86697e),
	.w2(32'hbb325467),
	.w3(32'hbb0ceeb6),
	.w4(32'hbaac96b4),
	.w5(32'hbb0eaf80),
	.w6(32'h3a29fad6),
	.w7(32'hba1fa1bd),
	.w8(32'hbb018daa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac712c),
	.w1(32'hbb1f5f6c),
	.w2(32'hbaffee8b),
	.w3(32'hbafad067),
	.w4(32'hbaa4bb27),
	.w5(32'hbb4cda96),
	.w6(32'hba272db0),
	.w7(32'hbb3cfe82),
	.w8(32'hbbc81956),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5794),
	.w1(32'hbb2ef735),
	.w2(32'hbb2e6cef),
	.w3(32'hbb1d245e),
	.w4(32'hbb311a25),
	.w5(32'hba666bae),
	.w6(32'hbb226a44),
	.w7(32'hba9ceacd),
	.w8(32'hba63ef3c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd3cfc),
	.w1(32'hba4a7c68),
	.w2(32'hba80df68),
	.w3(32'h399ae498),
	.w4(32'h392d436d),
	.w5(32'hbadcba0e),
	.w6(32'hba9403f3),
	.w7(32'hbab5be83),
	.w8(32'hbb1e3c2c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24b836),
	.w1(32'hbae99824),
	.w2(32'hbb24c88a),
	.w3(32'h38c8c1e4),
	.w4(32'hb9a8e646),
	.w5(32'hbb088a41),
	.w6(32'h3afb0155),
	.w7(32'hba1db085),
	.w8(32'hbb656386),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6a90e),
	.w1(32'hb7ddbd1d),
	.w2(32'hba5a5e6d),
	.w3(32'hb80b5a6f),
	.w4(32'h39c79d0b),
	.w5(32'h3aa8a694),
	.w6(32'h3ad0ebd1),
	.w7(32'h377399e2),
	.w8(32'h3a92a8be),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaee205),
	.w1(32'h3976cccf),
	.w2(32'hbb19a30d),
	.w3(32'h3aab6f34),
	.w4(32'hba1316ee),
	.w5(32'hba03a3f5),
	.w6(32'hb9f3d61b),
	.w7(32'hba68b79a),
	.w8(32'hba3a8865),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46cf8e),
	.w1(32'hbaa18420),
	.w2(32'hbb1316c2),
	.w3(32'hba71cce5),
	.w4(32'hbb084999),
	.w5(32'hba87fcec),
	.w6(32'hbad858b4),
	.w7(32'hbadc12c0),
	.w8(32'hb842429e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31b50c),
	.w1(32'h3a7b3685),
	.w2(32'hba9b7fdf),
	.w3(32'h3b8e14d3),
	.w4(32'h3ac1781c),
	.w5(32'hbb3cfb92),
	.w6(32'h3b62db72),
	.w7(32'h3a2900c4),
	.w8(32'hbb01e6c7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b7706),
	.w1(32'h3abc59c6),
	.w2(32'hba5bba57),
	.w3(32'hba53699e),
	.w4(32'hba241add),
	.w5(32'hb8da50df),
	.w6(32'h3b2e3bc6),
	.w7(32'hb91ad732),
	.w8(32'h3912a1eb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8831656),
	.w1(32'hba2890bc),
	.w2(32'hba3dd581),
	.w3(32'hba36ff93),
	.w4(32'h39117606),
	.w5(32'hbaa4e6ba),
	.w6(32'hb917ea9f),
	.w7(32'h3a8ce7e2),
	.w8(32'hbae87251),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f27bd),
	.w1(32'hbb1c0e6e),
	.w2(32'hbb2b6a7e),
	.w3(32'hba60cf60),
	.w4(32'hba98d310),
	.w5(32'hbaf47db9),
	.w6(32'h39f4fe3e),
	.w7(32'hbb147bc2),
	.w8(32'hba87e5be),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe1747),
	.w1(32'hbae31658),
	.w2(32'hbaf4ac8e),
	.w3(32'hbab13868),
	.w4(32'hbb1b2446),
	.w5(32'hbaffc1e2),
	.w6(32'hba6294f2),
	.w7(32'hbb178567),
	.w8(32'hb810a162),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d2e85),
	.w1(32'hba89becf),
	.w2(32'hbac26eec),
	.w3(32'hbb14bbf1),
	.w4(32'hbb16fcc6),
	.w5(32'h3a378cec),
	.w6(32'hba291ab5),
	.w7(32'hbadf6da1),
	.w8(32'hba3d8382),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dc7c7),
	.w1(32'hbae2b8f5),
	.w2(32'h39890757),
	.w3(32'hba11af1e),
	.w4(32'hbaa40e4a),
	.w5(32'hb9e3ba66),
	.w6(32'h3b43057a),
	.w7(32'h3a81e68e),
	.w8(32'hba5efc13),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e15a3d),
	.w1(32'h3a4a9b53),
	.w2(32'h3a6bfb87),
	.w3(32'h39bc5bf3),
	.w4(32'h3a74b2b0),
	.w5(32'hba3199a1),
	.w6(32'h3ab3a658),
	.w7(32'h3b05316f),
	.w8(32'hba9a452e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b19d09),
	.w1(32'hba06e26f),
	.w2(32'hb97954db),
	.w3(32'hba1cd003),
	.w4(32'hb9064a46),
	.w5(32'hbaa22910),
	.w6(32'hbaa9ea6c),
	.w7(32'hb9f1e2dc),
	.w8(32'h3874ee9a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392301),
	.w1(32'h38af3881),
	.w2(32'hbb42eecb),
	.w3(32'h39db0f7a),
	.w4(32'hb91877f7),
	.w5(32'hba77c2bb),
	.w6(32'hbb2778d3),
	.w7(32'hbb125917),
	.w8(32'hba1de749),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bc330),
	.w1(32'hb99885f9),
	.w2(32'hbaacace7),
	.w3(32'h3a9f6c14),
	.w4(32'h3a910803),
	.w5(32'hbb0df976),
	.w6(32'h3a1abbaf),
	.w7(32'h3a4823c7),
	.w8(32'hbb4ede12),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65e703),
	.w1(32'h3aa6993a),
	.w2(32'hbb127c0f),
	.w3(32'hbb02db48),
	.w4(32'h3a8018a0),
	.w5(32'hbb010f8e),
	.w6(32'hbada3bb9),
	.w7(32'hbae9f83a),
	.w8(32'hbabab0f4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2e95b),
	.w1(32'hba5775a1),
	.w2(32'hbad40b6a),
	.w3(32'hba2b6f2c),
	.w4(32'hba472c7a),
	.w5(32'hbae10cfd),
	.w6(32'h3b6e9856),
	.w7(32'h399dc603),
	.w8(32'hbab2377a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae411fc),
	.w1(32'hba94eb5d),
	.w2(32'hbb229fdd),
	.w3(32'h3a1faa5b),
	.w4(32'h3aeb4dbf),
	.w5(32'hb9fae78d),
	.w6(32'h3b0a2b92),
	.w7(32'h3b29d5cd),
	.w8(32'hb954d965),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9760bd),
	.w1(32'hba7a23e2),
	.w2(32'hbadeeb30),
	.w3(32'hbb181a55),
	.w4(32'hba9735a1),
	.w5(32'hba22439a),
	.w6(32'hbb16c0c5),
	.w7(32'h3a10a80c),
	.w8(32'h3b240084),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a116d6d),
	.w1(32'h3acfef21),
	.w2(32'h3a22e146),
	.w3(32'h3aecaad7),
	.w4(32'h3b0d0b8a),
	.w5(32'h39a1f40b),
	.w6(32'h3b4f7f89),
	.w7(32'hb876cc99),
	.w8(32'hbad046b0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d5971),
	.w1(32'hb98bbc8d),
	.w2(32'hb9da60ad),
	.w3(32'hb86ac9ee),
	.w4(32'hba49cf98),
	.w5(32'h3aef9982),
	.w6(32'h3a3d3c2d),
	.w7(32'hb9e6bdce),
	.w8(32'h3a4e54d4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fe670),
	.w1(32'h3b28fbb9),
	.w2(32'h3b2ea527),
	.w3(32'hbaf3f232),
	.w4(32'hba269f3a),
	.w5(32'h3b1c0ec1),
	.w6(32'h39dd8ae5),
	.w7(32'h3a42f39a),
	.w8(32'h3aaf9b18),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04642a),
	.w1(32'h3b097b18),
	.w2(32'h38ba3f9c),
	.w3(32'h3b168064),
	.w4(32'h3ab78c01),
	.w5(32'hbb2a33d6),
	.w6(32'h3ac89df7),
	.w7(32'h3a2415de),
	.w8(32'hb98ed1fd),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79c017),
	.w1(32'hbb1cbd06),
	.w2(32'hba0ea0ec),
	.w3(32'hbb0601be),
	.w4(32'hbb076261),
	.w5(32'hbaae8ccf),
	.w6(32'hbb01e96d),
	.w7(32'hbaaf695e),
	.w8(32'hbb06fb9d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a6c60),
	.w1(32'h39779f32),
	.w2(32'hba8f07a7),
	.w3(32'hb961935a),
	.w4(32'hbaaa2ebb),
	.w5(32'h37d7ec0c),
	.w6(32'h3a47ceb9),
	.w7(32'hbae285ae),
	.w8(32'h3a535a4a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc3c79),
	.w1(32'hb9d3429b),
	.w2(32'hbaa966ac),
	.w3(32'h3a71924a),
	.w4(32'h3a8883d1),
	.w5(32'hba56c8d3),
	.w6(32'h3a204e25),
	.w7(32'h3a0bbc84),
	.w8(32'hb89fa8bd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b017a),
	.w1(32'h3a6ba50d),
	.w2(32'h37bff5be),
	.w3(32'hb9695a27),
	.w4(32'hb950fd8b),
	.w5(32'h39d8c972),
	.w6(32'hb9e9e739),
	.w7(32'hba5ee486),
	.w8(32'h3a928c2a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1dfae),
	.w1(32'h3b2f7c45),
	.w2(32'h3a6231e1),
	.w3(32'h3b85e731),
	.w4(32'h3b10e729),
	.w5(32'hba980c57),
	.w6(32'h3b2a8bf6),
	.w7(32'hba907c79),
	.w8(32'hbab2eb58),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa848b3),
	.w1(32'hba8d4e3e),
	.w2(32'hbae064cf),
	.w3(32'hb9a3668e),
	.w4(32'hba91399e),
	.w5(32'hb9a076ba),
	.w6(32'h3ae4664c),
	.w7(32'h39505c06),
	.w8(32'hb9e476f5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08a7e7),
	.w1(32'h3928a967),
	.w2(32'hba1f32fa),
	.w3(32'hb94b3db4),
	.w4(32'h39f7181d),
	.w5(32'hbb13d59c),
	.w6(32'h3a269d8c),
	.w7(32'hbaae6b03),
	.w8(32'hba6fd214),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12da65),
	.w1(32'hba050e81),
	.w2(32'h3a5190be),
	.w3(32'hbb0911e8),
	.w4(32'hbb2d4393),
	.w5(32'h3a7b824e),
	.w6(32'hba78e388),
	.w7(32'h3aca8bfc),
	.w8(32'h3b5b09ba),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b358798),
	.w1(32'h3a50d9c6),
	.w2(32'hbaa7ea4e),
	.w3(32'h3a39ad1a),
	.w4(32'hb9246948),
	.w5(32'hbb1d6557),
	.w6(32'hbb88cc40),
	.w7(32'hbada2aba),
	.w8(32'hbb199547),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebf026),
	.w1(32'h3a8fee85),
	.w2(32'hb9776d7a),
	.w3(32'h3a15f1e9),
	.w4(32'h3a15c1ee),
	.w5(32'hb9057083),
	.w6(32'h3b17b1fb),
	.w7(32'h3a81942c),
	.w8(32'h390c59ef),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e40327),
	.w1(32'hba7824dd),
	.w2(32'hbad5c57c),
	.w3(32'hb99ff9e5),
	.w4(32'hba653ee0),
	.w5(32'hbb4d938e),
	.w6(32'h3b228e14),
	.w7(32'h3a80685e),
	.w8(32'hbb818643),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaf5c3),
	.w1(32'hbb352b8d),
	.w2(32'hbac0539e),
	.w3(32'hbb92aa38),
	.w4(32'hbb106fa8),
	.w5(32'hbb830156),
	.w6(32'h3a9f104e),
	.w7(32'hbb432d00),
	.w8(32'hbad109ff),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eeec8),
	.w1(32'hbae1444a),
	.w2(32'hb924ad1f),
	.w3(32'hbb9d978a),
	.w4(32'hbb40dc2a),
	.w5(32'h3a818740),
	.w6(32'hbba8989b),
	.w7(32'hbaedf519),
	.w8(32'hba23011a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba002b8e),
	.w1(32'hb9d43823),
	.w2(32'hbb0f5135),
	.w3(32'h3a2d8092),
	.w4(32'h37b181e1),
	.w5(32'hb9c447b7),
	.w6(32'h3a2791c5),
	.w7(32'hba1a270d),
	.w8(32'hba1f78a5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75f7b7),
	.w1(32'h38dd196f),
	.w2(32'h394079c2),
	.w3(32'h37b6b3bd),
	.w4(32'hb89338c8),
	.w5(32'h3a55e09f),
	.w6(32'hbae8cdca),
	.w7(32'hba24fd10),
	.w8(32'hbb0414b3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928a07c),
	.w1(32'h3a375b42),
	.w2(32'h3aa63435),
	.w3(32'h3af5ce65),
	.w4(32'h3b1ba6ea),
	.w5(32'hb9c9e329),
	.w6(32'h3aae4419),
	.w7(32'h3af6567c),
	.w8(32'h3a0c1d7e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3eb54),
	.w1(32'hbb33a9c5),
	.w2(32'hbb6330d0),
	.w3(32'hbb295140),
	.w4(32'hba8c01d0),
	.w5(32'hb8f910a7),
	.w6(32'hbaa858b9),
	.w7(32'hbac98a41),
	.w8(32'hba7703f1),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cbcee),
	.w1(32'h3912fc1c),
	.w2(32'h3a2efb4e),
	.w3(32'h3a908289),
	.w4(32'h3a15d98d),
	.w5(32'hbad00955),
	.w6(32'h39df1203),
	.w7(32'h39fb4a45),
	.w8(32'hbb53bba4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8b38d),
	.w1(32'hba384c7b),
	.w2(32'hba0af7c1),
	.w3(32'hbaede1dc),
	.w4(32'hbb1cf9b8),
	.w5(32'h3a7d3a26),
	.w6(32'hbaa647ae),
	.w7(32'hba4611e1),
	.w8(32'h3a28e6df),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad7d6c),
	.w1(32'hb7fecce0),
	.w2(32'hb97640d2),
	.w3(32'hb902a9b5),
	.w4(32'h3a72542e),
	.w5(32'hba37225e),
	.w6(32'h3a61da81),
	.w7(32'h39a71af6),
	.w8(32'hba78e161),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054026),
	.w1(32'hba3d2a20),
	.w2(32'hbb330a6a),
	.w3(32'hb9157c0f),
	.w4(32'hba87d951),
	.w5(32'hbacbf719),
	.w6(32'hba91659e),
	.w7(32'hba4663e3),
	.w8(32'hba66cf91),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80d699),
	.w1(32'hba46fa90),
	.w2(32'hbb436914),
	.w3(32'hbb4b38ea),
	.w4(32'hbaf4446e),
	.w5(32'hb9816b9f),
	.w6(32'hbb2bf8ef),
	.w7(32'hbb23c87e),
	.w8(32'hb85358ac),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366d6b43),
	.w1(32'hbaadef0d),
	.w2(32'hb950c9e6),
	.w3(32'h39647671),
	.w4(32'h397026c3),
	.w5(32'h38d567ac),
	.w6(32'h3ab28c22),
	.w7(32'h3ad209f7),
	.w8(32'h3ac84da1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7cf8e),
	.w1(32'h3a605f08),
	.w2(32'h3a2a5a15),
	.w3(32'h3ae565d7),
	.w4(32'h3b05ef49),
	.w5(32'h3a225747),
	.w6(32'h3b05090b),
	.w7(32'h3b0a55c3),
	.w8(32'h3abe4057),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a832cd6),
	.w1(32'h39d9a421),
	.w2(32'h39a184ba),
	.w3(32'h3b0706e4),
	.w4(32'h3b788142),
	.w5(32'hb8d8482e),
	.w6(32'h3afc8f3a),
	.w7(32'hb8119600),
	.w8(32'hbb24f194),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae52606),
	.w1(32'hb98f3f68),
	.w2(32'hba527b43),
	.w3(32'h374aac79),
	.w4(32'h3999e176),
	.w5(32'hba72fee9),
	.w6(32'h3a00f0a9),
	.w7(32'h3a51e5f2),
	.w8(32'hbb2c895d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c1894),
	.w1(32'hb9f99d41),
	.w2(32'hb9e39ba4),
	.w3(32'h3733e0eb),
	.w4(32'h389a5f64),
	.w5(32'hbab283ce),
	.w6(32'h39bad656),
	.w7(32'hb9b6a7cd),
	.w8(32'hbb03737f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea348c),
	.w1(32'hbba5d6b9),
	.w2(32'hbba49b8e),
	.w3(32'h39f39d04),
	.w4(32'hba6407aa),
	.w5(32'hbb5d295f),
	.w6(32'hbbb91bbe),
	.w7(32'hbb4a14a9),
	.w8(32'hbb73d2f1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd89da),
	.w1(32'h3abbed87),
	.w2(32'hba6bf3d2),
	.w3(32'hbabcdfc5),
	.w4(32'h3b31dd86),
	.w5(32'h3810d773),
	.w6(32'h3acddafe),
	.w7(32'h3a538d2a),
	.w8(32'hbad2f5d3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d3466),
	.w1(32'hb8350eb9),
	.w2(32'hbabbb424),
	.w3(32'h3a6156b5),
	.w4(32'hb914a0bb),
	.w5(32'hbb0f2e99),
	.w6(32'h3b26b744),
	.w7(32'hba1c1dbd),
	.w8(32'hbaad3d80),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37793b74),
	.w1(32'hba71baa5),
	.w2(32'hba54cb1c),
	.w3(32'hbb05b19d),
	.w4(32'hba9486fc),
	.w5(32'h391280b7),
	.w6(32'hb9ba648c),
	.w7(32'h370d0e34),
	.w8(32'h398e152a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa32397),
	.w1(32'h3920b50c),
	.w2(32'hba4bfe04),
	.w3(32'h3a586d00),
	.w4(32'h3abeaf4b),
	.w5(32'hba6749ad),
	.w6(32'hb98194a6),
	.w7(32'hb9ae47d3),
	.w8(32'hb922cb68),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888b9dc),
	.w1(32'hbada2346),
	.w2(32'hba20ea6a),
	.w3(32'hb99bbfdf),
	.w4(32'hba9e7e75),
	.w5(32'h3a85bd43),
	.w6(32'h3ab862b3),
	.w7(32'h38daf71d),
	.w8(32'h39742060),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36e96c),
	.w1(32'h39486c47),
	.w2(32'hbad63c31),
	.w3(32'h3b092897),
	.w4(32'hba424514),
	.w5(32'hbaaff2ab),
	.w6(32'h3aa470a7),
	.w7(32'h3a001b18),
	.w8(32'hbb17ba6d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafccc90),
	.w1(32'hbac0a3de),
	.w2(32'hbb79de22),
	.w3(32'h3aaf5742),
	.w4(32'hbb15a16f),
	.w5(32'hbb2754d8),
	.w6(32'h3aae6bcc),
	.w7(32'hbae9b421),
	.w8(32'hbb93766e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60e09d),
	.w1(32'hbb851c47),
	.w2(32'hbb6e3d7f),
	.w3(32'hbb83427d),
	.w4(32'hbb8b8cd3),
	.w5(32'hbaf234d2),
	.w6(32'hbb011b80),
	.w7(32'hbb2347b5),
	.w8(32'h3924dbee),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5c826),
	.w1(32'hbaf5700f),
	.w2(32'hba486f73),
	.w3(32'hb8ea4a46),
	.w4(32'hb9a99480),
	.w5(32'h3a271bd8),
	.w6(32'hba1affa9),
	.w7(32'h3a4cf406),
	.w8(32'h3aab3c2b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46f610),
	.w1(32'h39da56eb),
	.w2(32'hbb51d9ad),
	.w3(32'h38bf58cc),
	.w4(32'hbb0a90b4),
	.w5(32'hbb3bc0bc),
	.w6(32'h3b1bcfae),
	.w7(32'hbb7744ac),
	.w8(32'hbb8205c9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0f93d),
	.w1(32'hb9ff8f06),
	.w2(32'hba4c4702),
	.w3(32'hba11c64f),
	.w4(32'hba63882f),
	.w5(32'hb96b3d60),
	.w6(32'hba02d368),
	.w7(32'h3962e711),
	.w8(32'h3911a299),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98547ee),
	.w1(32'h3aad63a0),
	.w2(32'hb9fb9be9),
	.w3(32'hba180f4d),
	.w4(32'hba2c830d),
	.w5(32'hba4932a2),
	.w6(32'h398f0e77),
	.w7(32'hba6fa356),
	.w8(32'hbb5d688a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05322b),
	.w1(32'hbaebde8b),
	.w2(32'hbb370585),
	.w3(32'hba1d115f),
	.w4(32'h3896623d),
	.w5(32'h3a31d97e),
	.w6(32'hbb69bbf6),
	.w7(32'hba849719),
	.w8(32'h3a0ccc4b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a92127),
	.w1(32'h38a98d05),
	.w2(32'h385e2ddc),
	.w3(32'hb9a23435),
	.w4(32'hb98db879),
	.w5(32'h39c0aa81),
	.w6(32'h3a9d537e),
	.w7(32'hbaafaffa),
	.w8(32'h3ad17620),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c150c7),
	.w1(32'hba117def),
	.w2(32'hbb84a46d),
	.w3(32'h39fc7d50),
	.w4(32'hbb1dd5f2),
	.w5(32'hb9544539),
	.w6(32'h3ade3081),
	.w7(32'hbadfe4b8),
	.w8(32'h399cce5e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971be1f),
	.w1(32'h39f35397),
	.w2(32'hbab5739c),
	.w3(32'h3a370364),
	.w4(32'h39c09911),
	.w5(32'hb9ddb4fe),
	.w6(32'hb99ad0d5),
	.w7(32'hbaabc153),
	.w8(32'h39b61a2c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38629594),
	.w1(32'hba4339eb),
	.w2(32'hbaf556e3),
	.w3(32'hbab33c6f),
	.w4(32'hbaa56025),
	.w5(32'hbb02f183),
	.w6(32'hbb615f17),
	.w7(32'hbaa767e1),
	.w8(32'hba84b73e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed0e0c),
	.w1(32'h3acd5070),
	.w2(32'h3abfe1ee),
	.w3(32'hb9c7f7f9),
	.w4(32'h3798b823),
	.w5(32'h39c76778),
	.w6(32'h39d29ab7),
	.w7(32'h39258743),
	.w8(32'h3a457440),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1b3ff),
	.w1(32'h3a0c63fa),
	.w2(32'h3980e5d2),
	.w3(32'hba8a1b21),
	.w4(32'hba8e3f94),
	.w5(32'hbad343ff),
	.w6(32'hba731fd2),
	.w7(32'h3a4b96e2),
	.w8(32'hbad01811),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb875594d),
	.w1(32'hba97cb84),
	.w2(32'hbb2b5537),
	.w3(32'hbb01232a),
	.w4(32'hbaf2aa83),
	.w5(32'hb9cfe3f0),
	.w6(32'hba6e79f5),
	.w7(32'hbb3ca020),
	.w8(32'hba3be4da),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e170),
	.w1(32'hbb27d3fa),
	.w2(32'hbb55af21),
	.w3(32'hbb50ebd1),
	.w4(32'hbb2a51dd),
	.w5(32'hbb13f889),
	.w6(32'hbb811d7b),
	.w7(32'hba49e06a),
	.w8(32'hbab18203),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dc671),
	.w1(32'hb81acb12),
	.w2(32'hbac5b42c),
	.w3(32'hba960429),
	.w4(32'hbb074ee9),
	.w5(32'hbaf925fe),
	.w6(32'h392477bb),
	.w7(32'hbaff1681),
	.w8(32'hbb0a5d52),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c6aa),
	.w1(32'hbb14b6a0),
	.w2(32'hbaa1329b),
	.w3(32'hbac111b2),
	.w4(32'hba41dfec),
	.w5(32'h3b1f0ccf),
	.w6(32'hbb40748b),
	.w7(32'hba6039ad),
	.w8(32'h3b3ce813),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6ccd5),
	.w1(32'h3ad21a1c),
	.w2(32'hbb04f19a),
	.w3(32'h3bb38c2f),
	.w4(32'h39941a80),
	.w5(32'hba49189f),
	.w6(32'h3bab8d81),
	.w7(32'h3af81752),
	.w8(32'hba0c98ce),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389df9a1),
	.w1(32'hbb12e6b8),
	.w2(32'hbb0ef750),
	.w3(32'hba13d550),
	.w4(32'hba39f281),
	.w5(32'hba6861ae),
	.w6(32'hbb461bf3),
	.w7(32'hba82fdb3),
	.w8(32'hbaf56ec1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35019b),
	.w1(32'h3a1d216d),
	.w2(32'hbaa9dcc3),
	.w3(32'hba8e56f4),
	.w4(32'hba114078),
	.w5(32'hbb34c006),
	.w6(32'hb90a3df6),
	.w7(32'hb97319da),
	.w8(32'hbaf8482f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71eb05),
	.w1(32'hbb0bc2be),
	.w2(32'hbb0a3d6a),
	.w3(32'hba90e057),
	.w4(32'hb9bc0260),
	.w5(32'h3a757aa9),
	.w6(32'h3a57c061),
	.w7(32'hbb0bb158),
	.w8(32'hbac9dc03),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab469c9),
	.w1(32'hbaa7e438),
	.w2(32'hba7e5084),
	.w3(32'h39e42e83),
	.w4(32'hba97d522),
	.w5(32'hbb073505),
	.w6(32'h3a4ba0c3),
	.w7(32'hb89fd45d),
	.w8(32'hbb1cdc83),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09747b),
	.w1(32'hbb3584ac),
	.w2(32'hbb2ae463),
	.w3(32'hbb098b7d),
	.w4(32'hbb0bf392),
	.w5(32'hba830ab4),
	.w6(32'hba6cf786),
	.w7(32'hbb2cc1fa),
	.w8(32'h3979fec9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafb597),
	.w1(32'hb9c6d630),
	.w2(32'hba9f2828),
	.w3(32'h3ae110b8),
	.w4(32'h3ace0151),
	.w5(32'hba4011d5),
	.w6(32'h397493e1),
	.w7(32'h3b36d4d4),
	.w8(32'hba676007),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df6d7f),
	.w1(32'hbb3441e4),
	.w2(32'hbab81abf),
	.w3(32'h3a320975),
	.w4(32'hbb0be6f1),
	.w5(32'hba8df107),
	.w6(32'h39f0baca),
	.w7(32'hbaf864ee),
	.w8(32'hbb631726),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67aebe),
	.w1(32'h3afd3cc6),
	.w2(32'h3ad14160),
	.w3(32'h3b6dbdd6),
	.w4(32'hb9ab3f7a),
	.w5(32'h39e52f2d),
	.w6(32'h3bb06a72),
	.w7(32'h3a841b52),
	.w8(32'hb9a86460),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa6b47),
	.w1(32'h3a4e6298),
	.w2(32'h3b3b7f62),
	.w3(32'h39ab37df),
	.w4(32'h3b2b79fa),
	.w5(32'h3a44d118),
	.w6(32'h3b2b7d7b),
	.w7(32'h3ae68ee6),
	.w8(32'h3ac228be),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae300cd),
	.w1(32'h394c700a),
	.w2(32'hba3a8175),
	.w3(32'hba5c58c3),
	.w4(32'hba6aadb0),
	.w5(32'h3a09dd6a),
	.w6(32'hb9ad0a94),
	.w7(32'hb8cdb664),
	.w8(32'h3a5f87aa),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5196d),
	.w1(32'h39e0ebee),
	.w2(32'h394051ac),
	.w3(32'h39942f95),
	.w4(32'hb89bc4b7),
	.w5(32'h3a33a6f7),
	.w6(32'h39cae8d8),
	.w7(32'h3a0b59d4),
	.w8(32'h3af6db26),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe8280),
	.w1(32'hba18cf9d),
	.w2(32'hbae99658),
	.w3(32'h3aa36c57),
	.w4(32'hb9cf3a77),
	.w5(32'h3a8b54d1),
	.w6(32'h3b547692),
	.w7(32'h3abff4c4),
	.w8(32'h3a80dcc5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd5159),
	.w1(32'h3ab86cca),
	.w2(32'h3afa8b41),
	.w3(32'h3a70a857),
	.w4(32'h39b98f1a),
	.w5(32'hbb47b32c),
	.w6(32'hba7a5ba8),
	.w7(32'h39d5d794),
	.w8(32'hbafd520d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab28138),
	.w1(32'h390b712e),
	.w2(32'h3b192238),
	.w3(32'hbaa6fc48),
	.w4(32'hb9800adf),
	.w5(32'h3c427322),
	.w6(32'hba97a434),
	.w7(32'h3a2df590),
	.w8(32'h3a85f613),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad96118),
	.w1(32'h3af3b7a7),
	.w2(32'h3aec45da),
	.w3(32'h3c57d7a0),
	.w4(32'h3c3d06a8),
	.w5(32'h3ba3887a),
	.w6(32'h3a33d3d8),
	.w7(32'h3bc69ed0),
	.w8(32'hbaf9c0b4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21d244),
	.w1(32'h3b085af7),
	.w2(32'hbc080b86),
	.w3(32'hbc062cbf),
	.w4(32'hbbbaaa88),
	.w5(32'hba873dff),
	.w6(32'hbb640b2b),
	.w7(32'hbbfa90ec),
	.w8(32'hbc460bee),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd37c26),
	.w1(32'hbcb7b573),
	.w2(32'hbc50c3b4),
	.w3(32'h3ca5ab18),
	.w4(32'h3af23c8d),
	.w5(32'hbbf93a3b),
	.w6(32'h3b88b8f4),
	.w7(32'hbbb574e7),
	.w8(32'hb8dd2088),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a984ef6),
	.w1(32'hbb9562e9),
	.w2(32'hbad22745),
	.w3(32'hbc33c969),
	.w4(32'hbbd54e61),
	.w5(32'h3b1f7965),
	.w6(32'hbb026491),
	.w7(32'h3b39b2b6),
	.w8(32'h3b2de2b8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4c6e9),
	.w1(32'hba562758),
	.w2(32'hbaa0f6f3),
	.w3(32'h38c3432e),
	.w4(32'hbb13f030),
	.w5(32'h3a3f2c79),
	.w6(32'h3b5800b2),
	.w7(32'hbb1913fa),
	.w8(32'h3bed663c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d7811),
	.w1(32'h3ac985a9),
	.w2(32'hbae64d64),
	.w3(32'hbaf35fe1),
	.w4(32'hbc469ad5),
	.w5(32'hbbcec1d3),
	.w6(32'hba4e5fc4),
	.w7(32'hbbc67323),
	.w8(32'hbc889dc8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc880a6b),
	.w1(32'hbcb7e9ac),
	.w2(32'hbc5de20c),
	.w3(32'hb7b373a1),
	.w4(32'hbc2e11d4),
	.w5(32'hbb44a11e),
	.w6(32'hbc11d46e),
	.w7(32'hbc801f68),
	.w8(32'h3b4229b6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e6ddc),
	.w1(32'h3c00e8ee),
	.w2(32'h3a8f0ddf),
	.w3(32'hbc50fefa),
	.w4(32'hbc7bf23b),
	.w5(32'h3bae2522),
	.w6(32'hbb2cd294),
	.w7(32'hbbd407ab),
	.w8(32'hbbb6b513),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1e427),
	.w1(32'h3c085af9),
	.w2(32'hbc5a82d3),
	.w3(32'hbb2b35b2),
	.w4(32'hbc26263b),
	.w5(32'hbc023d76),
	.w6(32'hba8a768c),
	.w7(32'hbbebd09f),
	.w8(32'h3b964f1c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b110136),
	.w1(32'h3c0876ae),
	.w2(32'h3ade0bf6),
	.w3(32'hbc8aecbb),
	.w4(32'hbc1908a7),
	.w5(32'h3cc8b245),
	.w6(32'hbafd41d4),
	.w7(32'h39446ef6),
	.w8(32'h3bc5825b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f777),
	.w1(32'h3b452bc1),
	.w2(32'hbb95b03d),
	.w3(32'h3cbe2f9d),
	.w4(32'h3c8f78cc),
	.w5(32'hbbacebef),
	.w6(32'h39f91b21),
	.w7(32'h3b275f3d),
	.w8(32'hba3edb56),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d0222),
	.w1(32'h3c37c976),
	.w2(32'h3c3ac6de),
	.w3(32'hbc216da5),
	.w4(32'hbc3b5132),
	.w5(32'h3c163908),
	.w6(32'h39a8e065),
	.w7(32'h3b4a75d4),
	.w8(32'h3b82558e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5597f5),
	.w1(32'h3c0352b9),
	.w2(32'hbb4f9147),
	.w3(32'h3a7cf809),
	.w4(32'hbc3d6d6a),
	.w5(32'hbb757297),
	.w6(32'h3be5bdae),
	.w7(32'hbbba6ec7),
	.w8(32'hb94dc4d5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a31a7),
	.w1(32'h3b60154b),
	.w2(32'hbbac3a68),
	.w3(32'hbbe6390a),
	.w4(32'h3bdc13cb),
	.w5(32'h3ad3f979),
	.w6(32'h3b07b60d),
	.w7(32'h3bc0adfe),
	.w8(32'h3b844ab0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c464653),
	.w1(32'h3c5ffe53),
	.w2(32'h3c1b412e),
	.w3(32'hb90fd3fe),
	.w4(32'hb806fded),
	.w5(32'h39cf2457),
	.w6(32'h3c1310b4),
	.w7(32'h3b8f4d53),
	.w8(32'h3b15f5f3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850e90),
	.w1(32'hbb9ffcfb),
	.w2(32'hbb473f25),
	.w3(32'h3b1d44b7),
	.w4(32'hbae84cf7),
	.w5(32'hbc71ecd5),
	.w6(32'hba1a1965),
	.w7(32'hbb1bfe2f),
	.w8(32'hbba9ca91),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aa626),
	.w1(32'h3c290329),
	.w2(32'hbbb8a5a6),
	.w3(32'hbc00ba3b),
	.w4(32'h3be10cac),
	.w5(32'hba659e87),
	.w6(32'hbbb4e8f5),
	.w7(32'hb78006ed),
	.w8(32'hbad3ad9d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb0790),
	.w1(32'h3b952272),
	.w2(32'hbb9d9a53),
	.w3(32'hbbd04766),
	.w4(32'hbb913183),
	.w5(32'h3c636826),
	.w6(32'h3ad1b95f),
	.w7(32'h3b108205),
	.w8(32'hbac1a0fc),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8fc79),
	.w1(32'hbb69bcc8),
	.w2(32'h3baf279c),
	.w3(32'h3cce7d27),
	.w4(32'h3cb19287),
	.w5(32'hbc22a98c),
	.w6(32'h3bdfc479),
	.w7(32'h3c5a7887),
	.w8(32'hbc843b70),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84b7ca),
	.w1(32'hbc8cf8e2),
	.w2(32'hbc3a8991),
	.w3(32'hbba90b8e),
	.w4(32'hb9df0bf9),
	.w5(32'h3b9bdbed),
	.w6(32'hbc67a77d),
	.w7(32'hbc48a8d1),
	.w8(32'hbbfc171a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb386955),
	.w1(32'hbbc2ae4a),
	.w2(32'h3bce733d),
	.w3(32'h3bd077c1),
	.w4(32'h3c1d6793),
	.w5(32'h3a1fcdaf),
	.w6(32'hbc352c14),
	.w7(32'hbb1a43d1),
	.w8(32'hba04436b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb534906),
	.w1(32'h3af30ec0),
	.w2(32'hbb765735),
	.w3(32'h3a7526d0),
	.w4(32'hbbc149e4),
	.w5(32'hbb0d42b0),
	.w6(32'hbb0421a6),
	.w7(32'hbc1a1cd7),
	.w8(32'hbbf77f4d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b827177),
	.w1(32'h3b3955d9),
	.w2(32'h3a6d8d87),
	.w3(32'hbaf76723),
	.w4(32'h3a410468),
	.w5(32'h3a6cae53),
	.w6(32'hbbbd8376),
	.w7(32'h3b8fc7be),
	.w8(32'hba9883b6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba834fae),
	.w1(32'h3c607083),
	.w2(32'h3bd39586),
	.w3(32'hbbf73a16),
	.w4(32'hbc2bcb56),
	.w5(32'hbbb31bd2),
	.w6(32'h3acd56fe),
	.w7(32'hbc1d34c9),
	.w8(32'hbb21cf32),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0da93),
	.w1(32'h3a0e00a5),
	.w2(32'h3b177115),
	.w3(32'hbc6336ae),
	.w4(32'hbbbbdacb),
	.w5(32'h3af1b9c7),
	.w6(32'hbc0c604b),
	.w7(32'hbbf0d402),
	.w8(32'hba1d9ed8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e2550),
	.w1(32'h3bc4745f),
	.w2(32'h3ba91df5),
	.w3(32'hbc6379ce),
	.w4(32'hbbee27bf),
	.w5(32'hbb6e7137),
	.w6(32'hbac950fb),
	.w7(32'hbba0c2e0),
	.w8(32'hb9ce1282),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933713d),
	.w1(32'h3b8b6531),
	.w2(32'h3a64af3d),
	.w3(32'hbbee7cf5),
	.w4(32'hbb2cc248),
	.w5(32'h3a82950d),
	.w6(32'hbbc6d6cf),
	.w7(32'hbbe51768),
	.w8(32'h3bad584d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb438a8),
	.w1(32'hbafdd2df),
	.w2(32'hbab2fd0c),
	.w3(32'hbc0fce10),
	.w4(32'h3a32fba1),
	.w5(32'hb8ba584b),
	.w6(32'h3a130f14),
	.w7(32'hbab316ea),
	.w8(32'h3b2d972a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb337c0f),
	.w1(32'h3bedf759),
	.w2(32'h3c151583),
	.w3(32'hbb54dea4),
	.w4(32'hbb27d69c),
	.w5(32'hbc4c0975),
	.w6(32'h3c497f07),
	.w7(32'h3c0911eb),
	.w8(32'hbb2f6dbf),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4720d6),
	.w1(32'h3a10b54e),
	.w2(32'hbb21da87),
	.w3(32'hbb05c0fc),
	.w4(32'h3be3eb61),
	.w5(32'hbc09191b),
	.w6(32'hbb531036),
	.w7(32'h3b07025f),
	.w8(32'h3bc776eb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule