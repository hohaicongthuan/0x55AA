module layer_10_featuremap_33(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0571b),
	.w1(32'h3b775da9),
	.w2(32'h3c979ef5),
	.w3(32'h3b322379),
	.w4(32'h3ad69883),
	.w5(32'h3bb9ee54),
	.w6(32'h3b661d36),
	.w7(32'h3afdbbcc),
	.w8(32'h3b2b0579),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c2270),
	.w1(32'hbb01e8f1),
	.w2(32'h3c781cfb),
	.w3(32'hbcbaaa4e),
	.w4(32'hbbbeb6b8),
	.w5(32'h3c8fec10),
	.w6(32'hbcd5d516),
	.w7(32'hbb26fbe6),
	.w8(32'h3c0663dc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc522479),
	.w1(32'hbbee4e78),
	.w2(32'h3a50b748),
	.w3(32'hbc5046ac),
	.w4(32'hbb3f081c),
	.w5(32'hbaefd555),
	.w6(32'hbc0146f5),
	.w7(32'h3b72ead9),
	.w8(32'hbb6c1b54),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974a2b),
	.w1(32'hb833bec3),
	.w2(32'h3b44e83a),
	.w3(32'hbc6cb7b2),
	.w4(32'h3b8356f9),
	.w5(32'h3c691f44),
	.w6(32'hbbd635bd),
	.w7(32'h3c013d45),
	.w8(32'h3c81dff4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc379c05),
	.w1(32'hbcae2b4c),
	.w2(32'h3c9f2b93),
	.w3(32'hbc17d2ab),
	.w4(32'hbc66537a),
	.w5(32'h3b914cfc),
	.w6(32'hbb2414c9),
	.w7(32'hbc36dbbd),
	.w8(32'h3bd5c3a6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c501c6e),
	.w1(32'h3bf6bad8),
	.w2(32'h3ba630e1),
	.w3(32'h3c231590),
	.w4(32'hbbbfdf93),
	.w5(32'h3b16c3cd),
	.w6(32'hbbdfd4c3),
	.w7(32'hbc0a4620),
	.w8(32'h3ab179e9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a6dbf),
	.w1(32'hbb1493db),
	.w2(32'h39d0722b),
	.w3(32'h3a95a6c7),
	.w4(32'hbb95b205),
	.w5(32'h3ba898e2),
	.w6(32'hb911cec5),
	.w7(32'hbb1ed775),
	.w8(32'h3b8a936c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09f975),
	.w1(32'h3b472384),
	.w2(32'h3a70974d),
	.w3(32'h3c166f9b),
	.w4(32'hbb946dd2),
	.w5(32'hbb9e90a6),
	.w6(32'h3a92ddf6),
	.w7(32'h3b61d639),
	.w8(32'hbbb4025b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987d4c2),
	.w1(32'h3a94548e),
	.w2(32'h3b457d52),
	.w3(32'hbb31f601),
	.w4(32'hba960ff0),
	.w5(32'h3a8b6a63),
	.w6(32'hb8d57be4),
	.w7(32'hbc0040de),
	.w8(32'hba9a9c80),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13cdb9),
	.w1(32'hba9d8a3c),
	.w2(32'hbaffd8b7),
	.w3(32'h3989dd31),
	.w4(32'hbc092076),
	.w5(32'hbb33f150),
	.w6(32'hbc09a302),
	.w7(32'hbc256181),
	.w8(32'hbb0ac339),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a914d3d),
	.w1(32'h3b091bb3),
	.w2(32'h3b979576),
	.w3(32'h39a8fe7d),
	.w4(32'h3aa8de0b),
	.w5(32'hbab87adf),
	.w6(32'h3990ca5f),
	.w7(32'h3a65404d),
	.w8(32'hbb833cb8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11d142),
	.w1(32'hbb3b6952),
	.w2(32'h3b4de56d),
	.w3(32'hbbf6e147),
	.w4(32'h3c223b6e),
	.w5(32'hb9068fed),
	.w6(32'hbc135fba),
	.w7(32'h3bdbb64c),
	.w8(32'hba665e84),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49ab10),
	.w1(32'h3b3c4cb8),
	.w2(32'hbc4268bc),
	.w3(32'h3c3165b9),
	.w4(32'h3a707eb6),
	.w5(32'hbbf36d04),
	.w6(32'h3bd1cd83),
	.w7(32'h3ab72624),
	.w8(32'hbbf8c045),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28e57d),
	.w1(32'hbab60ba8),
	.w2(32'h3c8110b6),
	.w3(32'hb92d7f15),
	.w4(32'hba87f510),
	.w5(32'h3c4e7455),
	.w6(32'h3b75eb6e),
	.w7(32'hbbb73ac6),
	.w8(32'h3a7c4fc1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0890d7),
	.w1(32'hbc342c9b),
	.w2(32'hbad2118e),
	.w3(32'hbc5ff6b5),
	.w4(32'hbbe5fd35),
	.w5(32'h399652a5),
	.w6(32'hbc0a383c),
	.w7(32'h3b995dd9),
	.w8(32'h3b06bfbb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8389be),
	.w1(32'hbb77d8c9),
	.w2(32'h3b0dd2db),
	.w3(32'h3968032a),
	.w4(32'hbc1c01d6),
	.w5(32'h3ae71480),
	.w6(32'h3b16d169),
	.w7(32'hbbc478a2),
	.w8(32'h3aad8740),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d6cc7),
	.w1(32'h3b0e6a48),
	.w2(32'hbb14b4dd),
	.w3(32'h38bb251c),
	.w4(32'h3b0ee94d),
	.w5(32'h3b6b60e9),
	.w6(32'h3a8acc1c),
	.w7(32'h3b042f10),
	.w8(32'hba42e954),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1e2cf),
	.w1(32'hbb286936),
	.w2(32'hbad2d523),
	.w3(32'h3c13d504),
	.w4(32'hb99d24b5),
	.w5(32'hbc1848a0),
	.w6(32'h3bae9a79),
	.w7(32'hba0f43e1),
	.w8(32'hbb379fdf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf398a2),
	.w1(32'h3bdae983),
	.w2(32'hbbd9222c),
	.w3(32'h3bc183bb),
	.w4(32'h3b8557de),
	.w5(32'hbc82d81a),
	.w6(32'h3c29ce4b),
	.w7(32'h3c10cd79),
	.w8(32'hbc3008c1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9763dc),
	.w1(32'hbc44e0d1),
	.w2(32'h3b0c682a),
	.w3(32'hbcb3a55c),
	.w4(32'hbbb502b0),
	.w5(32'h3b956fb4),
	.w6(32'hbc072523),
	.w7(32'hba99e290),
	.w8(32'hba925a92),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba874cef),
	.w1(32'hbbcd066c),
	.w2(32'hbbba32aa),
	.w3(32'hbb23b0ec),
	.w4(32'hbc1fb0cf),
	.w5(32'hbc0c446e),
	.w6(32'hbc06fede),
	.w7(32'hbc08fa58),
	.w8(32'hbaa27a2d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d7f03),
	.w1(32'hba863a56),
	.w2(32'h3b856315),
	.w3(32'hbcc1fe8c),
	.w4(32'h3bfe9189),
	.w5(32'h3b34bbf7),
	.w6(32'hbc700002),
	.w7(32'h3c299d9c),
	.w8(32'h3ba4c7f9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23c993),
	.w1(32'h3b3c7d9d),
	.w2(32'h3bb9fe1d),
	.w3(32'h3b7e9fc6),
	.w4(32'h3ac4b507),
	.w5(32'hbbf0fb6b),
	.w6(32'h3c00f811),
	.w7(32'hbb38bcd3),
	.w8(32'hbbab7253),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca629f),
	.w1(32'hbaa9009c),
	.w2(32'hbbdc7ded),
	.w3(32'h3b6ba4db),
	.w4(32'hbb68221a),
	.w5(32'hbbb7e4fe),
	.w6(32'h3b2bed60),
	.w7(32'hbb3abf61),
	.w8(32'hbbd4f915),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be15666),
	.w1(32'hbab3a77f),
	.w2(32'h3b55658a),
	.w3(32'h3b3f6d0e),
	.w4(32'hbb9fdb4a),
	.w5(32'hbb890689),
	.w6(32'h3bd7a889),
	.w7(32'hbbb32cc7),
	.w8(32'hbc000fb3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca009f2),
	.w1(32'h3a8e242b),
	.w2(32'h3c659c59),
	.w3(32'hbcadd22d),
	.w4(32'h3aed9fcb),
	.w5(32'h3cdcca39),
	.w6(32'hbcaae3d4),
	.w7(32'h3b8897d9),
	.w8(32'h3cf075d1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0d435),
	.w1(32'hbc7edd9e),
	.w2(32'hb9ecd626),
	.w3(32'h3b9756d7),
	.w4(32'hbcd45fc6),
	.w5(32'hba108f04),
	.w6(32'h3c415f75),
	.w7(32'hbc872530),
	.w8(32'h39aa0f8b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa45bb4),
	.w1(32'h3b3fc321),
	.w2(32'h3bfad8a2),
	.w3(32'h3a6e4ec6),
	.w4(32'h3ad74794),
	.w5(32'h3c36f076),
	.w6(32'h3a2ab0fa),
	.w7(32'h3a297cb6),
	.w8(32'h3c4b0444),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34a288),
	.w1(32'h3c124a7c),
	.w2(32'hbb2d8236),
	.w3(32'hba91d2a6),
	.w4(32'hb8759ded),
	.w5(32'hb6e5c79e),
	.w6(32'hbb51bda7),
	.w7(32'hbad3f544),
	.w8(32'h3c30ce0b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4aeea1),
	.w1(32'h3c5759e9),
	.w2(32'hbb26111f),
	.w3(32'h3b4866a2),
	.w4(32'h3b781446),
	.w5(32'hbb713a37),
	.w6(32'hbad8d2ee),
	.w7(32'h3a544f88),
	.w8(32'hb8f849a0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ce0a),
	.w1(32'hbb05653b),
	.w2(32'hbbef4fbf),
	.w3(32'hbb74c7a8),
	.w4(32'hbafa5a1a),
	.w5(32'hbc9140e1),
	.w6(32'h39f348bf),
	.w7(32'h3ade1e04),
	.w8(32'hbc8ff28b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ef58b),
	.w1(32'hbc7c02da),
	.w2(32'h3aab1e3a),
	.w3(32'hbcbdaeef),
	.w4(32'hbc8b3130),
	.w5(32'h3bab5d29),
	.w6(32'hbcaf12e5),
	.w7(32'hbc9c06b4),
	.w8(32'h3ba69453),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e8e9),
	.w1(32'h3aaf0c9b),
	.w2(32'hb9c319fc),
	.w3(32'h3b72f88c),
	.w4(32'h3a985fe6),
	.w5(32'hbb80fbed),
	.w6(32'h3bb9f71c),
	.w7(32'h3b1a527f),
	.w8(32'hbb5cff3f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25f922),
	.w1(32'h3b3d5d3c),
	.w2(32'h3b6b8f7b),
	.w3(32'hbbdef367),
	.w4(32'hbb835d18),
	.w5(32'h3b328a5e),
	.w6(32'hbc1f6da9),
	.w7(32'hbbfdb111),
	.w8(32'hbc74e614),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebb2f4),
	.w1(32'hbc3da5fd),
	.w2(32'h3af916f9),
	.w3(32'hbb39d8d6),
	.w4(32'hbbca1c05),
	.w5(32'hbb1bb513),
	.w6(32'hbbe2ec39),
	.w7(32'hbb99224d),
	.w8(32'hbb636c5a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69eb40),
	.w1(32'hba9aa998),
	.w2(32'hbcab635f),
	.w3(32'hbb403641),
	.w4(32'hbbd696b4),
	.w5(32'hbc1a8153),
	.w6(32'hbc0b8686),
	.w7(32'hbc0c40b3),
	.w8(32'h3aaf8425),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c78e),
	.w1(32'h3b809663),
	.w2(32'h3b685538),
	.w3(32'h3b725e5d),
	.w4(32'h3ad8df04),
	.w5(32'hbb3c08bc),
	.w6(32'h3c88858e),
	.w7(32'h3bfd1922),
	.w8(32'hbbbcff08),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8882b9),
	.w1(32'h3c314e02),
	.w2(32'h3c5df4dc),
	.w3(32'hbc6044a0),
	.w4(32'hbaa82177),
	.w5(32'h3b94ba16),
	.w6(32'hbcb65a35),
	.w7(32'hbc0ecbac),
	.w8(32'hbc30effd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57bfe9),
	.w1(32'h3cbf0443),
	.w2(32'h3c853b10),
	.w3(32'hbbbf4b99),
	.w4(32'h3c412912),
	.w5(32'h3cc9e27d),
	.w6(32'hbcea34b0),
	.w7(32'hbc69a4af),
	.w8(32'h3caa8952),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8beabf8),
	.w1(32'hbb4dcec7),
	.w2(32'hba4f62e7),
	.w3(32'h3c0de5f4),
	.w4(32'hbb814fde),
	.w5(32'h3aa246c7),
	.w6(32'h3c20c516),
	.w7(32'h3bbef648),
	.w8(32'h3b01cd70),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5f0bf),
	.w1(32'h3bb11529),
	.w2(32'h3be46772),
	.w3(32'hbba9fde0),
	.w4(32'h3b09fd6d),
	.w5(32'h3c23bd68),
	.w6(32'hba480f99),
	.w7(32'h3ad181c9),
	.w8(32'h3be4d99b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c420c47),
	.w1(32'h3c191bcd),
	.w2(32'hbc5d9aa4),
	.w3(32'h3cd4c1f3),
	.w4(32'h3cad0f95),
	.w5(32'hbcb72f30),
	.w6(32'h3cb0bb8e),
	.w7(32'h3c56d82a),
	.w8(32'hbc64a341),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8b822),
	.w1(32'hbc7b690d),
	.w2(32'h3b8d0ad1),
	.w3(32'hbccda173),
	.w4(32'hbc94d3e8),
	.w5(32'hba43c537),
	.w6(32'hbcc5dd1e),
	.w7(32'hbc180bfb),
	.w8(32'hbb200d51),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33c772),
	.w1(32'h3b1213ab),
	.w2(32'hbc1cb216),
	.w3(32'h3a58f962),
	.w4(32'hbbab3b28),
	.w5(32'hbb8bd8cb),
	.w6(32'hbbf05df6),
	.w7(32'hbc10b9c3),
	.w8(32'hbb174cdf),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b249f17),
	.w1(32'hbbf3794c),
	.w2(32'hbc2061b0),
	.w3(32'h3b0f5fae),
	.w4(32'h37ac7ffb),
	.w5(32'hbc045221),
	.w6(32'h3c1963a4),
	.w7(32'h3a951e7b),
	.w8(32'hbbfed4bc),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7d986),
	.w1(32'h3b3bb32c),
	.w2(32'h3a9b6b12),
	.w3(32'h3ad23b4c),
	.w4(32'hba8ce031),
	.w5(32'hbb8886a3),
	.w6(32'h3a8ef985),
	.w7(32'hbbb70dda),
	.w8(32'hbba0f19f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b743786),
	.w1(32'h3b80122d),
	.w2(32'h3a8f5738),
	.w3(32'hba9b9aa1),
	.w4(32'h3b8ffcd5),
	.w5(32'hb92d0ede),
	.w6(32'h3b9a6269),
	.w7(32'h3be56e32),
	.w8(32'hbba50211),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bec22),
	.w1(32'h3b160cea),
	.w2(32'hba988b54),
	.w3(32'h3c40a6f9),
	.w4(32'h3c453940),
	.w5(32'hbc37b226),
	.w6(32'h3c7a98be),
	.w7(32'h3c5ef79e),
	.w8(32'hbc5668eb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b469c19),
	.w1(32'h3aabc0d8),
	.w2(32'h3bf652fb),
	.w3(32'hba888306),
	.w4(32'hbb11ad54),
	.w5(32'h3bc5f3e3),
	.w6(32'hbbd5d084),
	.w7(32'hbbadc6f7),
	.w8(32'h3b992d0c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab2e3e),
	.w1(32'h3b11c71d),
	.w2(32'h3c28833b),
	.w3(32'h3b7b6a4d),
	.w4(32'h3bd48a95),
	.w5(32'h3bb30bfa),
	.w6(32'hbbea5003),
	.w7(32'h39853244),
	.w8(32'h3bcfbc4c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e4b14),
	.w1(32'h3c1a5bf6),
	.w2(32'hbbf33db5),
	.w3(32'h3c8357e7),
	.w4(32'h3c262f2c),
	.w5(32'hbbb669d6),
	.w6(32'h3c142848),
	.w7(32'h3bb23126),
	.w8(32'h3b8db38b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b899c8e),
	.w1(32'h3c50b3b4),
	.w2(32'h3bf8a626),
	.w3(32'h3c95887d),
	.w4(32'h3c99930b),
	.w5(32'h3c1a2e68),
	.w6(32'h3cb088c9),
	.w7(32'h3c03bf42),
	.w8(32'h3c25fd49),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4aa8d7),
	.w1(32'h3c0a42aa),
	.w2(32'h3b4438be),
	.w3(32'h3bc70d43),
	.w4(32'h3ba151f8),
	.w5(32'hba94bb09),
	.w6(32'h3c29907f),
	.w7(32'h3c229d21),
	.w8(32'h3b1896ec),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b963352),
	.w1(32'hbaf9990a),
	.w2(32'hbb841e69),
	.w3(32'h3a72f061),
	.w4(32'hbc22c571),
	.w5(32'hbb47891b),
	.w6(32'h3c1a370b),
	.w7(32'hb9bde1c8),
	.w8(32'hbab6cb60),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f723e),
	.w1(32'h3bf6f81b),
	.w2(32'hbbb43904),
	.w3(32'h3c1a33da),
	.w4(32'h3b0be241),
	.w5(32'h3b4c136f),
	.w6(32'h3c4724dd),
	.w7(32'h3c034de6),
	.w8(32'hbaf00c69),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc317a48),
	.w1(32'hbc84a00d),
	.w2(32'h3c2084e8),
	.w3(32'hbc550c37),
	.w4(32'hbc890fc4),
	.w5(32'h3c11f28e),
	.w6(32'hbc72e744),
	.w7(32'hbc18d36f),
	.w8(32'h3bf9862c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b7b3d),
	.w1(32'h3c09a1b3),
	.w2(32'hb98d8f10),
	.w3(32'h3c2cb887),
	.w4(32'h3c4d7f68),
	.w5(32'h3a816f72),
	.w6(32'h3ba0a45e),
	.w7(32'h3ba81751),
	.w8(32'hb9c942ce),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b84fbf),
	.w1(32'hb932a402),
	.w2(32'hbad35643),
	.w3(32'hbb3abe6a),
	.w4(32'hbb942863),
	.w5(32'hbb3591ec),
	.w6(32'h388ff9f6),
	.w7(32'hbbff78c7),
	.w8(32'h3b12913f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dc5c8),
	.w1(32'h3c5cbede),
	.w2(32'h3c0c88f7),
	.w3(32'hbb12228a),
	.w4(32'h3c4ef6c1),
	.w5(32'h3c04447d),
	.w6(32'hbb7e191c),
	.w7(32'h3c118e81),
	.w8(32'h3b96bc2e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9f645),
	.w1(32'h3b78900b),
	.w2(32'h3a313c75),
	.w3(32'h3c83192e),
	.w4(32'h3c0c52fc),
	.w5(32'h3baaa9fd),
	.w6(32'h3b03c534),
	.w7(32'h3ae69979),
	.w8(32'h3c07a231),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c1141),
	.w1(32'hba87a2cf),
	.w2(32'hbc21bce5),
	.w3(32'h3c3f922c),
	.w4(32'h3c386f17),
	.w5(32'hbc9a7b5d),
	.w6(32'h3caa6d7e),
	.w7(32'h3c9ca623),
	.w8(32'hbb80d123),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d1599),
	.w1(32'h3c30b35b),
	.w2(32'h3c4243c9),
	.w3(32'hbb33f815),
	.w4(32'h3b8d07bc),
	.w5(32'h3c092fb5),
	.w6(32'h39e3339f),
	.w7(32'hbbefd1eb),
	.w8(32'h3a233cb6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bc2f5),
	.w1(32'hbaa07fb5),
	.w2(32'h3c00bc11),
	.w3(32'h3bcbe9b6),
	.w4(32'hbb72f491),
	.w5(32'h3bbd1b56),
	.w6(32'h3b86e532),
	.w7(32'h3a46a019),
	.w8(32'h3c0f3ab2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d02c0),
	.w1(32'h3c9e8748),
	.w2(32'hbc21e491),
	.w3(32'h3c8bc947),
	.w4(32'h3c94bfbc),
	.w5(32'hbc82975d),
	.w6(32'h3c28c4f5),
	.w7(32'h3c41929e),
	.w8(32'hbc48d9e5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9df400),
	.w1(32'hbc4f98ff),
	.w2(32'hbb0425d6),
	.w3(32'hbca89bac),
	.w4(32'hbc0b6b7f),
	.w5(32'hbbad9576),
	.w6(32'hbcaac20f),
	.w7(32'hbc3b52e9),
	.w8(32'hbb6fbab0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03ce90),
	.w1(32'h3b893e53),
	.w2(32'h3b9f71a3),
	.w3(32'hbb964b5e),
	.w4(32'hb9a8b561),
	.w5(32'h3b45e0d2),
	.w6(32'hbb3743ad),
	.w7(32'h3b1e7719),
	.w8(32'h3baab33c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ac71a),
	.w1(32'h3bc50f92),
	.w2(32'h3b94f530),
	.w3(32'h3be250ad),
	.w4(32'h3b82f906),
	.w5(32'h39db6eb5),
	.w6(32'h3b9f19eb),
	.w7(32'h3b30ae9e),
	.w8(32'h3b4b13fe),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91c214),
	.w1(32'h3b5d859a),
	.w2(32'hb9ce05bd),
	.w3(32'h3c083dc4),
	.w4(32'h3c39fae9),
	.w5(32'hbb6e767b),
	.w6(32'h3bd36ff3),
	.w7(32'h3b5b9181),
	.w8(32'hbb152d93),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedad5d),
	.w1(32'hbb5a8b74),
	.w2(32'h3b8ee640),
	.w3(32'hbaf0c361),
	.w4(32'hbc204590),
	.w5(32'h3ab52277),
	.w6(32'h3b6fabed),
	.w7(32'hbb50ccfe),
	.w8(32'h3aeecb3d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ab1d2),
	.w1(32'h3c4d85c8),
	.w2(32'hba081ed5),
	.w3(32'h3c42f176),
	.w4(32'h3c27822c),
	.w5(32'hbb60501c),
	.w6(32'h3c637cf5),
	.w7(32'h3c1b81a5),
	.w8(32'hbb6111f7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc021179),
	.w1(32'h3bb06c6f),
	.w2(32'hbba9f773),
	.w3(32'h3ae9f7a4),
	.w4(32'h3c5d8163),
	.w5(32'hba133efe),
	.w6(32'h3bab539f),
	.w7(32'h3c710e12),
	.w8(32'h3b903e31),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe278fd),
	.w1(32'hba86f74f),
	.w2(32'hbbc436c7),
	.w3(32'hbbb1016e),
	.w4(32'hbbb8f9b7),
	.w5(32'hbc2361f1),
	.w6(32'h3ba0581e),
	.w7(32'hbab977b7),
	.w8(32'hbb30cd34),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4bfa3),
	.w1(32'h39b28337),
	.w2(32'hbb209c0d),
	.w3(32'hbbe237b1),
	.w4(32'hbbfd4c1f),
	.w5(32'h3a809f0e),
	.w6(32'hbc23ea87),
	.w7(32'hbbb28dbe),
	.w8(32'h3bab436e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31eadf),
	.w1(32'hbb05c6a8),
	.w2(32'h3a880121),
	.w3(32'hbad7aa96),
	.w4(32'hbc027565),
	.w5(32'hbae12220),
	.w6(32'h3b46be38),
	.w7(32'hbac6dec0),
	.w8(32'hbb1979ba),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca4b5c),
	.w1(32'hbaaaf5d3),
	.w2(32'hb9763fed),
	.w3(32'hbb573e15),
	.w4(32'hbb4786f8),
	.w5(32'hba93a42e),
	.w6(32'hbb76130a),
	.w7(32'hbb3f733b),
	.w8(32'hbb28be78),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06c67c),
	.w1(32'hbc146b01),
	.w2(32'hbc3fd84c),
	.w3(32'hbb93bf73),
	.w4(32'hbc1467d8),
	.w5(32'hbc980f57),
	.w6(32'hbb991d57),
	.w7(32'hbc29b5d2),
	.w8(32'hbc8ed3bb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc083dc0),
	.w1(32'hbc6cd452),
	.w2(32'hbc823469),
	.w3(32'hbcb42024),
	.w4(32'hbcaed6cc),
	.w5(32'hbcc762a2),
	.w6(32'hbc27de56),
	.w7(32'hbbec9e36),
	.w8(32'hbc5f7600),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89f565),
	.w1(32'hbc7a36f9),
	.w2(32'h3bd6f3c7),
	.w3(32'hbd08dfeb),
	.w4(32'hbcbc4806),
	.w5(32'h3ab04df6),
	.w6(32'hbcbdb232),
	.w7(32'hbc8d2a4f),
	.w8(32'hbb8a07eb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86732f9),
	.w1(32'hbaba245d),
	.w2(32'hbb8b56d9),
	.w3(32'h3b86da6b),
	.w4(32'hbb45b758),
	.w5(32'hbb9c9385),
	.w6(32'h3c3e794d),
	.w7(32'h3c398383),
	.w8(32'hbb530037),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb358f8),
	.w1(32'h3a5d073f),
	.w2(32'h3a661396),
	.w3(32'hbbae1215),
	.w4(32'hb913f744),
	.w5(32'h3ad11104),
	.w6(32'hbac0cc8c),
	.w7(32'h3a2bc307),
	.w8(32'hbb099c9e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80298d1),
	.w1(32'h3b526ca2),
	.w2(32'hbc01d414),
	.w3(32'h3ac64ee5),
	.w4(32'h3b99b93b),
	.w5(32'hbc019d80),
	.w6(32'hbb439220),
	.w7(32'hb97771c4),
	.w8(32'hbb38e36a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a8f80),
	.w1(32'hbc0893e8),
	.w2(32'hbb35ab97),
	.w3(32'hbb3ef920),
	.w4(32'hbc07be13),
	.w5(32'hbbbf9a2f),
	.w6(32'hb9a2cbe3),
	.w7(32'hbbddc5f4),
	.w8(32'hbb0e7c16),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf30a39),
	.w1(32'h3bb862dc),
	.w2(32'hba9b2017),
	.w3(32'hba993940),
	.w4(32'hba89c6d0),
	.w5(32'h3a80c59d),
	.w6(32'hb843db14),
	.w7(32'hbb4ca2e2),
	.w8(32'h3be4d9e6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f1378),
	.w1(32'h3c50f509),
	.w2(32'h3b6eefc8),
	.w3(32'h3b2e786d),
	.w4(32'h3c1bc13b),
	.w5(32'h3c5ea68d),
	.w6(32'h3b8bf966),
	.w7(32'hbaba75b7),
	.w8(32'h3c43d64d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2395bc),
	.w1(32'h3c582a6a),
	.w2(32'h3b8efb72),
	.w3(32'h3c6e88f8),
	.w4(32'h3c5aa864),
	.w5(32'h3be4ff95),
	.w6(32'h3c0bd0be),
	.w7(32'h3b32a949),
	.w8(32'h3b48c65c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb030b),
	.w1(32'h3b528df3),
	.w2(32'h3b3587f3),
	.w3(32'h3c24daa3),
	.w4(32'h3b134c69),
	.w5(32'h3b9ed7a7),
	.w6(32'h3bb826f2),
	.w7(32'hbb2e8dc1),
	.w8(32'h3bced8f6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf047d),
	.w1(32'h3b8669eb),
	.w2(32'h3b65c58d),
	.w3(32'hbb9a6170),
	.w4(32'hbb430fa9),
	.w5(32'h3b5aabe4),
	.w6(32'hbbca309b),
	.w7(32'hbab66bbc),
	.w8(32'h3b82c1cb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be0f9e),
	.w1(32'h3b2125bd),
	.w2(32'h3c110f5e),
	.w3(32'h3b25403e),
	.w4(32'h3aded464),
	.w5(32'h3c2de600),
	.w6(32'h3ba38b34),
	.w7(32'h3ae75e13),
	.w8(32'h3bbb78a5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50a113),
	.w1(32'h3bcca3d2),
	.w2(32'hbbc2aaf4),
	.w3(32'h3c7bd522),
	.w4(32'h3bdbbe12),
	.w5(32'hbc569ded),
	.w6(32'h3be55a54),
	.w7(32'h3c2ec7b8),
	.w8(32'hbc1dd7cb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ac3dd),
	.w1(32'hbc78fafe),
	.w2(32'hbba46daf),
	.w3(32'hbcc719a0),
	.w4(32'hbc98c745),
	.w5(32'hbc9aff24),
	.w6(32'hbc340d0e),
	.w7(32'hbbc827b1),
	.w8(32'hbc309923),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef8368),
	.w1(32'h398845e2),
	.w2(32'h3c2c89d4),
	.w3(32'hbc88006f),
	.w4(32'hbbe1d15e),
	.w5(32'h3bd4bc49),
	.w6(32'hbc524e51),
	.w7(32'hbbcff977),
	.w8(32'h3bb18a37),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c609aa3),
	.w1(32'h3ca06cdc),
	.w2(32'hbb292658),
	.w3(32'h3c427903),
	.w4(32'h3c23e3e6),
	.w5(32'hbba95835),
	.w6(32'h3bdaf774),
	.w7(32'h3c3452e6),
	.w8(32'hbb98dcd3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29aa96),
	.w1(32'hbb923630),
	.w2(32'hbaddb653),
	.w3(32'h3a6efb1f),
	.w4(32'hbb118bc8),
	.w5(32'h3af33d9a),
	.w6(32'h3b04d327),
	.w7(32'hbac9f363),
	.w8(32'h3bab07da),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e375d),
	.w1(32'hbb7a7a19),
	.w2(32'hbb04b5eb),
	.w3(32'hba793cf1),
	.w4(32'hbb1471a1),
	.w5(32'hbbed021d),
	.w6(32'h3b62d7e7),
	.w7(32'hb84fe2e0),
	.w8(32'hbbf20a78),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a43b),
	.w1(32'hbb218466),
	.w2(32'h3b51cf1c),
	.w3(32'hbbdefba6),
	.w4(32'hbb20600a),
	.w5(32'hbbf9bd86),
	.w6(32'hbb32e9ef),
	.w7(32'hbbfba758),
	.w8(32'hbc1796d6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f4eb0),
	.w1(32'h3b8c0523),
	.w2(32'h3c0feb92),
	.w3(32'hbc65c64a),
	.w4(32'hbb609cbb),
	.w5(32'h3c8087e8),
	.w6(32'hbc87da38),
	.w7(32'h3a1a327e),
	.w8(32'h3b580e66),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b754e),
	.w1(32'h3a7e7491),
	.w2(32'h3c1db3d2),
	.w3(32'h3c31c284),
	.w4(32'h3bcdc1d5),
	.w5(32'h3c168a5a),
	.w6(32'h3be49b67),
	.w7(32'hbb4c442b),
	.w8(32'h3bf29594),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e0607),
	.w1(32'h3c23d6f9),
	.w2(32'h3b64bcf5),
	.w3(32'h3c46a19b),
	.w4(32'hbb005b46),
	.w5(32'hbc27a646),
	.w6(32'h3c610738),
	.w7(32'h3c04d77e),
	.w8(32'hbb88e944),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c220cee),
	.w1(32'h3c2228d1),
	.w2(32'hba3584d2),
	.w3(32'h3ba8b3f2),
	.w4(32'h3be81e66),
	.w5(32'hbb04da5c),
	.w6(32'h3b1ac53f),
	.w7(32'h3bb1a821),
	.w8(32'h3939ab5f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c98ca),
	.w1(32'h3ad48b6e),
	.w2(32'hbc651ea1),
	.w3(32'h3c3dfc1b),
	.w4(32'hba932a64),
	.w5(32'hbcd6642d),
	.w6(32'h3c0cb936),
	.w7(32'h3aa7ca74),
	.w8(32'hbc7b197d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1314da),
	.w1(32'hbc62ca9b),
	.w2(32'hbb790fed),
	.w3(32'hbd59fdf6),
	.w4(32'hbcbb2efa),
	.w5(32'hbc85909f),
	.w6(32'hbd42e861),
	.w7(32'hbcde808a),
	.w8(32'hbc572047),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0e034),
	.w1(32'hbca61acf),
	.w2(32'h3ac5343c),
	.w3(32'hbd2722f9),
	.w4(32'hbce7d13d),
	.w5(32'hb884c6d3),
	.w6(32'hbd049482),
	.w7(32'hbccb7476),
	.w8(32'hba79624c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f6f50),
	.w1(32'h3a21a076),
	.w2(32'hbbbdb7e8),
	.w3(32'h3c289538),
	.w4(32'hbb1d68e6),
	.w5(32'hbc16eb8a),
	.w6(32'h3be6f1bd),
	.w7(32'hba9c128c),
	.w8(32'hbba71374),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d1675),
	.w1(32'hbb3bf8a8),
	.w2(32'h3af831d6),
	.w3(32'hbc559597),
	.w4(32'hbb95a69b),
	.w5(32'hbb24bf4a),
	.w6(32'hbc223281),
	.w7(32'hbbc2ac5d),
	.w8(32'hbb7bcbd6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b729f69),
	.w1(32'h3b5786e4),
	.w2(32'hb7ad50d2),
	.w3(32'h3c59bb56),
	.w4(32'h3bd269dc),
	.w5(32'h3b294eb2),
	.w6(32'h3c71c47a),
	.w7(32'h3c233935),
	.w8(32'h3bde0195),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5e9d),
	.w1(32'h3c0e6375),
	.w2(32'h3a952d9a),
	.w3(32'h3c21b3db),
	.w4(32'h3b49f1f2),
	.w5(32'h3bc62c7d),
	.w6(32'h3c30d3d0),
	.w7(32'h3ba552f2),
	.w8(32'h3bd04248),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7526ca),
	.w1(32'h3b4913fd),
	.w2(32'h3b0d0127),
	.w3(32'hbac5086a),
	.w4(32'h3aa53836),
	.w5(32'h3b2db8cf),
	.w6(32'hba87e1ca),
	.w7(32'h3b0beed6),
	.w8(32'h3b291bb1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fb210),
	.w1(32'h3aad98af),
	.w2(32'h3b8e2af4),
	.w3(32'h3c1dec27),
	.w4(32'h398460cc),
	.w5(32'h3b016e86),
	.w6(32'h3c3b348c),
	.w7(32'h3bdc591d),
	.w8(32'h3bfb6123),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75842e),
	.w1(32'h3c1e965b),
	.w2(32'hbb40ee4d),
	.w3(32'h3c8401cb),
	.w4(32'h3be1090d),
	.w5(32'hbb03c56b),
	.w6(32'h3c1a45a3),
	.w7(32'h3b3ab327),
	.w8(32'hbba05503),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b202b05),
	.w1(32'hbc0629c2),
	.w2(32'hbac76e6d),
	.w3(32'hbc375789),
	.w4(32'hbc15f6cd),
	.w5(32'hbc6e8743),
	.w6(32'hbc5e6620),
	.w7(32'hbbc8a9c3),
	.w8(32'hbba26637),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306c34),
	.w1(32'hbc2be344),
	.w2(32'h39b47271),
	.w3(32'hbc6d3693),
	.w4(32'hbc8c91ab),
	.w5(32'hbbcf84ef),
	.w6(32'hbc2fbcf2),
	.w7(32'hbc48e26e),
	.w8(32'hbc05afed),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6feb2),
	.w1(32'hbc92deac),
	.w2(32'hb879172e),
	.w3(32'hbc0e2d9e),
	.w4(32'hbbaa0097),
	.w5(32'h3c474438),
	.w6(32'hbc537982),
	.w7(32'hbae38454),
	.w8(32'h3c18a5dd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9090e),
	.w1(32'h3b2c4383),
	.w2(32'hbb4490c3),
	.w3(32'h3c1bec8c),
	.w4(32'h3bd3e3c5),
	.w5(32'hbb79a0ea),
	.w6(32'h3bcc3e8d),
	.w7(32'h3b4c2444),
	.w8(32'hbbeba669),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc325c6f),
	.w1(32'hbc4c235a),
	.w2(32'h3af74a1e),
	.w3(32'hbb9c0d0c),
	.w4(32'hbbd5bc7a),
	.w5(32'h3b153e39),
	.w6(32'hbb94a3a4),
	.w7(32'hbb94dab2),
	.w8(32'h3c0751d5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27cd20),
	.w1(32'h3bafb9f4),
	.w2(32'h3b3a22ce),
	.w3(32'h3c7324a1),
	.w4(32'h3c8f3260),
	.w5(32'h3bbe1f3f),
	.w6(32'h3c953e6e),
	.w7(32'h3c9ca11d),
	.w8(32'h3b88ffed),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb91beb),
	.w1(32'h3a8916d1),
	.w2(32'hbbcefedf),
	.w3(32'h3c15551c),
	.w4(32'h3bb2960f),
	.w5(32'hbc5b8677),
	.w6(32'h3bc03929),
	.w7(32'h3b99f31e),
	.w8(32'hbb8a0ac8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc344f2f),
	.w1(32'h3b233c14),
	.w2(32'h3c34b9a7),
	.w3(32'hbc7c981d),
	.w4(32'hbc15c569),
	.w5(32'h3c22647a),
	.w6(32'h3a02f899),
	.w7(32'hb7f536c4),
	.w8(32'h3c1f4176),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07dbb5),
	.w1(32'h3bcee04a),
	.w2(32'h3b0221e0),
	.w3(32'h3c6248ba),
	.w4(32'h3c52ecc3),
	.w5(32'hbc4b246c),
	.w6(32'h3beb16b9),
	.w7(32'h3c038132),
	.w8(32'hbc71dff3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc353705),
	.w1(32'hbc60eeb4),
	.w2(32'hbc0e3eb7),
	.w3(32'hbcbfbe03),
	.w4(32'hbc94fb72),
	.w5(32'hbca5748f),
	.w6(32'hbcc8ee04),
	.w7(32'hbce04345),
	.w8(32'hbc69495e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca96925),
	.w1(32'hbc824c2d),
	.w2(32'hbb09c17e),
	.w3(32'hbd12c6bc),
	.w4(32'hbcd6988e),
	.w5(32'hbb58075b),
	.w6(32'hbcd1f647),
	.w7(32'hbc8d3ae6),
	.w8(32'h3ab8893a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc3697),
	.w1(32'hbb57a7b7),
	.w2(32'hba3353f5),
	.w3(32'hbbc0b896),
	.w4(32'hbbb175d3),
	.w5(32'h38f0a8d5),
	.w6(32'hbb2ee216),
	.w7(32'hbb722ed3),
	.w8(32'hb8439e31),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa351d9),
	.w1(32'h3a1bd2f2),
	.w2(32'hbad1df5b),
	.w3(32'h3abd02ba),
	.w4(32'h3afc7406),
	.w5(32'hbb0a0e38),
	.w6(32'h3afd323e),
	.w7(32'h3b54adda),
	.w8(32'h39e84096),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1aee0),
	.w1(32'hbb136946),
	.w2(32'h3b10cfd9),
	.w3(32'hbb849ae8),
	.w4(32'hba8a42f2),
	.w5(32'h3c4ed249),
	.w6(32'hbafcca21),
	.w7(32'hbb26ddc3),
	.w8(32'h3c75341c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b112f8e),
	.w1(32'h3c36a335),
	.w2(32'h3bd6b3aa),
	.w3(32'h3bb0f477),
	.w4(32'h396e95e3),
	.w5(32'h3c2a3108),
	.w6(32'hb7cad561),
	.w7(32'hbbed09a8),
	.w8(32'h3c1e5e67),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d22d0),
	.w1(32'h3b560462),
	.w2(32'h3b6d0a1c),
	.w3(32'h3bfc23eb),
	.w4(32'h3b51fcbb),
	.w5(32'h3c205693),
	.w6(32'h3c03db0f),
	.w7(32'h3bc71601),
	.w8(32'h3bf4c5ab),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23ad04),
	.w1(32'h3bedc1fa),
	.w2(32'hbc59aea9),
	.w3(32'h3c1a8e82),
	.w4(32'h3be96553),
	.w5(32'hbbc3bbb2),
	.w6(32'h3c0ca5cf),
	.w7(32'hbb6596c0),
	.w8(32'hbafc4bf9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb757457),
	.w1(32'h3b0ac465),
	.w2(32'hbb2e1008),
	.w3(32'hbc095c22),
	.w4(32'h3b04d07f),
	.w5(32'hbb84ba25),
	.w6(32'hba3cb040),
	.w7(32'h39ca8158),
	.w8(32'hbbc7fd19),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03d5e3),
	.w1(32'h3ba2a218),
	.w2(32'hbce5ae5c),
	.w3(32'hbc12d92c),
	.w4(32'h3a9aed6b),
	.w5(32'hbc81f91e),
	.w6(32'hbb4d8e5e),
	.w7(32'hbb00941c),
	.w8(32'hbbe86ece),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc943e11),
	.w1(32'hbb914620),
	.w2(32'hb72fe9e6),
	.w3(32'hbc2c9030),
	.w4(32'hbac077ef),
	.w5(32'hbba3c9c0),
	.w6(32'h3c081602),
	.w7(32'hbba7d3c0),
	.w8(32'hbaede821),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab83429),
	.w1(32'hba135fb9),
	.w2(32'hbb319cf1),
	.w3(32'h39a5b156),
	.w4(32'h3b3d826a),
	.w5(32'hb9b18fb5),
	.w6(32'hbac0a571),
	.w7(32'h3a5392d3),
	.w8(32'hb9b0d8c1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc469cc),
	.w1(32'h3c00452e),
	.w2(32'hbc182c52),
	.w3(32'hbbf32ac7),
	.w4(32'hbbb4b097),
	.w5(32'hbc69c151),
	.w6(32'hbac49b3a),
	.w7(32'hba8afffa),
	.w8(32'hbbb5fb4c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8901c3),
	.w1(32'hbc38ad46),
	.w2(32'hb99f4307),
	.w3(32'hbcb553e8),
	.w4(32'hbc9b16d0),
	.w5(32'hbc02c898),
	.w6(32'hbcaf0ac9),
	.w7(32'hbc935d9d),
	.w8(32'hbc34afed),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a5a68),
	.w1(32'hbc4aad65),
	.w2(32'hbc44efb6),
	.w3(32'hbc9ce35d),
	.w4(32'hbcad4261),
	.w5(32'hbc406188),
	.w6(32'hbc97eaa3),
	.w7(32'hbc74988e),
	.w8(32'hbc008738),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839134),
	.w1(32'hba56cd56),
	.w2(32'hbba881b8),
	.w3(32'hbbcffa6d),
	.w4(32'hbbc4e053),
	.w5(32'hbbd92f3a),
	.w6(32'hbb606fe0),
	.w7(32'hbbb04cf0),
	.w8(32'hbb35d0b0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4aaad),
	.w1(32'hba88692f),
	.w2(32'h3bfafd41),
	.w3(32'h3bad0bfc),
	.w4(32'hbb769e09),
	.w5(32'hbb835cf5),
	.w6(32'h3be5f65e),
	.w7(32'hba2c5dd6),
	.w8(32'h3a708093),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c113035),
	.w1(32'h3c61e375),
	.w2(32'hbb5b6720),
	.w3(32'h3b758cf9),
	.w4(32'h3c1920ae),
	.w5(32'hbb2f3916),
	.w6(32'hbb4a3972),
	.w7(32'h3bb3c456),
	.w8(32'hbb166f15),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a5a9f),
	.w1(32'hba6a153d),
	.w2(32'h3b7af673),
	.w3(32'hbc54c35b),
	.w4(32'hbbac8440),
	.w5(32'h3b20a916),
	.w6(32'hbb54aa59),
	.w7(32'h3b383fcb),
	.w8(32'h3995110d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36216c),
	.w1(32'h3b8bc4a1),
	.w2(32'hbbf210de),
	.w3(32'h3b443b4e),
	.w4(32'hbb791784),
	.w5(32'hbc104004),
	.w6(32'h3b7e5b11),
	.w7(32'hbb49f403),
	.w8(32'hbbc72406),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf90c),
	.w1(32'hbac1ea96),
	.w2(32'hbc1c949f),
	.w3(32'hba57b65d),
	.w4(32'h38ac4321),
	.w5(32'hbc2a188b),
	.w6(32'h3b1c87d6),
	.w7(32'h3a9f661a),
	.w8(32'hbc055ceb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85e437),
	.w1(32'hbbf8e360),
	.w2(32'hba914668),
	.w3(32'hbcc98b9a),
	.w4(32'hbc8e7a3d),
	.w5(32'hbb162ad1),
	.w6(32'hbc9769ca),
	.w7(32'hbc6d554e),
	.w8(32'hbb432dfb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2022c1),
	.w1(32'hbb817799),
	.w2(32'h3bf48bbd),
	.w3(32'hba523c65),
	.w4(32'hbb830ea0),
	.w5(32'h3bb72e5c),
	.w6(32'h3a4ce700),
	.w7(32'hbb1aba30),
	.w8(32'h3bdc488e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cce3871),
	.w1(32'h3c53877a),
	.w2(32'hbbdf7cf9),
	.w3(32'h3c640a99),
	.w4(32'h3c288f95),
	.w5(32'h3bb2e2ad),
	.w6(32'h3c10b421),
	.w7(32'h3c3e8eb9),
	.w8(32'h3b1f1612),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9daf7a),
	.w1(32'h3b2f0431),
	.w2(32'h3c12398a),
	.w3(32'h3b2a546b),
	.w4(32'h3b722425),
	.w5(32'h3b9c2be3),
	.w6(32'h3b60b47e),
	.w7(32'h3b887ce5),
	.w8(32'h3ba785f2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc65d7b),
	.w1(32'h3bd54188),
	.w2(32'hbae4c9c8),
	.w3(32'h3c0ac0ef),
	.w4(32'h3c442f86),
	.w5(32'h3a75a879),
	.w6(32'h3b9f6984),
	.w7(32'h3c13a8e1),
	.w8(32'h3b9aeb95),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48db6b),
	.w1(32'hbac4f8e9),
	.w2(32'h3baf127c),
	.w3(32'h3b0e8972),
	.w4(32'h3a8535f6),
	.w5(32'h3bbd47f0),
	.w6(32'h3be217e1),
	.w7(32'h3b90a46d),
	.w8(32'h3be64f4e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57910d),
	.w1(32'h3b9a32b5),
	.w2(32'h3c2b694b),
	.w3(32'h3bc489a1),
	.w4(32'h3bf46df2),
	.w5(32'h3c04c8e1),
	.w6(32'h3b089484),
	.w7(32'h3c179bd4),
	.w8(32'h3c1899ee),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57f2e0),
	.w1(32'h3c8e7005),
	.w2(32'h3c2dc8f3),
	.w3(32'h3c59e107),
	.w4(32'h3c44e8c4),
	.w5(32'h3c3a60e6),
	.w6(32'h3c4fd4de),
	.w7(32'h3c550681),
	.w8(32'h3beddcd4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bac67),
	.w1(32'h3c20f237),
	.w2(32'hbc18caa6),
	.w3(32'h3cad8a9c),
	.w4(32'h3902b166),
	.w5(32'hbc2375b6),
	.w6(32'h3c1f0b6c),
	.w7(32'h3c328334),
	.w8(32'hbbefbc98),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ee34),
	.w1(32'hbc05d6e9),
	.w2(32'h3c2a9c34),
	.w3(32'hbc0fc85c),
	.w4(32'hbbc909e9),
	.w5(32'h3c06c782),
	.w6(32'hbbb50511),
	.w7(32'hbb24b478),
	.w8(32'h3c2ce817),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e57c8),
	.w1(32'h3bf53cd1),
	.w2(32'hbc33388d),
	.w3(32'h3cb34249),
	.w4(32'h3ba29e01),
	.w5(32'hbc44c0a3),
	.w6(32'h3c26661a),
	.w7(32'h3b8bb133),
	.w8(32'hbbd3b806),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77893b),
	.w1(32'hbc33da04),
	.w2(32'hbb0baefc),
	.w3(32'hbbc5e040),
	.w4(32'hbc16bcf2),
	.w5(32'hbb7b7e2b),
	.w6(32'hbb8ff42f),
	.w7(32'hbc3143d3),
	.w8(32'hbb95930f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68cbb5),
	.w1(32'h3af41f54),
	.w2(32'h3c21a7aa),
	.w3(32'h3a4c7290),
	.w4(32'hbad81045),
	.w5(32'hbb85938f),
	.w6(32'h3ac49d86),
	.w7(32'hba31e57a),
	.w8(32'h3c02d7c2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbffab6),
	.w1(32'h3c6cafcb),
	.w2(32'h38ab8498),
	.w3(32'h3cb26630),
	.w4(32'h3be85685),
	.w5(32'hb99d8c1e),
	.w6(32'h3c5e5a2a),
	.w7(32'h3c2632cd),
	.w8(32'hbbd27e50),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5faf),
	.w1(32'hbbf91b22),
	.w2(32'hbb605273),
	.w3(32'hbc181500),
	.w4(32'hbc19e444),
	.w5(32'hbc955dd6),
	.w6(32'hbc82d996),
	.w7(32'hbc616f4e),
	.w8(32'hbc3584ad),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fc412),
	.w1(32'hbca91efa),
	.w2(32'h3a5fa8fb),
	.w3(32'hbd031190),
	.w4(32'hbcc17b5d),
	.w5(32'hbb434eae),
	.w6(32'hbcc28ac0),
	.w7(32'hbbd40ef1),
	.w8(32'hbaeec912),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93ae76),
	.w1(32'hb9906e40),
	.w2(32'h3b4b5ec6),
	.w3(32'hbc9b4fed),
	.w4(32'hbbf1fd39),
	.w5(32'h3b447071),
	.w6(32'hbc414d49),
	.w7(32'hbbba4c40),
	.w8(32'h3b4fd4e2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afad6e9),
	.w1(32'hbae124b3),
	.w2(32'h39769cde),
	.w3(32'h3bdc539c),
	.w4(32'h3acc1bf2),
	.w5(32'hbbb56bc0),
	.w6(32'h3b85852e),
	.w7(32'hbb4d4228),
	.w8(32'h3b13c8b7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1720b8),
	.w1(32'h3ba68c5b),
	.w2(32'hbc846197),
	.w3(32'hbbbd80e9),
	.w4(32'hbb955f2f),
	.w5(32'hbc434e14),
	.w6(32'h3bc11e01),
	.w7(32'h3b0068ea),
	.w8(32'hbc9462c2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ae61d),
	.w1(32'hbc85df84),
	.w2(32'hb9fc5bcf),
	.w3(32'hbbffedd8),
	.w4(32'hbc45888c),
	.w5(32'h3bac96e7),
	.w6(32'hbc6aaa68),
	.w7(32'hbc9f0a83),
	.w8(32'h3bac5a65),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399911e0),
	.w1(32'h3baeca21),
	.w2(32'hbb218079),
	.w3(32'h3bce22dd),
	.w4(32'h3bc089ea),
	.w5(32'h3ba9c8e0),
	.w6(32'h3be3773f),
	.w7(32'h3bee9192),
	.w8(32'h3c832302),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee75ec),
	.w1(32'h3a0bf2a2),
	.w2(32'hbc84c4e1),
	.w3(32'h3b481d3e),
	.w4(32'h3bb0eaa2),
	.w5(32'hbb6e7de5),
	.w6(32'h3c5ed3f8),
	.w7(32'h3bcf3b67),
	.w8(32'hbbe9a9e0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b27e),
	.w1(32'hbc4b9c84),
	.w2(32'h3c230755),
	.w3(32'h3ca0c546),
	.w4(32'h3bef1eab),
	.w5(32'h3b9c4d2c),
	.w6(32'h3c554bc4),
	.w7(32'hba35f722),
	.w8(32'h3a8ba591),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8a62b),
	.w1(32'h3aa823b2),
	.w2(32'hbbdd707e),
	.w3(32'h3b8a2292),
	.w4(32'h3b7179b7),
	.w5(32'hbbcd9c7c),
	.w6(32'h3b4e5323),
	.w7(32'h3aa67a2b),
	.w8(32'hbb214e1e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641f8b),
	.w1(32'hbb4d7805),
	.w2(32'hbb8c41ad),
	.w3(32'hbb38241a),
	.w4(32'hbb6e3bab),
	.w5(32'hbb700911),
	.w6(32'h37737266),
	.w7(32'h3b1cc6ca),
	.w8(32'h3bf5f6b4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a2d4a),
	.w1(32'hbb17d117),
	.w2(32'hbd204395),
	.w3(32'hbaf55e08),
	.w4(32'hbb2e4bdf),
	.w5(32'hbc9c2607),
	.w6(32'h3bc09a59),
	.w7(32'h3b24d8db),
	.w8(32'hbcc222db),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc931758),
	.w1(32'hbcdae1dc),
	.w2(32'hba57ef64),
	.w3(32'h3c0724e0),
	.w4(32'hbb92e9b1),
	.w5(32'hba16c0b6),
	.w6(32'h3a46b017),
	.w7(32'hbc4f3618),
	.w8(32'h3b5ddd3e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6d1d1),
	.w1(32'h3bccaa11),
	.w2(32'h3b1ef6f4),
	.w3(32'h3b907a25),
	.w4(32'h3b25420d),
	.w5(32'h3bc45416),
	.w6(32'h3bb6368d),
	.w7(32'h3c0cb09b),
	.w8(32'h3bc335aa),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba78db8),
	.w1(32'h3a8bafa6),
	.w2(32'h3b65b91f),
	.w3(32'h3b5cd39d),
	.w4(32'hb9976d0d),
	.w5(32'h3b9ce94f),
	.w6(32'h3ae69106),
	.w7(32'hb9d0b4dd),
	.w8(32'h3bb23994),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4836b),
	.w1(32'h3bf7d9b8),
	.w2(32'hba12a6f3),
	.w3(32'h3c0d4c7a),
	.w4(32'h3b5a6451),
	.w5(32'hbb7072ba),
	.w6(32'h3be47bb4),
	.w7(32'h3a5fe394),
	.w8(32'h3958198d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb979665e),
	.w1(32'h3b153407),
	.w2(32'h3c2e61ed),
	.w3(32'hb91f1550),
	.w4(32'hbaced2d4),
	.w5(32'h3c307877),
	.w6(32'h3bb90137),
	.w7(32'h3b29e1f8),
	.w8(32'h3bce67fd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c351ae6),
	.w1(32'h3c033eb8),
	.w2(32'hbc69343a),
	.w3(32'h3c567564),
	.w4(32'h3be2fcac),
	.w5(32'hbcf5024c),
	.w6(32'h3bcfa644),
	.w7(32'h3b111fa6),
	.w8(32'hbc9b722c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0ca26),
	.w1(32'hbc6090ac),
	.w2(32'h3ab983c8),
	.w3(32'hbd544a15),
	.w4(32'hbd1697dd),
	.w5(32'hb9c9d77e),
	.w6(32'hbd1c50f2),
	.w7(32'hbcb495f8),
	.w8(32'hbb5699e0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ef83a),
	.w1(32'h3b346eaf),
	.w2(32'h3b0251c8),
	.w3(32'h3c2ba460),
	.w4(32'h3ae6f634),
	.w5(32'hbb8b7c23),
	.w6(32'h3ba118b8),
	.w7(32'h3a9aeba1),
	.w8(32'hbbd289fa),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc81acb),
	.w1(32'h3b820dfa),
	.w2(32'h3b86ad4b),
	.w3(32'hbb7d99e0),
	.w4(32'hba82008a),
	.w5(32'h3ac40d14),
	.w6(32'hbbb86391),
	.w7(32'h3a2ff7bb),
	.w8(32'hbb425b68),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f5bfe),
	.w1(32'h3bf690d7),
	.w2(32'h3b9e0068),
	.w3(32'h3c197789),
	.w4(32'h3b77de59),
	.w5(32'hbb3f096c),
	.w6(32'h3bf57e85),
	.w7(32'h3bdf7019),
	.w8(32'h399411bc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f50c6),
	.w1(32'h3bce5479),
	.w2(32'hbb51ef40),
	.w3(32'h3beece57),
	.w4(32'hba83a18b),
	.w5(32'hbbc96f80),
	.w6(32'h3c65574d),
	.w7(32'hbb7d104c),
	.w8(32'hba24feca),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6529),
	.w1(32'hbbac4723),
	.w2(32'hbbfb4830),
	.w3(32'hbc0f02ff),
	.w4(32'hbc012b3c),
	.w5(32'hbc0b8dbc),
	.w6(32'hbb238584),
	.w7(32'hba66d37b),
	.w8(32'hbc11dada),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22a4ec),
	.w1(32'hbbf5e6f8),
	.w2(32'hbb03cd4c),
	.w3(32'hbc50870f),
	.w4(32'hbbadb6bf),
	.w5(32'h39c1760c),
	.w6(32'hbc128fb0),
	.w7(32'hbba913f4),
	.w8(32'h3baf1e2c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b472181),
	.w1(32'h3ab40467),
	.w2(32'h3b2c00b1),
	.w3(32'h3b0d7b8f),
	.w4(32'h39943f53),
	.w5(32'h3b9294d3),
	.w6(32'h3b70ad39),
	.w7(32'h3a880a60),
	.w8(32'hba9e2302),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad382),
	.w1(32'h3b0c64d3),
	.w2(32'h3858d77d),
	.w3(32'h3b96334d),
	.w4(32'h3b15b0ff),
	.w5(32'hbb22f8c9),
	.w6(32'hbbc0d49b),
	.w7(32'hbb60f667),
	.w8(32'h3a4577cb),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ed0b0),
	.w1(32'h3b792f62),
	.w2(32'h3b5f0fa1),
	.w3(32'hbae246c0),
	.w4(32'hbb92e3bf),
	.w5(32'h3bbee616),
	.w6(32'hbad9870b),
	.w7(32'hbb6a5d77),
	.w8(32'h399be55c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacfaf8),
	.w1(32'h3c20eb75),
	.w2(32'hbc221fb4),
	.w3(32'h3c1c91a9),
	.w4(32'h3c32e331),
	.w5(32'hbc6b0538),
	.w6(32'h3b11a999),
	.w7(32'h3b0e2136),
	.w8(32'hbc42cf3e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22d15a),
	.w1(32'hbb5cbe3c),
	.w2(32'h3aa68b92),
	.w3(32'hbc88e63e),
	.w4(32'hbc2bcb2b),
	.w5(32'hbaed9283),
	.w6(32'hbc65fe27),
	.w7(32'hbbdb24bf),
	.w8(32'hbb4e6596),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87101f),
	.w1(32'h3aa87c79),
	.w2(32'h3aff59c1),
	.w3(32'hbb012efa),
	.w4(32'h390184ab),
	.w5(32'h3bcaed61),
	.w6(32'hbb8135e1),
	.w7(32'h3b5e1071),
	.w8(32'h3bde7d8c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9168a0),
	.w1(32'h3b39e7c5),
	.w2(32'hbc11bfad),
	.w3(32'hba3ab4c4),
	.w4(32'hbb07d66a),
	.w5(32'hbbf20dcd),
	.w6(32'h3bb4ffc5),
	.w7(32'hbbabcd6b),
	.w8(32'hbb913aaf),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827413),
	.w1(32'h3c375939),
	.w2(32'hbaa111cf),
	.w3(32'hbb6d6e4a),
	.w4(32'h3c2864b9),
	.w5(32'h393fc667),
	.w6(32'h39f50933),
	.w7(32'h3c591a03),
	.w8(32'h3a8f7460),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc74f6),
	.w1(32'h3a37fa7b),
	.w2(32'hbba815bf),
	.w3(32'h39d63cea),
	.w4(32'hbb5e100c),
	.w5(32'h395c8b42),
	.w6(32'hba79c4fa),
	.w7(32'hbbbe756c),
	.w8(32'h3ba1d38e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa5603),
	.w1(32'h3c342257),
	.w2(32'hbc22dc3b),
	.w3(32'h3ccdfdae),
	.w4(32'h3c310510),
	.w5(32'hbc2ec08c),
	.w6(32'h3cb80730),
	.w7(32'h3ca356ba),
	.w8(32'hbc19bb31),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a397a99),
	.w1(32'h3c03f83f),
	.w2(32'h3bc89286),
	.w3(32'hba8b3376),
	.w4(32'h3bc02efc),
	.w5(32'h3a4f7cc2),
	.w6(32'hbaf96e8f),
	.w7(32'h3a3bb9f0),
	.w8(32'hba548a28),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b853508),
	.w1(32'h3bce4543),
	.w2(32'hbb03d12d),
	.w3(32'h3b2cc983),
	.w4(32'h3b454f7f),
	.w5(32'hbb38b96f),
	.w6(32'hbaa6dea3),
	.w7(32'h3b9c4e52),
	.w8(32'hbbb00618),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64404d),
	.w1(32'hba13b90d),
	.w2(32'h3aa3600d),
	.w3(32'hba3d4a79),
	.w4(32'hbade0c3e),
	.w5(32'h3a8cd845),
	.w6(32'h394f95e3),
	.w7(32'hba095f80),
	.w8(32'h3b888821),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b563b81),
	.w1(32'h3b777bea),
	.w2(32'h3ab21a1f),
	.w3(32'hba7e64ec),
	.w4(32'h3af9a5de),
	.w5(32'hbb7d41b0),
	.w6(32'h3b1338d3),
	.w7(32'h3bbd2419),
	.w8(32'hbb2bc974),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1d51),
	.w1(32'h3b0ae42e),
	.w2(32'h38ff5ca1),
	.w3(32'h3b4b3f93),
	.w4(32'h3b08d255),
	.w5(32'hba96de2a),
	.w6(32'hb9547355),
	.w7(32'h390970db),
	.w8(32'hba17b076),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a67b5e),
	.w1(32'hbadf662d),
	.w2(32'hbbb137cc),
	.w3(32'hba60d842),
	.w4(32'hbb2d37ee),
	.w5(32'hbc598cf9),
	.w6(32'hba8ca6fa),
	.w7(32'hbb438861),
	.w8(32'hbc0adca6),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec5820),
	.w1(32'hbbd99e11),
	.w2(32'hbbdf960e),
	.w3(32'hbceedbc4),
	.w4(32'hbcaa6e95),
	.w5(32'h399652e3),
	.w6(32'hbcb06468),
	.w7(32'hbc4321f1),
	.w8(32'hbacec86d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b529b),
	.w1(32'h3b6dcaab),
	.w2(32'hbb34b2cc),
	.w3(32'h3c4c32a4),
	.w4(32'h3c0b8165),
	.w5(32'h3a1dc6c9),
	.w6(32'h3beb6a6b),
	.w7(32'h3b1bfaaa),
	.w8(32'hba21cb70),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7da163),
	.w1(32'h3b614472),
	.w2(32'h3be4e182),
	.w3(32'h3b3784d2),
	.w4(32'h3b92735c),
	.w5(32'h3be86ba5),
	.w6(32'h3b2ecfb2),
	.w7(32'h3b942ccb),
	.w8(32'h3be6e4a5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55ff03),
	.w1(32'h3c1b4df2),
	.w2(32'h3c4b8748),
	.w3(32'h3c1b2236),
	.w4(32'h3bf2050c),
	.w5(32'h3c5da7f6),
	.w6(32'h3be2bf8c),
	.w7(32'h3bfeceb5),
	.w8(32'h3c7aba2a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43c64e),
	.w1(32'h3b3261d3),
	.w2(32'h3bc07071),
	.w3(32'h3caf3e27),
	.w4(32'h3b9b66af),
	.w5(32'h3bdef2a6),
	.w6(32'h3ca5f744),
	.w7(32'h3bccf9ec),
	.w8(32'h3b9a43a0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c149fbe),
	.w1(32'h3c14e9c3),
	.w2(32'h3a414f9c),
	.w3(32'h3c217e2f),
	.w4(32'h3c2cf429),
	.w5(32'h3b812e6d),
	.w6(32'h3b450f51),
	.w7(32'h3baae94b),
	.w8(32'h3b59aa50),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35f432),
	.w1(32'h3b961905),
	.w2(32'hbb95b4cf),
	.w3(32'h3c41a14f),
	.w4(32'h3b9daea5),
	.w5(32'hbc058ba7),
	.w6(32'h3c162287),
	.w7(32'h3b276a53),
	.w8(32'hbc0bbe90),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3735d),
	.w1(32'hbba9a423),
	.w2(32'hbc9365f8),
	.w3(32'hbbf5c6b3),
	.w4(32'hbbb3bf20),
	.w5(32'hbcc15a11),
	.w6(32'hbc00611c),
	.w7(32'hbc033310),
	.w8(32'hbca2e9b0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc598d70),
	.w1(32'hbbfc4675),
	.w2(32'h3c6732f4),
	.w3(32'hbcc638f8),
	.w4(32'hbc91d343),
	.w5(32'h3c8cc447),
	.w6(32'hbcbdfb26),
	.w7(32'hbc8e9b6f),
	.w8(32'h3c607cc7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1598c6),
	.w1(32'h3c0b17e0),
	.w2(32'h3a93ab57),
	.w3(32'h3c4faa6f),
	.w4(32'h3c337462),
	.w5(32'hb980a510),
	.w6(32'h3c03be5b),
	.w7(32'h3bfa69ac),
	.w8(32'h3b86f227),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baefacd),
	.w1(32'h3b288702),
	.w2(32'h3b65af69),
	.w3(32'h3a3255c6),
	.w4(32'h38d3cf4d),
	.w5(32'hbac2e365),
	.w6(32'h3a87826f),
	.w7(32'h3b8c74c3),
	.w8(32'hb93b52c5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b910e),
	.w1(32'h3c12aba1),
	.w2(32'h3b9ce6c0),
	.w3(32'h3a9569f2),
	.w4(32'h3bc563dd),
	.w5(32'h3c05edaa),
	.w6(32'h3b140c57),
	.w7(32'h3b4d133b),
	.w8(32'h3bdec9d7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd44458),
	.w1(32'h3b5b3afb),
	.w2(32'h3b4676d0),
	.w3(32'h3bade579),
	.w4(32'hbb2d631f),
	.w5(32'h3aac13fc),
	.w6(32'h3aeb4808),
	.w7(32'hbba1958b),
	.w8(32'hbbba985e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd83c1),
	.w1(32'hbb11c2b8),
	.w2(32'h3a3ef4fa),
	.w3(32'hbc33a8a6),
	.w4(32'hbbc713b9),
	.w5(32'hbb5c21dd),
	.w6(32'hbc26a9cb),
	.w7(32'hbbeec119),
	.w8(32'hb9f9a3e3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c783a2d),
	.w1(32'hbac34875),
	.w2(32'hbc4f67af),
	.w3(32'h3c6079d1),
	.w4(32'hbb9af5f7),
	.w5(32'hbca8dc80),
	.w6(32'h3bf6150a),
	.w7(32'hba976b12),
	.w8(32'hbca49cee),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc811a4e),
	.w1(32'hbc345de8),
	.w2(32'hbb4ac4cc),
	.w3(32'hbd1dfbb4),
	.w4(32'hbceb80e7),
	.w5(32'hbb9157bf),
	.w6(32'hbd1b1507),
	.w7(32'hbcce44dc),
	.w8(32'hbb5e624f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ec7e8),
	.w1(32'hbbcfbab9),
	.w2(32'h3c2cd65b),
	.w3(32'hbc37b99d),
	.w4(32'hbb48ff38),
	.w5(32'h3baa41fd),
	.w6(32'hbc0d57a2),
	.w7(32'hbb9d7f9c),
	.w8(32'h3bad16ea),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9db283),
	.w1(32'h3c5d4239),
	.w2(32'h3b517156),
	.w3(32'h3c3a15b5),
	.w4(32'h3c6b6121),
	.w5(32'hbac868f1),
	.w6(32'h3c04bb95),
	.w7(32'h3c1b38b0),
	.w8(32'hbb8a6706),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c414312),
	.w1(32'hbb0aedf7),
	.w2(32'h3bb46680),
	.w3(32'h3c5a9454),
	.w4(32'hbb5d9796),
	.w5(32'h3974ae59),
	.w6(32'h3c4681bb),
	.w7(32'hbad62e47),
	.w8(32'hbb1a1480),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c011043),
	.w1(32'h3b0f7be0),
	.w2(32'hbba971c7),
	.w3(32'hbb34c966),
	.w4(32'hbb443193),
	.w5(32'hbc0d4f0b),
	.w6(32'hbad43908),
	.w7(32'hbaab17d1),
	.w8(32'hbbd33c7a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b403911),
	.w1(32'h3a07c999),
	.w2(32'hbc8bb834),
	.w3(32'h3a9ff90e),
	.w4(32'hbb0ddf64),
	.w5(32'hbcb7abf2),
	.w6(32'h3a175214),
	.w7(32'hbb77697c),
	.w8(32'hbcac583f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadac9a),
	.w1(32'hbc9b6b5e),
	.w2(32'hbb7bf767),
	.w3(32'hbcfbb557),
	.w4(32'hbcdc58a8),
	.w5(32'h3af0a2c8),
	.w6(32'hbcf5b31c),
	.w7(32'hbcc91e4d),
	.w8(32'h3a734771),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c8916),
	.w1(32'h3adff99c),
	.w2(32'h3c1d750b),
	.w3(32'hbb007716),
	.w4(32'h3b25cd70),
	.w5(32'h3c337b2e),
	.w6(32'hbb2c5b49),
	.w7(32'hbbb9a141),
	.w8(32'hb965ddc0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c543d),
	.w1(32'h3c4f471b),
	.w2(32'hbc013d52),
	.w3(32'h3c942a78),
	.w4(32'h3c762a6b),
	.w5(32'hbbb757ab),
	.w6(32'h3bc85a2d),
	.w7(32'h3b42ae8b),
	.w8(32'hbb122077),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f439f),
	.w1(32'h3bd5abd7),
	.w2(32'hbc0f7566),
	.w3(32'h3c1ad80f),
	.w4(32'h3b25d4bf),
	.w5(32'hbbde493a),
	.w6(32'h3bd39da4),
	.w7(32'h3bd7b907),
	.w8(32'hbbe3961e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a39d5),
	.w1(32'h3c58a10c),
	.w2(32'h3b992acb),
	.w3(32'h3c6142bd),
	.w4(32'h3c4a16b1),
	.w5(32'h3abaf624),
	.w6(32'h3c4c0dde),
	.w7(32'h3bd30822),
	.w8(32'h3b35d6dd),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b309e32),
	.w1(32'h3c0db8dd),
	.w2(32'hb99bf9db),
	.w3(32'h39a86301),
	.w4(32'h3bb93a84),
	.w5(32'hbc393f02),
	.w6(32'h3b1d20a5),
	.w7(32'h3be0be02),
	.w8(32'hbc056562),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ebd1f),
	.w1(32'hbb090a5a),
	.w2(32'h3b06ac82),
	.w3(32'hbd06fbfc),
	.w4(32'hbca75061),
	.w5(32'h3a37f74d),
	.w6(32'hbcde9120),
	.w7(32'hbc6551d9),
	.w8(32'h3a86cc87),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877b05),
	.w1(32'h3b3a151e),
	.w2(32'hbb799c66),
	.w3(32'h3b652c64),
	.w4(32'h3ab7b437),
	.w5(32'hbc3d82fd),
	.w6(32'h3b0b6ff8),
	.w7(32'hba3ae790),
	.w8(32'hbc49e920),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dfcca),
	.w1(32'hbb6a28f7),
	.w2(32'h3a6ae2c0),
	.w3(32'hbc17cb89),
	.w4(32'hbb15454a),
	.w5(32'hbac84ff2),
	.w6(32'hbc14e36a),
	.w7(32'hbb7414fd),
	.w8(32'hbaf56385),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea631e),
	.w1(32'hbb433365),
	.w2(32'h3ae72659),
	.w3(32'h3a658cfd),
	.w4(32'hbb9eee66),
	.w5(32'h3b1b3a2d),
	.w6(32'hbac26530),
	.w7(32'hbbfdc405),
	.w8(32'h3a13c65b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f0063),
	.w1(32'h3b50d648),
	.w2(32'h3b9206f1),
	.w3(32'h3bb90bb8),
	.w4(32'h3a9fae46),
	.w5(32'h3b625052),
	.w6(32'hbac42ed9),
	.w7(32'h3ba9e801),
	.w8(32'h3b44873e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0b6a1),
	.w1(32'h3c2868ba),
	.w2(32'hbc3897d1),
	.w3(32'h3bc500ae),
	.w4(32'h3bd52729),
	.w5(32'hbbd83834),
	.w6(32'h3bc5e900),
	.w7(32'h3bf3ca57),
	.w8(32'hbc074c4d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1379be),
	.w1(32'h3b21d285),
	.w2(32'hb8d46333),
	.w3(32'h3b423702),
	.w4(32'h3b0baf7a),
	.w5(32'hbb88ba4a),
	.w6(32'hb7f4cd67),
	.w7(32'h3b79d5af),
	.w8(32'hbbedfb62),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ce4bf),
	.w1(32'h3c02aeff),
	.w2(32'h3b8ecc55),
	.w3(32'h3b11f348),
	.w4(32'h3b29317c),
	.w5(32'h3b6afa0b),
	.w6(32'h3b6eb29c),
	.w7(32'h3b762bd0),
	.w8(32'h3b4d9d7d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac446cd),
	.w1(32'h3b069568),
	.w2(32'h3ad245e7),
	.w3(32'h3bc42147),
	.w4(32'h3b64547f),
	.w5(32'h3b05b688),
	.w6(32'hba2e6c0c),
	.w7(32'h3b95baf0),
	.w8(32'h3bda51bf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c2dca),
	.w1(32'h3b853270),
	.w2(32'h3b854ca4),
	.w3(32'h3c358ff4),
	.w4(32'h3b13d240),
	.w5(32'hbb319d85),
	.w6(32'h3c26596b),
	.w7(32'h3bb0119f),
	.w8(32'hbaddbb4a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c362533),
	.w1(32'h3b5bac51),
	.w2(32'h3b746075),
	.w3(32'h3c2117cc),
	.w4(32'hb8e9e845),
	.w5(32'h3bd131a2),
	.w6(32'h3b86da62),
	.w7(32'hbad1ad08),
	.w8(32'h394d0f33),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a752e),
	.w1(32'h3ade35b7),
	.w2(32'h3a99db85),
	.w3(32'h3bf9d818),
	.w4(32'h3a459e7c),
	.w5(32'h3ac394c4),
	.w6(32'h3bd383e1),
	.w7(32'h3b101cf6),
	.w8(32'h3b4877d5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71d4a6),
	.w1(32'h3baed0ce),
	.w2(32'h3b195545),
	.w3(32'h3ba2b8ed),
	.w4(32'h3b453f5a),
	.w5(32'h3a47e88f),
	.w6(32'h3bb73b0c),
	.w7(32'h3bafb845),
	.w8(32'h3b3ecc3d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafc2d3),
	.w1(32'hbb24aac8),
	.w2(32'h39c93f3d),
	.w3(32'h3b9665a8),
	.w4(32'hbb13c3ed),
	.w5(32'h3b78f3a7),
	.w6(32'h3b991533),
	.w7(32'hba6b6a3a),
	.w8(32'h3b8f9782),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ae287),
	.w1(32'h3a0fcdfc),
	.w2(32'h3b425dca),
	.w3(32'h3c0bc3b9),
	.w4(32'h3b471c14),
	.w5(32'h3b3ac739),
	.w6(32'h3bda84f9),
	.w7(32'h3ba51551),
	.w8(32'h397610db),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a60f4),
	.w1(32'h3a5df95a),
	.w2(32'h3ae4cf25),
	.w3(32'h3b1c0fe2),
	.w4(32'hbb332a3c),
	.w5(32'hbaa679ff),
	.w6(32'h3ba211eb),
	.w7(32'hba29c996),
	.w8(32'h39c4a29f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fea874),
	.w1(32'h3b812025),
	.w2(32'h3bdf722b),
	.w3(32'h3b467324),
	.w4(32'h3a940b42),
	.w5(32'h38508d92),
	.w6(32'h3ade113e),
	.w7(32'h3b6d484f),
	.w8(32'hba13b9f1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a070c32),
	.w1(32'h3b406080),
	.w2(32'h3ba17330),
	.w3(32'h3b72d8f1),
	.w4(32'hbb35e187),
	.w5(32'h3be99068),
	.w6(32'hbac70fa4),
	.w7(32'h39fa5a9b),
	.w8(32'h3ba91936),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dd0c3),
	.w1(32'hbc3e73f9),
	.w2(32'hbbb3ce30),
	.w3(32'h3b9d21cf),
	.w4(32'hbbd335a3),
	.w5(32'hbb6ab7d2),
	.w6(32'hba775aee),
	.w7(32'hbc0e660b),
	.w8(32'hbb9781e9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987bb8),
	.w1(32'hb9b917d3),
	.w2(32'h3bf3d5df),
	.w3(32'h3c01c5e7),
	.w4(32'h3b7eca71),
	.w5(32'h3ba2301f),
	.w6(32'h3bbc5a0f),
	.w7(32'h3c57cef0),
	.w8(32'h3bbba977),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63b2ce),
	.w1(32'h3c0865b3),
	.w2(32'hbaf46cbe),
	.w3(32'h3c504fc3),
	.w4(32'h3b43f0f0),
	.w5(32'hbbc06851),
	.w6(32'h3c48c6cc),
	.w7(32'h3bc8fd90),
	.w8(32'hbbda4088),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53d4e9),
	.w1(32'hbb2abe13),
	.w2(32'hbb6b4f31),
	.w3(32'hbb1954e7),
	.w4(32'hbb4bff28),
	.w5(32'hbb4c4732),
	.w6(32'h3b0b6554),
	.w7(32'h3b5a0e07),
	.w8(32'hbaf82cb7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1ee16),
	.w1(32'hbb584ef1),
	.w2(32'h3b8913b9),
	.w3(32'hbafc2ee3),
	.w4(32'hba8a22b5),
	.w5(32'h3bf5d60e),
	.w6(32'hba395264),
	.w7(32'hba9e59bc),
	.w8(32'h3a67ddb1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c588fb2),
	.w1(32'h3c6bf4f7),
	.w2(32'h39a22bcc),
	.w3(32'h3c74ad43),
	.w4(32'h3c8b51a4),
	.w5(32'hbaf3c2f2),
	.w6(32'h3bb5271d),
	.w7(32'h3b640efa),
	.w8(32'h3b72e83f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13c98c),
	.w1(32'h3acf30e9),
	.w2(32'h3c2814b0),
	.w3(32'hba6b9c6b),
	.w4(32'hbb0b1341),
	.w5(32'h3bec04db),
	.w6(32'h3b81ad02),
	.w7(32'h3b01fae7),
	.w8(32'h3c0ef82e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2da6ad),
	.w1(32'h3c38f0ce),
	.w2(32'hbaaffdc0),
	.w3(32'h3c5554ab),
	.w4(32'h3c22af1a),
	.w5(32'h3ae48953),
	.w6(32'h3c1e5dc3),
	.w7(32'h3c46a802),
	.w8(32'hba93e442),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf267e0),
	.w1(32'h3975c1b0),
	.w2(32'hbbb9fc2e),
	.w3(32'h3a5a7916),
	.w4(32'h3b567de3),
	.w5(32'h3bae8dc6),
	.w6(32'h3bcfdd0f),
	.w7(32'h3ad76dac),
	.w8(32'h37d257a2),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4689c2),
	.w1(32'h39a84f36),
	.w2(32'hbc204276),
	.w3(32'h3b96fcbc),
	.w4(32'h3baf1b44),
	.w5(32'hbc02601f),
	.w6(32'h3ac45958),
	.w7(32'h386f8bc4),
	.w8(32'hbbe09c32),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c0182),
	.w1(32'hbbd85c55),
	.w2(32'hbbb25a64),
	.w3(32'hbae4b292),
	.w4(32'hba716843),
	.w5(32'hba0585bf),
	.w6(32'hba1d471e),
	.w7(32'hba86bc43),
	.w8(32'hbb8bcf6b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ed0ee),
	.w1(32'hba8379a0),
	.w2(32'h3b32076a),
	.w3(32'h3c07852d),
	.w4(32'h3b8a30cc),
	.w5(32'hba9fb746),
	.w6(32'h3b64713b),
	.w7(32'hba259838),
	.w8(32'h3a19eb4f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c272c03),
	.w1(32'h3c6d4382),
	.w2(32'hbb2e773e),
	.w3(32'h3c20d7d1),
	.w4(32'h3c16edef),
	.w5(32'hbb2287a4),
	.w6(32'h3bad071b),
	.w7(32'h3c3a3802),
	.w8(32'hba8d1359),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38853584),
	.w1(32'hbb819855),
	.w2(32'h3bc67c29),
	.w3(32'h394c154e),
	.w4(32'hbb4744d3),
	.w5(32'h3bc10a58),
	.w6(32'h388e6016),
	.w7(32'hbb59abb6),
	.w8(32'h3b184006),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c068a61),
	.w1(32'h3bae4304),
	.w2(32'h3b29e69b),
	.w3(32'h3bedfaf0),
	.w4(32'h3c23b2ff),
	.w5(32'h3a743aa9),
	.w6(32'h3c1f799b),
	.w7(32'h3c238dfe),
	.w8(32'hbaa154a3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be24734),
	.w1(32'h39d1251a),
	.w2(32'h3a460c26),
	.w3(32'h3c3a7bc1),
	.w4(32'h3b91806c),
	.w5(32'h3b34e077),
	.w6(32'h3b9f49f7),
	.w7(32'hb9cdeb65),
	.w8(32'h3b25f593),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70bc13),
	.w1(32'h3b672002),
	.w2(32'h3b823769),
	.w3(32'h3b723b12),
	.w4(32'hba75d90b),
	.w5(32'h3b63e9f5),
	.w6(32'h3b303554),
	.w7(32'h3aaf6fd3),
	.w8(32'h3b1b80c5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule