module layer_10_featuremap_480(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d7994),
	.w1(32'hbaa6e1b8),
	.w2(32'h3a60043c),
	.w3(32'hbb25982f),
	.w4(32'hba24e033),
	.w5(32'h3b76a2ba),
	.w6(32'hbaba181a),
	.w7(32'hbb844ac5),
	.w8(32'hbb730e23),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb504b65),
	.w1(32'hbbcd9ffc),
	.w2(32'hbb4084f0),
	.w3(32'hbc339bc3),
	.w4(32'hbb39aee1),
	.w5(32'hbc40e0b9),
	.w6(32'hbbe5c578),
	.w7(32'hbaed2a0a),
	.w8(32'hbaa5f27d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fc5ce),
	.w1(32'h3c048d31),
	.w2(32'h3b2808c4),
	.w3(32'h3b4d0567),
	.w4(32'h3a52aead),
	.w5(32'h3bab5234),
	.w6(32'h3b442409),
	.w7(32'hbbb81867),
	.w8(32'h3b101a46),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72363f),
	.w1(32'hbc0bca17),
	.w2(32'hbb5023b3),
	.w3(32'hbb34a55f),
	.w4(32'hbc445aa5),
	.w5(32'h3c2f3814),
	.w6(32'h3a321229),
	.w7(32'hbbb408c4),
	.w8(32'hbb51ab1f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e3bc7),
	.w1(32'h3b3cbccd),
	.w2(32'hbbd1082a),
	.w3(32'hbc76fa1b),
	.w4(32'h3bba094b),
	.w5(32'hbb8fcd2c),
	.w6(32'hbc277ad7),
	.w7(32'h3b8ac455),
	.w8(32'hbb61b28d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb60a85),
	.w1(32'hbb805bf8),
	.w2(32'hbabb522d),
	.w3(32'hbc2fd85d),
	.w4(32'h3b4404c3),
	.w5(32'hbc0bb072),
	.w6(32'hbc092fd4),
	.w7(32'hbb15b41c),
	.w8(32'h3b331267),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c0381),
	.w1(32'h3bed5a09),
	.w2(32'h3b2668e4),
	.w3(32'h3bff47b6),
	.w4(32'h3c77de67),
	.w5(32'h3b84753d),
	.w6(32'h3c524839),
	.w7(32'h3c309936),
	.w8(32'hbb7f48eb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab57e97),
	.w1(32'hbb88a0fe),
	.w2(32'h3b296e09),
	.w3(32'h3ab19057),
	.w4(32'hbc2e572a),
	.w5(32'hbaee6c94),
	.w6(32'h3b418d77),
	.w7(32'h3ac6e80e),
	.w8(32'h3b72bb29),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e066f),
	.w1(32'h3b74f995),
	.w2(32'h3b7dc3ce),
	.w3(32'h3c450544),
	.w4(32'h3bc82ddd),
	.w5(32'hb8137d17),
	.w6(32'h3c205c9f),
	.w7(32'h3bd514fd),
	.w8(32'h3b84a2be),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53b2ac),
	.w1(32'hba86fb58),
	.w2(32'hbbb93f60),
	.w3(32'h3b3a58dd),
	.w4(32'h3ac3f6a0),
	.w5(32'hba9bbb06),
	.w6(32'h3baee9bf),
	.w7(32'hb9b28b10),
	.w8(32'hbc2214c3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb527b1),
	.w1(32'hbc231b56),
	.w2(32'hbc029f5b),
	.w3(32'hbc569ae1),
	.w4(32'hbb1ccedd),
	.w5(32'hbb57b9c0),
	.w6(32'hbbf4bb0f),
	.w7(32'hbba8429e),
	.w8(32'hbb4ff9ef),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f82b64),
	.w1(32'h3bf00cdd),
	.w2(32'h3b0d428b),
	.w3(32'h3a3937e7),
	.w4(32'h3bccde14),
	.w5(32'hbba35846),
	.w6(32'h39388b8a),
	.w7(32'hbaa4c5a7),
	.w8(32'hbb8945cd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa604b9),
	.w1(32'h3bf2d821),
	.w2(32'h3b133864),
	.w3(32'hba65b5a0),
	.w4(32'h3c8ce17f),
	.w5(32'hbc4699c8),
	.w6(32'hbaad061f),
	.w7(32'h3c16fe11),
	.w8(32'h3b39e815),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84c297),
	.w1(32'h3b7a7932),
	.w2(32'hbba2ac50),
	.w3(32'h3cdb3264),
	.w4(32'h3b7c7c02),
	.w5(32'h3a8a3a31),
	.w6(32'h3cb8e460),
	.w7(32'h3bef45a1),
	.w8(32'h3c007c6f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75917d),
	.w1(32'hbc5df31d),
	.w2(32'h3a87c1ba),
	.w3(32'hbb2f8710),
	.w4(32'hbb6bed3b),
	.w5(32'hbc00d667),
	.w6(32'hbb5dfaa4),
	.w7(32'hbc22ac46),
	.w8(32'hb9e5eec7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06b185),
	.w1(32'hbae10ff0),
	.w2(32'hbba6d4b7),
	.w3(32'hbc4d6120),
	.w4(32'hbb945e6a),
	.w5(32'hbc963560),
	.w6(32'hbc71bc60),
	.w7(32'hbc50304c),
	.w8(32'hbc28777c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fbe85),
	.w1(32'hb9d2038e),
	.w2(32'hbae7904f),
	.w3(32'h3bf34798),
	.w4(32'hb9b13b91),
	.w5(32'hbab754b8),
	.w6(32'hbb6eba33),
	.w7(32'hbb7705e9),
	.w8(32'hbb35b833),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d6df8),
	.w1(32'hbac1441d),
	.w2(32'hbc195ad0),
	.w3(32'hbabfc36c),
	.w4(32'hbbcbed1f),
	.w5(32'hbc123232),
	.w6(32'h39d6a718),
	.w7(32'hbb90be0d),
	.w8(32'hba12ad95),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b993645),
	.w1(32'h3a2b8027),
	.w2(32'hbb669f79),
	.w3(32'h3ab05a57),
	.w4(32'h3b965f80),
	.w5(32'hbbfecb0c),
	.w6(32'h3b7c651d),
	.w7(32'hb975be88),
	.w8(32'hbaec6a1c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6076fc),
	.w1(32'h3b316c13),
	.w2(32'h3b4b3def),
	.w3(32'hbb2d8272),
	.w4(32'hba8c92a7),
	.w5(32'h3a8a01c2),
	.w6(32'hbba07b80),
	.w7(32'hbb4339f6),
	.w8(32'h3b1af383),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0a3a3),
	.w1(32'hbba42e84),
	.w2(32'hbb16d9c5),
	.w3(32'hbb8f00df),
	.w4(32'hbb6a59db),
	.w5(32'hbbad3887),
	.w6(32'hbbbb86aa),
	.w7(32'hbbafef14),
	.w8(32'hbb09fc52),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fc7ee),
	.w1(32'hbb5a1fd6),
	.w2(32'h3ad0983a),
	.w3(32'h3bf48d52),
	.w4(32'hbb211bb0),
	.w5(32'hba96109d),
	.w6(32'h3b88dc93),
	.w7(32'hbb8a7068),
	.w8(32'hbb872986),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdf0e7),
	.w1(32'h3beed9ca),
	.w2(32'hbb5604a8),
	.w3(32'h3aea4a9b),
	.w4(32'hbba7c94c),
	.w5(32'h3b878d44),
	.w6(32'h3a39ba6d),
	.w7(32'hbb133b33),
	.w8(32'h39d9f27c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1db082),
	.w1(32'h3c1a5752),
	.w2(32'h3ba84a2c),
	.w3(32'hbb822cea),
	.w4(32'h3bba6064),
	.w5(32'hbb081dbe),
	.w6(32'hbac4f654),
	.w7(32'h3abd86d0),
	.w8(32'hbad90bb8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8f61c),
	.w1(32'hbaaea3bb),
	.w2(32'hbaa121e1),
	.w3(32'hbc671f74),
	.w4(32'hbbdefb4e),
	.w5(32'h3c92dae1),
	.w6(32'hbc90e16a),
	.w7(32'hb8c7d0ab),
	.w8(32'h3b9a6d5a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f8de3),
	.w1(32'hba7264cd),
	.w2(32'hbb6ada22),
	.w3(32'hbc0d1b07),
	.w4(32'hbaf7d8fd),
	.w5(32'h3b3ef6d9),
	.w6(32'hbc1252a0),
	.w7(32'h3c0889b7),
	.w8(32'hbb19c2a8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb252807),
	.w1(32'hbab90de5),
	.w2(32'h3aedfeb3),
	.w3(32'hbc0f1caa),
	.w4(32'h3a644d9c),
	.w5(32'h3b77f433),
	.w6(32'hbbc9b32a),
	.w7(32'h3baca2ce),
	.w8(32'h390a836d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51529f),
	.w1(32'h3bcec08f),
	.w2(32'h3c3f0275),
	.w3(32'hbc4bbd49),
	.w4(32'hb7ed7668),
	.w5(32'h3cddabbc),
	.w6(32'hbbbddd13),
	.w7(32'h3b44f66a),
	.w8(32'h3c83568b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb4fc6),
	.w1(32'h3badb73a),
	.w2(32'h3c136898),
	.w3(32'h3c68617e),
	.w4(32'h3c1cebf4),
	.w5(32'h3bd1d116),
	.w6(32'h3b95886a),
	.w7(32'h3a00c9f2),
	.w8(32'hbb91007b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b038b14),
	.w1(32'hbb874766),
	.w2(32'hbb40c2fd),
	.w3(32'hbb41b09d),
	.w4(32'h3ae6d3a0),
	.w5(32'hbbf8e78d),
	.w6(32'hbaa46132),
	.w7(32'hbaa0ecb3),
	.w8(32'hbc042a83),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8098b7),
	.w1(32'h39d26c91),
	.w2(32'h3abea72b),
	.w3(32'h3c3cfcb1),
	.w4(32'h3af7f9f9),
	.w5(32'hbb833239),
	.w6(32'h3bf6603f),
	.w7(32'h3acf18b6),
	.w8(32'hbae89086),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbd25e),
	.w1(32'hb93bdadb),
	.w2(32'h3bda4694),
	.w3(32'hbb686687),
	.w4(32'hb94b01b5),
	.w5(32'h3c259829),
	.w6(32'h39eac5b6),
	.w7(32'hbb7d705d),
	.w8(32'h3b303546),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f361),
	.w1(32'h3c38c574),
	.w2(32'h3b5bf46c),
	.w3(32'hbb0c8ff2),
	.w4(32'h3bd2f68c),
	.w5(32'h3c3c348d),
	.w6(32'h3b1cf97e),
	.w7(32'hbb7fbd00),
	.w8(32'h3ac80c5f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2192f8),
	.w1(32'h3abf1a15),
	.w2(32'h3b8f6392),
	.w3(32'h3b709066),
	.w4(32'hbaf3dc61),
	.w5(32'h3c6253b3),
	.w6(32'h3a863261),
	.w7(32'h3ab0ea2e),
	.w8(32'h3bba8f5d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32f0c4),
	.w1(32'h3a6e21e5),
	.w2(32'h3b6d7ded),
	.w3(32'h3c4fac24),
	.w4(32'hbba1fabf),
	.w5(32'h3ba9817b),
	.w6(32'hba5b01c8),
	.w7(32'h3b8cddcb),
	.w8(32'h3be065d9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46d235),
	.w1(32'hbb833cc5),
	.w2(32'hbb0189fa),
	.w3(32'h3c2daf3f),
	.w4(32'hba9793eb),
	.w5(32'hbb49a8a7),
	.w6(32'h39ba2bdf),
	.w7(32'hbbcb24ed),
	.w8(32'hbad4ec5c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59ffda),
	.w1(32'hbc25ccfa),
	.w2(32'h3befd3f6),
	.w3(32'hbab9d5f9),
	.w4(32'h3b81b9d4),
	.w5(32'h3a64b36f),
	.w6(32'h3be6919a),
	.w7(32'hbb4b8bd0),
	.w8(32'hbc152bf5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc56e4),
	.w1(32'h3b25f82a),
	.w2(32'hbad48f65),
	.w3(32'hbc0f6530),
	.w4(32'h3c4d415a),
	.w5(32'h3b7ddfe5),
	.w6(32'hbbc5f07e),
	.w7(32'h3afaaa1b),
	.w8(32'h3a5c419e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819692),
	.w1(32'h3c956836),
	.w2(32'h3c82b331),
	.w3(32'h3bc5e2a0),
	.w4(32'h3c3b7097),
	.w5(32'h3cdc2f7f),
	.w6(32'h3ba933ae),
	.w7(32'h3bbcade5),
	.w8(32'h3c3c3bbf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c832f49),
	.w1(32'h3b2e12df),
	.w2(32'h3abf5a5d),
	.w3(32'h3c35b766),
	.w4(32'hbb1b1de1),
	.w5(32'h3c8618ec),
	.w6(32'h3c3a0676),
	.w7(32'h3adc2e9e),
	.w8(32'h3bab0c00),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdbcf5),
	.w1(32'h3a431ee2),
	.w2(32'hbb6bf6de),
	.w3(32'hbc45dd55),
	.w4(32'h3bdc6242),
	.w5(32'h3ac47b91),
	.w6(32'hbb63b212),
	.w7(32'h3acaab05),
	.w8(32'h3bc45bc5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabea762),
	.w1(32'hbb94b423),
	.w2(32'h3b71a2fa),
	.w3(32'h3bd84d51),
	.w4(32'hbb96ef8d),
	.w5(32'h3b08706d),
	.w6(32'h3b6c8f1d),
	.w7(32'hbb8c96d0),
	.w8(32'h3ad19df6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c340d),
	.w1(32'h3b20f4a2),
	.w2(32'h3ad7d356),
	.w3(32'hbc82a963),
	.w4(32'h3ab83b86),
	.w5(32'hbb4198d9),
	.w6(32'hbc6d7448),
	.w7(32'hba335527),
	.w8(32'h3ab37cb3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98294b),
	.w1(32'hb9ef4249),
	.w2(32'hbbc5b4b2),
	.w3(32'h3bd245d0),
	.w4(32'hbc8bb65e),
	.w5(32'h3c5a324c),
	.w6(32'h3c0db6e8),
	.w7(32'hbbbe3532),
	.w8(32'h3bc8b5de),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ef246),
	.w1(32'h39f7fc3b),
	.w2(32'h3a7440e2),
	.w3(32'hbb70cafb),
	.w4(32'h3aca97d5),
	.w5(32'hbb8db41c),
	.w6(32'hbba535bf),
	.w7(32'h3af9fd08),
	.w8(32'hbba56e2a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399aa574),
	.w1(32'h3998043a),
	.w2(32'hb934c61e),
	.w3(32'h3b30fdca),
	.w4(32'hb9d43545),
	.w5(32'hbbc4d2eb),
	.w6(32'hbb475057),
	.w7(32'hbb9bdf19),
	.w8(32'hbb09d7b5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b56c6),
	.w1(32'h3c4069af),
	.w2(32'h3c3f3d08),
	.w3(32'h3c1c197b),
	.w4(32'h3c3224c9),
	.w5(32'h3c68a0ab),
	.w6(32'hbbad3ff4),
	.w7(32'h3b7484ac),
	.w8(32'h3c532241),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb5754),
	.w1(32'h3c1f5208),
	.w2(32'h3b23432b),
	.w3(32'h3c8383b9),
	.w4(32'h3bcd397f),
	.w5(32'h3c536bc3),
	.w6(32'h3c90ebcd),
	.w7(32'h3c038360),
	.w8(32'h3c0190be),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44b869),
	.w1(32'h3b0da19d),
	.w2(32'h3b394016),
	.w3(32'h3b9dbf74),
	.w4(32'hb8952bfd),
	.w5(32'h3ae12ba0),
	.w6(32'hbae963aa),
	.w7(32'h3b9e9df5),
	.w8(32'h3c2412f1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63eb6f),
	.w1(32'hbba35a18),
	.w2(32'h3bd4ce4f),
	.w3(32'h3c117b65),
	.w4(32'hbb6a56d5),
	.w5(32'h3b7a7cab),
	.w6(32'h3c117111),
	.w7(32'hbbdaba35),
	.w8(32'h3b8cddcc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1f7f2),
	.w1(32'h3be26a39),
	.w2(32'hbb11353d),
	.w3(32'hbacbb962),
	.w4(32'h3beee39c),
	.w5(32'hbbc55034),
	.w6(32'h3c0134d8),
	.w7(32'h3bc48c15),
	.w8(32'hbbb0292a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91dc50),
	.w1(32'hba085f9f),
	.w2(32'hbb9e32d1),
	.w3(32'hbc030462),
	.w4(32'hbbabf146),
	.w5(32'h3bd87714),
	.w6(32'hbb8f0927),
	.w7(32'hbbb321bd),
	.w8(32'hba8ae18c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09965d),
	.w1(32'hbb627339),
	.w2(32'h3947cb6b),
	.w3(32'hbbe98943),
	.w4(32'hbb26e588),
	.w5(32'hbbb351c8),
	.w6(32'hbb8e2b5e),
	.w7(32'h3ae6c563),
	.w8(32'h3b20122b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b1bd),
	.w1(32'h3b07971c),
	.w2(32'hbb6b3bc7),
	.w3(32'h3b935bd9),
	.w4(32'h397cf52a),
	.w5(32'h3c105acc),
	.w6(32'h3c1486cb),
	.w7(32'hbba5ae21),
	.w8(32'hbb18dcd8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b790a3c),
	.w1(32'h3b69eefb),
	.w2(32'hbba20be6),
	.w3(32'hb9f7a254),
	.w4(32'hbb40e672),
	.w5(32'hbb302ebd),
	.w6(32'hbbb14214),
	.w7(32'hbaa24b85),
	.w8(32'hbbabf95b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf84fa6),
	.w1(32'hbb33bb7a),
	.w2(32'hbb4122db),
	.w3(32'hbbfc51f3),
	.w4(32'h3ae7d656),
	.w5(32'hbbc57f8e),
	.w6(32'hbadb6c45),
	.w7(32'h3b2556dd),
	.w8(32'hbb150021),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17db7a),
	.w1(32'hbc04b062),
	.w2(32'hbb627b3a),
	.w3(32'h3b82f355),
	.w4(32'hbbb44b46),
	.w5(32'hbb9c3156),
	.w6(32'h3b7cb188),
	.w7(32'hbc04a13e),
	.w8(32'hbbc6a4ba),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb016ef7),
	.w1(32'hbbc063e1),
	.w2(32'h3abd1c61),
	.w3(32'hbb7e665e),
	.w4(32'hbbcb955d),
	.w5(32'h39cd1006),
	.w6(32'hbba86f99),
	.w7(32'h3b2a37e4),
	.w8(32'hbac3eeb0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba775e85),
	.w1(32'h39666ee3),
	.w2(32'h3b7a2b52),
	.w3(32'h3a4e1f5f),
	.w4(32'hbb9e4092),
	.w5(32'h3c430a09),
	.w6(32'hba5bddc6),
	.w7(32'hbb1adfd8),
	.w8(32'h3986dca5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b689494),
	.w1(32'h3b020961),
	.w2(32'h3ab1aa8d),
	.w3(32'h3b0bebff),
	.w4(32'hbc0cc353),
	.w5(32'h3bcd7359),
	.w6(32'h3bfa0bc3),
	.w7(32'hb9a6b2e8),
	.w8(32'hbbbb6e51),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3f42),
	.w1(32'h3a01c6ec),
	.w2(32'hbb3cd3ba),
	.w3(32'h3b53933f),
	.w4(32'hbaf93be4),
	.w5(32'hbaf14260),
	.w6(32'h3ae474ae),
	.w7(32'h3b354403),
	.w8(32'h38ab6083),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96e981),
	.w1(32'h3c1e5575),
	.w2(32'h3c2e2fe0),
	.w3(32'h3b175ae5),
	.w4(32'h3b8df7d6),
	.w5(32'h3b1a3517),
	.w6(32'hbad318b0),
	.w7(32'h3b5efe60),
	.w8(32'h3c31eaab),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3245d),
	.w1(32'h3b44f10a),
	.w2(32'hbad71a2a),
	.w3(32'h3b9b9864),
	.w4(32'hbbb66099),
	.w5(32'h3b92ce90),
	.w6(32'h3922dd9d),
	.w7(32'hbade95d7),
	.w8(32'hbafc3500),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba85636),
	.w1(32'h3b28546b),
	.w2(32'hbb8b091a),
	.w3(32'hba6bcf92),
	.w4(32'h3abc9e3e),
	.w5(32'hbbdd2bc0),
	.w6(32'hbb1b6293),
	.w7(32'hbbb6da51),
	.w8(32'hbba55f1f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ebe9d),
	.w1(32'h3a762751),
	.w2(32'h3b7650b9),
	.w3(32'hbad0b1c1),
	.w4(32'h3bc7abdf),
	.w5(32'h3b81c0b5),
	.w6(32'h3b14511e),
	.w7(32'h3b38c016),
	.w8(32'h3b7fd71c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b035f),
	.w1(32'h3c0ec813),
	.w2(32'h3c5449f8),
	.w3(32'h3b23e5a5),
	.w4(32'h3a372399),
	.w5(32'h3c37109d),
	.w6(32'h3bc928fd),
	.w7(32'h3acdda3f),
	.w8(32'h3becb987),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5138c1),
	.w1(32'hbc2a629e),
	.w2(32'hbc398fea),
	.w3(32'hbbd3f181),
	.w4(32'hbcab981d),
	.w5(32'hbbf8ba76),
	.w6(32'h3a937a36),
	.w7(32'hbc53d075),
	.w8(32'hbc38e621),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf63c1d),
	.w1(32'h3b880496),
	.w2(32'h3b066929),
	.w3(32'h3bf40a3f),
	.w4(32'hbbb939cd),
	.w5(32'hbc5c477c),
	.w6(32'h3c14e7da),
	.w7(32'hbaa88cff),
	.w8(32'h3aa8002b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33428c),
	.w1(32'h3b7ea7ce),
	.w2(32'hbc1e0387),
	.w3(32'h3cba2ae8),
	.w4(32'h3b858820),
	.w5(32'h3b0ebfbe),
	.w6(32'h3c80fe9f),
	.w7(32'hbab510a3),
	.w8(32'hbb9da83c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba673356),
	.w1(32'hbacb87a8),
	.w2(32'hb9a29f18),
	.w3(32'hbc541627),
	.w4(32'hb9d91066),
	.w5(32'h3a518196),
	.w6(32'hbc7aafcf),
	.w7(32'hbc189557),
	.w8(32'hbbf124ee),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb260926),
	.w1(32'hbb8efafa),
	.w2(32'hbb4102ef),
	.w3(32'hbb4034d2),
	.w4(32'hbb6d5017),
	.w5(32'hbad2ffd9),
	.w6(32'hbb62420d),
	.w7(32'hba2f58a0),
	.w8(32'h3a619694),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb876340d),
	.w1(32'hba8486be),
	.w2(32'hbac6a240),
	.w3(32'h3aeb95e6),
	.w4(32'h357dc135),
	.w5(32'hbae0c52d),
	.w6(32'h3b49cb1c),
	.w7(32'h3aff32eb),
	.w8(32'h3999735a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb89aa),
	.w1(32'h380ebee0),
	.w2(32'hb9de6494),
	.w3(32'hb9e388d8),
	.w4(32'hbac1587a),
	.w5(32'hba254f50),
	.w6(32'h3a81b978),
	.w7(32'hba9be6c8),
	.w8(32'hbac29f7f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a755a7d),
	.w1(32'hb924b3a6),
	.w2(32'hbb128da8),
	.w3(32'h3b1c386d),
	.w4(32'h3aaffc6e),
	.w5(32'hba8e08a2),
	.w6(32'h3b29596c),
	.w7(32'h3ae239a4),
	.w8(32'hb99fa61a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3fa39),
	.w1(32'hbb3bf68c),
	.w2(32'hbb751587),
	.w3(32'hbada9ec4),
	.w4(32'hbb54bb8f),
	.w5(32'hbba445c3),
	.w6(32'hbac56696),
	.w7(32'hbb21fef6),
	.w8(32'hbbda9f77),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98db45),
	.w1(32'hbb3d1500),
	.w2(32'hbb843ec1),
	.w3(32'hbad1d016),
	.w4(32'hbb423734),
	.w5(32'hbb62744d),
	.w6(32'hbadb73ef),
	.w7(32'hbb12c58a),
	.w8(32'hbb8f09a2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926de68),
	.w1(32'hbb0a0374),
	.w2(32'hbb132b66),
	.w3(32'hba6f22a1),
	.w4(32'hbbb86ab4),
	.w5(32'hbb8cc3b9),
	.w6(32'h3b189623),
	.w7(32'hbb9d21a2),
	.w8(32'hbbb6a481),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099aff),
	.w1(32'h3a4504ba),
	.w2(32'h3a15c221),
	.w3(32'hbb51d344),
	.w4(32'hba031f86),
	.w5(32'hba9b11bd),
	.w6(32'hbbb0a4da),
	.w7(32'hbb2fdc83),
	.w8(32'hbb7c089c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7af9373),
	.w1(32'hbb3e74ab),
	.w2(32'hbb9a49a1),
	.w3(32'h3a9b80a5),
	.w4(32'hbb6334d2),
	.w5(32'hbb42e55b),
	.w6(32'h3a975118),
	.w7(32'hbb120007),
	.w8(32'hbb53831d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2b6e1),
	.w1(32'h3acf555c),
	.w2(32'hbae19f4c),
	.w3(32'h3a81865c),
	.w4(32'hbb94e02b),
	.w5(32'hbafca6af),
	.w6(32'h3b9fc039),
	.w7(32'hba83039f),
	.w8(32'hbb85ff16),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6238d7),
	.w1(32'h3b43e8ba),
	.w2(32'h3a998952),
	.w3(32'hbb79aae7),
	.w4(32'h3b66cbfc),
	.w5(32'h3a8a78c3),
	.w6(32'hbb706cf9),
	.w7(32'hba1ae51a),
	.w8(32'hbaddc1ca),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3aa91),
	.w1(32'hb7e1826e),
	.w2(32'hba6fcde1),
	.w3(32'h3b1e4cde),
	.w4(32'hb8aefd08),
	.w5(32'hb98cbd3a),
	.w6(32'h39e94c84),
	.w7(32'h3a5dc492),
	.w8(32'h3a20c8c0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbababa56),
	.w1(32'h39ad8b25),
	.w2(32'h3993a859),
	.w3(32'hbaa14919),
	.w4(32'hba29c5f1),
	.w5(32'hbaa6fcae),
	.w6(32'hba8b4346),
	.w7(32'h3ac7659b),
	.w8(32'h3aec9005),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a8383),
	.w1(32'hba1a2ebe),
	.w2(32'hbb7d71e1),
	.w3(32'hbaaf7ff8),
	.w4(32'hbb1677fb),
	.w5(32'hbb8367fa),
	.w6(32'h37a86832),
	.w7(32'hbaf60459),
	.w8(32'hba12bc76),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf4a3),
	.w1(32'h3a067d82),
	.w2(32'h37d396de),
	.w3(32'hba4b7b69),
	.w4(32'h3a3356a7),
	.w5(32'h3a6d8888),
	.w6(32'h39c4866d),
	.w7(32'h3a58e13a),
	.w8(32'h3aeb320c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39974ba3),
	.w1(32'hbb63a31c),
	.w2(32'hbba29524),
	.w3(32'h3a3def19),
	.w4(32'hbb8fd483),
	.w5(32'hbc0573f0),
	.w6(32'h3b38ec4e),
	.w7(32'hbb48cd14),
	.w8(32'hbbeaf7c2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93c864),
	.w1(32'h3a3cbeee),
	.w2(32'h3ab9303d),
	.w3(32'hbc0b65e5),
	.w4(32'h3ad10a6e),
	.w5(32'h3a51eed3),
	.w6(32'hbbdc80a8),
	.w7(32'hba1017a0),
	.w8(32'hbab287ba),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90004a),
	.w1(32'h3b8f6ef4),
	.w2(32'h3a4d528c),
	.w3(32'h39fbac76),
	.w4(32'h3b25481f),
	.w5(32'hbb4bed0a),
	.w6(32'h3aa6ec07),
	.w7(32'h3b4484f5),
	.w8(32'hbabcd8ca),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38980a),
	.w1(32'hbb64587a),
	.w2(32'hbb082902),
	.w3(32'hba8acb95),
	.w4(32'hbb69100f),
	.w5(32'hb9f245c3),
	.w6(32'hba7ef424),
	.w7(32'hbbd3cb68),
	.w8(32'hbb5c712e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959f80a),
	.w1(32'hbaed8d2e),
	.w2(32'hbbaee385),
	.w3(32'h3af4dfc4),
	.w4(32'hbb7c26d6),
	.w5(32'hbb731c88),
	.w6(32'h3ada5b23),
	.w7(32'hbb497902),
	.w8(32'hbb16889c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d8a92),
	.w1(32'hbb7778d7),
	.w2(32'hbb0d5cf7),
	.w3(32'hba3c4ae6),
	.w4(32'h3986d602),
	.w5(32'h3ae4b098),
	.w6(32'hba9d51f6),
	.w7(32'hbb47cf1b),
	.w8(32'hba8474d9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe0ff6),
	.w1(32'h3b0693c1),
	.w2(32'hbbb049cf),
	.w3(32'hbace2379),
	.w4(32'hb9a7b80f),
	.w5(32'hbbdb5036),
	.w6(32'hba1ff219),
	.w7(32'hbc06a520),
	.w8(32'hbc627ac5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ad8c2),
	.w1(32'h392fc43c),
	.w2(32'h3b217d09),
	.w3(32'hbacf6ec4),
	.w4(32'h3b55d529),
	.w5(32'h3ac5dc5b),
	.w6(32'hbbccb4ce),
	.w7(32'h3a6ec6f4),
	.w8(32'h3a581614),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90aa30f),
	.w1(32'hbb1e2662),
	.w2(32'hbbe7fd0f),
	.w3(32'hbb8269ae),
	.w4(32'hbc2bd3c0),
	.w5(32'hbc2430fa),
	.w6(32'hb99503b0),
	.w7(32'hbc008eb2),
	.w8(32'hbc0fbdae),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50e95b),
	.w1(32'hbb34c905),
	.w2(32'hbbd05375),
	.w3(32'hbb32fbe6),
	.w4(32'hbbdf554c),
	.w5(32'hbbf351bf),
	.w6(32'hbae741ec),
	.w7(32'hbbc474a1),
	.w8(32'hbc0810af),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7685e4),
	.w1(32'h3980f444),
	.w2(32'h3a6c61f2),
	.w3(32'hbbcd9bf6),
	.w4(32'hba8d5fc3),
	.w5(32'h3a1bcf31),
	.w6(32'hbb9613dd),
	.w7(32'hb945970a),
	.w8(32'hbafaf404),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1e45e),
	.w1(32'h3ac385c0),
	.w2(32'h3a3e79b3),
	.w3(32'hbb003180),
	.w4(32'h3a450fe0),
	.w5(32'h39898db0),
	.w6(32'hba7028c7),
	.w7(32'h3b14ee82),
	.w8(32'h3ab466ca),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88c1e1),
	.w1(32'hbb3677cd),
	.w2(32'hbbba192d),
	.w3(32'h39a327f4),
	.w4(32'hbb6a1c4d),
	.w5(32'hbb380013),
	.w6(32'h3b7fc90c),
	.w7(32'hbb570ea1),
	.w8(32'hbb15be13),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a8d95),
	.w1(32'h3b84b8f5),
	.w2(32'h3ade7e5a),
	.w3(32'hbb568152),
	.w4(32'h3bd7d970),
	.w5(32'h3c1a3f0f),
	.w6(32'h3a92538e),
	.w7(32'hbb2dbde0),
	.w8(32'hbbd44c0c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f83f5),
	.w1(32'hbc2f7197),
	.w2(32'hbc1f4ce7),
	.w3(32'h36c0d21a),
	.w4(32'hbc80d872),
	.w5(32'hbc32f175),
	.w6(32'hbbf095c8),
	.w7(32'hbc0d742b),
	.w8(32'hbbdb670b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe39566),
	.w1(32'hb895e415),
	.w2(32'h3b2bac32),
	.w3(32'hbb96db74),
	.w4(32'h3b5b8a9c),
	.w5(32'h3bd56b27),
	.w6(32'hbbe2cef1),
	.w7(32'hb9dddfb0),
	.w8(32'h3b86d153),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb0239),
	.w1(32'h3a1e9e24),
	.w2(32'h3aea046d),
	.w3(32'hbb132860),
	.w4(32'h3abd1ad5),
	.w5(32'h3adba75f),
	.w6(32'hbbb78ef9),
	.w7(32'hb9921138),
	.w8(32'h3a494561),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb959198),
	.w1(32'h3ab7049a),
	.w2(32'h3a7b311e),
	.w3(32'h3b89c22a),
	.w4(32'h393fcaa7),
	.w5(32'hbb80bf33),
	.w6(32'h3c244a2b),
	.w7(32'hba86f72d),
	.w8(32'hbb954121),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad071a4),
	.w1(32'h3b572c22),
	.w2(32'h3ad83700),
	.w3(32'hbb27832b),
	.w4(32'h3b958e6b),
	.w5(32'h3b04c6f3),
	.w6(32'hbae81852),
	.w7(32'h3baf6a9f),
	.w8(32'h3b8951d1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43c0fe),
	.w1(32'hbb92778c),
	.w2(32'h3a2db4f1),
	.w3(32'hbb5e3975),
	.w4(32'hbbe5b54e),
	.w5(32'hbbe547e8),
	.w6(32'h3c14cf0a),
	.w7(32'h3a621f98),
	.w8(32'hbc04f479),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46491e),
	.w1(32'hbaf64d69),
	.w2(32'h3add5e49),
	.w3(32'h3b89dfd6),
	.w4(32'h3af47187),
	.w5(32'h3aacf429),
	.w6(32'h3b1e408b),
	.w7(32'h3b02a5cf),
	.w8(32'h3a1149ed),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03704f),
	.w1(32'hbae50aab),
	.w2(32'hbb14ba20),
	.w3(32'hba743bdb),
	.w4(32'hba308cb8),
	.w5(32'hbaf9bf3d),
	.w6(32'hb734a0e6),
	.w7(32'h3a320dad),
	.w8(32'hb9b745d4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5696ef),
	.w1(32'hba951e28),
	.w2(32'hbb05619e),
	.w3(32'hbb60bdba),
	.w4(32'hbb50854e),
	.w5(32'hbb05bb1c),
	.w6(32'hbb698ecc),
	.w7(32'hbbb26597),
	.w8(32'hbbd3c67f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1510a3),
	.w1(32'h3aa9e90f),
	.w2(32'hba6c2c93),
	.w3(32'hbb36e2a0),
	.w4(32'h3abd1204),
	.w5(32'hb9f78102),
	.w6(32'hbb40c0a8),
	.w7(32'hb9fe9efb),
	.w8(32'hb8e0a392),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00facc),
	.w1(32'h3b2571ca),
	.w2(32'h3ae1e886),
	.w3(32'hbb221176),
	.w4(32'h3b0e17ac),
	.w5(32'h3abc7b80),
	.w6(32'hbae2a2c5),
	.w7(32'hbb09c95d),
	.w8(32'hbb02a373),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1f736),
	.w1(32'hbb98c045),
	.w2(32'hbb33dfc5),
	.w3(32'h3adbd788),
	.w4(32'hbaafb4e5),
	.w5(32'hba047da1),
	.w6(32'hba46fa92),
	.w7(32'hbbc1e3fb),
	.w8(32'hbb9a9581),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5aad2),
	.w1(32'hbad77671),
	.w2(32'h3a225e0a),
	.w3(32'hbbad90b8),
	.w4(32'hbb2cde32),
	.w5(32'h38e5d96a),
	.w6(32'hbbc83e4f),
	.w7(32'hbb8acb74),
	.w8(32'hbabd1c7a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b421b55),
	.w1(32'h3b84c148),
	.w2(32'h3b1d9399),
	.w3(32'hba69cb13),
	.w4(32'h3b943d2d),
	.w5(32'h3b8d4672),
	.w6(32'hba9f4bdb),
	.w7(32'h3b528b5c),
	.w8(32'h3b33073a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14106c),
	.w1(32'hbb8e98cc),
	.w2(32'hbc22eba9),
	.w3(32'hbb78475a),
	.w4(32'hbc1672b9),
	.w5(32'hbc0eab0a),
	.w6(32'hba18ce70),
	.w7(32'hbbb74c0a),
	.w8(32'hbb8c7ad4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084bee),
	.w1(32'hb976b380),
	.w2(32'hba6b2d7b),
	.w3(32'hb9fb1247),
	.w4(32'h391a3819),
	.w5(32'hbaa6e973),
	.w6(32'hbb37ce24),
	.w7(32'hba4621a9),
	.w8(32'hba73d602),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99112d),
	.w1(32'hbb3a80a8),
	.w2(32'hba0a9843),
	.w3(32'hba8fecf2),
	.w4(32'hbb64fe7c),
	.w5(32'hbacacf36),
	.w6(32'hba976fdf),
	.w7(32'hbabb9b11),
	.w8(32'hba687cf1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803e41),
	.w1(32'hbb18babf),
	.w2(32'hbb783036),
	.w3(32'hbb1691e8),
	.w4(32'hba7a2dcb),
	.w5(32'hba0cfc2d),
	.w6(32'hb9a31ac4),
	.w7(32'hb937a8ce),
	.w8(32'hba37fde3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb583527),
	.w1(32'hb9d4b125),
	.w2(32'h3ad31b6d),
	.w3(32'hbb2c8a89),
	.w4(32'hb769cbd7),
	.w5(32'h3b1f92b6),
	.w6(32'hba82c777),
	.w7(32'hba01dcb1),
	.w8(32'h3a9ded6f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed0ce9),
	.w1(32'h3b03392c),
	.w2(32'h39e3d1f3),
	.w3(32'hba0ca1dd),
	.w4(32'h3b282366),
	.w5(32'hbad35c23),
	.w6(32'hbaa4f84d),
	.w7(32'h3b518e7d),
	.w8(32'h385126e0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2521e2),
	.w1(32'h3b41b4e2),
	.w2(32'h3ae19e1a),
	.w3(32'h3ae4d810),
	.w4(32'h3b8171bc),
	.w5(32'h3b59ec91),
	.w6(32'h3a89ae01),
	.w7(32'h3b217739),
	.w8(32'h3ac6bdb8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cc053),
	.w1(32'hbbc28140),
	.w2(32'hbbc309d7),
	.w3(32'hba99150f),
	.w4(32'hbbd5db9b),
	.w5(32'hbba54861),
	.w6(32'h3a215cb2),
	.w7(32'hbbfafe6a),
	.w8(32'hbbcc5bce),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfab94a),
	.w1(32'hbb02ded3),
	.w2(32'hba9bd36f),
	.w3(32'hbb8e8d5a),
	.w4(32'hba02d911),
	.w5(32'hbad52c03),
	.w6(32'hbb9e3500),
	.w7(32'hbbab3f07),
	.w8(32'hbb4c348f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b0507),
	.w1(32'hbb006635),
	.w2(32'hbafc2b56),
	.w3(32'hbbb503cb),
	.w4(32'hbb79e4b9),
	.w5(32'hbb6be6c5),
	.w6(32'hbc1d141b),
	.w7(32'hbb8c870c),
	.w8(32'hbb9276ea),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba177f3e),
	.w1(32'hbad26a8c),
	.w2(32'hbb4c2b68),
	.w3(32'hba6f847c),
	.w4(32'hba928f86),
	.w5(32'hbae75f2a),
	.w6(32'hba92454d),
	.w7(32'hba87dc6a),
	.w8(32'hbad96375),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1599df),
	.w1(32'h3afddb67),
	.w2(32'hb9b8e9d7),
	.w3(32'hbb003cbf),
	.w4(32'h3b174dcd),
	.w5(32'hba03b3f4),
	.w6(32'hbaeb0cc6),
	.w7(32'h3b2ef3ba),
	.w8(32'h3971eb66),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e12e6),
	.w1(32'hba53da61),
	.w2(32'h382b9396),
	.w3(32'hba50f349),
	.w4(32'h3a459c20),
	.w5(32'hb939c80c),
	.w6(32'h3a8da20d),
	.w7(32'hb88afac5),
	.w8(32'hb95503fa),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d679a),
	.w1(32'hbc0d0618),
	.w2(32'hbc3df13a),
	.w3(32'h3a806ae4),
	.w4(32'hbc4b1bc2),
	.w5(32'hbc6836a1),
	.w6(32'hb9bf27c7),
	.w7(32'hbc1b7a76),
	.w8(32'hbc3b37df),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba698822),
	.w1(32'h3befee87),
	.w2(32'hb77c8e04),
	.w3(32'hbbbba126),
	.w4(32'h3b4dcb73),
	.w5(32'h3a045f6b),
	.w6(32'hbb53f5ec),
	.w7(32'hba1e8706),
	.w8(32'hbb793e75),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098668),
	.w1(32'h3aa5c8e6),
	.w2(32'hbb1d0bf3),
	.w3(32'hba3d6787),
	.w4(32'hbada1447),
	.w5(32'h39fa0a4c),
	.w6(32'hba3d4090),
	.w7(32'hbb60fdfa),
	.w8(32'hbaef4142),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b1b08),
	.w1(32'hbaef1d13),
	.w2(32'hba823863),
	.w3(32'h3a264c77),
	.w4(32'hbb190037),
	.w5(32'hba3fabbd),
	.w6(32'h398fdc35),
	.w7(32'hbaaa2f04),
	.w8(32'h389c2cf5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e03c),
	.w1(32'hbb36354c),
	.w2(32'hba979e4f),
	.w3(32'hbafbc90c),
	.w4(32'hba1a93b8),
	.w5(32'hbb11e5c7),
	.w6(32'h3a50c36d),
	.w7(32'hbaa85222),
	.w8(32'hba8460ca),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad193c6),
	.w1(32'h3aa0bb8d),
	.w2(32'h3a445fbb),
	.w3(32'hba49dd17),
	.w4(32'h39fdc883),
	.w5(32'h39cde5e8),
	.w6(32'hba626a86),
	.w7(32'h39df7cc4),
	.w8(32'hb88d5026),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdb6d2),
	.w1(32'hbba7cd52),
	.w2(32'hbb836ead),
	.w3(32'h3a3a9248),
	.w4(32'hbbb4212a),
	.w5(32'hbb4a41fe),
	.w6(32'h3a9b5670),
	.w7(32'hbb9e9ec5),
	.w8(32'hbb463b98),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6abb6b),
	.w1(32'hbb339cd0),
	.w2(32'hbbb8453b),
	.w3(32'hbbc653b4),
	.w4(32'hbbbe2a6c),
	.w5(32'hbbd17b43),
	.w6(32'hbb752d60),
	.w7(32'hbba7dd50),
	.w8(32'hbbed7170),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb211679),
	.w1(32'h3aaecb6e),
	.w2(32'hbb98d134),
	.w3(32'hbacccaa1),
	.w4(32'h3ad29a8c),
	.w5(32'hba8a16a1),
	.w6(32'h3b2bde84),
	.w7(32'h3b007b47),
	.w8(32'hba94a359),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949915a),
	.w1(32'hbaad509f),
	.w2(32'h3b12fdb6),
	.w3(32'hb971ef2f),
	.w4(32'hb9c12036),
	.w5(32'h3a9d33d2),
	.w6(32'h3a80da19),
	.w7(32'hbb632406),
	.w8(32'hbaeadaf6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa90568),
	.w1(32'h3a34ee77),
	.w2(32'hbb871ec2),
	.w3(32'hba876b44),
	.w4(32'hbaaf4ff6),
	.w5(32'hbb4e926d),
	.w6(32'hbb30b705),
	.w7(32'hb9c070cc),
	.w8(32'hbb6b5fbb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb303d84),
	.w1(32'hbb976adb),
	.w2(32'hbc0e7e13),
	.w3(32'hb84a847a),
	.w4(32'hbb7f3dc2),
	.w5(32'hbbc47b0f),
	.w6(32'h3ab183f6),
	.w7(32'hba5d1b80),
	.w8(32'hbae3a2c1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5546de),
	.w1(32'h396198cf),
	.w2(32'h39c60ab2),
	.w3(32'hbb1b1a3c),
	.w4(32'hbabecdfe),
	.w5(32'h38f5f9ce),
	.w6(32'hbb1a4a76),
	.w7(32'hbb1cd561),
	.w8(32'hba8a93e6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e97033),
	.w1(32'hbb0c2fee),
	.w2(32'hbb05e1b7),
	.w3(32'h39b7baa3),
	.w4(32'hbb9a17e4),
	.w5(32'hbb23bd13),
	.w6(32'h3b283da9),
	.w7(32'hbb3169e9),
	.w8(32'hbb497e68),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadac76),
	.w1(32'h384d339c),
	.w2(32'h3ac3444f),
	.w3(32'hbac0ce48),
	.w4(32'hba50afab),
	.w5(32'h394ae133),
	.w6(32'hbb086b34),
	.w7(32'h3ad59e9e),
	.w8(32'h39623719),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf250d),
	.w1(32'h3aa3dd5b),
	.w2(32'h3b03b575),
	.w3(32'h3b20fa40),
	.w4(32'hba5c79f6),
	.w5(32'hbb0f2145),
	.w6(32'hba4bcac8),
	.w7(32'hba96fbbb),
	.w8(32'hb92dffc9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b438034),
	.w1(32'hba93491f),
	.w2(32'hba90b110),
	.w3(32'hba9b7979),
	.w4(32'hb9cd0f3e),
	.w5(32'h3a39771d),
	.w6(32'h398b2a66),
	.w7(32'hba2c0534),
	.w8(32'h3a0cc6c6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391732ea),
	.w1(32'h3a1f1c42),
	.w2(32'hba0666df),
	.w3(32'hba677901),
	.w4(32'hb9d381df),
	.w5(32'hba78c67c),
	.w6(32'h3ab89fcb),
	.w7(32'h38ded19d),
	.w8(32'hbad5b9fd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba839edf),
	.w1(32'hbad7186d),
	.w2(32'hbb09b6ab),
	.w3(32'hbb0ff337),
	.w4(32'hbacc3fb3),
	.w5(32'hbaf0437f),
	.w6(32'hbac484ca),
	.w7(32'hbb4aff66),
	.w8(32'hbb65f96d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f51c),
	.w1(32'hb9cb60bb),
	.w2(32'h3b14a618),
	.w3(32'hbaf46c9a),
	.w4(32'h3a2fb502),
	.w5(32'h3b4175b7),
	.w6(32'hbb4406c0),
	.w7(32'hba43d2f0),
	.w8(32'h3a6e1547),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94a809),
	.w1(32'hba9535f7),
	.w2(32'h3a8c67b8),
	.w3(32'h39d27814),
	.w4(32'h3b0dc0e2),
	.w5(32'h3b1f21b9),
	.w6(32'hbabd15cc),
	.w7(32'hb8d97e8e),
	.w8(32'h39116418),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c0985),
	.w1(32'hbb2cd7e0),
	.w2(32'hbbc3b02c),
	.w3(32'hb9b84369),
	.w4(32'hbb2acbc6),
	.w5(32'hbbc99667),
	.w6(32'h3ac78ae0),
	.w7(32'hbaaf82e4),
	.w8(32'hbbb04cb7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11fbda),
	.w1(32'h3ae92893),
	.w2(32'h3a063aeb),
	.w3(32'hbb4a08a8),
	.w4(32'h3ab3df53),
	.w5(32'h39930764),
	.w6(32'hba56b095),
	.w7(32'h3b475b36),
	.w8(32'h3b2ef016),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09223a),
	.w1(32'hba333976),
	.w2(32'hbbb2f332),
	.w3(32'h39b0c0ba),
	.w4(32'h3ab2ce0a),
	.w5(32'hbb6b38c2),
	.w6(32'h3af303f9),
	.w7(32'h3ab117d1),
	.w8(32'hbb458d46),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b78a3),
	.w1(32'hbb628eff),
	.w2(32'hbbb5b582),
	.w3(32'hbb99f95e),
	.w4(32'hbb7d685d),
	.w5(32'hbb241df7),
	.w6(32'hbb6cb5a1),
	.w7(32'hba8f0b50),
	.w8(32'hba80f676),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39d0ce),
	.w1(32'hb9318ab1),
	.w2(32'hbb71e8e1),
	.w3(32'h3b6474e0),
	.w4(32'h38fb783c),
	.w5(32'hbba8eac4),
	.w6(32'h3b5a7c9a),
	.w7(32'hbba00b7b),
	.w8(32'hbbaac3ea),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab97f1d),
	.w1(32'h39222a2c),
	.w2(32'hb8576c88),
	.w3(32'h3b4d8be6),
	.w4(32'hbb32f08e),
	.w5(32'hbaf1a568),
	.w6(32'hbb8b2c52),
	.w7(32'hbc00a466),
	.w8(32'hbbee05ed),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0035c),
	.w1(32'hbb59dc15),
	.w2(32'hbbaba7b2),
	.w3(32'hbbb9190d),
	.w4(32'hbb9cff84),
	.w5(32'hbc0ac1ec),
	.w6(32'hbb9580fb),
	.w7(32'hbb8d32b8),
	.w8(32'hbbc34f6a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaceeb1),
	.w1(32'h3ab1d650),
	.w2(32'hb906703c),
	.w3(32'hbbc9d179),
	.w4(32'hba89217f),
	.w5(32'hbba13bc5),
	.w6(32'hbbca539d),
	.w7(32'hbb07168e),
	.w8(32'hbbd0ace9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a100206),
	.w1(32'hbb1ddc20),
	.w2(32'h3b0a70f4),
	.w3(32'hbb3dda1c),
	.w4(32'hba4b531e),
	.w5(32'h3b59383e),
	.w6(32'hbba32b54),
	.w7(32'hbad32c35),
	.w8(32'h3b0c78e6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840ac5),
	.w1(32'hbb454345),
	.w2(32'hbade1106),
	.w3(32'hbac8b5aa),
	.w4(32'hbb1bf92c),
	.w5(32'hba54fb41),
	.w6(32'hbab94f05),
	.w7(32'hbbaadd40),
	.w8(32'hbbb38c2a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb101939),
	.w1(32'hbaed5202),
	.w2(32'hb7f7b654),
	.w3(32'hbbb0b3a5),
	.w4(32'hbb3d0289),
	.w5(32'hbab19a13),
	.w6(32'hbbca09e9),
	.w7(32'hbb0503f8),
	.w8(32'hbaabc056),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6bf31),
	.w1(32'hbbb741fc),
	.w2(32'hbb9995ea),
	.w3(32'h3a66eb99),
	.w4(32'hbb0d72cd),
	.w5(32'hba0af8ad),
	.w6(32'h3a036d89),
	.w7(32'hbb8c3aa0),
	.w8(32'hbb949173),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ad7f),
	.w1(32'h39ef07b5),
	.w2(32'h3a3dbdcc),
	.w3(32'hb9e9f01e),
	.w4(32'h3ad45a4d),
	.w5(32'h3ad5f5b4),
	.w6(32'hbb854702),
	.w7(32'h3ac2dfe6),
	.w8(32'h3b00ead3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae267dd),
	.w1(32'h3b974850),
	.w2(32'hb938f572),
	.w3(32'h3ad37fa2),
	.w4(32'h3a1862d2),
	.w5(32'hba21a6ff),
	.w6(32'h3b94a9ba),
	.w7(32'hbaf3b2e6),
	.w8(32'hbb2b5aff),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913f0da),
	.w1(32'h3accf777),
	.w2(32'h39fd24be),
	.w3(32'h3b5d2671),
	.w4(32'h3b57b5df),
	.w5(32'h3a1d3e29),
	.w6(32'h39b41a2e),
	.w7(32'h3abc924b),
	.w8(32'h3a04fb22),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e7823),
	.w1(32'hba564c97),
	.w2(32'hba703119),
	.w3(32'hbafceb72),
	.w4(32'hba67b517),
	.w5(32'h38ba394d),
	.w6(32'hbb411906),
	.w7(32'hb9b5cc66),
	.w8(32'h3b06a7f8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64cc55),
	.w1(32'h3a1aebcb),
	.w2(32'hbaae3ccc),
	.w3(32'hbb44fbae),
	.w4(32'h3a88622b),
	.w5(32'h3a817c55),
	.w6(32'h39a59a1f),
	.w7(32'h38fdf5f7),
	.w8(32'hba9c0142),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b336219),
	.w1(32'h3b36fcbc),
	.w2(32'hba09bd8d),
	.w3(32'h3b7bef3f),
	.w4(32'hba25439e),
	.w5(32'h3a7822e9),
	.w6(32'h3b2a955b),
	.w7(32'h3a224a48),
	.w8(32'hbae6fcb6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0a439),
	.w1(32'hb99467cc),
	.w2(32'hba7ee9e5),
	.w3(32'hba7c1f18),
	.w4(32'h39d68a3c),
	.w5(32'h391a5151),
	.w6(32'hb9fa4407),
	.w7(32'h3a0ffb22),
	.w8(32'hb9740f59),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac93cb),
	.w1(32'h3ab8c3ab),
	.w2(32'h3b07c3c0),
	.w3(32'hba923ea5),
	.w4(32'h39721c22),
	.w5(32'h3b215264),
	.w6(32'h3a263e19),
	.w7(32'h3846fee9),
	.w8(32'hb949a7d1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af245ee),
	.w1(32'hba97b5ba),
	.w2(32'hba33dc5c),
	.w3(32'h3a50bd35),
	.w4(32'hbac5790b),
	.w5(32'hba3094ca),
	.w6(32'h3a54dec4),
	.w7(32'hbb2ee0ea),
	.w8(32'hbae850bb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f86ec),
	.w1(32'h3aa25cec),
	.w2(32'h3b33d557),
	.w3(32'h3b3566d1),
	.w4(32'hba5583c3),
	.w5(32'h3ad64df9),
	.w6(32'h3aaf4799),
	.w7(32'h3a707188),
	.w8(32'h3b67bf86),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaacb99),
	.w1(32'hba84205d),
	.w2(32'hba95c161),
	.w3(32'h3a1b2bcb),
	.w4(32'hbb0f6ba8),
	.w5(32'hba9fc651),
	.w6(32'h396c178a),
	.w7(32'hba97a136),
	.w8(32'hba1dc5b5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98c8f4),
	.w1(32'h3b106189),
	.w2(32'h3b0a582a),
	.w3(32'hbb5d3e2d),
	.w4(32'h3b41cdcc),
	.w5(32'h3b4a6f74),
	.w6(32'hbb0c5cca),
	.w7(32'h3b6d5d9d),
	.w8(32'h3b102ba8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af75010),
	.w1(32'h3ab30601),
	.w2(32'hb962f43e),
	.w3(32'h3a43c4f8),
	.w4(32'hbac30e82),
	.w5(32'hb944df08),
	.w6(32'h3b1b57bb),
	.w7(32'hba989f8c),
	.w8(32'h39409b02),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0374b),
	.w1(32'hbaea9920),
	.w2(32'hbbff6255),
	.w3(32'hbb52f85d),
	.w4(32'hbb523eb6),
	.w5(32'hbb55c15a),
	.w6(32'h3a13ebcb),
	.w7(32'hbb014d35),
	.w8(32'hbb6892c3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa251e8),
	.w1(32'hbaa2ee88),
	.w2(32'hbb19ec98),
	.w3(32'hba90a7c0),
	.w4(32'hbb3b873f),
	.w5(32'hbb1c65bb),
	.w6(32'h3af536c4),
	.w7(32'hbab63545),
	.w8(32'hbaf14247),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bbb76f),
	.w1(32'h3a2af971),
	.w2(32'hbb8b5ab5),
	.w3(32'h3ac1599f),
	.w4(32'hb9a0f57c),
	.w5(32'hbb9f2c6b),
	.w6(32'h3b424b70),
	.w7(32'hb97e7d0f),
	.w8(32'hbb6abf0d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8636ff),
	.w1(32'h3aca77c7),
	.w2(32'h3a51989e),
	.w3(32'hb98e3a96),
	.w4(32'h3a6fa5d0),
	.w5(32'h3a16d2e3),
	.w6(32'hbab5a6cf),
	.w7(32'h3a69cdc2),
	.w8(32'hb9a63b84),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a379e),
	.w1(32'h3a8cce21),
	.w2(32'hbb61b6e3),
	.w3(32'hbb946575),
	.w4(32'h3a9ced1e),
	.w5(32'hbaaef750),
	.w6(32'hbace2251),
	.w7(32'h3b0de2b6),
	.w8(32'hba157713),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cab81),
	.w1(32'hbaa50484),
	.w2(32'hba5b341c),
	.w3(32'h3ab8cd66),
	.w4(32'hba2fcd33),
	.w5(32'h3b0e6591),
	.w6(32'h3a68abfe),
	.w7(32'h3985d944),
	.w8(32'h3abb4093),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae023d),
	.w1(32'hbb2662ce),
	.w2(32'h3ab377bb),
	.w3(32'h3b33c427),
	.w4(32'hbb1e0294),
	.w5(32'h3a658b6c),
	.w6(32'h3a7f181b),
	.w7(32'hbb777f2d),
	.w8(32'h3a0e80ef),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdadc8),
	.w1(32'h3b2afa67),
	.w2(32'hbb04d4b1),
	.w3(32'hbaf01bf2),
	.w4(32'h3b15a302),
	.w5(32'hbb3920b1),
	.w6(32'hbb235b86),
	.w7(32'h3b64d6e8),
	.w8(32'hba5511f3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f38c0a),
	.w1(32'hba2b1ee2),
	.w2(32'hbba8e809),
	.w3(32'hbb00dfc0),
	.w4(32'hbb49ef99),
	.w5(32'hbb9d1718),
	.w6(32'h3af10ddf),
	.w7(32'hbb336d1f),
	.w8(32'hbb9d838d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba708a75),
	.w1(32'h3b054ed0),
	.w2(32'h3b0d43e9),
	.w3(32'hba0f2a4d),
	.w4(32'h3aa48652),
	.w5(32'h3a184024),
	.w6(32'hba92112d),
	.w7(32'h39e9456c),
	.w8(32'h3a350a2d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5410a3),
	.w1(32'hbb3736cd),
	.w2(32'hba880c4c),
	.w3(32'hb9a0de87),
	.w4(32'hbb2f0cc0),
	.w5(32'hba5c22cc),
	.w6(32'h395b5ee4),
	.w7(32'hbb6ef66b),
	.w8(32'hbb44dd76),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b0535),
	.w1(32'h3a8fb83e),
	.w2(32'h39dbf26f),
	.w3(32'hba8782ef),
	.w4(32'h3a625513),
	.w5(32'h3ae90705),
	.w6(32'hbaaa868f),
	.w7(32'h38a27f91),
	.w8(32'h3abccaa7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e237),
	.w1(32'hbb500411),
	.w2(32'hbb825cb5),
	.w3(32'hb9f7bfb8),
	.w4(32'hbba09961),
	.w5(32'hbb357ef7),
	.w6(32'h3b991283),
	.w7(32'hbb15bc70),
	.w8(32'hbbf147e8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaedfaa),
	.w1(32'hbc10b59f),
	.w2(32'hbb06ddd0),
	.w3(32'hbadf16a9),
	.w4(32'hbbb28140),
	.w5(32'hbb5d5357),
	.w6(32'h3a3ccd91),
	.w7(32'hbb8a9392),
	.w8(32'hbba5d767),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba460de),
	.w1(32'h3b1a0b57),
	.w2(32'h3b04e579),
	.w3(32'hbbbc0842),
	.w4(32'h3aed73de),
	.w5(32'h3959a5aa),
	.w6(32'hbbaf0a9b),
	.w7(32'h3b078e08),
	.w8(32'h38a035a9),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26f75a),
	.w1(32'hb98ab1ed),
	.w2(32'hbba1179b),
	.w3(32'hb8e8e383),
	.w4(32'hbb9cc785),
	.w5(32'hbbbe037f),
	.w6(32'h3b5d0e06),
	.w7(32'hbb2b9586),
	.w8(32'hbbfd84f1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0be25e),
	.w1(32'h3b3f2a64),
	.w2(32'h3896613e),
	.w3(32'hbbbfe891),
	.w4(32'hbb1b6858),
	.w5(32'hbaff091c),
	.w6(32'hbc157d89),
	.w7(32'hbc383de9),
	.w8(32'hbc3bd7f3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4612e5),
	.w1(32'h3af6f518),
	.w2(32'h3b0debdd),
	.w3(32'hbb28bfb9),
	.w4(32'h3b252aa5),
	.w5(32'h3b6aaef9),
	.w6(32'hbbcabbdc),
	.w7(32'h3a87bb42),
	.w8(32'h3a034e00),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0db6b),
	.w1(32'h3a5677a9),
	.w2(32'hba60e456),
	.w3(32'h38e10a65),
	.w4(32'h38eb8d9f),
	.w5(32'hba84e2a9),
	.w6(32'h3a36644e),
	.w7(32'h3a461a8e),
	.w8(32'h37a56777),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba762f48),
	.w1(32'hbac44189),
	.w2(32'h3997e011),
	.w3(32'hbac34423),
	.w4(32'hba848653),
	.w5(32'h3aae4473),
	.w6(32'h37c0b21e),
	.w7(32'hbadb4a09),
	.w8(32'hba69aba3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba577f59),
	.w1(32'h3ae69435),
	.w2(32'h3ae12045),
	.w3(32'hba510ca6),
	.w4(32'h3b09b93d),
	.w5(32'h3b0d2732),
	.w6(32'hbb16cdf3),
	.w7(32'h39348be7),
	.w8(32'h39d8b5d5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a139349),
	.w1(32'h3b3e500e),
	.w2(32'h38ab7de8),
	.w3(32'h3b766bf8),
	.w4(32'h3a5624eb),
	.w5(32'hba5cdbf3),
	.w6(32'h3ac3434a),
	.w7(32'h3aedf3ef),
	.w8(32'hbb1f9a38),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de56ae),
	.w1(32'hba1c728b),
	.w2(32'hbb199f3f),
	.w3(32'h39976be9),
	.w4(32'hb78bce75),
	.w5(32'hbb555037),
	.w6(32'h3ac7b729),
	.w7(32'h3aed2342),
	.w8(32'h3abb1cc5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ecc76),
	.w1(32'hbbe2b6c4),
	.w2(32'hbb3e4051),
	.w3(32'hbbb4c5fd),
	.w4(32'hbbc9e87d),
	.w5(32'hba91573c),
	.w6(32'hbae75c9f),
	.w7(32'hbc011442),
	.w8(32'hbb630650),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb838b85),
	.w1(32'hbb5d9fba),
	.w2(32'hbb464d8a),
	.w3(32'hbaeb1bf5),
	.w4(32'hbb88d6da),
	.w5(32'hbaf0776c),
	.w6(32'hbb50c3c9),
	.w7(32'hbba24ce0),
	.w8(32'hbb461000),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c98e1),
	.w1(32'h3bf5fbbf),
	.w2(32'h3b5b1ef1),
	.w3(32'hbb507400),
	.w4(32'h3c0b4451),
	.w5(32'hbb21dac2),
	.w6(32'hbada60a8),
	.w7(32'h3c1780b6),
	.w8(32'hbb285a49),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a4875),
	.w1(32'hbafe87e6),
	.w2(32'hba83e086),
	.w3(32'hbb90682b),
	.w4(32'hbaa201b0),
	.w5(32'h3afc92b3),
	.w6(32'hbac1571a),
	.w7(32'hbc19e12e),
	.w8(32'hbbd85e56),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f624c),
	.w1(32'hbbb57168),
	.w2(32'hbb8a4f0c),
	.w3(32'hbb9383e7),
	.w4(32'h3950f8da),
	.w5(32'h3cc494a6),
	.w6(32'hbb38912b),
	.w7(32'h3bd0c832),
	.w8(32'h3b42421d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbcb38),
	.w1(32'hbbe20102),
	.w2(32'hbc2262e8),
	.w3(32'h3c81e999),
	.w4(32'hbbc03028),
	.w5(32'hbc4b2d29),
	.w6(32'hbbc63d65),
	.w7(32'hbbc305f3),
	.w8(32'hbaf1f19c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37da12),
	.w1(32'h3a3fe842),
	.w2(32'h3b209e44),
	.w3(32'hba1691a4),
	.w4(32'hbb993702),
	.w5(32'hbb279ec4),
	.w6(32'hb9bcdb1b),
	.w7(32'h3a29f489),
	.w8(32'h3b89dbb2),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebf290),
	.w1(32'h3bbe3334),
	.w2(32'hbbb57388),
	.w3(32'hbbab29a3),
	.w4(32'h38b2327d),
	.w5(32'hbace059b),
	.w6(32'h399a166b),
	.w7(32'hbaf7de6e),
	.w8(32'hbc211722),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9849f68),
	.w1(32'hb9b25927),
	.w2(32'h3b94b9a9),
	.w3(32'hbb48944a),
	.w4(32'h3970e886),
	.w5(32'h3a988883),
	.w6(32'hbc1aa9f1),
	.w7(32'hbbce8604),
	.w8(32'hbbd6a301),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a55e),
	.w1(32'h3b9940c9),
	.w2(32'h3bc5986d),
	.w3(32'hba68537e),
	.w4(32'h3bd2c1ef),
	.w5(32'hbba5589e),
	.w6(32'hbb53bdb4),
	.w7(32'h3bc81793),
	.w8(32'h3b88996d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d8800),
	.w1(32'h3afe94e6),
	.w2(32'h3b27914d),
	.w3(32'hba3274cc),
	.w4(32'h3ab14b12),
	.w5(32'hbc0a695a),
	.w6(32'h3b8e7d25),
	.w7(32'h3b984c09),
	.w8(32'hbb1de968),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6df6d1),
	.w1(32'h3b646ec1),
	.w2(32'hbaa675f2),
	.w3(32'hbaa9ca18),
	.w4(32'h3affb13f),
	.w5(32'h3c17aa2a),
	.w6(32'hb9fca27c),
	.w7(32'h390ab94c),
	.w8(32'h3b145c39),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b4ac5),
	.w1(32'h3b31930c),
	.w2(32'h3bbdd778),
	.w3(32'h3bdb46f6),
	.w4(32'h3b695874),
	.w5(32'h3b18394b),
	.w6(32'h3b014a9a),
	.w7(32'hbaff7830),
	.w8(32'hbb08f1c9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd3f18),
	.w1(32'h3be61db0),
	.w2(32'h3b9e7c7a),
	.w3(32'h3beb430d),
	.w4(32'h3b2a03e8),
	.w5(32'hb8921398),
	.w6(32'hbad315f4),
	.w7(32'h3c0e7512),
	.w8(32'h3b199dfe),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24d681),
	.w1(32'h39db804e),
	.w2(32'hba42cfe3),
	.w3(32'h3bae79a4),
	.w4(32'h3897ea4f),
	.w5(32'hba65e27b),
	.w6(32'h3b663eba),
	.w7(32'hba20d8dd),
	.w8(32'hbb432c4c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50ce7d),
	.w1(32'hbbb30132),
	.w2(32'hbb178aab),
	.w3(32'hbbd4fab0),
	.w4(32'hbb18327a),
	.w5(32'h3c98a452),
	.w6(32'hbb32abd0),
	.w7(32'h3be4ab31),
	.w8(32'h3baf7045),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89d03d),
	.w1(32'h3c00eb23),
	.w2(32'h3c597d6c),
	.w3(32'h3c9efc54),
	.w4(32'h3c2dd426),
	.w5(32'h3c44cdc9),
	.w6(32'h384501ab),
	.w7(32'h3bfd1faf),
	.w8(32'h3bc50f24),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd91454),
	.w1(32'hbb4ae60a),
	.w2(32'hbc0e8be9),
	.w3(32'h3c09a55e),
	.w4(32'h3a646c1e),
	.w5(32'hbb415a9d),
	.w6(32'h3c13d302),
	.w7(32'hba113ec1),
	.w8(32'hbc2ce56e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80a5d3),
	.w1(32'h3ad61484),
	.w2(32'hbb70e472),
	.w3(32'hb98cba50),
	.w4(32'hbb3db405),
	.w5(32'h3be30508),
	.w6(32'h3a4b06d7),
	.w7(32'h3b0c5dfc),
	.w8(32'hbb11480e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa17fc),
	.w1(32'h3b0ed91a),
	.w2(32'hbc0a7ff5),
	.w3(32'h3845d029),
	.w4(32'hbbae1f46),
	.w5(32'hbc5bc68c),
	.w6(32'h3c39311d),
	.w7(32'hbc320713),
	.w8(32'hbc360252),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba881d4),
	.w1(32'h3ae4f1df),
	.w2(32'hbaa5df08),
	.w3(32'hbc0a4985),
	.w4(32'h3aa53259),
	.w5(32'h3b1835e5),
	.w6(32'hbb94c2e0),
	.w7(32'hba0707e5),
	.w8(32'h3b105a3b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba939c43),
	.w1(32'h3b06312a),
	.w2(32'hba3578cc),
	.w3(32'hbb1efe9c),
	.w4(32'h3ad59507),
	.w5(32'hbb11b4d7),
	.w6(32'hb9cdbd9c),
	.w7(32'h39a29b32),
	.w8(32'hbb79d8f5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf4a82),
	.w1(32'h3c032b4d),
	.w2(32'h3c601163),
	.w3(32'h3bd25b75),
	.w4(32'h3c34081c),
	.w5(32'h3bd1c519),
	.w6(32'hba02d7d1),
	.w7(32'h3b005df5),
	.w8(32'h3c2e042b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4321de),
	.w1(32'hb98c8fda),
	.w2(32'h3a9269b9),
	.w3(32'h3bd0d316),
	.w4(32'hbbb1bc8b),
	.w5(32'hbb965323),
	.w6(32'h3c1990ee),
	.w7(32'hbb268665),
	.w8(32'hbb8666b9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5749ae),
	.w1(32'h3bafa543),
	.w2(32'h3a87a88d),
	.w3(32'hba3f4928),
	.w4(32'hbb434ff1),
	.w5(32'hbc1d7a7e),
	.w6(32'h3b8b3dae),
	.w7(32'h3b1c1a2d),
	.w8(32'h3b65bf92),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab7857),
	.w1(32'h39130d9a),
	.w2(32'h3b8806c4),
	.w3(32'hbb576d32),
	.w4(32'hbae4cb01),
	.w5(32'h3c844e97),
	.w6(32'hbaabfc86),
	.w7(32'h3b5d4435),
	.w8(32'hbb269f5c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad1b98),
	.w1(32'h3b4bc66b),
	.w2(32'hbb286b50),
	.w3(32'h3bbfe192),
	.w4(32'hbb6ecdb0),
	.w5(32'hbc09a9a3),
	.w6(32'hbc427e0c),
	.w7(32'hbb284888),
	.w8(32'hbb271c01),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcce1ee),
	.w1(32'hbb0c922f),
	.w2(32'hbb0f18b3),
	.w3(32'hbc008992),
	.w4(32'h3b5b633e),
	.w5(32'h3c023754),
	.w6(32'hbb3f830b),
	.w7(32'hbbbc8a0a),
	.w8(32'hbc351514),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4b80b),
	.w1(32'hbb9618e2),
	.w2(32'h3ad9c451),
	.w3(32'h3c27a247),
	.w4(32'hbb2304e0),
	.w5(32'hbae15d13),
	.w6(32'h3b8183a8),
	.w7(32'h3b8996ad),
	.w8(32'h3c014037),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf30e08),
	.w1(32'h3b532ef7),
	.w2(32'h3a9ab2ad),
	.w3(32'h39e348dd),
	.w4(32'h3aa72a76),
	.w5(32'h3b569b87),
	.w6(32'hbb8653a0),
	.w7(32'h3a5274e6),
	.w8(32'h3b9356d2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafab086),
	.w1(32'hbbb5dc58),
	.w2(32'hbb7137b5),
	.w3(32'hbaecf888),
	.w4(32'hbbb19458),
	.w5(32'hbb7b650e),
	.w6(32'h3bc14a29),
	.w7(32'hbbf8229b),
	.w8(32'h3ab431e7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b728637),
	.w1(32'h3a8effec),
	.w2(32'h3ab50ad8),
	.w3(32'h3b2f269b),
	.w4(32'hb8b094eb),
	.w5(32'hbb851b90),
	.w6(32'h390747d2),
	.w7(32'hbb028eea),
	.w8(32'hbbeec7d5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add540e),
	.w1(32'h3b81d3f8),
	.w2(32'h3bd95509),
	.w3(32'hbbe8c5a4),
	.w4(32'hbaeca4bb),
	.w5(32'hbae58272),
	.w6(32'h37ce1ebb),
	.w7(32'hbc074f3a),
	.w8(32'hbb91d537),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e94bc),
	.w1(32'h3b431a39),
	.w2(32'h3b17765e),
	.w3(32'h3b287296),
	.w4(32'hba47f515),
	.w5(32'hb8e6a700),
	.w6(32'h3b1e7df0),
	.w7(32'h39f8b009),
	.w8(32'h3b2b52c2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a3d1c),
	.w1(32'hbaeae57a),
	.w2(32'hbc197c8b),
	.w3(32'hbbbd9a80),
	.w4(32'hbb838395),
	.w5(32'hbc2bacbd),
	.w6(32'h3b143133),
	.w7(32'hbb8ff002),
	.w8(32'hbbe6159e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc016ef2),
	.w1(32'hbb7a0437),
	.w2(32'hbc13c22d),
	.w3(32'h3a8be66a),
	.w4(32'h3a4f882f),
	.w5(32'h3c885a1f),
	.w6(32'h3b39bbe2),
	.w7(32'h3c3c2dc4),
	.w8(32'h3b44d2ff),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b379504),
	.w1(32'hbbb515ec),
	.w2(32'hbb8032a0),
	.w3(32'h3c0c9f2e),
	.w4(32'hbba7f211),
	.w5(32'hbc0b985e),
	.w6(32'h3a274f41),
	.w7(32'hbace354a),
	.w8(32'hbbc9fa91),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16fb27),
	.w1(32'hbbd05d2c),
	.w2(32'hbbd51ed1),
	.w3(32'hb970a4c5),
	.w4(32'hbbe1f852),
	.w5(32'h3c94f805),
	.w6(32'h3b9019a2),
	.w7(32'hbbd9f823),
	.w8(32'hbb4762df),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb973503f),
	.w1(32'hba5a20aa),
	.w2(32'hbb9ef82e),
	.w3(32'h3bf73551),
	.w4(32'hba28f4f1),
	.w5(32'h3ba63a9d),
	.w6(32'hbb33f342),
	.w7(32'h392c0ed7),
	.w8(32'h3b229f54),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaa543),
	.w1(32'h3bdffcc8),
	.w2(32'h3b4a88ff),
	.w3(32'h3ae0de87),
	.w4(32'h3ba8b24e),
	.w5(32'h3b86b2bf),
	.w6(32'hba1c5f30),
	.w7(32'h39abc6cf),
	.w8(32'hbb35a0a7),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79ee32),
	.w1(32'hbac8093f),
	.w2(32'h3a3764b7),
	.w3(32'h3b187d6e),
	.w4(32'h3b33ec61),
	.w5(32'h38ed853a),
	.w6(32'h3a9f9cb2),
	.w7(32'h3ad44943),
	.w8(32'hbb8be501),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61a964),
	.w1(32'h3ac69fa5),
	.w2(32'hb9be61a8),
	.w3(32'hbb0b43a8),
	.w4(32'h3b6a55d5),
	.w5(32'h3c5ca663),
	.w6(32'h3b0ce714),
	.w7(32'h3be906d8),
	.w8(32'h3b050fb6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab35c68),
	.w1(32'hb9238773),
	.w2(32'hbb97cd55),
	.w3(32'h3bdb3aeb),
	.w4(32'hbbf4cbad),
	.w5(32'hbbe95544),
	.w6(32'hbb3132b5),
	.w7(32'hbaeeab88),
	.w8(32'hbb4721fe),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba81f97),
	.w1(32'hbb5d49ae),
	.w2(32'hbb14feaa),
	.w3(32'h3a840bb3),
	.w4(32'hbb477c7d),
	.w5(32'h3bb89309),
	.w6(32'hba695a5c),
	.w7(32'hba98acfd),
	.w8(32'h3b80e1e8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32cdb5),
	.w1(32'h3c0d0d38),
	.w2(32'hbba3bb6e),
	.w3(32'h3bf825d0),
	.w4(32'hba5964db),
	.w5(32'hbb5e55ff),
	.w6(32'h3bcb98e7),
	.w7(32'hbb0fd641),
	.w8(32'hbaa40a85),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe096e),
	.w1(32'hba889c0b),
	.w2(32'hbb71bf40),
	.w3(32'h3bc89365),
	.w4(32'hbbb1984d),
	.w5(32'hbab3cdea),
	.w6(32'h3b129ee5),
	.w7(32'hbb321773),
	.w8(32'h39b50ee2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937567),
	.w1(32'h3baf768e),
	.w2(32'h3b99009a),
	.w3(32'hbb95327d),
	.w4(32'h3b64c6b9),
	.w5(32'hbc749c7d),
	.w6(32'h3b8dccb8),
	.w7(32'hbb82cede),
	.w8(32'hbc3c3f77),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6c0f8),
	.w1(32'hbac52589),
	.w2(32'h3bb3fcbb),
	.w3(32'hbc698fe7),
	.w4(32'h3bda1637),
	.w5(32'h3c1a7d43),
	.w6(32'hba5f1be0),
	.w7(32'h3b1c33bd),
	.w8(32'h3b5e6f39),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b913b7c),
	.w1(32'h3b3fcb0d),
	.w2(32'h3b5349eb),
	.w3(32'h3c1f6398),
	.w4(32'h3b41c1e1),
	.w5(32'h3b5bbef3),
	.w6(32'hbafef708),
	.w7(32'h3b7261e1),
	.w8(32'h3b66058f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82cc48),
	.w1(32'hbb3048bd),
	.w2(32'h3b57ab34),
	.w3(32'hbb8c1b5e),
	.w4(32'h3b551193),
	.w5(32'h3b0e64d2),
	.w6(32'h3a565203),
	.w7(32'h3a6741f3),
	.w8(32'h3b99aa00),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc012cb),
	.w1(32'h3be4ffbc),
	.w2(32'hba0fee82),
	.w3(32'h3abe3853),
	.w4(32'h3b1635a7),
	.w5(32'hb9afe744),
	.w6(32'hbbb8bae8),
	.w7(32'h3b5587a0),
	.w8(32'h3ae9bc2c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4be6b),
	.w1(32'hbbf68b46),
	.w2(32'hbba7fd5a),
	.w3(32'hbbbef89d),
	.w4(32'hbc454f47),
	.w5(32'hbbe275b6),
	.w6(32'hbb2fb8c4),
	.w7(32'hb9fb4a84),
	.w8(32'hbb427e09),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad22a42),
	.w1(32'hbbbb972e),
	.w2(32'hbbc95b2e),
	.w3(32'hbb2e68c0),
	.w4(32'hbb805725),
	.w5(32'h3c34119a),
	.w6(32'h3b378a63),
	.w7(32'h3b7233b5),
	.w8(32'h3c055883),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae87dd),
	.w1(32'h3bf3875d),
	.w2(32'h3bba4a13),
	.w3(32'h3c261492),
	.w4(32'h3b82da06),
	.w5(32'h3b4c8bac),
	.w6(32'h3b2146c4),
	.w7(32'h3b89ac80),
	.w8(32'h3b7ddf15),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ece5e),
	.w1(32'hbb6fc120),
	.w2(32'hbb274ce7),
	.w3(32'hba9790a0),
	.w4(32'h3b9ec0a2),
	.w5(32'h3b62eb7e),
	.w6(32'h39cd6a0b),
	.w7(32'h3a9bcd1c),
	.w8(32'hba7e24bb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe317e),
	.w1(32'hbae92fc5),
	.w2(32'hbaa53c63),
	.w3(32'hbbeb3731),
	.w4(32'hb9c2e827),
	.w5(32'h3c58b52c),
	.w6(32'h3a6519cc),
	.w7(32'hbb9ce750),
	.w8(32'hb9b70003),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81404c),
	.w1(32'h3a404cbf),
	.w2(32'hbb8a8cb2),
	.w3(32'hba0fe000),
	.w4(32'hbba301fc),
	.w5(32'hbc439997),
	.w6(32'h3aa01ae1),
	.w7(32'hbbe9c914),
	.w8(32'hbbe0d650),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd79481),
	.w1(32'hb99e8907),
	.w2(32'hbb9cd272),
	.w3(32'hbbea8203),
	.w4(32'hbb8e0b91),
	.w5(32'h3baf91f7),
	.w6(32'hb9f31dab),
	.w7(32'hbb92907a),
	.w8(32'hbc429b8f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc214e7c),
	.w1(32'h395dda92),
	.w2(32'hbc032d41),
	.w3(32'hbc0479e6),
	.w4(32'hbbfdef95),
	.w5(32'h3c43695c),
	.w6(32'hbc5ce4dc),
	.w7(32'hbc0825a6),
	.w8(32'hbbc14080),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeecfd),
	.w1(32'hbb025e57),
	.w2(32'h3a845d83),
	.w3(32'h3b8340b1),
	.w4(32'h3acd7807),
	.w5(32'hbaf5f3b1),
	.w6(32'h3a999362),
	.w7(32'hbabf5d34),
	.w8(32'hbba9f1fc),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea4ed9),
	.w1(32'h3b846e35),
	.w2(32'hbbc1ac14),
	.w3(32'hbb80ab95),
	.w4(32'h38e4d416),
	.w5(32'h394dcdfd),
	.w6(32'hbbf2f5a9),
	.w7(32'hbba78dba),
	.w8(32'hbc249cc1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule