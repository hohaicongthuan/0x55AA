module layer_10_featuremap_464(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0ab05),
	.w1(32'h3b4162b5),
	.w2(32'h3b0e98b1),
	.w3(32'h3b5b1d21),
	.w4(32'h3b125aee),
	.w5(32'h3ae7d1f6),
	.w6(32'hbafeebf2),
	.w7(32'h39544a37),
	.w8(32'h3a2899e8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeb65e),
	.w1(32'hba5771e8),
	.w2(32'h3c1058d3),
	.w3(32'h3b1925c7),
	.w4(32'hbbb639a3),
	.w5(32'h3b179804),
	.w6(32'h382897e1),
	.w7(32'hbbf050c6),
	.w8(32'h3b787295),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb741023),
	.w1(32'hbc1bfc12),
	.w2(32'hbaa0773d),
	.w3(32'h3a28861c),
	.w4(32'h3b0c3681),
	.w5(32'hbb075fbb),
	.w6(32'hba9dd063),
	.w7(32'hb8fd4ac1),
	.w8(32'h3bed336d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1eaef5),
	.w1(32'hbb260b74),
	.w2(32'hbb3152f3),
	.w3(32'hbbb1f330),
	.w4(32'h3b43a39d),
	.w5(32'hbc0424e5),
	.w6(32'hb9c95515),
	.w7(32'h3b3d4dec),
	.w8(32'hbacbed83),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2742f6),
	.w1(32'hbae06b89),
	.w2(32'hbb4dd619),
	.w3(32'hbb9ac76c),
	.w4(32'h3ae0ca19),
	.w5(32'h3c3c65ff),
	.w6(32'h3ac08ecf),
	.w7(32'hbbc508ff),
	.w8(32'hba96f8b2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e6190),
	.w1(32'h3acf3a45),
	.w2(32'h3b8ced8d),
	.w3(32'h3b3f681a),
	.w4(32'hba5a58ac),
	.w5(32'hba9fc2f0),
	.w6(32'h3bcafd77),
	.w7(32'hbb4e4ea7),
	.w8(32'hbb878aa3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d0ebb),
	.w1(32'h3aef1ee5),
	.w2(32'h3bc4cce6),
	.w3(32'hbaf167b5),
	.w4(32'h3bbc393d),
	.w5(32'h3bb2f356),
	.w6(32'h39997b18),
	.w7(32'h3b75b950),
	.w8(32'h3a66e93e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf6036),
	.w1(32'h3baddd96),
	.w2(32'h3c3aeab1),
	.w3(32'h3c76dc2e),
	.w4(32'h3bcc3886),
	.w5(32'hbbb90fa6),
	.w6(32'h3bdf1945),
	.w7(32'h3bda05cb),
	.w8(32'h3b589023),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f05ba),
	.w1(32'hbba72001),
	.w2(32'hbc039338),
	.w3(32'h3ae2258e),
	.w4(32'hba625276),
	.w5(32'h3aa231c3),
	.w6(32'hbb8ef97e),
	.w7(32'h3b3183ae),
	.w8(32'hbbca6c9e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ced3),
	.w1(32'h379876e3),
	.w2(32'hbb2f9228),
	.w3(32'h39e6cb2c),
	.w4(32'h3c06ffc5),
	.w5(32'h3bdf412e),
	.w6(32'hbba53afe),
	.w7(32'h3b37ac56),
	.w8(32'hba06bb94),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b191d09),
	.w1(32'h39643552),
	.w2(32'hbbd7de4e),
	.w3(32'h3949c3d1),
	.w4(32'hbbb58cfa),
	.w5(32'h3b80db7b),
	.w6(32'hbadbee96),
	.w7(32'hbb7b3664),
	.w8(32'hbbbdaa16),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b23e0),
	.w1(32'hbb82ff95),
	.w2(32'h3b8af300),
	.w3(32'hba8fad8d),
	.w4(32'h3b4bc566),
	.w5(32'h3bdd5037),
	.w6(32'hbbb58b53),
	.w7(32'h3b8112e1),
	.w8(32'h3b4f5f99),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aad617),
	.w1(32'hbb5c2c25),
	.w2(32'h3b16b632),
	.w3(32'h3b322d80),
	.w4(32'h3b566941),
	.w5(32'hbc206172),
	.w6(32'h3b578bcf),
	.w7(32'h3b33b8f3),
	.w8(32'h3bdd3c5d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb5646),
	.w1(32'h3b77c2c9),
	.w2(32'hbbb381f9),
	.w3(32'hbb90dbfb),
	.w4(32'h3c28c1a3),
	.w5(32'h3cdb413c),
	.w6(32'hbba144d1),
	.w7(32'hbbdb41c4),
	.w8(32'h3b23dc80),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf10438),
	.w1(32'h3a37c9d3),
	.w2(32'hbbd246c3),
	.w3(32'hb93424d2),
	.w4(32'hbb29a7f5),
	.w5(32'h3c2d919d),
	.w6(32'h3c403117),
	.w7(32'hbb349f03),
	.w8(32'hbb0831c5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f017b),
	.w1(32'h3994a29e),
	.w2(32'hbb086a7f),
	.w3(32'h3bcdbdc6),
	.w4(32'h3a8c7ad8),
	.w5(32'hbb97ecf0),
	.w6(32'h3c1afe04),
	.w7(32'h3b8fa145),
	.w8(32'h3b6343f3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a89b3),
	.w1(32'h3c34bef8),
	.w2(32'h3a987eae),
	.w3(32'hbb4fbe92),
	.w4(32'h3c069abf),
	.w5(32'h3c6d361f),
	.w6(32'hbb3bd450),
	.w7(32'h3933246c),
	.w8(32'h388680da),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9816110),
	.w1(32'h3c09ce8f),
	.w2(32'h3bd33b50),
	.w3(32'h3c1423b1),
	.w4(32'h397efaaf),
	.w5(32'h3b8f1c34),
	.w6(32'h3c0d31e9),
	.w7(32'h3ba5a7a2),
	.w8(32'h3bf4d554),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcea58a),
	.w1(32'h3b3a84d0),
	.w2(32'h3b08846f),
	.w3(32'hbb047fc3),
	.w4(32'hbaa63fa8),
	.w5(32'h3babf92b),
	.w6(32'hbb6cb619),
	.w7(32'hb9f71100),
	.w8(32'hba89b7bd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a090b),
	.w1(32'h3cd07417),
	.w2(32'h3c6fcd30),
	.w3(32'h3ae71387),
	.w4(32'h3b9c68e2),
	.w5(32'h3ca43c2d),
	.w6(32'hbaadf006),
	.w7(32'hba1be1ed),
	.w8(32'hbb3e538a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc389e2),
	.w1(32'h3babae40),
	.w2(32'h3bbe39b7),
	.w3(32'h3c610a24),
	.w4(32'hbb27ae79),
	.w5(32'hbb5e8a65),
	.w6(32'h3be2e168),
	.w7(32'hba64f85d),
	.w8(32'hba8fcbd9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9bfac),
	.w1(32'h38ce7259),
	.w2(32'h3b78b1b5),
	.w3(32'h3aa511c8),
	.w4(32'hbb85df9a),
	.w5(32'hba8771c6),
	.w6(32'hba4f20d7),
	.w7(32'hbb38a18e),
	.w8(32'h3a6028bc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c3dd9),
	.w1(32'h3bf17f27),
	.w2(32'h3c22121b),
	.w3(32'h3b5b8384),
	.w4(32'h3a99ccda),
	.w5(32'h3c2f71d5),
	.w6(32'h3c1bb53f),
	.w7(32'h3ba4e460),
	.w8(32'h3c19d451),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beda1d1),
	.w1(32'hba3490d6),
	.w2(32'hbb9e8afd),
	.w3(32'h3bd33508),
	.w4(32'hb85891d8),
	.w5(32'hbbc753a0),
	.w6(32'h3ad1a48a),
	.w7(32'h3b9a8d64),
	.w8(32'h3b5c7423),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c5e7d),
	.w1(32'hbb451b3f),
	.w2(32'hbb95d264),
	.w3(32'h3b12d8fa),
	.w4(32'hbbb40e03),
	.w5(32'h3b521999),
	.w6(32'h3c045139),
	.w7(32'h3b0cfa1d),
	.w8(32'h3982d06b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac28980),
	.w1(32'h3b61b5ff),
	.w2(32'h3b3258a7),
	.w3(32'hbc0c84a9),
	.w4(32'h3b39f0cb),
	.w5(32'hba217d4a),
	.w6(32'hbacf2993),
	.w7(32'h3aab71a5),
	.w8(32'h3b23cedd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990d1a5),
	.w1(32'hb9388fea),
	.w2(32'hbafa8e45),
	.w3(32'h3b2ba68a),
	.w4(32'hbb628c5f),
	.w5(32'hbb427b0c),
	.w6(32'h3b742821),
	.w7(32'h399ee91c),
	.w8(32'hb98cfece),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00c6fb),
	.w1(32'h3b10d022),
	.w2(32'h3b288182),
	.w3(32'hbbd87fda),
	.w4(32'h3b80da53),
	.w5(32'h3b58b8e9),
	.w6(32'hbc05f263),
	.w7(32'h3ba56210),
	.w8(32'hba444a4d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e7987),
	.w1(32'h3b867ac3),
	.w2(32'h3c46e3ea),
	.w3(32'hbbef8b23),
	.w4(32'h3bdea99a),
	.w5(32'h3c2a9397),
	.w6(32'hbbe25732),
	.w7(32'hbb9955c3),
	.w8(32'h3912d5b7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4ad99),
	.w1(32'hbbdadfff),
	.w2(32'hbb1bacb1),
	.w3(32'h3bcc2150),
	.w4(32'h3a349165),
	.w5(32'hbbff8970),
	.w6(32'hba93cd89),
	.w7(32'h3b2dedf7),
	.w8(32'h3b87e673),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb23a79),
	.w1(32'h3ab2c144),
	.w2(32'hbc32f55e),
	.w3(32'h3bb1e8b5),
	.w4(32'hbaafa491),
	.w5(32'hbaac0e36),
	.w6(32'hba89cc54),
	.w7(32'hb99b5a6c),
	.w8(32'hbad272c7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e1be8),
	.w1(32'hbb8352b1),
	.w2(32'h3a379738),
	.w3(32'h3b71f866),
	.w4(32'h3a10c6c8),
	.w5(32'hbb348d23),
	.w6(32'h3ac19f57),
	.w7(32'h39c1e5e8),
	.w8(32'hba76c8d0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ce298),
	.w1(32'hba9b47ab),
	.w2(32'hba844915),
	.w3(32'h3b4aab32),
	.w4(32'h3c38204d),
	.w5(32'hba91cc40),
	.w6(32'hbada5e1b),
	.w7(32'h3b9363e2),
	.w8(32'h3b86688e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabe33c),
	.w1(32'hbb1d74b5),
	.w2(32'hbae6a83b),
	.w3(32'hbb2270fc),
	.w4(32'h3b5da824),
	.w5(32'h3ac45eda),
	.w6(32'h3b90c494),
	.w7(32'h3b9fe646),
	.w8(32'hb928e719),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0be238),
	.w1(32'h3ba5ee73),
	.w2(32'hba9f3c57),
	.w3(32'h3aa81631),
	.w4(32'h3962954f),
	.w5(32'hbbb585e9),
	.w6(32'hbb7740fb),
	.w7(32'h3bf516db),
	.w8(32'h3b03570a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87d834),
	.w1(32'h3b654b13),
	.w2(32'h3b7ebb51),
	.w3(32'hbb77d3b5),
	.w4(32'h3b120504),
	.w5(32'h3b4c36d7),
	.w6(32'hbad6296d),
	.w7(32'h3b82d610),
	.w8(32'h3baa2171),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14479f),
	.w1(32'h3b953d50),
	.w2(32'hbb603f47),
	.w3(32'h3ba814da),
	.w4(32'hbb5b00cc),
	.w5(32'h3b08a052),
	.w6(32'h3bae2bd0),
	.w7(32'hbc109209),
	.w8(32'hbbba0fda),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb53687),
	.w1(32'hbc25ba21),
	.w2(32'h3c16c022),
	.w3(32'h3b646d57),
	.w4(32'hbbfcbf83),
	.w5(32'h3b0cc877),
	.w6(32'h3bb61da3),
	.w7(32'hbbacc0ac),
	.w8(32'h3c352a9a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc618819),
	.w1(32'hbc098817),
	.w2(32'hbb247aa2),
	.w3(32'hbba70a47),
	.w4(32'hbb78d932),
	.w5(32'h3cb151e5),
	.w6(32'hbc1e2ce1),
	.w7(32'h3a815bb7),
	.w8(32'h3bd5cd36),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01eadb),
	.w1(32'hba3a0fef),
	.w2(32'h3b26cd65),
	.w3(32'hbaa07c27),
	.w4(32'hbb3639a3),
	.w5(32'hbb8d02a0),
	.w6(32'hbaac86db),
	.w7(32'h3ac2fa65),
	.w8(32'h3b5da14c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83f37f),
	.w1(32'hbbc478b8),
	.w2(32'hbb1fde4c),
	.w3(32'hbad929c7),
	.w4(32'hba8eebe4),
	.w5(32'hbbe8b194),
	.w6(32'hbaf340e5),
	.w7(32'hbc068253),
	.w8(32'hbb97a230),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99e2ef),
	.w1(32'h3a48e389),
	.w2(32'hbaadda98),
	.w3(32'hb97afe09),
	.w4(32'hba443ab7),
	.w5(32'hbacf87bc),
	.w6(32'h3bb3e3b0),
	.w7(32'h3a9ded51),
	.w8(32'hbb882474),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb82a0),
	.w1(32'h3b8103d4),
	.w2(32'h3bdd2af8),
	.w3(32'hbbcca7fa),
	.w4(32'h3c0a369e),
	.w5(32'hbb861ebb),
	.w6(32'hbb4c33b9),
	.w7(32'h3bb446b2),
	.w8(32'h3b709df1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5350e5),
	.w1(32'h3b2825ef),
	.w2(32'h3ab89c1c),
	.w3(32'h3af3b553),
	.w4(32'hbb749b04),
	.w5(32'hbc0c4e50),
	.w6(32'h3ab2104a),
	.w7(32'h3b5faa45),
	.w8(32'h3b47ae58),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b832ac5),
	.w1(32'hb96c2b70),
	.w2(32'h3a9c5402),
	.w3(32'hbb1151a4),
	.w4(32'hbb1751f9),
	.w5(32'hba3e92f3),
	.w6(32'h3b3a4a54),
	.w7(32'h3be91300),
	.w8(32'h3b73b065),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86d014),
	.w1(32'hbb8b7c3a),
	.w2(32'hbbfef3f3),
	.w3(32'hba8ad22b),
	.w4(32'hbb3867b3),
	.w5(32'hbb56f377),
	.w6(32'h3b060eb3),
	.w7(32'h3ba10892),
	.w8(32'hba100292),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b4fac),
	.w1(32'hbb3d583d),
	.w2(32'hbb8f0f3b),
	.w3(32'h3b0cb895),
	.w4(32'hbbacdb85),
	.w5(32'h3c1750c2),
	.w6(32'h3b1b7166),
	.w7(32'hba067d72),
	.w8(32'hbb205ecb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb680edc),
	.w1(32'h3b944a2e),
	.w2(32'h3b1f6b6c),
	.w3(32'hbb6e2b69),
	.w4(32'h3a4c942f),
	.w5(32'h3c1147a5),
	.w6(32'hbb3b733f),
	.w7(32'h3a99a2fa),
	.w8(32'h3c2bdf2e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd706e4),
	.w1(32'hba94cd41),
	.w2(32'hbb7f6c0f),
	.w3(32'hbb3304d3),
	.w4(32'hbac20c31),
	.w5(32'h3b12444c),
	.w6(32'h3ace0a94),
	.w7(32'h3b47ad75),
	.w8(32'hbb3d88bd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9355d6),
	.w1(32'hbb181862),
	.w2(32'hbad6013a),
	.w3(32'hbb12d0d0),
	.w4(32'h3acf7232),
	.w5(32'hbb0bf64a),
	.w6(32'hbadd2860),
	.w7(32'h3bbc0887),
	.w8(32'h3bb01911),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95670a),
	.w1(32'hbb46656c),
	.w2(32'h3bc8f07b),
	.w3(32'hba862d39),
	.w4(32'hbbac4b84),
	.w5(32'h3ab323d3),
	.w6(32'h3b20f37c),
	.w7(32'hbb923a81),
	.w8(32'hba848c82),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb323787),
	.w1(32'h3ba13434),
	.w2(32'h3ade4bfd),
	.w3(32'hba9059ab),
	.w4(32'hbb7a3ee0),
	.w5(32'h3bcf4a7f),
	.w6(32'h3b7aa1cd),
	.w7(32'hbba27a31),
	.w8(32'hba58dff4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc0e8d),
	.w1(32'h3a83f0cc),
	.w2(32'h3b47ef93),
	.w3(32'hba86b06d),
	.w4(32'h3a0ff56d),
	.w5(32'hbbee2921),
	.w6(32'h399bce16),
	.w7(32'h3b4cb969),
	.w8(32'hb9f23f37),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a5bf8),
	.w1(32'h3af1a4f4),
	.w2(32'h3c1b0408),
	.w3(32'h3b568aa5),
	.w4(32'hb9f984aa),
	.w5(32'hbb390211),
	.w6(32'h3a4e6761),
	.w7(32'h3bcbc74e),
	.w8(32'h3c1f395d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58dc1a),
	.w1(32'hba216dea),
	.w2(32'h3c02c39f),
	.w3(32'hbb1950f5),
	.w4(32'hbb849b7e),
	.w5(32'hb94be497),
	.w6(32'hbb8d34e3),
	.w7(32'hbaa2790b),
	.w8(32'h3ac5a6c0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabe82d),
	.w1(32'h3b8f65fe),
	.w2(32'h3c337065),
	.w3(32'h3b384783),
	.w4(32'h3aea59f2),
	.w5(32'h3be8a820),
	.w6(32'hbaacc039),
	.w7(32'hbb02d68e),
	.w8(32'h3c2ed892),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70054b),
	.w1(32'hbb04f7cd),
	.w2(32'h3aab8665),
	.w3(32'h3b3b794f),
	.w4(32'h39292ff1),
	.w5(32'hbaf5ac45),
	.w6(32'hbb32521d),
	.w7(32'hbab53595),
	.w8(32'hba6617c6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae65670),
	.w1(32'h3bb8c79d),
	.w2(32'hbbd9c2db),
	.w3(32'h3b5c7afd),
	.w4(32'h3bc4c87f),
	.w5(32'h3ba14787),
	.w6(32'h3a89ae5f),
	.w7(32'hbbd5ab26),
	.w8(32'h3bb70dc8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd015c),
	.w1(32'h39cd5763),
	.w2(32'h3bcf3278),
	.w3(32'hbb7e5bc5),
	.w4(32'h3a17f82e),
	.w5(32'h3bad5544),
	.w6(32'h3bd12575),
	.w7(32'h3a3f6ec3),
	.w8(32'h3bcd20fd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7106),
	.w1(32'hbafd49f0),
	.w2(32'hbc1126be),
	.w3(32'h3af6fcf6),
	.w4(32'hb96213ca),
	.w5(32'h3c4e8a96),
	.w6(32'h3bcfa675),
	.w7(32'hbab51bb8),
	.w8(32'h3b89a18f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc20f20),
	.w1(32'hb7b4a13e),
	.w2(32'hba6eb62a),
	.w3(32'hb964239c),
	.w4(32'hb9b6b1f3),
	.w5(32'h3bbde5d3),
	.w6(32'h3b24277f),
	.w7(32'h3b970cf4),
	.w8(32'h3bb4ef42),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2a16d),
	.w1(32'h3b8c9851),
	.w2(32'h3bb11d37),
	.w3(32'h3b0ffb18),
	.w4(32'h3b486e27),
	.w5(32'h3c32d40f),
	.w6(32'hbaa75e47),
	.w7(32'h3bca9101),
	.w8(32'h3b2d199c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b957f39),
	.w1(32'h3bbb4532),
	.w2(32'h3b4b6a40),
	.w3(32'h3bcde42c),
	.w4(32'h3b3f0940),
	.w5(32'hbbf4a602),
	.w6(32'h3b980cc1),
	.w7(32'h3bbdfd8b),
	.w8(32'h3b95e0e1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcee03),
	.w1(32'h3a457091),
	.w2(32'h3ad70e7e),
	.w3(32'hbbc222d7),
	.w4(32'h3ac63f67),
	.w5(32'hb7e3176f),
	.w6(32'hba6a7867),
	.w7(32'h399d877b),
	.w8(32'h3a739e15),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa71ab3),
	.w1(32'h3af33ea3),
	.w2(32'h3b644f24),
	.w3(32'h3ab2a45b),
	.w4(32'h3af737ba),
	.w5(32'hbb42c603),
	.w6(32'h3b4cc2ee),
	.w7(32'h3ba6bb84),
	.w8(32'h3b39cb44),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd6b2b),
	.w1(32'h3b08338d),
	.w2(32'hbb72dfeb),
	.w3(32'h3bb19dc7),
	.w4(32'hbae0c0e6),
	.w5(32'h3bc2e573),
	.w6(32'h3adac5ca),
	.w7(32'h3ba800be),
	.w8(32'hbb349550),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b960639),
	.w1(32'h3b35ef06),
	.w2(32'h3c2b55dd),
	.w3(32'h3b86df79),
	.w4(32'hbb7078ff),
	.w5(32'h39d785ca),
	.w6(32'h3b5f53f3),
	.w7(32'h3a919393),
	.w8(32'h3b29c81b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95634c),
	.w1(32'h39d2db4c),
	.w2(32'hb94b83c0),
	.w3(32'h39af752e),
	.w4(32'hbab6bf2e),
	.w5(32'h3ba56d0a),
	.w6(32'h3b8e2b51),
	.w7(32'h3b161835),
	.w8(32'h3b88d701),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39e32b),
	.w1(32'h3b1425b5),
	.w2(32'h3c241ac0),
	.w3(32'hb9125c30),
	.w4(32'hbb60cc35),
	.w5(32'h3c04423c),
	.w6(32'h3b0384d1),
	.w7(32'hba964b6f),
	.w8(32'h3c0064bb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28291c),
	.w1(32'h3b8b5ed9),
	.w2(32'h3bcc0ca2),
	.w3(32'hba9977e6),
	.w4(32'h3b451e8c),
	.w5(32'h3bdae85c),
	.w6(32'h3b4555fc),
	.w7(32'h3bf00e0b),
	.w8(32'h3c464caf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc3dc4),
	.w1(32'h3b526e61),
	.w2(32'hba502829),
	.w3(32'hbbd01fb5),
	.w4(32'h3c166ddb),
	.w5(32'h3bc9c9e8),
	.w6(32'h3b9e0742),
	.w7(32'h3b3d1869),
	.w8(32'hbb49367e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81c522),
	.w1(32'h3b97f515),
	.w2(32'h3b0924ab),
	.w3(32'h3b253aea),
	.w4(32'hbb413e17),
	.w5(32'hbac79590),
	.w6(32'hbb1f13de),
	.w7(32'hbbb4ef04),
	.w8(32'hba82af20),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98e336),
	.w1(32'h3aa0c510),
	.w2(32'h3c3b0546),
	.w3(32'h3a56b0bf),
	.w4(32'hbaddbb38),
	.w5(32'h3c65b695),
	.w6(32'h3c261092),
	.w7(32'h3b87d477),
	.w8(32'h3c16fd70),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01316b),
	.w1(32'h3b3d6483),
	.w2(32'hba0d16c0),
	.w3(32'hba9f6566),
	.w4(32'hbae30780),
	.w5(32'hba13aeba),
	.w6(32'h3c0423b9),
	.w7(32'h3ad1e76d),
	.w8(32'h3b55a8ef),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f55ca6),
	.w1(32'hbbc81fa8),
	.w2(32'hbbd68fcc),
	.w3(32'h3b92b627),
	.w4(32'hbbe9f142),
	.w5(32'hba83213c),
	.w6(32'hbb4f3913),
	.w7(32'hbb42582c),
	.w8(32'hbb82751b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de2e88),
	.w1(32'h3b2386e2),
	.w2(32'h3bac873b),
	.w3(32'hbb03dd69),
	.w4(32'h3bbaab0e),
	.w5(32'h3bc20bf2),
	.w6(32'h3bd695a3),
	.w7(32'h3bf7fb07),
	.w8(32'h3bde6f24),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b926a47),
	.w1(32'h3af484d3),
	.w2(32'h3b060e22),
	.w3(32'hb9055083),
	.w4(32'h3b94a7e9),
	.w5(32'hba214ac2),
	.w6(32'h3b0e600f),
	.w7(32'h3a560f62),
	.w8(32'hb9e6f0d0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b055402),
	.w1(32'h3b92c168),
	.w2(32'h39b6a5b5),
	.w3(32'h3b55d9b5),
	.w4(32'h3b65afbf),
	.w5(32'h3b9d2dea),
	.w6(32'h3bc2f188),
	.w7(32'h38a395bd),
	.w8(32'h3c26e6d8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ec1b6),
	.w1(32'hba53be04),
	.w2(32'h3b42eaf0),
	.w3(32'hbb3a93e2),
	.w4(32'hbb050eb1),
	.w5(32'h3bee456f),
	.w6(32'h3bcc7593),
	.w7(32'h3ae65c3f),
	.w8(32'h3bb23cae),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45d030),
	.w1(32'h3b646bec),
	.w2(32'h3b36f5d6),
	.w3(32'hbb91f2e5),
	.w4(32'h3be1150a),
	.w5(32'hbb526e0a),
	.w6(32'hba67b7ef),
	.w7(32'h3bd1c636),
	.w8(32'h3a2b58ba),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02bd41),
	.w1(32'h3b6fe37b),
	.w2(32'hb9b0f47b),
	.w3(32'h3bd3d62c),
	.w4(32'h39fbd90f),
	.w5(32'hbc14e6b5),
	.w6(32'hbb95f5f1),
	.w7(32'h3b205581),
	.w8(32'hbb7f7f21),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b949aa1),
	.w1(32'h3b8d4d97),
	.w2(32'h3b0f5264),
	.w3(32'h3ba603a3),
	.w4(32'h3bc721cb),
	.w5(32'h3b62ad0b),
	.w6(32'h398b1452),
	.w7(32'h3bad2c96),
	.w8(32'h3bdf785c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9beec),
	.w1(32'hbb488675),
	.w2(32'hba0b74b6),
	.w3(32'hbb6ea55e),
	.w4(32'hbc068cfb),
	.w5(32'h39d9e9ff),
	.w6(32'hbb695fc6),
	.w7(32'hbb027947),
	.w8(32'h3aad9106),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74a004),
	.w1(32'h3b56534a),
	.w2(32'hba5be041),
	.w3(32'h3bc1bb6e),
	.w4(32'h3bca2a8d),
	.w5(32'h3caa0e63),
	.w6(32'hba0463ac),
	.w7(32'h3becb481),
	.w8(32'h3be3b6ab),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fe34c),
	.w1(32'h3ba90314),
	.w2(32'h3b9a2579),
	.w3(32'h3c0d50d2),
	.w4(32'h3b8c1d70),
	.w5(32'h3ba4d67e),
	.w6(32'h3b099ef4),
	.w7(32'hb86e0490),
	.w8(32'h3b6dba7f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba418f10),
	.w1(32'hbbec2f41),
	.w2(32'h3b12f1c9),
	.w3(32'h3a304bf4),
	.w4(32'hbb1d87ab),
	.w5(32'h395e89ad),
	.w6(32'h3b8302e7),
	.w7(32'hbb50bfde),
	.w8(32'hbb0137df),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9468c2),
	.w1(32'hbb6ca27b),
	.w2(32'hbb6df66f),
	.w3(32'h3be8b816),
	.w4(32'h3b60a151),
	.w5(32'h3a9e93df),
	.w6(32'h3bd828a5),
	.w7(32'h3c09d917),
	.w8(32'h3a9adaed),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4f8db),
	.w1(32'hbba48f60),
	.w2(32'hbba5d123),
	.w3(32'h3b9d6d18),
	.w4(32'hbbba5987),
	.w5(32'hbb1b8dd5),
	.w6(32'hba99a487),
	.w7(32'h3a2d4ee6),
	.w8(32'hbb344eec),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb88911),
	.w1(32'h3af99b64),
	.w2(32'hbb828aee),
	.w3(32'hbabb8d6c),
	.w4(32'h3b06476b),
	.w5(32'h3bca5a05),
	.w6(32'h3b886100),
	.w7(32'h3b9f38b4),
	.w8(32'h3c060313),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa6867),
	.w1(32'hbba05e4e),
	.w2(32'hbb3d2b2f),
	.w3(32'h3c9dc6f9),
	.w4(32'hb9977688),
	.w5(32'h3ac4c033),
	.w6(32'h3b934e10),
	.w7(32'h3bb77612),
	.w8(32'h3b790b85),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c361b),
	.w1(32'hbb27b8a8),
	.w2(32'hbb9886c2),
	.w3(32'hbb44c8b9),
	.w4(32'hbb64cc51),
	.w5(32'h3a3a9349),
	.w6(32'hbb8ad083),
	.w7(32'hba0c5151),
	.w8(32'h3b9d2dbd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc05507),
	.w1(32'h3b975827),
	.w2(32'h3bd113e7),
	.w3(32'h3c4e0d73),
	.w4(32'h3ba1a1c0),
	.w5(32'h3c10dd03),
	.w6(32'h3b789068),
	.w7(32'hbb771231),
	.w8(32'h3b14b5b4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4e4b6),
	.w1(32'hbc002c16),
	.w2(32'hbb1d3755),
	.w3(32'h3a895543),
	.w4(32'hbb3146b8),
	.w5(32'hbb154a56),
	.w6(32'h3b03c494),
	.w7(32'hbb88710f),
	.w8(32'hbba9b9cd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26ac82),
	.w1(32'h3b7b23f6),
	.w2(32'h3bacb0cb),
	.w3(32'h3b5c463f),
	.w4(32'h39b2a95f),
	.w5(32'hbaf4800e),
	.w6(32'h3bc1e63a),
	.w7(32'h3abda051),
	.w8(32'h3a0ceea8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44791e),
	.w1(32'hbad3dcc1),
	.w2(32'hbbb739d8),
	.w3(32'h3b0a6a3e),
	.w4(32'h3b9e7019),
	.w5(32'h3c4689e5),
	.w6(32'h386422d9),
	.w7(32'h3a912735),
	.w8(32'h3ad8cc84),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07c87e),
	.w1(32'h3b637312),
	.w2(32'hbb172a84),
	.w3(32'h3c0491f1),
	.w4(32'hbb44e4a1),
	.w5(32'hbc27cef4),
	.w6(32'h3a6db7f7),
	.w7(32'h3b0ecd27),
	.w8(32'h3b9fe8e2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eb9a8),
	.w1(32'hbb2cd66a),
	.w2(32'hba6054e6),
	.w3(32'h3c43fa17),
	.w4(32'h39c6d262),
	.w5(32'h3b9f064f),
	.w6(32'h3ba278b3),
	.w7(32'h3a8c533c),
	.w8(32'h39cb9d60),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff8db),
	.w1(32'h3ba18926),
	.w2(32'hba63818a),
	.w3(32'h3a0ac318),
	.w4(32'h3c390659),
	.w5(32'hbb905a85),
	.w6(32'h3aae2f40),
	.w7(32'h3c46141f),
	.w8(32'h3bd1bed0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeeb93),
	.w1(32'h3ba0040f),
	.w2(32'h3bebd501),
	.w3(32'h3bdac63a),
	.w4(32'h3c23052f),
	.w5(32'h3c0d75f8),
	.w6(32'h3c2d75b4),
	.w7(32'h3c3db8b8),
	.w8(32'h3c2e64a9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c449d88),
	.w1(32'h3c0afffe),
	.w2(32'h3b3f2dcc),
	.w3(32'h3bb629a7),
	.w4(32'h3a74e7ce),
	.w5(32'hbb222e55),
	.w6(32'h3c2d7521),
	.w7(32'h3aa79c0f),
	.w8(32'hb9821a33),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2166d2),
	.w1(32'hbc08b9f8),
	.w2(32'hb7d6112c),
	.w3(32'h3b79547f),
	.w4(32'hbb9c91d9),
	.w5(32'h3b4a3bbf),
	.w6(32'h3b6e7a6e),
	.w7(32'hbb4d82a4),
	.w8(32'hbb7fad26),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f536a),
	.w1(32'hbbf129a6),
	.w2(32'h3758fe29),
	.w3(32'h3b6a5e32),
	.w4(32'hbbcd4e97),
	.w5(32'h3c10a988),
	.w6(32'hbb347879),
	.w7(32'hba781a6f),
	.w8(32'h3bc52f9a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a52fb),
	.w1(32'h3b9e8c01),
	.w2(32'hbac0e124),
	.w3(32'h3a04e551),
	.w4(32'h3a5d5d77),
	.w5(32'hbba435d9),
	.w6(32'h388de5cb),
	.w7(32'hbaef4068),
	.w8(32'hbb0cfe89),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8587ca),
	.w1(32'hbb86167a),
	.w2(32'hbaaa37d8),
	.w3(32'hbb121571),
	.w4(32'hbb0c774e),
	.w5(32'h39af617e),
	.w6(32'hbb6c4627),
	.w7(32'hbaa5a01f),
	.w8(32'h3b946609),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe363b),
	.w1(32'hb92e334d),
	.w2(32'h3c054d48),
	.w3(32'hbb364f45),
	.w4(32'h3a9224bf),
	.w5(32'h3c51b9f1),
	.w6(32'hbaa47b25),
	.w7(32'h3be9d0f4),
	.w8(32'h3bafd140),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06cf15),
	.w1(32'hbacf5638),
	.w2(32'h3b88ab1d),
	.w3(32'h39e8de87),
	.w4(32'h3b5e0f0c),
	.w5(32'h3c31f75c),
	.w6(32'hbc0360e2),
	.w7(32'h3b798c15),
	.w8(32'h3aab961f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5abe67),
	.w1(32'hba82c93f),
	.w2(32'h3aa07393),
	.w3(32'hbb965c60),
	.w4(32'hbb837ea8),
	.w5(32'hba39aa99),
	.w6(32'hbbb212cc),
	.w7(32'h37ef0005),
	.w8(32'h3b22eee5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd9ea8),
	.w1(32'h3b18188c),
	.w2(32'h3b269005),
	.w3(32'h3a94b164),
	.w4(32'h3bae8bf7),
	.w5(32'hbb2e1223),
	.w6(32'h3b9db201),
	.w7(32'h3b1f9ebd),
	.w8(32'h3ac5f1d8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01bfd7),
	.w1(32'h3a32a7a4),
	.w2(32'h3bb587d4),
	.w3(32'hbba15325),
	.w4(32'hba325ae3),
	.w5(32'h3b27694a),
	.w6(32'hba964512),
	.w7(32'h3bb37460),
	.w8(32'h3a056183),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d1afc),
	.w1(32'hbc44d0bf),
	.w2(32'hbbbdce7d),
	.w3(32'hba422f4d),
	.w4(32'hba457e37),
	.w5(32'h3b55837d),
	.w6(32'hba280474),
	.w7(32'h3a7795fc),
	.w8(32'h3b6a3409),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2f6a1),
	.w1(32'hba903b6a),
	.w2(32'h3a60f98f),
	.w3(32'h3b9085eb),
	.w4(32'h3920a0e9),
	.w5(32'hbb71ad6e),
	.w6(32'hbbb7c039),
	.w7(32'hbad1971c),
	.w8(32'h3ac0ef7c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb721c71),
	.w1(32'h3b0690a2),
	.w2(32'hbbbf85f2),
	.w3(32'hb992a20f),
	.w4(32'hbad0c19d),
	.w5(32'hbba23745),
	.w6(32'h3b01ad1f),
	.w7(32'h3aa73de0),
	.w8(32'hbb60070e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9ee8b),
	.w1(32'h3b2dff6a),
	.w2(32'hbb34e21a),
	.w3(32'h39b407e5),
	.w4(32'hbb9198fb),
	.w5(32'hbb2fbb0b),
	.w6(32'h3a3276cc),
	.w7(32'h39f3df90),
	.w8(32'h3c148082),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddced7),
	.w1(32'h3be178e5),
	.w2(32'h3b3cb938),
	.w3(32'h3bef3056),
	.w4(32'h3c193bf2),
	.w5(32'hbbe07e8b),
	.w6(32'hba9f377d),
	.w7(32'h3bc184e1),
	.w8(32'h3b1d9914),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7588ed),
	.w1(32'hbb9627cd),
	.w2(32'hbbc34070),
	.w3(32'hba15e891),
	.w4(32'hbba11d1f),
	.w5(32'hbb60b459),
	.w6(32'h3b753dd7),
	.w7(32'hbb596079),
	.w8(32'hbb0e1538),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98568eb),
	.w1(32'h3b48e051),
	.w2(32'h3c02f7a0),
	.w3(32'h3ab89ce6),
	.w4(32'h3c39b026),
	.w5(32'h3c3678e9),
	.w6(32'hba9e8af7),
	.w7(32'h3bfab8ca),
	.w8(32'h3bad1217),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0afbab),
	.w1(32'hb964d4c4),
	.w2(32'hbb21dcd5),
	.w3(32'hbb4e7e9c),
	.w4(32'hba481f97),
	.w5(32'h396a603a),
	.w6(32'hba2f5446),
	.w7(32'h3bb38974),
	.w8(32'h3b909fd6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef896e),
	.w1(32'h3b855a96),
	.w2(32'h3b902726),
	.w3(32'h3b2d24d2),
	.w4(32'hbbc2d4ae),
	.w5(32'hbb120f72),
	.w6(32'hbb60c6f7),
	.w7(32'hbba5c8d0),
	.w8(32'hbba191c3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b204384),
	.w1(32'hb9c07084),
	.w2(32'hbb8368de),
	.w3(32'h3ba8d9c6),
	.w4(32'hbbb45e2f),
	.w5(32'hbbbcc0f9),
	.w6(32'h3a4de1ee),
	.w7(32'hbb66c699),
	.w8(32'hbba3efc6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fb17c),
	.w1(32'h3baac0e6),
	.w2(32'hbbb12510),
	.w3(32'h3aaabb9d),
	.w4(32'h3bbcd0e3),
	.w5(32'hbc106eb7),
	.w6(32'hba5704cc),
	.w7(32'h3be7e8bb),
	.w8(32'h3b25307a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dcb3ad),
	.w1(32'h3ae116b9),
	.w2(32'h3bb1c9bd),
	.w3(32'hba0fa61f),
	.w4(32'hba3c2607),
	.w5(32'h3c13b41f),
	.w6(32'hbb2445b9),
	.w7(32'hbb1ea7dd),
	.w8(32'h3c1acfeb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb80a5),
	.w1(32'hbab5877b),
	.w2(32'hba354475),
	.w3(32'h3bd6447c),
	.w4(32'hbb2e2f88),
	.w5(32'hbb92e378),
	.w6(32'h3b95cde8),
	.w7(32'h3b2af8f5),
	.w8(32'h394b6b36),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad233a6),
	.w1(32'h3a711de6),
	.w2(32'h3af88fee),
	.w3(32'hbb2f4d89),
	.w4(32'h3b219b3e),
	.w5(32'h3c6cc761),
	.w6(32'hbc24a00f),
	.w7(32'h3bf97b70),
	.w8(32'h3c19f425),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a8f46),
	.w1(32'hbbbd466c),
	.w2(32'hbaa1058b),
	.w3(32'h3bc1421f),
	.w4(32'hbc10fb7c),
	.w5(32'h3b1a0937),
	.w6(32'hbab8937c),
	.w7(32'hba771d8b),
	.w8(32'h3a9a3e0c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904850),
	.w1(32'h3b96b674),
	.w2(32'h3be2cdf8),
	.w3(32'hbbd0d2f1),
	.w4(32'h3aae4b4e),
	.w5(32'h3c11b592),
	.w6(32'hbc00ccf1),
	.w7(32'h3a50fc43),
	.w8(32'h3a817456),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb42dd),
	.w1(32'hbae2ce6c),
	.w2(32'hba3f9a4d),
	.w3(32'hbae6c098),
	.w4(32'hbaae4fd1),
	.w5(32'h3b44360e),
	.w6(32'h3aba4f76),
	.w7(32'hba6f397a),
	.w8(32'h3a0f9e23),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6f2a1),
	.w1(32'h3a9fec66),
	.w2(32'hbc07c996),
	.w3(32'hbb95fc8d),
	.w4(32'hba83ecd7),
	.w5(32'hbb314782),
	.w6(32'hbb4984c6),
	.w7(32'hbbf72a22),
	.w8(32'hbc2e796e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ec81a),
	.w1(32'hb9721bc8),
	.w2(32'h3be085fd),
	.w3(32'hbb845d48),
	.w4(32'h3c5adc59),
	.w5(32'h3c82ae78),
	.w6(32'hbbd435f7),
	.w7(32'h3c00630e),
	.w8(32'h3be9bc74),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c601a),
	.w1(32'h3b8a01e9),
	.w2(32'hbb5aef2d),
	.w3(32'h3b5c6829),
	.w4(32'h3b7732c7),
	.w5(32'h3a61cc84),
	.w6(32'h3b6d7ea3),
	.w7(32'hb943a768),
	.w8(32'hbad16d7f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c8920),
	.w1(32'hbb676029),
	.w2(32'hbbf819d3),
	.w3(32'h3bd8c291),
	.w4(32'hbbea9884),
	.w5(32'hbbdcaff9),
	.w6(32'h3bb8808b),
	.w7(32'hbbb1368e),
	.w8(32'hbb280b8a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfe205),
	.w1(32'hbb84288e),
	.w2(32'hbb4b270a),
	.w3(32'hbbbf93e8),
	.w4(32'h3a9e673f),
	.w5(32'hba0c2c4b),
	.w6(32'hbbc06603),
	.w7(32'h3b7f4bbf),
	.w8(32'hbbb37f9c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e41791),
	.w1(32'h3ba2d643),
	.w2(32'h3a268a7d),
	.w3(32'h3b1dd745),
	.w4(32'h3c2e5d64),
	.w5(32'hbbfebc04),
	.w6(32'hbb2108a5),
	.w7(32'h3b34eafd),
	.w8(32'h3b1896a7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c046b90),
	.w1(32'h3b15796b),
	.w2(32'h3b505b79),
	.w3(32'h3b81fe95),
	.w4(32'hbb5c22a2),
	.w5(32'h3ac62599),
	.w6(32'h3bc95a77),
	.w7(32'hbaab06bc),
	.w8(32'h3b03f09e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affdc03),
	.w1(32'h3b0a81a5),
	.w2(32'hbaa39813),
	.w3(32'h3808b8c8),
	.w4(32'hbba54752),
	.w5(32'h3bb4310d),
	.w6(32'h39e50fe9),
	.w7(32'hbb61665d),
	.w8(32'h3b87f454),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e4f52),
	.w1(32'h3c20b244),
	.w2(32'h3a30b1bc),
	.w3(32'h3a2da5b5),
	.w4(32'h3bbcf12c),
	.w5(32'hba714d09),
	.w6(32'hbab7a6c5),
	.w7(32'h3b431843),
	.w8(32'h3ba54397),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac04fe0),
	.w1(32'h3bdc11a1),
	.w2(32'h3b2e1c46),
	.w3(32'h3bbee3da),
	.w4(32'h3a86f50a),
	.w5(32'hbbcbfc12),
	.w6(32'h3c0554a5),
	.w7(32'hb9f7f325),
	.w8(32'hbc0080fc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f8283),
	.w1(32'h3b035452),
	.w2(32'h3ae84832),
	.w3(32'h3bad6027),
	.w4(32'h3a8307d5),
	.w5(32'h39397f6a),
	.w6(32'hb7f25c42),
	.w7(32'h3a11927b),
	.w8(32'h3c1c6e2a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3574d2),
	.w1(32'h3a047011),
	.w2(32'hbb42d4a7),
	.w3(32'h3ba6dfe9),
	.w4(32'hba9bdbe8),
	.w5(32'hbb986b44),
	.w6(32'h3b42fd7e),
	.w7(32'hbb93c8e3),
	.w8(32'hbb096c01),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3789e033),
	.w1(32'h3b567755),
	.w2(32'hbafdfd8d),
	.w3(32'h39f33d00),
	.w4(32'h3989484c),
	.w5(32'hbb7b5e61),
	.w6(32'hba8d8777),
	.w7(32'h3aa3c9a1),
	.w8(32'h3b2bccac),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02392b),
	.w1(32'hbb1ef376),
	.w2(32'h3b0cba52),
	.w3(32'h3b6778fd),
	.w4(32'h3ab0b7fe),
	.w5(32'h3b82291e),
	.w6(32'h3a19fe6a),
	.w7(32'hb9faf069),
	.w8(32'hbb48307a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7c0ea),
	.w1(32'hbb203ae1),
	.w2(32'h39c58306),
	.w3(32'hbbaff108),
	.w4(32'h3b9479c7),
	.w5(32'hb93bb395),
	.w6(32'hbb7dae09),
	.w7(32'hbb91ed62),
	.w8(32'h3b45c514),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e035a),
	.w1(32'hbb4372c0),
	.w2(32'hb9c0281c),
	.w3(32'hbc07e85a),
	.w4(32'hbae81ef4),
	.w5(32'h3c29bca7),
	.w6(32'hbc10629d),
	.w7(32'h3a9fe271),
	.w8(32'h3b0f0f49),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b2f6),
	.w1(32'h3bd67369),
	.w2(32'h3c0dbffb),
	.w3(32'h3be1d0cd),
	.w4(32'h3bdb03c7),
	.w5(32'h3be99933),
	.w6(32'h3b6df8f4),
	.w7(32'h3b14c9b1),
	.w8(32'h3c335810),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db7ae),
	.w1(32'h3c180243),
	.w2(32'h3c297087),
	.w3(32'h3ac36699),
	.w4(32'h3c578937),
	.w5(32'h3c31ce9f),
	.w6(32'h3b88f8ce),
	.w7(32'h3b06893a),
	.w8(32'h3a9ee925),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81ac3f),
	.w1(32'h3b50ed63),
	.w2(32'hba8b068e),
	.w3(32'hbb5dbd15),
	.w4(32'h3af022d0),
	.w5(32'h3b313a5f),
	.w6(32'h3af48a09),
	.w7(32'h3b14824d),
	.w8(32'h3c08e224),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf7419),
	.w1(32'hbb4e99ec),
	.w2(32'hbc04451f),
	.w3(32'hbaa970d2),
	.w4(32'hbb7b35b6),
	.w5(32'hbc1d41b4),
	.w6(32'h3b251f17),
	.w7(32'hbb999ffa),
	.w8(32'hbc1aa8d4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c1d9d),
	.w1(32'h3bb24b67),
	.w2(32'h3a05d37b),
	.w3(32'h3b8ad3e8),
	.w4(32'h3b938e14),
	.w5(32'hba83b0d6),
	.w6(32'h3c167171),
	.w7(32'h3bd6ac3f),
	.w8(32'h3bdabdf5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62ebd4),
	.w1(32'h3c0f66bc),
	.w2(32'h3bceecb3),
	.w3(32'hbabd5bb8),
	.w4(32'h3cb8090b),
	.w5(32'h3c9e2264),
	.w6(32'hbb7d4120),
	.w7(32'h3aabf10d),
	.w8(32'h3c3bc487),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb877c0d),
	.w1(32'hbb07167f),
	.w2(32'hbc08d86e),
	.w3(32'h3bb35e6f),
	.w4(32'hbbe1cbdf),
	.w5(32'hbc0bc010),
	.w6(32'h39bdcbc1),
	.w7(32'hbbc20a66),
	.w8(32'hbaccdf27),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b939dd2),
	.w1(32'hba63cd35),
	.w2(32'h3b8237ad),
	.w3(32'h3b1354ac),
	.w4(32'h3aade180),
	.w5(32'h3c21b3f5),
	.w6(32'h3aab6e91),
	.w7(32'hbc0fa869),
	.w8(32'h3c2be5dc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44cf75),
	.w1(32'hbb3b99ec),
	.w2(32'hba6af764),
	.w3(32'hbaaf576b),
	.w4(32'h3a0fbf90),
	.w5(32'h3b650fdc),
	.w6(32'h3a460330),
	.w7(32'h3b8c329b),
	.w8(32'h3b2c4f1d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ac2a6),
	.w1(32'h3c0667bb),
	.w2(32'h3b18eb42),
	.w3(32'hbb1c1d8f),
	.w4(32'h3b4767bf),
	.w5(32'hba08e0a1),
	.w6(32'h39f045bc),
	.w7(32'h3bc188d9),
	.w8(32'h3acfb600),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2ce9),
	.w1(32'h3ae5968a),
	.w2(32'hbb88831e),
	.w3(32'hbb71a573),
	.w4(32'hbbb111d5),
	.w5(32'h3b8b637e),
	.w6(32'hbbb4fb6d),
	.w7(32'h3ad9525d),
	.w8(32'h3c1aab27),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1977b7),
	.w1(32'hbb408bb2),
	.w2(32'hb944463e),
	.w3(32'h3bc20da3),
	.w4(32'hbb6554d8),
	.w5(32'hbbc94070),
	.w6(32'hbc065551),
	.w7(32'h3b0a160c),
	.w8(32'hbbd4d5bf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02ec89),
	.w1(32'hba9de48e),
	.w2(32'h3a8aa2bc),
	.w3(32'hbb7ee33d),
	.w4(32'h3a7c63ae),
	.w5(32'h3858cdd6),
	.w6(32'hbbc51d6a),
	.w7(32'h3b30c7ce),
	.w8(32'h3a1f5789),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7f182),
	.w1(32'hbbd1506d),
	.w2(32'hbbd7be72),
	.w3(32'h3c0672cb),
	.w4(32'hbc1de71c),
	.w5(32'hbbc0c334),
	.w6(32'h3bb9a245),
	.w7(32'hba2cc2d1),
	.w8(32'h3aa07930),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b689),
	.w1(32'h3c340be8),
	.w2(32'hbaa4284d),
	.w3(32'h3b207cb6),
	.w4(32'hbb676bd3),
	.w5(32'hbba1e827),
	.w6(32'hbaf6fd62),
	.w7(32'h3b5b46db),
	.w8(32'h3bba3b6b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1953a5),
	.w1(32'hbbb41c2f),
	.w2(32'hbb90b658),
	.w3(32'h3bf59bac),
	.w4(32'hbb89239b),
	.w5(32'hbbdb1f11),
	.w6(32'h3c0c4166),
	.w7(32'hbb1441a7),
	.w8(32'hbb3821fa),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bf439),
	.w1(32'h3c037633),
	.w2(32'h3aca20a8),
	.w3(32'hbb98f52e),
	.w4(32'h3bde6993),
	.w5(32'hbabeefb2),
	.w6(32'hbae127d8),
	.w7(32'h3bb4d319),
	.w8(32'h391e1b07),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843a84),
	.w1(32'h3a6eb3dd),
	.w2(32'h3a0b5836),
	.w3(32'h3969a404),
	.w4(32'h3b607d5f),
	.w5(32'h3b7b69ec),
	.w6(32'h38f0468e),
	.w7(32'h3b9773e0),
	.w8(32'h3c080af2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddcad4),
	.w1(32'h39d92909),
	.w2(32'hbb8ebe92),
	.w3(32'h3b6d706f),
	.w4(32'h3a79857e),
	.w5(32'hbb07c786),
	.w6(32'h3bf80fc2),
	.w7(32'h3b4f8d68),
	.w8(32'hbafd1cb8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89094e),
	.w1(32'h3b420773),
	.w2(32'hbb3fdc71),
	.w3(32'h3ba18ab7),
	.w4(32'hb999ea67),
	.w5(32'hba8cb6f2),
	.w6(32'hba5bc099),
	.w7(32'h394f42f0),
	.w8(32'hbb80cbbe),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a105b),
	.w1(32'h3a3d91db),
	.w2(32'h3a6a060c),
	.w3(32'h3a70df33),
	.w4(32'h3b8a9114),
	.w5(32'hbba8d8a9),
	.w6(32'h3af09cc1),
	.w7(32'hb9be4112),
	.w8(32'hbaa8afc2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a85a6),
	.w1(32'hba04efca),
	.w2(32'h3a8840f6),
	.w3(32'hb90f025d),
	.w4(32'h3b274050),
	.w5(32'hbb839e5f),
	.w6(32'h3b7fe58c),
	.w7(32'h3aa70756),
	.w8(32'hbb5dc781),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba138bc3),
	.w1(32'h3a62df48),
	.w2(32'hbbd35729),
	.w3(32'hbb095e74),
	.w4(32'h3b33145c),
	.w5(32'hbb3f3f3b),
	.w6(32'hb963caea),
	.w7(32'hbaa10316),
	.w8(32'h39f8e5bd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf569de),
	.w1(32'hbbac6e45),
	.w2(32'hba802492),
	.w3(32'hbb51c9c7),
	.w4(32'hbc28cc3f),
	.w5(32'h3b93778e),
	.w6(32'hbb4d3f0c),
	.w7(32'hbc0e60f6),
	.w8(32'h3b6a40b9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba470),
	.w1(32'h3b9518e0),
	.w2(32'hbb834ccc),
	.w3(32'hbb7c1ad2),
	.w4(32'h3ba2d652),
	.w5(32'hbbd3c3e0),
	.w6(32'hbb30aae4),
	.w7(32'h3b766fb7),
	.w8(32'h39b883bc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e50e0),
	.w1(32'h39b4ae3c),
	.w2(32'h373af9d3),
	.w3(32'h3b083d78),
	.w4(32'hba04bd6d),
	.w5(32'hbba7f32f),
	.w6(32'hbae5c5d5),
	.w7(32'h3802a145),
	.w8(32'hb9f0e8e5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c061b71),
	.w1(32'hb90457a4),
	.w2(32'hb9df7d9b),
	.w3(32'h3c36cb8e),
	.w4(32'hbb286dd9),
	.w5(32'hba771056),
	.w6(32'h3c109886),
	.w7(32'hbb2b7ffe),
	.w8(32'hbadc2008),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98cb75),
	.w1(32'hbc0b0006),
	.w2(32'hbaca0d1c),
	.w3(32'h3b2c53c0),
	.w4(32'hbb988e8e),
	.w5(32'h3b25a698),
	.w6(32'hbb01fe91),
	.w7(32'hba835174),
	.w8(32'h3b0ba419),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae35e4d),
	.w1(32'hbb85a1c3),
	.w2(32'hbbc38d82),
	.w3(32'hbb2eb554),
	.w4(32'h3b725b4a),
	.w5(32'hbb47fb5b),
	.w6(32'hbac7fa37),
	.w7(32'hba5c2e42),
	.w8(32'h3a6dad3e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3801e09b),
	.w1(32'h3c248852),
	.w2(32'hbaf16880),
	.w3(32'hbb661530),
	.w4(32'h3c06bc49),
	.w5(32'hbb8a3626),
	.w6(32'h38333687),
	.w7(32'h3a39b54d),
	.w8(32'hbb296aa2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99a6b2),
	.w1(32'h3b9f685b),
	.w2(32'h3be97b45),
	.w3(32'h3c84291c),
	.w4(32'h3bdcf462),
	.w5(32'h3ab02a46),
	.w6(32'h3c8ffe16),
	.w7(32'h3bdaeacc),
	.w8(32'h3bf38daf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b620153),
	.w1(32'h3c1a4b4d),
	.w2(32'h3c53e090),
	.w3(32'h399f62f8),
	.w4(32'h3cce9592),
	.w5(32'h3c75beee),
	.w6(32'h3890114e),
	.w7(32'h3bf96828),
	.w8(32'h39feffd5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ddb78),
	.w1(32'hbbde2385),
	.w2(32'h37cac593),
	.w3(32'hba4545c9),
	.w4(32'hbb4cc035),
	.w5(32'h3b50736a),
	.w6(32'h3c1338cd),
	.w7(32'hbb8057dd),
	.w8(32'h3ad3e806),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eb577),
	.w1(32'h3b95f3aa),
	.w2(32'hbb4268f1),
	.w3(32'hbbaca922),
	.w4(32'hb9c5f1da),
	.w5(32'hbbb3d396),
	.w6(32'hbb9146be),
	.w7(32'hba3bed11),
	.w8(32'hbbb43bc9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfa67f),
	.w1(32'h3b6bfe02),
	.w2(32'hbb6a1f89),
	.w3(32'h3b4b27d0),
	.w4(32'h3b029d3e),
	.w5(32'hbbd42810),
	.w6(32'h3bdd6526),
	.w7(32'hbac50c0a),
	.w8(32'h3b69c63c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81fe75),
	.w1(32'hb9da389d),
	.w2(32'h3b5657fc),
	.w3(32'h3b66b2bd),
	.w4(32'h39520e98),
	.w5(32'hbae1819f),
	.w6(32'h3be299ef),
	.w7(32'h3bd3d811),
	.w8(32'h3af913c0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc977b2),
	.w1(32'h3b89b073),
	.w2(32'hba0590f0),
	.w3(32'h3aaa53e8),
	.w4(32'hbbdae4d7),
	.w5(32'hbab7e501),
	.w6(32'h3bcad73c),
	.w7(32'h3b825b19),
	.w8(32'h3af083ec),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f85bc),
	.w1(32'hb9824501),
	.w2(32'hbbc6727d),
	.w3(32'hbbd765e6),
	.w4(32'h3c3face6),
	.w5(32'hbc0275d5),
	.w6(32'hbc0d9d86),
	.w7(32'h3bb5b245),
	.w8(32'hb867a87e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3176b0),
	.w1(32'h3b4fde8d),
	.w2(32'h3b04b4ba),
	.w3(32'h3bcb6c2f),
	.w4(32'hbb26e490),
	.w5(32'hbb6f2525),
	.w6(32'h3c2f35a2),
	.w7(32'h3a12c49c),
	.w8(32'hba77c4f2),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac06241),
	.w1(32'hbb5f5f3c),
	.w2(32'hbb42502e),
	.w3(32'h3a35ce68),
	.w4(32'h3ae778d5),
	.w5(32'hbab87e21),
	.w6(32'hb9b07842),
	.w7(32'h3b635e5b),
	.w8(32'h3a246b16),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b065bcc),
	.w1(32'h3baf6947),
	.w2(32'h3b238d67),
	.w3(32'h3b1d001e),
	.w4(32'h3c03eb6d),
	.w5(32'h3bb0a9da),
	.w6(32'h3bc67a4c),
	.w7(32'h3a3dba8b),
	.w8(32'h3b685485),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd8456),
	.w1(32'hba2c1050),
	.w2(32'hbb1496ed),
	.w3(32'h3b9d9197),
	.w4(32'hbba3400f),
	.w5(32'h3b987a09),
	.w6(32'h3b66f36c),
	.w7(32'h3ae8e03c),
	.w8(32'h3b0496a3),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e263e),
	.w1(32'h3b5a0055),
	.w2(32'h3bb668e5),
	.w3(32'hbabe2e85),
	.w4(32'h3b5d5099),
	.w5(32'h3b83d4f2),
	.w6(32'h3b90c352),
	.w7(32'h3b0cd947),
	.w8(32'hbac5c323),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98bdc9),
	.w1(32'hbaadafe1),
	.w2(32'h3beca9a1),
	.w3(32'hbb4b14bb),
	.w4(32'h3b9154b3),
	.w5(32'h3c1ac5ce),
	.w6(32'hbbc2d2e0),
	.w7(32'h3b05289c),
	.w8(32'h3c0fe904),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f2561),
	.w1(32'hb97dbcd8),
	.w2(32'h3be8758d),
	.w3(32'hb9b01a22),
	.w4(32'h3b9d7c23),
	.w5(32'h3c16bad2),
	.w6(32'h3b2addd1),
	.w7(32'hbb954513),
	.w8(32'hbab24127),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a11e0),
	.w1(32'h3c5b5d5d),
	.w2(32'h3b90e762),
	.w3(32'hbbb9c189),
	.w4(32'h3c92bfa3),
	.w5(32'h3c102034),
	.w6(32'h3b9f8018),
	.w7(32'h3c46dcdb),
	.w8(32'h3c368599),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7720fb),
	.w1(32'hb9cec7ee),
	.w2(32'h3c1068bb),
	.w3(32'hbad327e8),
	.w4(32'hbaad29bf),
	.w5(32'hbaa3df01),
	.w6(32'hbbed49fc),
	.w7(32'h3b17af29),
	.w8(32'h3bb7c13f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9b807),
	.w1(32'h3bdc150d),
	.w2(32'hbaf47720),
	.w3(32'h3a5b41ad),
	.w4(32'h3bb342ae),
	.w5(32'hbb968c1f),
	.w6(32'h3b64e5b7),
	.w7(32'h3bf7e908),
	.w8(32'h3b6502e1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873a0a),
	.w1(32'hbbadf028),
	.w2(32'hbbad797a),
	.w3(32'h3c40d856),
	.w4(32'hbb2167fe),
	.w5(32'hbafc93fd),
	.w6(32'h3b533b37),
	.w7(32'hbba39472),
	.w8(32'h3b03b2aa),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a607cea),
	.w1(32'h3ac5a922),
	.w2(32'h3c15149b),
	.w3(32'h3afa76e8),
	.w4(32'h3bfd9c7b),
	.w5(32'h3c73bfca),
	.w6(32'h3b3982bd),
	.w7(32'h3bfde2a1),
	.w8(32'h3b0f42e1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567db6),
	.w1(32'h3ac78e30),
	.w2(32'h3ac8b09b),
	.w3(32'hbc01db05),
	.w4(32'h3b58504a),
	.w5(32'hb9c8f60f),
	.w6(32'hbc0f7916),
	.w7(32'h3bb3cfc0),
	.w8(32'h39d395d5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b851685),
	.w1(32'hbb0a7d7a),
	.w2(32'h3ab47c69),
	.w3(32'h3bf14516),
	.w4(32'hba930283),
	.w5(32'hba7c553e),
	.w6(32'h3b479f8e),
	.w7(32'h3b1bcbae),
	.w8(32'hbacb3614),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc28d5),
	.w1(32'hba86cd13),
	.w2(32'hbbe0b475),
	.w3(32'h3bdac87f),
	.w4(32'h39d85681),
	.w5(32'hbad36611),
	.w6(32'h3ba2b927),
	.w7(32'hba4b4168),
	.w8(32'hbc0daef4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2796ff),
	.w1(32'hbc07c81a),
	.w2(32'hbbcd8790),
	.w3(32'h3a883d2f),
	.w4(32'hbb72a842),
	.w5(32'hbbfe6853),
	.w6(32'hbafac516),
	.w7(32'h3c099ccb),
	.w8(32'h3c2dcace),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b552a27),
	.w1(32'h3c14f81e),
	.w2(32'hbc16ed60),
	.w3(32'h3c496332),
	.w4(32'hbba4536e),
	.w5(32'hbc2ddba9),
	.w6(32'h3c1adcc9),
	.w7(32'hbb8e0bc5),
	.w8(32'hbb8a3c7d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf98b90),
	.w1(32'h3b5049c2),
	.w2(32'h3c16d1f8),
	.w3(32'h3bfe2978),
	.w4(32'hbb424436),
	.w5(32'h3c560f04),
	.w6(32'h3c2bb4a5),
	.w7(32'hbb23dcd9),
	.w8(32'h3c0b4edf),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8cf86),
	.w1(32'h3b8133fc),
	.w2(32'hb86e9f5c),
	.w3(32'h3ac0a772),
	.w4(32'h3bd4c516),
	.w5(32'h3b35325c),
	.w6(32'h3b355247),
	.w7(32'h3ba99c91),
	.w8(32'hbaa9e55a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b4311),
	.w1(32'h3b0b98c6),
	.w2(32'h39e4fb68),
	.w3(32'h3a621dc9),
	.w4(32'hbaa9cc7e),
	.w5(32'hbb8c2a5f),
	.w6(32'h3ba1a897),
	.w7(32'hbb78cf1c),
	.w8(32'h3b929b44),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2c0a),
	.w1(32'h3bbd30d3),
	.w2(32'h3c150776),
	.w3(32'hbb816cd3),
	.w4(32'h39caafba),
	.w5(32'h3c1fc076),
	.w6(32'h3a89db60),
	.w7(32'h3a1c7368),
	.w8(32'h3bf4ac52),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386217b6),
	.w1(32'hbbdb6823),
	.w2(32'h3b5ba521),
	.w3(32'h3b0e3f4f),
	.w4(32'hbad40e8b),
	.w5(32'h3c45e14c),
	.w6(32'h3ad88e3e),
	.w7(32'h3b84dcfe),
	.w8(32'hba8ff4c3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b449d38),
	.w1(32'h3ac321ee),
	.w2(32'h3c111371),
	.w3(32'hbbbb7eb9),
	.w4(32'hba0a137b),
	.w5(32'hbbae04b4),
	.w6(32'hbc2cb030),
	.w7(32'h3c0ab32e),
	.w8(32'h3c305691),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce26eb),
	.w1(32'hbba8f9ff),
	.w2(32'h3bce7213),
	.w3(32'h3b05bee0),
	.w4(32'hbc069eaa),
	.w5(32'h3c06aaf2),
	.w6(32'h3c0a4c63),
	.w7(32'h3b5a2d85),
	.w8(32'h3bff4323),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67bdb5),
	.w1(32'h3aba08dc),
	.w2(32'h3b201a3b),
	.w3(32'hba8f08ab),
	.w4(32'hbb6c6e18),
	.w5(32'h3b59928d),
	.w6(32'hbb21fafe),
	.w7(32'hbb26b49d),
	.w8(32'h3c04ef03),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af043fe),
	.w1(32'hbc2cf792),
	.w2(32'hbbd65387),
	.w3(32'h3b327fc7),
	.w4(32'hbbb543f3),
	.w5(32'hbb2a4961),
	.w6(32'h3b3d6664),
	.w7(32'h3b8fbd8d),
	.w8(32'hbc4c2dbe),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36e020),
	.w1(32'h3bc48b21),
	.w2(32'h3bed1dac),
	.w3(32'h3bef339f),
	.w4(32'h3bab4a05),
	.w5(32'h3cdfe111),
	.w6(32'hbabc2827),
	.w7(32'h37034f45),
	.w8(32'h3c752631),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11d869),
	.w1(32'h39a0aff0),
	.w2(32'hbb8ba390),
	.w3(32'hbb057768),
	.w4(32'h3b282ac4),
	.w5(32'hbb051981),
	.w6(32'h3b32eaff),
	.w7(32'h3b4a9578),
	.w8(32'hbaee4c12),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80bced),
	.w1(32'h3bead431),
	.w2(32'h3c093f00),
	.w3(32'hbb8dd944),
	.w4(32'h3bc572d0),
	.w5(32'h3bf9f87e),
	.w6(32'h3ab91e4c),
	.w7(32'h3bde662c),
	.w8(32'h3c6ca5f5),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5f20b),
	.w1(32'hbb58a33a),
	.w2(32'hbba0b37b),
	.w3(32'hba509781),
	.w4(32'hbb16dc03),
	.w5(32'hbbf699a6),
	.w6(32'h3bdc5afc),
	.w7(32'hba8e311a),
	.w8(32'hbbfa4d87),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55694b),
	.w1(32'h3a09e6ee),
	.w2(32'h3a983933),
	.w3(32'hbbdfbf0d),
	.w4(32'hbc18561a),
	.w5(32'hbc0e8360),
	.w6(32'hbbe8f666),
	.w7(32'hbc63d1b7),
	.w8(32'h3bdd5370),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11f2cb),
	.w1(32'h3b17d530),
	.w2(32'h3baea5c2),
	.w3(32'h3c68cb21),
	.w4(32'h3aec1908),
	.w5(32'h3b22acb6),
	.w6(32'h3cc1f9ea),
	.w7(32'h3a39f80b),
	.w8(32'h3b3856ff),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e1e39),
	.w1(32'hbb3096db),
	.w2(32'hbbb67c8a),
	.w3(32'h3aeb9e2e),
	.w4(32'hbb4a10c0),
	.w5(32'h3baaaefe),
	.w6(32'h3c49e2f2),
	.w7(32'hbaf352cc),
	.w8(32'h3c0e05ac),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdee4d0),
	.w1(32'h3b573023),
	.w2(32'hbb919ac3),
	.w3(32'hbc4845ca),
	.w4(32'hba5940b3),
	.w5(32'hbad019db),
	.w6(32'hb9f467d0),
	.w7(32'h3b4155bf),
	.w8(32'h3b63ce95),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc793bf),
	.w1(32'hbb3bebf7),
	.w2(32'hbb1d1e29),
	.w3(32'hba4e5843),
	.w4(32'h3bd197c5),
	.w5(32'h3bddfbc1),
	.w6(32'h3a2afea3),
	.w7(32'h3989cfbe),
	.w8(32'hba27e815),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba426f2c),
	.w1(32'hbbe7199c),
	.w2(32'h3b1be84b),
	.w3(32'hbb3350b6),
	.w4(32'h3a5c65d8),
	.w5(32'hb98a6caf),
	.w6(32'hbbe29cc2),
	.w7(32'hbb07593b),
	.w8(32'h3ba4edcd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9f4d),
	.w1(32'hbab03d5d),
	.w2(32'hbbba0d58),
	.w3(32'hbb539e45),
	.w4(32'hbc15ed4e),
	.w5(32'hbafe3a2f),
	.w6(32'hbb675530),
	.w7(32'hbbb6d373),
	.w8(32'h39d3463a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e9cca),
	.w1(32'hbb9259ea),
	.w2(32'hbb02cd32),
	.w3(32'h393cbb39),
	.w4(32'hba88330b),
	.w5(32'hbad10c96),
	.w6(32'h3b4985df),
	.w7(32'hba167855),
	.w8(32'hbbb197cc),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977086),
	.w1(32'h3aeada46),
	.w2(32'h3b418dc1),
	.w3(32'h3aa1701d),
	.w4(32'h3ad091f8),
	.w5(32'h3c271ee0),
	.w6(32'h3ac47930),
	.w7(32'h3b108eb1),
	.w8(32'h3baa178c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bc5b4),
	.w1(32'h3bd7dc9a),
	.w2(32'h3b0616e8),
	.w3(32'hbaa2af15),
	.w4(32'h3b9cb88c),
	.w5(32'h392ccc61),
	.w6(32'h3b85e14e),
	.w7(32'h3bb81aab),
	.w8(32'h3b47d6d8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72ce4e),
	.w1(32'hbbfdf3e5),
	.w2(32'hbbd0e464),
	.w3(32'h3aea8490),
	.w4(32'hbb7b65d6),
	.w5(32'h3a943fc3),
	.w6(32'h39a869b7),
	.w7(32'hba7d07ec),
	.w8(32'h3b8d7f7f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ed44f),
	.w1(32'hbba062a9),
	.w2(32'h3ae33858),
	.w3(32'h3b147b45),
	.w4(32'hba0f616b),
	.w5(32'hbb483e57),
	.w6(32'h3b5f19f1),
	.w7(32'h3c048c75),
	.w8(32'h39c72e6f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949d811),
	.w1(32'hba5639b8),
	.w2(32'hbaefe4f4),
	.w3(32'hbbb094dd),
	.w4(32'hbb955f7a),
	.w5(32'hbb76aacb),
	.w6(32'hbbfd0b13),
	.w7(32'hba3e7628),
	.w8(32'hbb3aec3f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6356c8),
	.w1(32'hbadd66ac),
	.w2(32'h3b91d020),
	.w3(32'hbb39d991),
	.w4(32'hbb8e5ee3),
	.w5(32'h3b20bdc6),
	.w6(32'hba1cea4f),
	.w7(32'hbb207787),
	.w8(32'h3ba5d0d0),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ead92),
	.w1(32'hbad2061f),
	.w2(32'hbb20d9a6),
	.w3(32'h3c1f68ab),
	.w4(32'hb98e0408),
	.w5(32'h3c285345),
	.w6(32'h3c4ad1e3),
	.w7(32'h3afad021),
	.w8(32'hba38aa1b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba942a15),
	.w1(32'h3aaddcfc),
	.w2(32'h3b719a0b),
	.w3(32'hbbe9e4cd),
	.w4(32'hb823f76c),
	.w5(32'h3b47316d),
	.w6(32'h3b864946),
	.w7(32'h3c0e554f),
	.w8(32'h3b2b6d7b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e91e0),
	.w1(32'h3b61d36f),
	.w2(32'hbab4162a),
	.w3(32'hbba95b15),
	.w4(32'hbb108d7f),
	.w5(32'h39e4e26c),
	.w6(32'hbbea9996),
	.w7(32'hbb1d5985),
	.w8(32'h3b3901ab),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fd9ca),
	.w1(32'h3bd41081),
	.w2(32'h3ac5df04),
	.w3(32'hbb229e7a),
	.w4(32'h3ab52d3a),
	.w5(32'h3b7124d7),
	.w6(32'h3b2bc86e),
	.w7(32'h3becd797),
	.w8(32'h3b19168f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801f1c),
	.w1(32'hbb35ddf4),
	.w2(32'hbb7dd56a),
	.w3(32'h3b1daca8),
	.w4(32'hbbac07d8),
	.w5(32'hbb24e408),
	.w6(32'hbbd9b5fd),
	.w7(32'h3b5d854a),
	.w8(32'hbba5b21c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb64b5b),
	.w1(32'h3bb84b68),
	.w2(32'h3b1b60e3),
	.w3(32'hbc5064cc),
	.w4(32'h3c21bfb2),
	.w5(32'h3bce9874),
	.w6(32'hbc04dab7),
	.w7(32'h3bb5fa00),
	.w8(32'h3bddfdd0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84588e),
	.w1(32'hbbc543a4),
	.w2(32'h3c5d8f81),
	.w3(32'h3a25b353),
	.w4(32'hbb31b45e),
	.w5(32'h3b9ff0a2),
	.w6(32'h3a9b31e5),
	.w7(32'hbc7d2d73),
	.w8(32'h3c42c704),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9ab75),
	.w1(32'hbb815c2a),
	.w2(32'hbc32fb56),
	.w3(32'h39647fbc),
	.w4(32'h3c22ddb2),
	.w5(32'h3d514c6a),
	.w6(32'hbb31775e),
	.w7(32'hbc8136f0),
	.w8(32'h3bf3c5b6),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8700e0),
	.w1(32'h3bdd0110),
	.w2(32'hba3ac527),
	.w3(32'hbc998f1c),
	.w4(32'hbadad489),
	.w5(32'h3bbc5512),
	.w6(32'hbc1b73f2),
	.w7(32'hbb8477a9),
	.w8(32'h3ba0cff0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae32325),
	.w1(32'h3bf0881b),
	.w2(32'h3b9beb2b),
	.w3(32'h3bcc2d87),
	.w4(32'h3ba1660e),
	.w5(32'h3bee41b3),
	.w6(32'h3c0e0ca9),
	.w7(32'h3ad8f001),
	.w8(32'h3b076c55),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27e537),
	.w1(32'hbb97044c),
	.w2(32'h3b542c8c),
	.w3(32'h3b313afe),
	.w4(32'hbbe681c0),
	.w5(32'h3b822e62),
	.w6(32'h3aba22b1),
	.w7(32'hbb2975be),
	.w8(32'hb8c1cf8a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2f76b),
	.w1(32'hbb182c5f),
	.w2(32'h3ab55889),
	.w3(32'h3c326419),
	.w4(32'hbb74181f),
	.w5(32'h3b11a268),
	.w6(32'h3b1bafd2),
	.w7(32'hbb532376),
	.w8(32'hbb6342f3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40f91d),
	.w1(32'h3b66fa7f),
	.w2(32'h3b0974c0),
	.w3(32'hbbb2d106),
	.w4(32'h3a7f2b1d),
	.w5(32'hbb864188),
	.w6(32'hbbc05ff7),
	.w7(32'h397b9912),
	.w8(32'hbaef6c80),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92e623),
	.w1(32'h3ac40b03),
	.w2(32'h3c1cb405),
	.w3(32'hbb8968bc),
	.w4(32'hbb0d6e46),
	.w5(32'h3bffd155),
	.w6(32'h3ab53232),
	.w7(32'hbb500a0e),
	.w8(32'hbb566e8e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc6a6e),
	.w1(32'h38af6576),
	.w2(32'hbb66c325),
	.w3(32'h3b884352),
	.w4(32'hbba801e6),
	.w5(32'h39881c37),
	.w6(32'h3b3aa199),
	.w7(32'hbc0bde63),
	.w8(32'hbb31e78c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf58ac3),
	.w1(32'h3b4f25f6),
	.w2(32'h392835ac),
	.w3(32'h3b88bcb9),
	.w4(32'h39c14805),
	.w5(32'h3b8e6282),
	.w6(32'h3c0bea2e),
	.w7(32'h3b299ff9),
	.w8(32'h3b8d585e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce1c87),
	.w1(32'h3bc01c88),
	.w2(32'hbbad840a),
	.w3(32'h3b349839),
	.w4(32'h3b24518c),
	.w5(32'hbc2cc24a),
	.w6(32'h3b09677b),
	.w7(32'h3b3bcfd2),
	.w8(32'hb8b7cb6e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4f44),
	.w1(32'hbc893761),
	.w2(32'h3bae1b52),
	.w3(32'hbae6c321),
	.w4(32'hbcf0fc0d),
	.w5(32'h3d08eec0),
	.w6(32'h3b4a9d2b),
	.w7(32'hbbee1de0),
	.w8(32'hbbc6a6eb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34d62d),
	.w1(32'hbafa2479),
	.w2(32'hbb859552),
	.w3(32'h3c22a6a9),
	.w4(32'h37e3e98c),
	.w5(32'h3aacecc0),
	.w6(32'hbbbdb4d2),
	.w7(32'hbbf68138),
	.w8(32'hbb0c3380),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5c8f4),
	.w1(32'h3c084c96),
	.w2(32'h3ae3fd18),
	.w3(32'hb7de51c2),
	.w4(32'h3b629654),
	.w5(32'hbb521763),
	.w6(32'hbabcbd47),
	.w7(32'h3ad43d60),
	.w8(32'hbbc3b136),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6c10f),
	.w1(32'h3a638f56),
	.w2(32'h3b37db91),
	.w3(32'h3bc408b5),
	.w4(32'h3b8b4617),
	.w5(32'h3a8caa65),
	.w6(32'h3c0797d0),
	.w7(32'h3a0d75a8),
	.w8(32'h38ada367),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b425b46),
	.w1(32'hbb164839),
	.w2(32'hbb0af3ca),
	.w3(32'h3c1b435f),
	.w4(32'h3ba6c81a),
	.w5(32'h3b96ac7c),
	.w6(32'hb9263a98),
	.w7(32'h3c193d27),
	.w8(32'hba619060),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08cb9b),
	.w1(32'hbb6b9776),
	.w2(32'h3b8e006e),
	.w3(32'h3b8b3609),
	.w4(32'hbb8b5b69),
	.w5(32'h3b7873bd),
	.w6(32'h39a8b8d5),
	.w7(32'h3a3f16d4),
	.w8(32'h3bffd114),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e67501),
	.w1(32'h3b0ae281),
	.w2(32'h3c3e6642),
	.w3(32'h3a72acfc),
	.w4(32'h3c0d37ea),
	.w5(32'h3c667162),
	.w6(32'h3a5d6433),
	.w7(32'h3abe4b7f),
	.w8(32'h3bb3d6b9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7de2c2),
	.w1(32'h3b74032d),
	.w2(32'h3b1bcc28),
	.w3(32'h3c1b1fac),
	.w4(32'hbb60d08a),
	.w5(32'h3b783169),
	.w6(32'hbb911949),
	.w7(32'hbacb6db5),
	.w8(32'h3bddaf2c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514d4d),
	.w1(32'h3b2ae3b2),
	.w2(32'h393cafc7),
	.w3(32'h3b0cab01),
	.w4(32'h3ba22f08),
	.w5(32'h3b50b618),
	.w6(32'h3b82fbb4),
	.w7(32'h3a1b90e5),
	.w8(32'h3b2a20db),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b589f8a),
	.w1(32'hb9a13a62),
	.w2(32'h3bff2f80),
	.w3(32'h3a6b6f62),
	.w4(32'h3b3b09cb),
	.w5(32'h3b8a91de),
	.w6(32'h3bb45a75),
	.w7(32'h3a616958),
	.w8(32'h3bb5532a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beadc12),
	.w1(32'hb9d48039),
	.w2(32'hbb79f014),
	.w3(32'h3c32dc6b),
	.w4(32'hba17a42f),
	.w5(32'hbb5362b3),
	.w6(32'h3c32b000),
	.w7(32'h3b520c38),
	.w8(32'h3b9ec576),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba594fd1),
	.w1(32'hbb8a3326),
	.w2(32'h39ab67e4),
	.w3(32'hbb1b6b44),
	.w4(32'hbb0fe0b8),
	.w5(32'hbb253599),
	.w6(32'h3b15024f),
	.w7(32'hbb7a8bd8),
	.w8(32'h3a2cf1ab),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988f75f),
	.w1(32'h3b7eddce),
	.w2(32'h3bdd6a0f),
	.w3(32'h3a60eded),
	.w4(32'hbaa8ceaf),
	.w5(32'h3c287b1e),
	.w6(32'h3a8db054),
	.w7(32'h3a4d1664),
	.w8(32'h3c1ce243),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be82a),
	.w1(32'hbb180944),
	.w2(32'hbba3194c),
	.w3(32'h3c453ac0),
	.w4(32'hbc043152),
	.w5(32'hbbade0b1),
	.w6(32'h3bc42bb0),
	.w7(32'hba794230),
	.w8(32'hbbbf9e2d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa0115),
	.w1(32'hbb8a0345),
	.w2(32'hbace91fc),
	.w3(32'hbb2ba180),
	.w4(32'h3a64e217),
	.w5(32'hba38bcb5),
	.w6(32'h3ae589ad),
	.w7(32'h3a504564),
	.w8(32'h3adf0329),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule