module layer_10_featuremap_487(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a143ec6),
	.w1(32'hb8dac835),
	.w2(32'hba163503),
	.w3(32'h39794ddf),
	.w4(32'hba16d5fa),
	.w5(32'h3a008d94),
	.w6(32'h3a663dd5),
	.w7(32'hb9e233f1),
	.w8(32'hba321c8e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ed685),
	.w1(32'h3a9a7200),
	.w2(32'h39ee0bbf),
	.w3(32'h3a2ed69a),
	.w4(32'hba2a6814),
	.w5(32'hbaa13095),
	.w6(32'h3923edd5),
	.w7(32'hbb2beb80),
	.w8(32'hbacf6c6c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6baac),
	.w1(32'hba433c6d),
	.w2(32'hbad5392b),
	.w3(32'h396359e9),
	.w4(32'hb9f9feee),
	.w5(32'hbad03754),
	.w6(32'hb7b32bbe),
	.w7(32'h3a4bec15),
	.w8(32'hba2e3456),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f468b),
	.w1(32'h3a2a2f84),
	.w2(32'h39791f4e),
	.w3(32'hba506666),
	.w4(32'h3a2d69f2),
	.w5(32'h3b09623a),
	.w6(32'hb7e0ea35),
	.w7(32'h39f867a8),
	.w8(32'h3a360825),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba204b32),
	.w1(32'h3a528bf0),
	.w2(32'h3a0a8312),
	.w3(32'hb998a776),
	.w4(32'h3a824bb7),
	.w5(32'h3a0986c6),
	.w6(32'hb94afc4b),
	.w7(32'h39f6f602),
	.w8(32'h394eb966),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5a899),
	.w1(32'hb9c4cd81),
	.w2(32'h39c71e86),
	.w3(32'h39b3b284),
	.w4(32'hb99938e6),
	.w5(32'hbaabd2d9),
	.w6(32'hba0fc1a8),
	.w7(32'hb9d48d1a),
	.w8(32'h38fe15c4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bf725),
	.w1(32'hbb09088d),
	.w2(32'hbb24ecb9),
	.w3(32'h3b8e11f6),
	.w4(32'h38b33f08),
	.w5(32'h3ac56e00),
	.w6(32'h3a8adf83),
	.w7(32'hbaa5eaf9),
	.w8(32'hba6e8d8c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeb67f),
	.w1(32'hbc24adf0),
	.w2(32'hbc031333),
	.w3(32'hbbfcc84b),
	.w4(32'hbb328784),
	.w5(32'h3a6e7471),
	.w6(32'hbbded433),
	.w7(32'hbbbc5c4b),
	.w8(32'h3abccdbf),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2897a6),
	.w1(32'h3adf9678),
	.w2(32'h39a6f9ac),
	.w3(32'h3aafcf0d),
	.w4(32'h3aabb485),
	.w5(32'hb9fa0540),
	.w6(32'h3b6ef9e2),
	.w7(32'h3b4140c0),
	.w8(32'hb9ae644a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba29df),
	.w1(32'hba42eec3),
	.w2(32'hbab78d76),
	.w3(32'h3ac97df2),
	.w4(32'hb85190ed),
	.w5(32'hba23738c),
	.w6(32'hbb0fd970),
	.w7(32'h3b3d3a3b),
	.w8(32'hb985f141),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3f07c),
	.w1(32'hb8bd192b),
	.w2(32'h399d1876),
	.w3(32'h39c3175e),
	.w4(32'h3a148b38),
	.w5(32'h398621c1),
	.w6(32'hb995de0d),
	.w7(32'hb94d5b57),
	.w8(32'hb9cbf6f7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c2705),
	.w1(32'hb9c17380),
	.w2(32'h38f2f580),
	.w3(32'h3bc4b75a),
	.w4(32'h3aef045f),
	.w5(32'h3b538e41),
	.w6(32'h3b0d1842),
	.w7(32'hb91b17c2),
	.w8(32'h3a812fd9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae71cd0),
	.w1(32'hbb00a2af),
	.w2(32'hbb38a688),
	.w3(32'h3aec53fe),
	.w4(32'hba0099a1),
	.w5(32'hbac2f02b),
	.w6(32'h3a67d0cf),
	.w7(32'h37e41e2e),
	.w8(32'hba65f493),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397235d3),
	.w1(32'hba7f747f),
	.w2(32'hbad57379),
	.w3(32'hba890820),
	.w4(32'hbb05bc11),
	.w5(32'hbacaba44),
	.w6(32'hb9a23a8b),
	.w7(32'hbac53f98),
	.w8(32'hba951e9b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40db02),
	.w1(32'h3afca23c),
	.w2(32'hba0f1bf1),
	.w3(32'h3a262840),
	.w4(32'h3ae81be0),
	.w5(32'hba2b35a0),
	.w6(32'h39bbd485),
	.w7(32'h3ab74ea7),
	.w8(32'h3ac77bec),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bd194),
	.w1(32'h39faf461),
	.w2(32'hbab16b7d),
	.w3(32'hbb18ba15),
	.w4(32'hbaa1e82b),
	.w5(32'hba8107de),
	.w6(32'hbb50057d),
	.w7(32'h3a86c9bc),
	.w8(32'h398ae512),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a653782),
	.w1(32'hbaf31663),
	.w2(32'hbad006b6),
	.w3(32'hb9a44080),
	.w4(32'hbabd8a78),
	.w5(32'hbb321542),
	.w6(32'hb890b905),
	.w7(32'hba9e5370),
	.w8(32'hbac6b2be),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1331b),
	.w1(32'hbc173a59),
	.w2(32'hbbe6e82d),
	.w3(32'hbbf82b3a),
	.w4(32'hbbd66554),
	.w5(32'hbb2aa3eb),
	.w6(32'hbbbbd5c2),
	.w7(32'hbb5b360f),
	.w8(32'hbb01a932),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6df513),
	.w1(32'hbba06123),
	.w2(32'hbb106c06),
	.w3(32'hbb2693a0),
	.w4(32'hbb0b78fa),
	.w5(32'hb9bfcaf0),
	.w6(32'hbaea98fc),
	.w7(32'hb948713d),
	.w8(32'h39f52a12),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11660c),
	.w1(32'hba037fb0),
	.w2(32'h3abef173),
	.w3(32'h398b1655),
	.w4(32'h393eb21f),
	.w5(32'hb9f22331),
	.w6(32'h39096ddb),
	.w7(32'h393ffddb),
	.w8(32'h3b34ad8e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa32f4),
	.w1(32'h3a4ba3b8),
	.w2(32'h3b04dd85),
	.w3(32'hb921a4a9),
	.w4(32'h3aaaac2b),
	.w5(32'h3a3d33a8),
	.w6(32'h3a5ed211),
	.w7(32'h38532cd5),
	.w8(32'hba29dc58),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b135900),
	.w1(32'h3a52c205),
	.w2(32'h3ad325d3),
	.w3(32'h3ae0c20f),
	.w4(32'h3a4c61f8),
	.w5(32'hb9b7332f),
	.w6(32'h39ed35d1),
	.w7(32'hba89b8b3),
	.w8(32'hb96068e0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc434ff2),
	.w1(32'hbc1e981c),
	.w2(32'hbb8f5db9),
	.w3(32'hbbcc613c),
	.w4(32'hbbc9c188),
	.w5(32'hba58b365),
	.w6(32'hbc415045),
	.w7(32'hbb85b622),
	.w8(32'h3b0bd8a4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad66e22),
	.w1(32'h3a6c9b22),
	.w2(32'hbb060fff),
	.w3(32'h3b4e5223),
	.w4(32'h396a642e),
	.w5(32'hbb37f507),
	.w6(32'h3acb0c2d),
	.w7(32'h39fe7ed3),
	.w8(32'hbb5373cc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8625f5),
	.w1(32'h3bb28cff),
	.w2(32'h3b182148),
	.w3(32'hb8647868),
	.w4(32'h39634b77),
	.w5(32'hbaa7b62a),
	.w6(32'hbb09d659),
	.w7(32'hbb693743),
	.w8(32'hbbb5e56e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdb14f),
	.w1(32'h3aeec67e),
	.w2(32'h3b04b996),
	.w3(32'h3a9c1697),
	.w4(32'h3a0e5367),
	.w5(32'h3ab44138),
	.w6(32'hbb28a76b),
	.w7(32'h3a89bef9),
	.w8(32'h3a85e849),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a82e1),
	.w1(32'h3b3da69a),
	.w2(32'h3b67c726),
	.w3(32'h3b0da112),
	.w4(32'h3b835f2d),
	.w5(32'h3b61cfb7),
	.w6(32'h3aa4efcf),
	.w7(32'h3b0eac35),
	.w8(32'h3ad499c2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6118d7),
	.w1(32'h3ab842a6),
	.w2(32'h39fae57f),
	.w3(32'h3b1c592a),
	.w4(32'h3a9428c9),
	.w5(32'hbb6c76b7),
	.w6(32'h3b2c3fd5),
	.w7(32'h3b856d08),
	.w8(32'hbafff23f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d98ec),
	.w1(32'h3a4d1808),
	.w2(32'hb913f504),
	.w3(32'h3accdbb3),
	.w4(32'h3acc697f),
	.w5(32'h3aec4a3c),
	.w6(32'h3abaf344),
	.w7(32'h3abddcc3),
	.w8(32'h3a92da91),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b0973),
	.w1(32'h3be503e6),
	.w2(32'h3b583fc5),
	.w3(32'h3b281a92),
	.w4(32'h3a94eb16),
	.w5(32'hba8e0eb6),
	.w6(32'h3b3d0b17),
	.w7(32'h3b38ce44),
	.w8(32'hbad5be4f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399433d9),
	.w1(32'hb9d6f433),
	.w2(32'hba1b615f),
	.w3(32'h3a62e2e1),
	.w4(32'hbadbd244),
	.w5(32'hbb23881d),
	.w6(32'h3a0fd9c1),
	.w7(32'hb9e870ad),
	.w8(32'hba171931),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba841a6c),
	.w1(32'h3a3eb88b),
	.w2(32'hba2270ea),
	.w3(32'hbb4be83a),
	.w4(32'h3aabb8fe),
	.w5(32'hb9fb3111),
	.w6(32'hba2737fa),
	.w7(32'h3a9a21c7),
	.w8(32'h39f825b8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a232ff),
	.w1(32'hb99a6100),
	.w2(32'hb7f192b3),
	.w3(32'h3a5ba0d0),
	.w4(32'h389daa42),
	.w5(32'h3b09e7ca),
	.w6(32'hb7451d4c),
	.w7(32'h3a67a1a3),
	.w8(32'h3ae83e36),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8abb67),
	.w1(32'h3a6bca6c),
	.w2(32'hba74f1d7),
	.w3(32'h39b9f7d0),
	.w4(32'hba60db0b),
	.w5(32'h3a0d1b76),
	.w6(32'hba1afb64),
	.w7(32'hbafd4cbc),
	.w8(32'hbab5eded),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a69763),
	.w1(32'h3a8ec70e),
	.w2(32'h3a5322f2),
	.w3(32'hba3ca99f),
	.w4(32'hba98b553),
	.w5(32'h3a8e51b3),
	.w6(32'h39460322),
	.w7(32'hb7ef937a),
	.w8(32'h39a103f7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af962fe),
	.w1(32'hba18dbe4),
	.w2(32'hb9f47b04),
	.w3(32'h3ab8a92f),
	.w4(32'hba09ab77),
	.w5(32'h3a3507cf),
	.w6(32'hb9f6d490),
	.w7(32'h3a6411a7),
	.w8(32'h39e04423),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4be80a),
	.w1(32'hbc098744),
	.w2(32'h39ef4214),
	.w3(32'hb9941c6c),
	.w4(32'hbb907e02),
	.w5(32'h3b1c5422),
	.w6(32'hbaa41b02),
	.w7(32'hbc107b50),
	.w8(32'h3b0edaa7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e33c1),
	.w1(32'h3bd54cd3),
	.w2(32'hba2d06e7),
	.w3(32'h3b7b6fe3),
	.w4(32'h3b4aa965),
	.w5(32'hbb3b77dd),
	.w6(32'h3b2e3557),
	.w7(32'hbb706f76),
	.w8(32'hbb9b9547),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6c3e6),
	.w1(32'h3bc04cab),
	.w2(32'hba195cdf),
	.w3(32'h3bd8a152),
	.w4(32'h3b3dac65),
	.w5(32'hbba0b1cc),
	.w6(32'h3c162c48),
	.w7(32'h3b0e2f9c),
	.w8(32'hbb35b0c8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9fd8a),
	.w1(32'h3ab09868),
	.w2(32'hba6ef969),
	.w3(32'h3ad1a30c),
	.w4(32'hb93872ae),
	.w5(32'hba83b509),
	.w6(32'h3acff853),
	.w7(32'h393d8308),
	.w8(32'hba62798c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c111b),
	.w1(32'h3a0a735d),
	.w2(32'h3838d98a),
	.w3(32'hba2ae08b),
	.w4(32'h3a097e57),
	.w5(32'h39bf24ef),
	.w6(32'h3824380f),
	.w7(32'hb9f4c2d3),
	.w8(32'hb9a6c019),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60dafc),
	.w1(32'hba4c099e),
	.w2(32'h39cdab23),
	.w3(32'hba006eab),
	.w4(32'h38d8fdfb),
	.w5(32'h3a581af9),
	.w6(32'h3a3ddf4a),
	.w7(32'hb9e32fce),
	.w8(32'h3a9373a8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a276fdd),
	.w1(32'h3aa0b819),
	.w2(32'h3a6afdeb),
	.w3(32'h39f76849),
	.w4(32'h39e94be2),
	.w5(32'h3a269431),
	.w6(32'hb9edb597),
	.w7(32'h3a32e203),
	.w8(32'h39c35c5b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc79085),
	.w1(32'hba9f67b7),
	.w2(32'hbb118eb0),
	.w3(32'hbb4bc418),
	.w4(32'h3a02c312),
	.w5(32'h3a304834),
	.w6(32'hbb3dc8dd),
	.w7(32'h3b95bf02),
	.w8(32'h3b455812),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39591949),
	.w1(32'h3b1b6473),
	.w2(32'hb9563a2d),
	.w3(32'h3a8c569e),
	.w4(32'h3b1dc47f),
	.w5(32'h3a2b56ce),
	.w6(32'h3a84ac4b),
	.w7(32'h3af897b8),
	.w8(32'hba3a7f6d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a6dae),
	.w1(32'h3b20dd05),
	.w2(32'hb922ccaf),
	.w3(32'h3b343b68),
	.w4(32'h3b054daa),
	.w5(32'h3a7b844e),
	.w6(32'hba1fa203),
	.w7(32'h3a9b1e10),
	.w8(32'hba3901be),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de0ab5),
	.w1(32'h3a3b30fb),
	.w2(32'hba0b74d3),
	.w3(32'hb7e12b6f),
	.w4(32'hb8ee2b14),
	.w5(32'hb9ce222d),
	.w6(32'hbb15ecd5),
	.w7(32'h39ad5273),
	.w8(32'hbaa0ec54),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42aa59),
	.w1(32'hbc230a46),
	.w2(32'hbc02b629),
	.w3(32'hbb2e508a),
	.w4(32'hbb719933),
	.w5(32'hbaaa6ea7),
	.w6(32'hbbb29a85),
	.w7(32'hba73e181),
	.w8(32'h3ae816bf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd534d),
	.w1(32'h3a20e920),
	.w2(32'h398bd990),
	.w3(32'hb9285c4c),
	.w4(32'h3a7d69b4),
	.w5(32'hb8a61726),
	.w6(32'hb89171c4),
	.w7(32'h396c2c92),
	.w8(32'hba417872),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987acb3),
	.w1(32'h3aa48743),
	.w2(32'h3ade65ac),
	.w3(32'hba06d081),
	.w4(32'h3a592915),
	.w5(32'h39f5e580),
	.w6(32'hba0636ae),
	.w7(32'h3a752b96),
	.w8(32'h39a89ef2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a297f8b),
	.w1(32'hb9fc9f31),
	.w2(32'hbab2aaac),
	.w3(32'h39dcc110),
	.w4(32'h39e2de70),
	.w5(32'hba8d4e5f),
	.w6(32'h3af0d6ae),
	.w7(32'h393254b4),
	.w8(32'hba5152c1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34db27),
	.w1(32'hbabed579),
	.w2(32'hbb41dff3),
	.w3(32'hba90d5a4),
	.w4(32'h3a03a8c9),
	.w5(32'hbb3497ed),
	.w6(32'hbaec3628),
	.w7(32'hbaf07ca6),
	.w8(32'hba953ce0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f0ae1),
	.w1(32'hbadf93ac),
	.w2(32'hbb0f6a1c),
	.w3(32'hba9b0f13),
	.w4(32'hba9e4346),
	.w5(32'hba1c0373),
	.w6(32'hbac56910),
	.w7(32'hba87e140),
	.w8(32'hba5dc623),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaa6cc),
	.w1(32'hbc0f6b0b),
	.w2(32'hbbafed5f),
	.w3(32'hbb2fa531),
	.w4(32'hbb5b1f94),
	.w5(32'h39cda9cd),
	.w6(32'hbb4a2919),
	.w7(32'h3adb5b34),
	.w8(32'h3b5d016b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe93aa),
	.w1(32'hba95885b),
	.w2(32'hbb804de9),
	.w3(32'h36ea02e4),
	.w4(32'hb9aaf3c6),
	.w5(32'hbb21c54d),
	.w6(32'h3a7e23c2),
	.w7(32'h399cd583),
	.w8(32'hbabb4c0b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefcd78),
	.w1(32'h3af62db7),
	.w2(32'h3aaa0395),
	.w3(32'hbb017b49),
	.w4(32'h363ce2df),
	.w5(32'hba667609),
	.w6(32'hbaa881ff),
	.w7(32'hb9a14f20),
	.w8(32'h3aa39ef6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa012b6),
	.w1(32'h39468334),
	.w2(32'h3a3c3cb4),
	.w3(32'h3a63bd47),
	.w4(32'hba4661df),
	.w5(32'h39824b2d),
	.w6(32'h3a6643d0),
	.w7(32'hba891b23),
	.w8(32'hba714c08),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a384190),
	.w1(32'hbacd64e2),
	.w2(32'hb9abf594),
	.w3(32'h39a4cd3f),
	.w4(32'hba9fc1d7),
	.w5(32'hba4103b5),
	.w6(32'hba1e77c6),
	.w7(32'hba256eba),
	.w8(32'h394e2c87),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9034a87),
	.w1(32'hba12d3d6),
	.w2(32'hba8614c1),
	.w3(32'h3a547efb),
	.w4(32'h3a6c4b31),
	.w5(32'hba12613f),
	.w6(32'h3a269148),
	.w7(32'hb8e9d5f6),
	.w8(32'h39c208ec),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921268c),
	.w1(32'hbb48ad4d),
	.w2(32'hbb24187c),
	.w3(32'h3a20c6a3),
	.w4(32'hbb8086df),
	.w5(32'hbb95a824),
	.w6(32'h39edd4f7),
	.w7(32'hba225522),
	.w8(32'hbb249472),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb471e99),
	.w1(32'hbb03e315),
	.w2(32'hbb3ccf59),
	.w3(32'hbb1eccf2),
	.w4(32'hbadd634e),
	.w5(32'hbb449d89),
	.w6(32'hbb271a1a),
	.w7(32'h3a2348a0),
	.w8(32'hba59727e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c1813),
	.w1(32'hbb2a5f46),
	.w2(32'hbabccdc1),
	.w3(32'hbc0143d0),
	.w4(32'hbb019ed8),
	.w5(32'hbb512eb3),
	.w6(32'hbb91f9ce),
	.w7(32'hba734e21),
	.w8(32'hb9bc247f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba344f37),
	.w1(32'hba87e061),
	.w2(32'hba8d8b14),
	.w3(32'hba03db24),
	.w4(32'hbaea9102),
	.w5(32'hbaddf26d),
	.w6(32'h385a286e),
	.w7(32'hbab60323),
	.w8(32'hbac4c860),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed7eb7),
	.w1(32'hba23213f),
	.w2(32'h393fb545),
	.w3(32'hbb0b9f8a),
	.w4(32'hba616f98),
	.w5(32'hb9ff3723),
	.w6(32'hbafd5d7d),
	.w7(32'hba6cb5bc),
	.w8(32'hbaa94034),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed41b8),
	.w1(32'h3b10968f),
	.w2(32'h3b1f2ef9),
	.w3(32'hba57bd04),
	.w4(32'h3b0136ff),
	.w5(32'h3af3f323),
	.w6(32'hb9938b97),
	.w7(32'h3b144176),
	.w8(32'h3aeda14f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b222d64),
	.w1(32'h3ac3470f),
	.w2(32'h37c52b32),
	.w3(32'h3b046cb2),
	.w4(32'h3ac9d628),
	.w5(32'h39c72dba),
	.w6(32'h3b5c34bb),
	.w7(32'h39bec6c2),
	.w8(32'h3a569a8b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fe6f0),
	.w1(32'hbb8e89c0),
	.w2(32'hbac67a8f),
	.w3(32'h3b8cf3d0),
	.w4(32'hbb0156ab),
	.w5(32'hba9c36d5),
	.w6(32'hba867fb6),
	.w7(32'h384fe66d),
	.w8(32'hbaf47771),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b554ef4),
	.w1(32'h3b09cf17),
	.w2(32'hbb291336),
	.w3(32'h38e19cac),
	.w4(32'h3aa173bf),
	.w5(32'hba1b68b4),
	.w6(32'hbbc3ddc6),
	.w7(32'h38fec864),
	.w8(32'hbaa61c50),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7d2cf),
	.w1(32'hbb3402b2),
	.w2(32'hbb10fa30),
	.w3(32'hbb783c73),
	.w4(32'hba37b243),
	.w5(32'h3a675071),
	.w6(32'hbb73bb7e),
	.w7(32'hbac24b9a),
	.w8(32'hba557d42),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82aa08),
	.w1(32'h3b9313c3),
	.w2(32'hbc95f20a),
	.w3(32'h3b8e475d),
	.w4(32'hbb53d178),
	.w5(32'hbca9c760),
	.w6(32'h393b1e6a),
	.w7(32'hbc677cac),
	.w8(32'hbcaa8c4f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af84b4f),
	.w1(32'hba0d2d5e),
	.w2(32'h3abca616),
	.w3(32'h3c002cbe),
	.w4(32'h3a6c2eee),
	.w5(32'hbaa2be73),
	.w6(32'h3b4b93b2),
	.w7(32'hba59e791),
	.w8(32'h3b802441),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b414299),
	.w1(32'hb99ad260),
	.w2(32'hbb6e9886),
	.w3(32'hba0c7a85),
	.w4(32'h3a0c9da5),
	.w5(32'hbb8d94ee),
	.w6(32'h3c0fed07),
	.w7(32'hb9aa48d1),
	.w8(32'h3b935886),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfba20),
	.w1(32'hbb62489f),
	.w2(32'hbb46be03),
	.w3(32'h3c0bf230),
	.w4(32'hb9b13fcb),
	.w5(32'hbbf097b3),
	.w6(32'hbbd2ca92),
	.w7(32'hbb03d991),
	.w8(32'hbb84b53e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be036e1),
	.w1(32'hbbb07a75),
	.w2(32'hbbe7003a),
	.w3(32'h3c136ec8),
	.w4(32'hbb5ae5da),
	.w5(32'hbb4f2206),
	.w6(32'h3b2f1078),
	.w7(32'h3b93d566),
	.w8(32'h3b08ecca),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb243316),
	.w1(32'h3b308806),
	.w2(32'h3b3e1fbe),
	.w3(32'h39b2edbb),
	.w4(32'h3c210bbe),
	.w5(32'hbc0fec9a),
	.w6(32'h3aaac1ec),
	.w7(32'h3ba3a3fa),
	.w8(32'hbbe362ef),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be938f4),
	.w1(32'hbc25fc1c),
	.w2(32'hba804f7c),
	.w3(32'h3b75f7f2),
	.w4(32'hbbb9f636),
	.w5(32'hbb307c9a),
	.w6(32'hba3714d9),
	.w7(32'h3ba62de4),
	.w8(32'hbb1e2c8b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39547c),
	.w1(32'hbb51cbb2),
	.w2(32'hbb2c2553),
	.w3(32'hbc276ed6),
	.w4(32'h3b35b572),
	.w5(32'h3c58b028),
	.w6(32'hbc48672c),
	.w7(32'hbb90f7f5),
	.w8(32'h3b149fd1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bd37e),
	.w1(32'hbbba0c53),
	.w2(32'hbc2a8337),
	.w3(32'h3bf1fff0),
	.w4(32'hbbc112c5),
	.w5(32'hbc6fd23f),
	.w6(32'h3a99673d),
	.w7(32'hbb912ef8),
	.w8(32'hbbe2db51),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fe7d7),
	.w1(32'h3a692e0c),
	.w2(32'hba024554),
	.w3(32'hbc18be97),
	.w4(32'h3bdd5ac1),
	.w5(32'hba77256f),
	.w6(32'h3ab204b9),
	.w7(32'h3bd6d9a1),
	.w8(32'h3ad5a372),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e0f26),
	.w1(32'hbb9bf65d),
	.w2(32'h3be225a5),
	.w3(32'hbbbbbbd7),
	.w4(32'h3a1fe402),
	.w5(32'hbc5547c9),
	.w6(32'h3adb045e),
	.w7(32'h3b81e5ed),
	.w8(32'hbbeeca31),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba73b27),
	.w1(32'h3bd1b714),
	.w2(32'hbb662599),
	.w3(32'h3bece2ea),
	.w4(32'h3c15b617),
	.w5(32'hbbe61b08),
	.w6(32'h3aab9144),
	.w7(32'h3c0e1bee),
	.w8(32'hbbd97b36),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104410),
	.w1(32'hbaad8a82),
	.w2(32'hbb4c2c9c),
	.w3(32'hbc8407a8),
	.w4(32'h3af09a14),
	.w5(32'h3b903a80),
	.w6(32'hbb87dc90),
	.w7(32'h3b448558),
	.w8(32'h3a6ab8a6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed671c),
	.w1(32'hbb3f70ce),
	.w2(32'hbb8b3135),
	.w3(32'hbc0622b8),
	.w4(32'h39cd6dd7),
	.w5(32'hbb0296db),
	.w6(32'hbbcb310a),
	.w7(32'h3b0c380b),
	.w8(32'h3ad6e7b5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3cf8a),
	.w1(32'hbc05a9ce),
	.w2(32'hbbe70873),
	.w3(32'h3a0e559f),
	.w4(32'hbba24cc4),
	.w5(32'hbb2f12d1),
	.w6(32'hbb8b29c2),
	.w7(32'hbbadf532),
	.w8(32'h3ba062a1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96550b),
	.w1(32'h3a231ceb),
	.w2(32'h3a619c57),
	.w3(32'h3a864921),
	.w4(32'h3b6fb45a),
	.w5(32'h3b89400d),
	.w6(32'h3c517b90),
	.w7(32'hbb2d7f44),
	.w8(32'hbb4788de),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c371795),
	.w1(32'hbb8e8447),
	.w2(32'hbc111908),
	.w3(32'h3b3cb5eb),
	.w4(32'hbc642bab),
	.w5(32'hbb7f5a27),
	.w6(32'h3b8d94f5),
	.w7(32'hbc6f491c),
	.w8(32'hbc8e72ec),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc458b98),
	.w1(32'hbb623faa),
	.w2(32'h3b367d76),
	.w3(32'hbc6f86f5),
	.w4(32'h3b5a1b2a),
	.w5(32'h3a0226ea),
	.w6(32'hbc923875),
	.w7(32'hbbc9f80a),
	.w8(32'hbb8bd48b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b168aee),
	.w1(32'h38c85db6),
	.w2(32'h3b6cd7c3),
	.w3(32'h3bbe05f3),
	.w4(32'hb834f317),
	.w5(32'h3ba10d72),
	.w6(32'h3b230e9f),
	.w7(32'hbbb52ce5),
	.w8(32'hbbba9973),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35d75c),
	.w1(32'hbb87e78f),
	.w2(32'h3af0c849),
	.w3(32'hbb8dc63b),
	.w4(32'h39f23ce6),
	.w5(32'h3c15a041),
	.w6(32'hbc609b76),
	.w7(32'hbbb0e381),
	.w8(32'hbaa8f591),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccf88e),
	.w1(32'hbbe4d2d4),
	.w2(32'hbbd9518f),
	.w3(32'hbc24d4e9),
	.w4(32'hbbc9d3de),
	.w5(32'h3a4a648e),
	.w6(32'hbc1a9229),
	.w7(32'h3b0dec89),
	.w8(32'h3ba28498),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc621186),
	.w1(32'hbae19c38),
	.w2(32'hbc0997e0),
	.w3(32'hbc6a75b9),
	.w4(32'h3b976cb6),
	.w5(32'h3bcd1f5e),
	.w6(32'hbb7611df),
	.w7(32'h396ac3d9),
	.w8(32'h3b5cd786),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1090e1),
	.w1(32'hbbc48a9f),
	.w2(32'hbb1fb1b1),
	.w3(32'hb9a3fee6),
	.w4(32'hbc026788),
	.w5(32'hbc2734cf),
	.w6(32'hbb23d912),
	.w7(32'h39d4d6da),
	.w8(32'h3b324f43),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3f9e8),
	.w1(32'h3bf54c4c),
	.w2(32'h3b374447),
	.w3(32'hbc403d00),
	.w4(32'h3c5f6dee),
	.w5(32'h3c402a8f),
	.w6(32'h3ad7c1cf),
	.w7(32'h3b3adea7),
	.w8(32'hba98656e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbed509),
	.w1(32'h3b110748),
	.w2(32'h39b4a7aa),
	.w3(32'hba8839ea),
	.w4(32'h3b329357),
	.w5(32'h3bb22fac),
	.w6(32'hbb827010),
	.w7(32'h3af58189),
	.w8(32'h3ae1e3c9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e66e6),
	.w1(32'hbb5e9ab1),
	.w2(32'h39c05762),
	.w3(32'hbbc6586a),
	.w4(32'hbb5b4b99),
	.w5(32'hbc777ad3),
	.w6(32'hbb358c7b),
	.w7(32'h3bae3d43),
	.w8(32'hbbc15271),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe32933),
	.w1(32'hbc6accf9),
	.w2(32'hbc79f480),
	.w3(32'hbb85a1e0),
	.w4(32'hbc3e5351),
	.w5(32'hbc6df08a),
	.w6(32'h3a8b6fa5),
	.w7(32'hbb9e08b0),
	.w8(32'hb902b9ee),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ae84a),
	.w1(32'h3bf60801),
	.w2(32'h3b0d320e),
	.w3(32'h3bdf966c),
	.w4(32'h3bbb7b94),
	.w5(32'h3c23d041),
	.w6(32'h3b3e4e14),
	.w7(32'hbaffa88e),
	.w8(32'hbc07ea42),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a973),
	.w1(32'h3ae0ca33),
	.w2(32'hbb0d1332),
	.w3(32'h3b498a80),
	.w4(32'h3bb25cd3),
	.w5(32'h3b2a5c08),
	.w6(32'hbc259a71),
	.w7(32'h3c764d88),
	.w8(32'h3b9ab4dd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3520f7),
	.w1(32'hbb988d93),
	.w2(32'hbb21b7c4),
	.w3(32'hbb8c94a8),
	.w4(32'hbb7f5629),
	.w5(32'hbbc88adf),
	.w6(32'hbb1e84d6),
	.w7(32'hbbbb8c9c),
	.w8(32'hbbbc2a94),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0339a1),
	.w1(32'hbc6aaff1),
	.w2(32'hbc51ebba),
	.w3(32'hbc421faf),
	.w4(32'hbc870b94),
	.w5(32'hbc82d761),
	.w6(32'hbc3394ce),
	.w7(32'hbbd450c7),
	.w8(32'h3b849af9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbace695),
	.w1(32'h3b85b926),
	.w2(32'h3b98afc0),
	.w3(32'hbc7bcce4),
	.w4(32'h3b950f82),
	.w5(32'h3be5c81d),
	.w6(32'hbba640e8),
	.w7(32'h3b8ab191),
	.w8(32'h363b4c88),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc21752),
	.w1(32'h3b6ee894),
	.w2(32'h3b837830),
	.w3(32'h3c28061a),
	.w4(32'h3b857bb4),
	.w5(32'h3bfc2bb9),
	.w6(32'h3b7feca1),
	.w7(32'h3b808e9b),
	.w8(32'h3bf361f9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eef9b),
	.w1(32'hbc8e739b),
	.w2(32'h3b024b54),
	.w3(32'h3a5c88cd),
	.w4(32'hbbb41fb4),
	.w5(32'hba8defe9),
	.w6(32'hbb1324b4),
	.w7(32'h3a96cf0f),
	.w8(32'h3c338e0f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bb3f7),
	.w1(32'h3b8fea69),
	.w2(32'h3b2fbd85),
	.w3(32'h3c06e118),
	.w4(32'h3a773754),
	.w5(32'h3afe2f52),
	.w6(32'h3c45f0f8),
	.w7(32'hba8a0ad1),
	.w8(32'h3bc0c7cc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c2b0f),
	.w1(32'hbbcc941f),
	.w2(32'hbc258710),
	.w3(32'hbc4223c4),
	.w4(32'h3abda578),
	.w5(32'hbae8fd6c),
	.w6(32'hbadf8d73),
	.w7(32'hbb8fc1e4),
	.w8(32'hbb8fc3e9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40057c),
	.w1(32'h3bd84540),
	.w2(32'h38b43bb3),
	.w3(32'h3ae50b8b),
	.w4(32'h3c02724d),
	.w5(32'h3bc9fbf7),
	.w6(32'hbbe2ef1d),
	.w7(32'hbb503725),
	.w8(32'hbc4ee6c3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba81303),
	.w1(32'hb9e29dd5),
	.w2(32'hbb2b1d68),
	.w3(32'hbc24b685),
	.w4(32'hbbb87bf8),
	.w5(32'h3b0f72c9),
	.w6(32'hbc86c549),
	.w7(32'hbabff7c4),
	.w8(32'hbb343cfc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f9ca5),
	.w1(32'hbc1e020f),
	.w2(32'hbc6915f1),
	.w3(32'hbba8e72b),
	.w4(32'hbc53e2ce),
	.w5(32'hbc79a160),
	.w6(32'hbad44118),
	.w7(32'hbc94b705),
	.w8(32'hbca5674c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6b4f),
	.w1(32'h3b50ee55),
	.w2(32'hba3a1864),
	.w3(32'h3ae46b79),
	.w4(32'h3b8aef40),
	.w5(32'h3b07103f),
	.w6(32'hbc327c7d),
	.w7(32'h3b8fa953),
	.w8(32'h3c0adae0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1406b2),
	.w1(32'h3a4cb63a),
	.w2(32'h3b120617),
	.w3(32'h3a454e58),
	.w4(32'h3b13a40a),
	.w5(32'hbc24b954),
	.w6(32'h3b97fa28),
	.w7(32'hbc0baea6),
	.w8(32'hbc3512fa),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918a52b),
	.w1(32'h3c4117b0),
	.w2(32'h3b87f4a4),
	.w3(32'hba173f30),
	.w4(32'hbb97e53f),
	.w5(32'hbbc86635),
	.w6(32'hbc024056),
	.w7(32'hbc234073),
	.w8(32'hbc35c08a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ea1f5),
	.w1(32'hbc1e1714),
	.w2(32'hbc86c98d),
	.w3(32'hbc75cd7d),
	.w4(32'hbaa4b214),
	.w5(32'hbb9703d1),
	.w6(32'hbc8bd0d9),
	.w7(32'h3aabfca8),
	.w8(32'hbb0e01ac),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69f5de),
	.w1(32'hbb63fafb),
	.w2(32'h3b70fe92),
	.w3(32'hbc37777f),
	.w4(32'hbb559ddd),
	.w5(32'h3bd69e5e),
	.w6(32'hbc442302),
	.w7(32'hba0a700a),
	.w8(32'hbad0cd61),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02de82),
	.w1(32'h3a0e02fc),
	.w2(32'h3bbe620e),
	.w3(32'h3b6c9d7b),
	.w4(32'hbb8ac93d),
	.w5(32'hbbc1ea19),
	.w6(32'h3a3c2eaf),
	.w7(32'h3bbcff1d),
	.w8(32'h3b63d6ed),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ef9fc),
	.w1(32'hbb18f381),
	.w2(32'hbc53a643),
	.w3(32'hbb3e0fab),
	.w4(32'hbb8a76bf),
	.w5(32'hbcaf24de),
	.w6(32'h3b48d09d),
	.w7(32'hbbc71cac),
	.w8(32'hbc8182ab),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1482d3),
	.w1(32'h3aebce51),
	.w2(32'hbbc1db71),
	.w3(32'hbc75e332),
	.w4(32'hb9bd9973),
	.w5(32'hbc19ec8e),
	.w6(32'hbc37c2bf),
	.w7(32'hbbf02cd8),
	.w8(32'hbc5da931),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3f2e3),
	.w1(32'h394d2d1b),
	.w2(32'hbc22088a),
	.w3(32'hbc5c39c6),
	.w4(32'hbbe33e10),
	.w5(32'hbbd0814c),
	.w6(32'hbc15fa3b),
	.w7(32'hba583cd4),
	.w8(32'hbb1c913e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37afa8),
	.w1(32'hbaf064f3),
	.w2(32'h3b2e36ef),
	.w3(32'hbc94eb58),
	.w4(32'hbaa81986),
	.w5(32'h3bf6859f),
	.w6(32'hbbc9e2df),
	.w7(32'hb9bb8682),
	.w8(32'h3b97aafb),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad02af4),
	.w1(32'hbb8868ca),
	.w2(32'hbb4b7808),
	.w3(32'h3bfa321f),
	.w4(32'h3b4b66cc),
	.w5(32'hbbecc18c),
	.w6(32'hb9a7dbf9),
	.w7(32'h3b8c6400),
	.w8(32'hbb31ad2d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f1d5e),
	.w1(32'h3ba7c8ef),
	.w2(32'h3ba2f49a),
	.w3(32'hbb65edaf),
	.w4(32'hba35e60b),
	.w5(32'hbbb700c9),
	.w6(32'hbaf8d448),
	.w7(32'h3c19da31),
	.w8(32'h3bce9d1f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83efca),
	.w1(32'hba44ee0d),
	.w2(32'h3bc74f41),
	.w3(32'h3c435881),
	.w4(32'hbae81d35),
	.w5(32'h3b5d2fc2),
	.w6(32'h3c2b7c79),
	.w7(32'hbb3ee10d),
	.w8(32'h3bb2123a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd26412),
	.w1(32'hbc67cd51),
	.w2(32'hbc93141f),
	.w3(32'h3a5d84be),
	.w4(32'hbc80b63c),
	.w5(32'hbc919df9),
	.w6(32'h3b86e1fa),
	.w7(32'hbc6db0ed),
	.w8(32'hbc14647b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf98bb),
	.w1(32'h3a734822),
	.w2(32'h3b109f62),
	.w3(32'hbc9aa192),
	.w4(32'hbab87683),
	.w5(32'hbb3c700c),
	.w6(32'h3c162570),
	.w7(32'hbbf11f49),
	.w8(32'hbc31f516),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58fb12),
	.w1(32'h3a2e3e69),
	.w2(32'hbbcded65),
	.w3(32'hb78cc73d),
	.w4(32'h3b15826c),
	.w5(32'hbb3e3ad1),
	.w6(32'hbbb4039c),
	.w7(32'h3b109e1c),
	.w8(32'hbb218dd0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030202),
	.w1(32'hbba3d176),
	.w2(32'hbb909ed6),
	.w3(32'hbc68f7ee),
	.w4(32'hbb3fbacb),
	.w5(32'hbc177312),
	.w6(32'hbc05727e),
	.w7(32'hbb0476a6),
	.w8(32'h3c1585a4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6407d1),
	.w1(32'h3b2d3a71),
	.w2(32'h3b76d127),
	.w3(32'h3b82fdbe),
	.w4(32'h3ae47bce),
	.w5(32'hbb0587e2),
	.w6(32'h3bdd21d6),
	.w7(32'hba9420e8),
	.w8(32'h3bd19c2f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1944ba),
	.w1(32'hbc205078),
	.w2(32'hbbbc1e57),
	.w3(32'h3c442332),
	.w4(32'hbc4d660c),
	.w5(32'hbc8097a3),
	.w6(32'h3be41034),
	.w7(32'hbc37a41f),
	.w8(32'hbb303ece),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5819),
	.w1(32'h3bc1f19a),
	.w2(32'h3b4e6e7e),
	.w3(32'h3bbb1dcd),
	.w4(32'h3b0c5a14),
	.w5(32'hbb057405),
	.w6(32'hbb636ac2),
	.w7(32'hbb5472e1),
	.w8(32'h3a97e0f6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3fbfa),
	.w1(32'hbbaf1b54),
	.w2(32'h3b674f43),
	.w3(32'h3b440eda),
	.w4(32'hbbbc4089),
	.w5(32'hbb66a30a),
	.w6(32'hbad7f46c),
	.w7(32'hbbb37f08),
	.w8(32'h3b3bdc28),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27818b),
	.w1(32'hba8df2c2),
	.w2(32'hbb6dd09b),
	.w3(32'h3c2af263),
	.w4(32'h3a91b5b5),
	.w5(32'hbb03c644),
	.w6(32'h3c184498),
	.w7(32'h3ba81531),
	.w8(32'h3af564c8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c505d),
	.w1(32'hbb408224),
	.w2(32'h3bddeda0),
	.w3(32'hbc3799fb),
	.w4(32'hbafb6965),
	.w5(32'h3b3c8eba),
	.w6(32'hbc403664),
	.w7(32'hbbd3509f),
	.w8(32'hbc023b57),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9311c9),
	.w1(32'hbb55fe12),
	.w2(32'hbb1b5720),
	.w3(32'h3bcf84b5),
	.w4(32'hbad33994),
	.w5(32'hbbe2cc5e),
	.w6(32'h3afed078),
	.w7(32'h3a933b25),
	.w8(32'hbb3827d3),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9325fb),
	.w1(32'hbaaea74d),
	.w2(32'hb9f91a11),
	.w3(32'hba000d33),
	.w4(32'h3a51262e),
	.w5(32'hba15219b),
	.w6(32'hbb205080),
	.w7(32'h3b76b24f),
	.w8(32'h3ac531e7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ebf21),
	.w1(32'hbbddb6f2),
	.w2(32'hbc8d56fd),
	.w3(32'hbc687a82),
	.w4(32'hbc21669e),
	.w5(32'hbcc88d13),
	.w6(32'hbbc4803c),
	.w7(32'h3b09dde5),
	.w8(32'hbc184104),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bb6e4),
	.w1(32'hbc564714),
	.w2(32'hbc25731f),
	.w3(32'hbcaed5d8),
	.w4(32'h3ad3d4c3),
	.w5(32'h372d8bcd),
	.w6(32'hbc7ed567),
	.w7(32'h3b86d1c7),
	.w8(32'h3bcd99d3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab2969),
	.w1(32'h39d9bd2e),
	.w2(32'h39aaaf0e),
	.w3(32'h3bbfe060),
	.w4(32'hbadbc630),
	.w5(32'h3bf5f24c),
	.w6(32'h3b305c5a),
	.w7(32'hbacffd14),
	.w8(32'h3b297a2e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ab39e),
	.w1(32'hbb565bcf),
	.w2(32'hb9d22803),
	.w3(32'hba908d97),
	.w4(32'hbbaa01f5),
	.w5(32'hb969a7ab),
	.w6(32'h3bdb0e33),
	.w7(32'h3afa641c),
	.w8(32'h3ba63f11),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3b015),
	.w1(32'hbb06a4e9),
	.w2(32'hbba31a0f),
	.w3(32'h3bcaca8d),
	.w4(32'h3b8a0d2f),
	.w5(32'h3b4d2e26),
	.w6(32'h3c12c1c3),
	.w7(32'h3b97d947),
	.w8(32'h3c698db3),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a4aee),
	.w1(32'hba51fd04),
	.w2(32'hbc25f10c),
	.w3(32'h3bd5788b),
	.w4(32'h3c0935ef),
	.w5(32'h3be28064),
	.w6(32'h3c32e6df),
	.w7(32'h3c27aa3c),
	.w8(32'h3c3c32c8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89e930),
	.w1(32'h3bf8cbc4),
	.w2(32'h3c19adc6),
	.w3(32'hbba6aacb),
	.w4(32'h3c71030d),
	.w5(32'h3c3d44ed),
	.w6(32'h3a6fa13d),
	.w7(32'h3b42ba52),
	.w8(32'h3b884d33),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe410a),
	.w1(32'h3baed240),
	.w2(32'hbad8bb7a),
	.w3(32'hbc3dc417),
	.w4(32'hba2a081f),
	.w5(32'hbae41b06),
	.w6(32'hbc3bada9),
	.w7(32'hbc0a7056),
	.w8(32'hbc350372),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17acee),
	.w1(32'h3b8de41a),
	.w2(32'h3ba283b5),
	.w3(32'hbc5d2dc3),
	.w4(32'h3b653be2),
	.w5(32'hbba62f2d),
	.w6(32'hbc692dd2),
	.w7(32'hbbcd6e78),
	.w8(32'hbbda06e9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81bf8b),
	.w1(32'hbbb317bc),
	.w2(32'hbbf5f000),
	.w3(32'hbbf346cf),
	.w4(32'hbb256603),
	.w5(32'hbc0ab8d3),
	.w6(32'hbc3fa0f7),
	.w7(32'h3ac79231),
	.w8(32'h3b373129),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25f4a1),
	.w1(32'h3b7cce77),
	.w2(32'h3bba9c03),
	.w3(32'h3a8491fb),
	.w4(32'hba15d445),
	.w5(32'h3ae9b50b),
	.w6(32'h3b3ac388),
	.w7(32'hbbb4ac34),
	.w8(32'h38608443),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2859bc),
	.w1(32'hbbaf4ce8),
	.w2(32'hbc495761),
	.w3(32'h3bc8f38a),
	.w4(32'hba3d79c2),
	.w5(32'hbb809c60),
	.w6(32'h3bf8c1a2),
	.w7(32'h3bdf8fac),
	.w8(32'h3bf8544e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d9145),
	.w1(32'hbc949dd5),
	.w2(32'hbb9d6f6b),
	.w3(32'hbb98632f),
	.w4(32'hbc92886f),
	.w5(32'hbb8bd022),
	.w6(32'h3b461df7),
	.w7(32'hbc0da50e),
	.w8(32'h3b92d33e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2854a9),
	.w1(32'h3aee0eca),
	.w2(32'hbae37344),
	.w3(32'h3ce047a6),
	.w4(32'h3af6cd01),
	.w5(32'h3bb78422),
	.w6(32'h3cbabf06),
	.w7(32'hbb3b3f79),
	.w8(32'hba779df0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae225a8),
	.w1(32'hbc8cf989),
	.w2(32'hbb9f1b93),
	.w3(32'hbabe80d3),
	.w4(32'hbb46ae2a),
	.w5(32'hbb8cd493),
	.w6(32'hb9f2fc2b),
	.w7(32'hbb744104),
	.w8(32'hbc0ebd14),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc700de),
	.w1(32'hbb3a1375),
	.w2(32'hbc0f8cfa),
	.w3(32'hbbf67d17),
	.w4(32'hbb88fe00),
	.w5(32'hbc17dcb0),
	.w6(32'hbb8e88bd),
	.w7(32'h3a9cb7fd),
	.w8(32'hbbeafd89),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27d12b),
	.w1(32'hba7efb13),
	.w2(32'hbc55ffc3),
	.w3(32'hbc706b5c),
	.w4(32'h3ba33d28),
	.w5(32'hbc40d188),
	.w6(32'hbc0cfade),
	.w7(32'h3b7f7f03),
	.w8(32'hbc2f6594),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d551d2),
	.w1(32'hbb0476df),
	.w2(32'hbc911199),
	.w3(32'hbb2f9e4b),
	.w4(32'hbc2cccce),
	.w5(32'hbcd2000e),
	.w6(32'hba9ada88),
	.w7(32'hbbde39d4),
	.w8(32'hbb81ec24),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab9fb6),
	.w1(32'hbbdd8cb8),
	.w2(32'h3b721f6a),
	.w3(32'hbb8fc61c),
	.w4(32'h3b827c3d),
	.w5(32'h3cad64b3),
	.w6(32'hbaf250e5),
	.w7(32'hbaee1b0c),
	.w8(32'h3c9029ca),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947276),
	.w1(32'hbc38d4f1),
	.w2(32'hbba8f0e3),
	.w3(32'h3c0cef4f),
	.w4(32'hbc56fcff),
	.w5(32'hbb9ab566),
	.w6(32'h3afb4189),
	.w7(32'hbc80683c),
	.w8(32'hbb2d800d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebfc34),
	.w1(32'h3b6bc62e),
	.w2(32'hbc255d76),
	.w3(32'h3c6d9880),
	.w4(32'hbb6da857),
	.w5(32'hbbfd7f22),
	.w6(32'h3c05f709),
	.w7(32'h3b75427d),
	.w8(32'hbc37323e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12e05f),
	.w1(32'h3bd4865b),
	.w2(32'h3c2d2ae1),
	.w3(32'hbbf7a707),
	.w4(32'h3a946de2),
	.w5(32'h3c7bb68b),
	.w6(32'h3b0c4c1b),
	.w7(32'hbb37306e),
	.w8(32'h3bb5c405),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba310ae8),
	.w1(32'hbacc122b),
	.w2(32'hbbe96888),
	.w3(32'hba1b98be),
	.w4(32'hbb66c5a3),
	.w5(32'hbbfbbc27),
	.w6(32'hbbe2b3ec),
	.w7(32'hba1ba125),
	.w8(32'h3bf4cb0b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f25de),
	.w1(32'h3bc7775d),
	.w2(32'hbbe4ba9a),
	.w3(32'h3c9f0f3e),
	.w4(32'hbba7595a),
	.w5(32'hbc8f88df),
	.w6(32'h3cd5027b),
	.w7(32'hbbbb65f2),
	.w8(32'hbaeb025c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc299f9b),
	.w1(32'h3c202d0b),
	.w2(32'h3bf3635c),
	.w3(32'h3ab5f483),
	.w4(32'h3c0b4c1a),
	.w5(32'h3c387fc2),
	.w6(32'h3c6aabce),
	.w7(32'h3bf68fc0),
	.w8(32'h3b874206),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc128277),
	.w1(32'h3b47f86c),
	.w2(32'h3b908c9b),
	.w3(32'hbc4e2f63),
	.w4(32'hbb3d35c8),
	.w5(32'h39f970b4),
	.w6(32'hbc099e51),
	.w7(32'hbba04399),
	.w8(32'h3a91e245),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0585e8),
	.w1(32'h3c2e3819),
	.w2(32'h3c31bad8),
	.w3(32'h3c195435),
	.w4(32'h3ac1aca6),
	.w5(32'h3b083181),
	.w6(32'h3af60af7),
	.w7(32'h3bee39b7),
	.w8(32'h3b3bde7f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41e3e4),
	.w1(32'hbbf1d7b5),
	.w2(32'hbc2ed751),
	.w3(32'hba373ae9),
	.w4(32'h3a1d4e9a),
	.w5(32'hbba879e3),
	.w6(32'h3baabe63),
	.w7(32'h3bd83681),
	.w8(32'h3be36fe2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc731142),
	.w1(32'hbbe39e89),
	.w2(32'hbc564608),
	.w3(32'hbc2b98f9),
	.w4(32'hbbca1043),
	.w5(32'hbc527246),
	.w6(32'hba30e432),
	.w7(32'hbb0ddffa),
	.w8(32'hb9c499ec),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc225780),
	.w1(32'hbb8ae0a8),
	.w2(32'h3bb330ea),
	.w3(32'hbbc5152b),
	.w4(32'h3b15e42e),
	.w5(32'h3c4d7572),
	.w6(32'h3b70eda2),
	.w7(32'hbb18a3c4),
	.w8(32'h3ba36812),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a15ce),
	.w1(32'h39b910d5),
	.w2(32'h3b76c745),
	.w3(32'h3b92cedf),
	.w4(32'h3b556309),
	.w5(32'hbb6e78ca),
	.w6(32'hbb0d544d),
	.w7(32'h3b232867),
	.w8(32'h3b3ab622),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d57c3),
	.w1(32'h3a9cdeb2),
	.w2(32'hbacb9dad),
	.w3(32'h3b97cccd),
	.w4(32'h3aa2dd82),
	.w5(32'hba99beaf),
	.w6(32'h3c196e70),
	.w7(32'h3b62076f),
	.w8(32'hbb682a09),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d8193),
	.w1(32'h3c1e9d50),
	.w2(32'h3b7a5640),
	.w3(32'hbc842195),
	.w4(32'h3c074324),
	.w5(32'h3b5c74b3),
	.w6(32'hbc6f9314),
	.w7(32'h3bfb7591),
	.w8(32'h3b2b0552),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aa32e),
	.w1(32'hba842a9b),
	.w2(32'h3aaa3c77),
	.w3(32'hbc41b816),
	.w4(32'hb9820487),
	.w5(32'hbbe54b46),
	.w6(32'hbbed637a),
	.w7(32'hbbaf6474),
	.w8(32'hbb25b143),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bc2af),
	.w1(32'hba651115),
	.w2(32'hbb78124c),
	.w3(32'h3c816ac4),
	.w4(32'hbb61f2be),
	.w5(32'hbc4440e1),
	.w6(32'h3c1a4b98),
	.w7(32'hbb4bf1db),
	.w8(32'hbbd23964),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbf6b2),
	.w1(32'h3a86888a),
	.w2(32'hbba0aa6c),
	.w3(32'h3aaf25c8),
	.w4(32'h3acc0464),
	.w5(32'hbca92444),
	.w6(32'hbb7e4567),
	.w7(32'h3b7eb8cc),
	.w8(32'hbaf9ff33),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba629813),
	.w1(32'hbb3a6c1d),
	.w2(32'hbb17c7e9),
	.w3(32'hba1ed332),
	.w4(32'hbb522af9),
	.w5(32'h3a823dd9),
	.w6(32'hbb91a7e9),
	.w7(32'h3a58e06d),
	.w8(32'hbb0d302e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae72b5f),
	.w1(32'h3c2c2af6),
	.w2(32'h3b545057),
	.w3(32'hbba82ec7),
	.w4(32'h3c1cfa3c),
	.w5(32'hbb84a590),
	.w6(32'hbc3b2f5a),
	.w7(32'h3bd26543),
	.w8(32'hbbdc8e4f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc041f15),
	.w1(32'hbc0a2c74),
	.w2(32'hb7e8288d),
	.w3(32'hbc336eb1),
	.w4(32'hbbb54026),
	.w5(32'hbaccdfe6),
	.w6(32'hbc25ec29),
	.w7(32'hbaf2c0e5),
	.w8(32'h3bcca1ba),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99de31),
	.w1(32'h3a1cc5c9),
	.w2(32'hbbb7b2e2),
	.w3(32'h3b3d3504),
	.w4(32'hb8a72ef6),
	.w5(32'hbc0ac453),
	.w6(32'h3c006b85),
	.w7(32'hba602ed3),
	.w8(32'hbbd354e9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf421ba),
	.w1(32'h3bd0a968),
	.w2(32'h3c45c988),
	.w3(32'hbbb5a67d),
	.w4(32'h3b7146b5),
	.w5(32'h3c20f066),
	.w6(32'hbb137ac5),
	.w7(32'h3b06210c),
	.w8(32'h3c2d971d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816092),
	.w1(32'h395d8894),
	.w2(32'hbb09e0ac),
	.w3(32'h3c24473f),
	.w4(32'hbb7d9cc1),
	.w5(32'hbc173aa1),
	.w6(32'h3bfb0a0b),
	.w7(32'hbc4537c2),
	.w8(32'hbc862bd7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70c555),
	.w1(32'hbb8ab883),
	.w2(32'hbb2d1dcb),
	.w3(32'hbc303a9f),
	.w4(32'hbbd61b97),
	.w5(32'hbbc5fdcf),
	.w6(32'hbc9afba8),
	.w7(32'hbb9e3fa4),
	.w8(32'h3b96c8b6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19e17b),
	.w1(32'hb9e97887),
	.w2(32'hbad62de5),
	.w3(32'h3ca440dc),
	.w4(32'h3ba17418),
	.w5(32'h3b196ffa),
	.w6(32'h3c88d8dd),
	.w7(32'h3b8b6992),
	.w8(32'h38aa333c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae736fa),
	.w1(32'h39f938e3),
	.w2(32'hbacf608b),
	.w3(32'hbc660f77),
	.w4(32'h3b6e7158),
	.w5(32'hbac34b38),
	.w6(32'hbacdc25d),
	.w7(32'h3c102c5c),
	.w8(32'h3ba6e4e4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fa5f7),
	.w1(32'hb8f1b68a),
	.w2(32'hbc2d2244),
	.w3(32'hbb30430c),
	.w4(32'hbaba795d),
	.w5(32'hbbccb3a3),
	.w6(32'h3b31c438),
	.w7(32'hbb0fc831),
	.w8(32'hbb29db46),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b3a53),
	.w1(32'hbb9567a3),
	.w2(32'hba879b8e),
	.w3(32'h3b0e02a2),
	.w4(32'hbb834551),
	.w5(32'hb9974d51),
	.w6(32'hbb5b485f),
	.w7(32'hbb11f20f),
	.w8(32'h37855297),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e71c5),
	.w1(32'h3bf65eed),
	.w2(32'h3b2b5365),
	.w3(32'hbc1bfec8),
	.w4(32'h3b9192ef),
	.w5(32'hbb8dd4a2),
	.w6(32'hbc68a243),
	.w7(32'h3bc12129),
	.w8(32'h3b162134),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a181e10),
	.w1(32'h3ac37077),
	.w2(32'h3ba6ccbe),
	.w3(32'hbb215ae7),
	.w4(32'h3abe4d25),
	.w5(32'h3bf574cf),
	.w6(32'h3b4fd357),
	.w7(32'hba8951c9),
	.w8(32'hbb1dca69),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cce1a),
	.w1(32'h3b9a0a24),
	.w2(32'h3b3d1f07),
	.w3(32'hbb422f16),
	.w4(32'h3be5ec90),
	.w5(32'h3b08236e),
	.w6(32'hbba3b1e9),
	.w7(32'h3a3004f7),
	.w8(32'hbb8bf1c7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dc88b),
	.w1(32'h39dbb700),
	.w2(32'h3bffff75),
	.w3(32'h3b74ee49),
	.w4(32'hbae480cb),
	.w5(32'h3a4f7f9e),
	.w6(32'hbb619e55),
	.w7(32'hbb144d8f),
	.w8(32'hbae0e229),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beac40f),
	.w1(32'h3ba4488d),
	.w2(32'hbb910dce),
	.w3(32'h3c4b1551),
	.w4(32'h3b60bd9f),
	.w5(32'hba96b15a),
	.w6(32'h3bef0b63),
	.w7(32'h3b08c30a),
	.w8(32'hbadb97a6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb22a37),
	.w1(32'hbcb16c39),
	.w2(32'hbc8ee4d1),
	.w3(32'hbc1d7d4e),
	.w4(32'hbc86dbb1),
	.w5(32'hbc67dd3b),
	.w6(32'hbbf8a5ce),
	.w7(32'hbb98b6c8),
	.w8(32'hbc0da721),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64b086),
	.w1(32'h3ae06864),
	.w2(32'h38a817af),
	.w3(32'hbbdd2759),
	.w4(32'h3ad395c6),
	.w5(32'h3a61ed2d),
	.w6(32'hbb9a1161),
	.w7(32'h3a8cf80c),
	.w8(32'h3b539d66),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc4a88),
	.w1(32'hbc65c7dd),
	.w2(32'hbbfc83cf),
	.w3(32'hbaebfe8b),
	.w4(32'hbc641d21),
	.w5(32'hbcc24095),
	.w6(32'hbb7897b2),
	.w7(32'hbc4502b7),
	.w8(32'hbcbf0c6f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87e1f9),
	.w1(32'h3a05c844),
	.w2(32'hbb68b5af),
	.w3(32'h3bca285d),
	.w4(32'hbba22968),
	.w5(32'hbc10ee4c),
	.w6(32'hbc7a74f7),
	.w7(32'h3ad6759c),
	.w8(32'hbb9654f6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85671c),
	.w1(32'h3b97bda4),
	.w2(32'h3aca5863),
	.w3(32'hbba15d9f),
	.w4(32'h3b9cc88a),
	.w5(32'h3a91baec),
	.w6(32'hba464302),
	.w7(32'h3bad8042),
	.w8(32'h3a61c4f1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db1f9),
	.w1(32'hbc5372bf),
	.w2(32'hbb705411),
	.w3(32'hbb03466f),
	.w4(32'hbc4f0da8),
	.w5(32'hbaae60a1),
	.w6(32'hbb2bdfb4),
	.w7(32'hbc20482a),
	.w8(32'h3bcf6344),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b698a6a),
	.w1(32'h3c52da06),
	.w2(32'h3bc2f76b),
	.w3(32'h3c9c6457),
	.w4(32'h3c3d72cf),
	.w5(32'h3bd64f15),
	.w6(32'h3c4cf143),
	.w7(32'hba7472eb),
	.w8(32'hbc0da875),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb142ea2),
	.w1(32'hbb1c04d0),
	.w2(32'hbb7ab3e2),
	.w3(32'hbc39b60d),
	.w4(32'h3a8aa315),
	.w5(32'hbb20f74d),
	.w6(32'hbc3cdf75),
	.w7(32'h3b78692a),
	.w8(32'hbafc13f5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57bee0),
	.w1(32'h3b4a555c),
	.w2(32'h3bc7782f),
	.w3(32'hba8e3c3b),
	.w4(32'h3c11570e),
	.w5(32'h3c1a7131),
	.w6(32'h3a8d1463),
	.w7(32'h3bbf7f68),
	.w8(32'h3bf5bd1b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4fb62),
	.w1(32'hbc2c8c57),
	.w2(32'hbc8c1d85),
	.w3(32'hbaa289c1),
	.w4(32'hbc9c07b8),
	.w5(32'hbc8d87f2),
	.w6(32'hbb43cf91),
	.w7(32'hbc605020),
	.w8(32'hbc9779d4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5ce3d),
	.w1(32'hbb6c9534),
	.w2(32'hbbf2bda3),
	.w3(32'hbc064bd7),
	.w4(32'hbc182632),
	.w5(32'hbb98e610),
	.w6(32'hbc289b64),
	.w7(32'hbb889581),
	.w8(32'hbb6aeae6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16d7e6),
	.w1(32'h3b5a0f9d),
	.w2(32'h3bdbf470),
	.w3(32'h3b19dc50),
	.w4(32'h3b9ebcb7),
	.w5(32'hbc3d9383),
	.w6(32'h3be4c956),
	.w7(32'h3bf97a9c),
	.w8(32'h3ac9461a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a8701),
	.w1(32'hbb2725c6),
	.w2(32'hbb56db69),
	.w3(32'h3c66714b),
	.w4(32'h3b125a00),
	.w5(32'hbab07e59),
	.w6(32'h3bc38594),
	.w7(32'h3a2184ca),
	.w8(32'hbb19581e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f22301),
	.w1(32'hbb061777),
	.w2(32'hbaf0040e),
	.w3(32'hbad9397f),
	.w4(32'hbb0fa33d),
	.w5(32'hba9876e2),
	.w6(32'hbb1a8a6a),
	.w7(32'hbaaca75b),
	.w8(32'hbb0de058),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0c0d9),
	.w1(32'h3a419e9e),
	.w2(32'h3b066d81),
	.w3(32'hba8949a7),
	.w4(32'h3ad316c0),
	.w5(32'h3a93101b),
	.w6(32'hba9b8a37),
	.w7(32'hbb1a580b),
	.w8(32'hbb554ff0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1aaf9e),
	.w1(32'hbb577407),
	.w2(32'hbb592a48),
	.w3(32'hbac5de21),
	.w4(32'hba14b3d8),
	.w5(32'hba83b932),
	.w6(32'hbaa61f12),
	.w7(32'hb943e219),
	.w8(32'h3a478f1f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4380f5),
	.w1(32'h371dea11),
	.w2(32'hb9effe36),
	.w3(32'hbb3dfdf0),
	.w4(32'h39e5e9ac),
	.w5(32'h3a328f14),
	.w6(32'hba6753fd),
	.w7(32'hb99ee6ac),
	.w8(32'hba3d57ef),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88ecf4),
	.w1(32'hba4db792),
	.w2(32'hba6de061),
	.w3(32'h39971983),
	.w4(32'h3a4fd348),
	.w5(32'h39c491a1),
	.w6(32'hba631d65),
	.w7(32'h3b9d06c7),
	.w8(32'h3b4e034c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e283d7),
	.w1(32'h3b7b91fe),
	.w2(32'h3b51010e),
	.w3(32'h3b335239),
	.w4(32'h3ade7af7),
	.w5(32'h3a94aee5),
	.w6(32'h3abf1f0b),
	.w7(32'h39e33953),
	.w8(32'h3945f091),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b182478),
	.w1(32'h3adbfcc4),
	.w2(32'hbb3deb34),
	.w3(32'h3b12ae55),
	.w4(32'h3b001507),
	.w5(32'hbb508a52),
	.w6(32'h3ac11736),
	.w7(32'h3a3f421a),
	.w8(32'hbb538d6d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8399eb),
	.w1(32'hbb17ced8),
	.w2(32'hbb016a79),
	.w3(32'hbb5d86ef),
	.w4(32'hbbb7c42a),
	.w5(32'hbb872304),
	.w6(32'hbaddad94),
	.w7(32'hbb9004bf),
	.w8(32'hbb88b573),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3719b8),
	.w1(32'h3b640220),
	.w2(32'h3a06a5ad),
	.w3(32'h3a887eb4),
	.w4(32'h3b1bbc7a),
	.w5(32'h3a47e3b6),
	.w6(32'hbad1b653),
	.w7(32'h3b313faa),
	.w8(32'h399b27b9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a810895),
	.w1(32'hbb171c28),
	.w2(32'hba1f0a4b),
	.w3(32'h3a932bf9),
	.w4(32'hbac204af),
	.w5(32'hba5ad161),
	.w6(32'h39589d05),
	.w7(32'h3aa20485),
	.w8(32'hbac5c957),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43963f),
	.w1(32'h3b6c3b6d),
	.w2(32'h3b8440b5),
	.w3(32'h3913e1c7),
	.w4(32'h3b87880a),
	.w5(32'h3b5dc73d),
	.w6(32'hbad5faf5),
	.w7(32'h3b4886c6),
	.w8(32'h3b42429e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbafb34),
	.w1(32'hb97acdf6),
	.w2(32'h3a258e4d),
	.w3(32'h3b9f29d3),
	.w4(32'hba58b97c),
	.w5(32'hb9dcd1aa),
	.w6(32'h3bb6fb4c),
	.w7(32'hbafbb877),
	.w8(32'hbad73d42),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8995c1),
	.w1(32'h390d1a9b),
	.w2(32'h3a9e1503),
	.w3(32'hb98c446a),
	.w4(32'h39795bac),
	.w5(32'h3a9618a3),
	.w6(32'h3a7fc994),
	.w7(32'hba291d97),
	.w8(32'h3a9a72d3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7ebd9),
	.w1(32'hb87f44d8),
	.w2(32'hba0989e2),
	.w3(32'h3b2ae4aa),
	.w4(32'h3a313f8b),
	.w5(32'h3b214b8d),
	.w6(32'h3b214140),
	.w7(32'hba646a5a),
	.w8(32'hbaa9b7e4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978e6a4),
	.w1(32'hbb325f03),
	.w2(32'hbb78f140),
	.w3(32'hb8817292),
	.w4(32'hbb57326e),
	.w5(32'hbabeaabe),
	.w6(32'hbb4dbbc4),
	.w7(32'hba9ffdb3),
	.w8(32'hbad21744),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980e4dc),
	.w1(32'h3b51b0a7),
	.w2(32'hba474b6c),
	.w3(32'hb9a45d5f),
	.w4(32'h3b86bf9a),
	.w5(32'h3ba0e857),
	.w6(32'h38e9bd69),
	.w7(32'h3b37673d),
	.w8(32'hba769a56),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f5681),
	.w1(32'hbb36021f),
	.w2(32'h3af005f7),
	.w3(32'h3b4c900e),
	.w4(32'hba01b455),
	.w5(32'h3ab9f8e2),
	.w6(32'h3b59c4bb),
	.w7(32'h3b004b3b),
	.w8(32'h3a96b276),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144c99),
	.w1(32'h36a51a4b),
	.w2(32'hb89738d5),
	.w3(32'hb8c1a6f4),
	.w4(32'hbabdc1e6),
	.w5(32'h3a85b120),
	.w6(32'hbab51323),
	.w7(32'hb8ace251),
	.w8(32'hba874017),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f19d8),
	.w1(32'h3a9d7774),
	.w2(32'h391570da),
	.w3(32'h3a80323f),
	.w4(32'hb9c2b892),
	.w5(32'h3982b33c),
	.w6(32'hbae28682),
	.w7(32'h380537f1),
	.w8(32'h3923b9fc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab7655),
	.w1(32'hba5935f9),
	.w2(32'hbb1d5f1f),
	.w3(32'h3a149dcc),
	.w4(32'hba5b1e2e),
	.w5(32'h38b697c0),
	.w6(32'hbb27e50e),
	.w7(32'hba676352),
	.w8(32'hbaaa69ba),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27fd8a),
	.w1(32'hbbf00f0b),
	.w2(32'hbb3312f4),
	.w3(32'hbb02fef3),
	.w4(32'hbb726b74),
	.w5(32'h3a68a246),
	.w6(32'hbaf535dc),
	.w7(32'hbb9d63eb),
	.w8(32'hbb15ee20),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7a065),
	.w1(32'hbbc641f2),
	.w2(32'hbb952582),
	.w3(32'hbadd1546),
	.w4(32'hbb0794c8),
	.w5(32'h3a9bc8b6),
	.w6(32'hbbc39220),
	.w7(32'hbb2a5ec7),
	.w8(32'h3aaad94f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa08ddf),
	.w1(32'h3b93f28d),
	.w2(32'h3b30a05b),
	.w3(32'hbabbeb39),
	.w4(32'h3b3151a9),
	.w5(32'h3ae07ec0),
	.w6(32'h3a4ac1c8),
	.w7(32'hb6782597),
	.w8(32'h39b7f72e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae73d27),
	.w1(32'h3b90114c),
	.w2(32'h3accc6cb),
	.w3(32'h3adc4c56),
	.w4(32'h3b315b61),
	.w5(32'h3a8c71e9),
	.w6(32'h3b2b1d93),
	.w7(32'hbb1d670a),
	.w8(32'hbaf145fd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a836611),
	.w1(32'hb96b591a),
	.w2(32'hb9a5a785),
	.w3(32'h3a119e75),
	.w4(32'hbb27a313),
	.w5(32'hb9ddcf66),
	.w6(32'h3853fe33),
	.w7(32'h3abe0701),
	.w8(32'hba800bf4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba704e5a),
	.w1(32'h3a6f6ae6),
	.w2(32'h3aadaffa),
	.w3(32'hb9bc3899),
	.w4(32'h3ae8c23d),
	.w5(32'h3aa7862e),
	.w6(32'h3a91276b),
	.w7(32'h3a17a00e),
	.w8(32'hba908df4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ac130),
	.w1(32'hbad95c69),
	.w2(32'hbb1d9362),
	.w3(32'hb85c25f7),
	.w4(32'hbb2b8fcd),
	.w5(32'h39c891cd),
	.w6(32'h3983a160),
	.w7(32'hbb0980a1),
	.w8(32'hbb5b9a3d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06a36e),
	.w1(32'h39fc4f52),
	.w2(32'h39e24e89),
	.w3(32'hbb084aaa),
	.w4(32'h39604294),
	.w5(32'h38a5f591),
	.w6(32'hbac0cb00),
	.w7(32'h3acbd2c2),
	.w8(32'hbaa0c4d4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65a48d),
	.w1(32'hba6afd25),
	.w2(32'hbaef688a),
	.w3(32'h3a10ca77),
	.w4(32'hba504cc6),
	.w5(32'hbaff5ba8),
	.w6(32'h3950e0b2),
	.w7(32'hbb1ce033),
	.w8(32'hbb486a90),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7c7e1),
	.w1(32'hbb3c9c5b),
	.w2(32'hbb3cc08c),
	.w3(32'hbb584002),
	.w4(32'hbb82d32f),
	.w5(32'hbb5b20d4),
	.w6(32'hbbb8343f),
	.w7(32'h3a2eea46),
	.w8(32'h3a2a2e71),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63ed86),
	.w1(32'h398f1c21),
	.w2(32'hba3c64d5),
	.w3(32'hbad6e464),
	.w4(32'hbabfd65c),
	.w5(32'hba3e2d24),
	.w6(32'hbad30d0a),
	.w7(32'hbaadaa10),
	.w8(32'hbb69c0d4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390121de),
	.w1(32'hba990605),
	.w2(32'hbb1320ba),
	.w3(32'hba132ba0),
	.w4(32'hbb4f6722),
	.w5(32'hbb82661c),
	.w6(32'hbb088219),
	.w7(32'hbb01b640),
	.w8(32'hbb34bfc5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedddd8),
	.w1(32'hbc1c6fee),
	.w2(32'hbb9735d9),
	.w3(32'hbb4ebf39),
	.w4(32'hbb864dfd),
	.w5(32'h3aca7afd),
	.w6(32'hbbd3b54b),
	.w7(32'hbb428d85),
	.w8(32'h39557447),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22fab5),
	.w1(32'hbb8a6edf),
	.w2(32'hba2c3574),
	.w3(32'hbb8ac21b),
	.w4(32'hbb4ce303),
	.w5(32'hbb3233cc),
	.w6(32'hbb6ef6ec),
	.w7(32'hb9ac9f90),
	.w8(32'hbaaa232d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df63b8),
	.w1(32'h3b0ef17a),
	.w2(32'h3acc1f31),
	.w3(32'hbb293640),
	.w4(32'h3ab9db86),
	.w5(32'h3b32b8ac),
	.w6(32'hba9f35cf),
	.w7(32'h38d3df16),
	.w8(32'h3a783121),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4b8fd),
	.w1(32'hbb265a91),
	.w2(32'hbadecf6c),
	.w3(32'h3abab353),
	.w4(32'hba5aa230),
	.w5(32'h38ae9ef3),
	.w6(32'hb9bac20d),
	.w7(32'hba5ac863),
	.w8(32'h38c0e537),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3056f7),
	.w1(32'h3ab26a76),
	.w2(32'h3b0bb035),
	.w3(32'hb8d2e407),
	.w4(32'h3a909346),
	.w5(32'h3ac75e72),
	.w6(32'h3a3ab379),
	.w7(32'h3a9f09b5),
	.w8(32'h3b14bdf9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f9577),
	.w1(32'hbaca7f90),
	.w2(32'hbb7dff8f),
	.w3(32'h3b39cf35),
	.w4(32'hba71825b),
	.w5(32'hbb0044dd),
	.w6(32'h3b424196),
	.w7(32'hbaa9743e),
	.w8(32'h3907b56b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0514aa),
	.w1(32'hbaa1caa7),
	.w2(32'hb9602cd9),
	.w3(32'hbb3b0454),
	.w4(32'hbb850f21),
	.w5(32'hbb5bc6be),
	.w6(32'hbaf0ee3d),
	.w7(32'hbb5493a1),
	.w8(32'hbb1b127a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b58378),
	.w1(32'hb80caf60),
	.w2(32'hbaa16d31),
	.w3(32'hba91b540),
	.w4(32'hbb319ed1),
	.w5(32'hbb72ff64),
	.w6(32'hb89d0256),
	.w7(32'hbb2445dc),
	.w8(32'hbb714b78),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c148b),
	.w1(32'h3a8c2a09),
	.w2(32'h3a59c431),
	.w3(32'hba857835),
	.w4(32'h39c29df5),
	.w5(32'hba52e50c),
	.w6(32'hbb689244),
	.w7(32'hb99c90ef),
	.w8(32'hba08d47e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aaf0a),
	.w1(32'hbb04e19a),
	.w2(32'hbabf3ae8),
	.w3(32'h39ba736a),
	.w4(32'hbb2acad0),
	.w5(32'hbb5ba756),
	.w6(32'hba50f495),
	.w7(32'h3aac4cfc),
	.w8(32'hbacae825),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b32a0),
	.w1(32'hbb4205ca),
	.w2(32'hbb117881),
	.w3(32'hbb17691a),
	.w4(32'h3a7a30c5),
	.w5(32'h3a35239e),
	.w6(32'hbb1304d1),
	.w7(32'h3b8b5d8d),
	.w8(32'h3acec25e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba49a3d),
	.w1(32'hbba9dbca),
	.w2(32'hbb8f09a7),
	.w3(32'h39264d5f),
	.w4(32'hbb1ff806),
	.w5(32'h3afc0a7f),
	.w6(32'hba99f347),
	.w7(32'hbb08427e),
	.w8(32'hba9384cd),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e1be88),
	.w1(32'hba489abd),
	.w2(32'hb90ea80b),
	.w3(32'h3a951f45),
	.w4(32'h392251dc),
	.w5(32'h398c003a),
	.w6(32'hbad65987),
	.w7(32'h38ebb2f8),
	.w8(32'hba3b8f7a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f409a),
	.w1(32'hbadb7491),
	.w2(32'h3930eea4),
	.w3(32'h38a43a38),
	.w4(32'hbb374fbf),
	.w5(32'h39386f38),
	.w6(32'hb9522282),
	.w7(32'hbb2bb9fd),
	.w8(32'hba0d6663),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba242a3f),
	.w1(32'hba3d6631),
	.w2(32'hb962dc2d),
	.w3(32'hbad510b6),
	.w4(32'hbadc774c),
	.w5(32'hbacd236c),
	.w6(32'hba3a8428),
	.w7(32'hba11a22e),
	.w8(32'h3a6632af),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393da7ef),
	.w1(32'h3a5caed0),
	.w2(32'hba4d6039),
	.w3(32'h3ad1aedc),
	.w4(32'h3a8c994a),
	.w5(32'hbad0b55e),
	.w6(32'h3ac6afef),
	.w7(32'hbb3f9f8d),
	.w8(32'hbb3058b6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706d61),
	.w1(32'hba64dc7a),
	.w2(32'hba000f49),
	.w3(32'hbb9f2c09),
	.w4(32'hba283e8c),
	.w5(32'h3a895c60),
	.w6(32'hbb3dcc35),
	.w7(32'hba2acd44),
	.w8(32'h3a33dabc),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a958c07),
	.w1(32'hbb3a4fa1),
	.w2(32'hb98d15b4),
	.w3(32'h3a83a42f),
	.w4(32'hba451869),
	.w5(32'hb8df8a61),
	.w6(32'h3a68bc55),
	.w7(32'h3ac8d509),
	.w8(32'h3a04f38b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac638cb),
	.w1(32'h3b02d6dd),
	.w2(32'h3a75cf4b),
	.w3(32'hb9253624),
	.w4(32'h3b27f62a),
	.w5(32'h3b129b21),
	.w6(32'h3a6f56d8),
	.w7(32'h3ae13075),
	.w8(32'h3a60aa41),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e354e),
	.w1(32'hb9aac04b),
	.w2(32'hb9ecfae1),
	.w3(32'hbad3ed66),
	.w4(32'hb8632f21),
	.w5(32'hb5806fa6),
	.w6(32'h39b5ddb1),
	.w7(32'h389adfe3),
	.w8(32'h3b6ad131),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae03ce5),
	.w1(32'h39a1615e),
	.w2(32'h3ac20f31),
	.w3(32'h3a8cae0a),
	.w4(32'hbb1a841d),
	.w5(32'h3a8c1b65),
	.w6(32'h3ae9dfbb),
	.w7(32'hba994e32),
	.w8(32'hba581a9f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a311422),
	.w1(32'h3a07309d),
	.w2(32'hb9f70560),
	.w3(32'h3a0af83b),
	.w4(32'h38e799c7),
	.w5(32'hb9ddaa4b),
	.w6(32'h3a99d2b1),
	.w7(32'h39acf5a6),
	.w8(32'h39eb6698),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa75c8e),
	.w1(32'h3682ac1b),
	.w2(32'h3aa51166),
	.w3(32'h3af4c6ec),
	.w4(32'hbb203855),
	.w5(32'hbab8501d),
	.w6(32'h3b844b48),
	.w7(32'hbb553910),
	.w8(32'hba4400dc),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6c49b),
	.w1(32'hbb37d200),
	.w2(32'hbaba49d7),
	.w3(32'hbaaeecf7),
	.w4(32'hba963cdd),
	.w5(32'hba42f2eb),
	.w6(32'hbb1be5fe),
	.w7(32'hbb3b9bdd),
	.w8(32'hba3c8516),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84e3c46),
	.w1(32'hbbbb9e38),
	.w2(32'hbc17ef8d),
	.w3(32'hba6beb67),
	.w4(32'hbb42b34c),
	.w5(32'hbb3e2366),
	.w6(32'hba89fc10),
	.w7(32'h394159fc),
	.w8(32'h39ba8c2a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46b862),
	.w1(32'h38e95c84),
	.w2(32'hbadfa626),
	.w3(32'hbc17bbef),
	.w4(32'h39470d44),
	.w5(32'h3ae75a6c),
	.w6(32'hbb4b8c6e),
	.w7(32'h3b09a782),
	.w8(32'hb85afd40),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule