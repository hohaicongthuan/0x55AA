module layer_8_featuremap_245(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed54b),
	.w1(32'hbca5e1ea),
	.w2(32'hbcdfdee6),
	.w3(32'h3bb49138),
	.w4(32'hbac3acc5),
	.w5(32'hbc17f8c5),
	.w6(32'hbc355047),
	.w7(32'hbcbcecdc),
	.w8(32'hbc1b45cc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80261e),
	.w1(32'h3b96f8fa),
	.w2(32'h3afdc305),
	.w3(32'hbc54b69c),
	.w4(32'h3b8c7faa),
	.w5(32'h3b34e442),
	.w6(32'h3b87a86a),
	.w7(32'h3b291ed7),
	.w8(32'h3bb4d3ff),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac25e5d),
	.w1(32'h3c53f07c),
	.w2(32'h3c7c007d),
	.w3(32'hba1b0253),
	.w4(32'h3bc913a7),
	.w5(32'h3b2c31d3),
	.w6(32'h3c431835),
	.w7(32'h3c0cd32c),
	.w8(32'h3c6aeac7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb52c07),
	.w1(32'h3b6c8c4c),
	.w2(32'h3bfed00c),
	.w3(32'h3c4edc52),
	.w4(32'hbb4b36fe),
	.w5(32'hb995b2dd),
	.w6(32'h3c6dce22),
	.w7(32'h3c43279d),
	.w8(32'h3c8430e9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb09878),
	.w1(32'hba2619d8),
	.w2(32'hbb209017),
	.w3(32'h3be3d181),
	.w4(32'h3a43e911),
	.w5(32'h3b6d99fe),
	.w6(32'h3a7c5d6b),
	.w7(32'hba9943cc),
	.w8(32'h393f33bb),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae23cf3),
	.w1(32'h3a777320),
	.w2(32'h3bbb1395),
	.w3(32'hbb1f952d),
	.w4(32'h3b43b225),
	.w5(32'hbb1a672b),
	.w6(32'hbab9949b),
	.w7(32'h3c0e0c04),
	.w8(32'h3c49cbaf),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbd368),
	.w1(32'h3bc5da5e),
	.w2(32'h3bfb844a),
	.w3(32'hbc536b69),
	.w4(32'h3b67d021),
	.w5(32'h3bc3b61a),
	.w6(32'h3bec3963),
	.w7(32'h3c33b02a),
	.w8(32'h3bbe9521),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf424ea),
	.w1(32'hbc4b81a2),
	.w2(32'hbc8e4404),
	.w3(32'h3b823707),
	.w4(32'hbb872582),
	.w5(32'hbb32e443),
	.w6(32'hbc7b058c),
	.w7(32'hbc2e00c0),
	.w8(32'h3b929cf3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ad5fd),
	.w1(32'h3bd76c28),
	.w2(32'h3946fcdc),
	.w3(32'hb90f4619),
	.w4(32'h3c47f229),
	.w5(32'h3c1175fc),
	.w6(32'h3bb70a87),
	.w7(32'hbb8a0314),
	.w8(32'hbaecfef6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac21f10),
	.w1(32'h3ba1ba8c),
	.w2(32'hb8c85ff7),
	.w3(32'hbb2c7732),
	.w4(32'h3c3b24e7),
	.w5(32'h3bfd58d7),
	.w6(32'h3b520cb9),
	.w7(32'h3ac39a6d),
	.w8(32'h3b92fa8b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36cf19),
	.w1(32'hbb252b34),
	.w2(32'hbc413054),
	.w3(32'h3bee3641),
	.w4(32'hbba93f90),
	.w5(32'hbc71bf92),
	.w6(32'h3c265a6f),
	.w7(32'h3b92cad8),
	.w8(32'h3bf02e84),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb903a7f),
	.w1(32'hbb16ec5d),
	.w2(32'hbbb0b2da),
	.w3(32'hbb885e54),
	.w4(32'hb96f740e),
	.w5(32'hbb12520c),
	.w6(32'hbbed5e19),
	.w7(32'hbb8801a3),
	.w8(32'hbbc14358),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf24045),
	.w1(32'h3c9c9dc7),
	.w2(32'h3ca9b3ce),
	.w3(32'hbb846b3d),
	.w4(32'h3c5eef3b),
	.w5(32'h3bf4f4a8),
	.w6(32'h3c58a5ac),
	.w7(32'h3be36465),
	.w8(32'h3b823948),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68ebf0),
	.w1(32'h3b338b6a),
	.w2(32'h3c40dceb),
	.w3(32'h3c5fa8d5),
	.w4(32'h3bdcea0d),
	.w5(32'h3c26a013),
	.w6(32'h3b752526),
	.w7(32'h3b76221b),
	.w8(32'h3c05e078),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c531398),
	.w1(32'h3b974337),
	.w2(32'hbb487c1a),
	.w3(32'h3c175aa4),
	.w4(32'h3b1b44bc),
	.w5(32'hbbd88f39),
	.w6(32'h3bd7eb8f),
	.w7(32'h3a78440f),
	.w8(32'hba677e6a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7a3c0),
	.w1(32'h3bbf6b61),
	.w2(32'hbc72bfd8),
	.w3(32'hba2a39e5),
	.w4(32'h3a89918d),
	.w5(32'hbc9932c8),
	.w6(32'h3c64dc2b),
	.w7(32'hbc3c85d7),
	.w8(32'hbccb5e27),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8f455),
	.w1(32'hbb84c493),
	.w2(32'hbc73c48f),
	.w3(32'hbce6824e),
	.w4(32'hbc08c53c),
	.w5(32'hbbc069b7),
	.w6(32'hbb1c09ae),
	.w7(32'hbc251439),
	.w8(32'hbb68d6ae),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39f9d3),
	.w1(32'hbbcea916),
	.w2(32'hbbea8d4f),
	.w3(32'h3b82c238),
	.w4(32'hbcbe5830),
	.w5(32'hbc934d00),
	.w6(32'h3b883bfa),
	.w7(32'h3c35c008),
	.w8(32'hbabd7f00),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb597b),
	.w1(32'hbbd13d3d),
	.w2(32'hbc5e3a44),
	.w3(32'hbca4829c),
	.w4(32'h3b468a6d),
	.w5(32'hbc99dcde),
	.w6(32'h3bad16e3),
	.w7(32'h3baf38de),
	.w8(32'hbb2dce52),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87ab67),
	.w1(32'h3bb7b3d7),
	.w2(32'h3b7bd920),
	.w3(32'hbcc5d479),
	.w4(32'h3bb2c655),
	.w5(32'h3b079eee),
	.w6(32'h3bb951a1),
	.w7(32'h3bc37448),
	.w8(32'h3b6367ef),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a72a8),
	.w1(32'h3c39625f),
	.w2(32'h3be3d673),
	.w3(32'h3b495733),
	.w4(32'h3c887880),
	.w5(32'h3c4b8174),
	.w6(32'h3b83663f),
	.w7(32'h3c3607e2),
	.w8(32'h3c1122cd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45d4b9),
	.w1(32'h3b55b8cf),
	.w2(32'h3bfadcfc),
	.w3(32'h3b5a69d8),
	.w4(32'hba6bb6b8),
	.w5(32'hbc40c7f9),
	.w6(32'hbab821d9),
	.w7(32'h3c1ca2d2),
	.w8(32'h3b9903aa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9272fc),
	.w1(32'hbb277799),
	.w2(32'hbc6df842),
	.w3(32'hbc2ab8b2),
	.w4(32'hbbae786b),
	.w5(32'hbcc4792e),
	.w6(32'hbae7d2a3),
	.w7(32'h3a34e297),
	.w8(32'h3bc00755),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc260860),
	.w1(32'hbb885366),
	.w2(32'h3b20b48d),
	.w3(32'hbc23e28e),
	.w4(32'h3b380ccc),
	.w5(32'hba8c8b3e),
	.w6(32'h3b9487ac),
	.w7(32'h38ec0b3a),
	.w8(32'hbae49ff0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab75a09),
	.w1(32'h3b7befd9),
	.w2(32'h3bf3144c),
	.w3(32'hbb7ce7f9),
	.w4(32'hbbc45bbf),
	.w5(32'hbba24c59),
	.w6(32'h3b90d911),
	.w7(32'h3c0987a4),
	.w8(32'h3c412fc4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6bf37),
	.w1(32'hbca0b9a0),
	.w2(32'hbc2964df),
	.w3(32'hba5a445c),
	.w4(32'hbb2ae9f8),
	.w5(32'hbb699861),
	.w6(32'hbb691552),
	.w7(32'h391676de),
	.w8(32'hbbdf3170),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16cd3a),
	.w1(32'hbb9cc6a6),
	.w2(32'hbbe6d5b3),
	.w3(32'hbbf040b2),
	.w4(32'hbbf5ab2b),
	.w5(32'hbc5689bc),
	.w6(32'h39055c15),
	.w7(32'h3bf8c750),
	.w8(32'h3a0b95ca),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18d218),
	.w1(32'h3b123dcb),
	.w2(32'hbb2c3cd3),
	.w3(32'hbc08e3d7),
	.w4(32'hbab49be2),
	.w5(32'hbb79ca21),
	.w6(32'h3c1b0dad),
	.w7(32'h3c620bcf),
	.w8(32'h3c0e7490),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b573546),
	.w1(32'h3bb5ae3e),
	.w2(32'h3b2ea973),
	.w3(32'hbbeab718),
	.w4(32'h3bbc5906),
	.w5(32'hbb16e790),
	.w6(32'h3c5ac29a),
	.w7(32'h3c32b0e5),
	.w8(32'h3b4754a4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb356e90),
	.w1(32'hba9c3806),
	.w2(32'hbb91dfdb),
	.w3(32'hbb97d03e),
	.w4(32'h3c659b57),
	.w5(32'h3c2e1d8a),
	.w6(32'hbab07144),
	.w7(32'hbb655980),
	.w8(32'h39d2021f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f65cbe),
	.w1(32'hbbc2219c),
	.w2(32'hbbf58a72),
	.w3(32'h3c3aa7c5),
	.w4(32'hbb84bda4),
	.w5(32'hbc0389a7),
	.w6(32'h3b5d20ff),
	.w7(32'hba49e2eb),
	.w8(32'h3c295d1b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bb6e5),
	.w1(32'h3c2fcdf2),
	.w2(32'h3ba30e08),
	.w3(32'hbb5259de),
	.w4(32'h3c5b6c01),
	.w5(32'h39cbac36),
	.w6(32'h3b431c35),
	.w7(32'h3ab68ec4),
	.w8(32'hbb3087a7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a069e),
	.w1(32'hbc1c97d6),
	.w2(32'hbcc10a17),
	.w3(32'h3985aa19),
	.w4(32'hbc36bbfb),
	.w5(32'hbc47d933),
	.w6(32'hbb4b165f),
	.w7(32'hbbc86dcb),
	.w8(32'hbb3abf6b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddc7d1),
	.w1(32'h3bf29f88),
	.w2(32'h3ba4c22e),
	.w3(32'hbc412b6c),
	.w4(32'h3c6a1bb0),
	.w5(32'h3c712853),
	.w6(32'hbba8ac34),
	.w7(32'hbbb74cf4),
	.w8(32'h37f2155c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d140f),
	.w1(32'h3c01640e),
	.w2(32'h3c09e826),
	.w3(32'h3bc40a61),
	.w4(32'h3bc1477d),
	.w5(32'h3bf23401),
	.w6(32'hba46d760),
	.w7(32'h3a51cdd9),
	.w8(32'h3b34b8bf),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b527065),
	.w1(32'hbb9801f7),
	.w2(32'hbb536eb6),
	.w3(32'h3a8ee081),
	.w4(32'hbc1c9619),
	.w5(32'hbb8cadb7),
	.w6(32'h3a2d951f),
	.w7(32'hbc053215),
	.w8(32'hbbfac268),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9a92d),
	.w1(32'h3af1cf63),
	.w2(32'h3bb9c248),
	.w3(32'hbb117801),
	.w4(32'hb9c3eac5),
	.w5(32'h3adea8ad),
	.w6(32'h3a343616),
	.w7(32'h3b84e10d),
	.w8(32'h3b55ba03),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0d8a1),
	.w1(32'h3b7efd4c),
	.w2(32'hbb2d35ee),
	.w3(32'h3b35b042),
	.w4(32'h3b190a8a),
	.w5(32'hb80f5724),
	.w6(32'h3b8c61b0),
	.w7(32'hbb142a27),
	.w8(32'h3ab03bc4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fefc2),
	.w1(32'h3c7624d6),
	.w2(32'h3cbe41d7),
	.w3(32'h3b4eacdb),
	.w4(32'h3c1a5363),
	.w5(32'hba242467),
	.w6(32'h3c66c829),
	.w7(32'h3ce5d85e),
	.w8(32'h3c4ddd0a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26148c),
	.w1(32'hbc060cd0),
	.w2(32'hbc57a2d8),
	.w3(32'hbb68d1ca),
	.w4(32'hbb8ec202),
	.w5(32'hbb498f5c),
	.w6(32'hbb17d8f1),
	.w7(32'hbc11ac1a),
	.w8(32'hbaa44762),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b1fdd),
	.w1(32'hbc1a4207),
	.w2(32'hbbcef975),
	.w3(32'hb9e07e74),
	.w4(32'hbb5f7276),
	.w5(32'hba20f64b),
	.w6(32'hbc5806a7),
	.w7(32'hbc39fd29),
	.w8(32'hbc21c170),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc629aa),
	.w1(32'h3ad193d5),
	.w2(32'hbaef12c4),
	.w3(32'hbab1f3ea),
	.w4(32'hb9c95184),
	.w5(32'hbc08686c),
	.w6(32'h3c19a8e9),
	.w7(32'h3bf04fba),
	.w8(32'h3b8025f8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7701b),
	.w1(32'h3b0d6a90),
	.w2(32'h3b04d878),
	.w3(32'hbbaaa0d4),
	.w4(32'hbb5d4506),
	.w5(32'hbba91949),
	.w6(32'h3bd8ae4a),
	.w7(32'h3c05ef2e),
	.w8(32'h3b43e10b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b4f8c),
	.w1(32'h3a7a76d8),
	.w2(32'h3c76d1ce),
	.w3(32'h3b182924),
	.w4(32'hbbbaa98c),
	.w5(32'hbbb55a09),
	.w6(32'h3c9b9461),
	.w7(32'h3cb6e6f6),
	.w8(32'h3b9d4e2a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b8b1b),
	.w1(32'hbce203ba),
	.w2(32'hbd44720d),
	.w3(32'hbb99a110),
	.w4(32'hbbc93185),
	.w5(32'hbcbbc7a1),
	.w6(32'hbcde7bf2),
	.w7(32'hbd234b62),
	.w8(32'hbca3a06e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb9593),
	.w1(32'hbb948eb8),
	.w2(32'hbbacc22c),
	.w3(32'hbb012529),
	.w4(32'hbba0b9a4),
	.w5(32'hbbf0a617),
	.w6(32'hbb59bb82),
	.w7(32'hbb84368c),
	.w8(32'hba7cba2f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82af3b),
	.w1(32'h3bec48bd),
	.w2(32'hbc327d07),
	.w3(32'hbb0f4caa),
	.w4(32'h3a3285b1),
	.w5(32'hbc89c565),
	.w6(32'h3c063aee),
	.w7(32'h3c1195e5),
	.w8(32'h3b590494),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3670ca),
	.w1(32'hbb17e293),
	.w2(32'hbc1f1db6),
	.w3(32'hbc28ff40),
	.w4(32'hbbcf7d7b),
	.w5(32'hbbe2535c),
	.w6(32'h3b8bb308),
	.w7(32'h3b5ac5e0),
	.w8(32'h3ad5dbb6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae6da8),
	.w1(32'h3ba35260),
	.w2(32'h3b8c28e0),
	.w3(32'hbb0f80f6),
	.w4(32'hbc089844),
	.w5(32'hbc5960b5),
	.w6(32'h3c4a2754),
	.w7(32'h3c64a0bf),
	.w8(32'h3c310f0d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba3029),
	.w1(32'h3c0c4862),
	.w2(32'h3c0f3068),
	.w3(32'hbbe71c84),
	.w4(32'h3b6cb631),
	.w5(32'h3ad4f784),
	.w6(32'h3c6ae66e),
	.w7(32'h3c1f5f83),
	.w8(32'h3c08baf0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3fc3),
	.w1(32'hbc03e6b3),
	.w2(32'hbb1c78a9),
	.w3(32'hbc02d83d),
	.w4(32'hbba73291),
	.w5(32'h3906f05e),
	.w6(32'hbbba415c),
	.w7(32'h3b0cc1a1),
	.w8(32'hbb8db1e3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0325b5),
	.w1(32'h3ad6a54b),
	.w2(32'h3bacb982),
	.w3(32'hbb3cba84),
	.w4(32'hbb21203c),
	.w5(32'hbb323b95),
	.w6(32'h3b9b7e32),
	.w7(32'h3c21554e),
	.w8(32'h3c2a1270),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a105fa1),
	.w1(32'h3b395ec4),
	.w2(32'hbb45de6b),
	.w3(32'hbbc40920),
	.w4(32'hb9102935),
	.w5(32'hbaf336c7),
	.w6(32'h3b8d1dbb),
	.w7(32'hb9392c9f),
	.w8(32'h3b758561),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea5066),
	.w1(32'h3b868f24),
	.w2(32'h3c1d2ad8),
	.w3(32'h3b00d861),
	.w4(32'hb93b4a02),
	.w5(32'hba40ef47),
	.w6(32'hbb77ff7b),
	.w7(32'h3c4a5306),
	.w8(32'h3b1fc8e1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955414),
	.w1(32'h3a1c356d),
	.w2(32'hbc92ef1c),
	.w3(32'hbc0757ba),
	.w4(32'hba97a993),
	.w5(32'hbcaadb20),
	.w6(32'h3bcc70b8),
	.w7(32'hbb1d7221),
	.w8(32'hbc0799b4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3feafd),
	.w1(32'h3bc96cb5),
	.w2(32'h3ba55e20),
	.w3(32'hbc7c7056),
	.w4(32'hbba851d2),
	.w5(32'hbb957628),
	.w6(32'h3c48f642),
	.w7(32'h3bed9257),
	.w8(32'h3c464235),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81914a),
	.w1(32'hbb9e3823),
	.w2(32'hbc4c8491),
	.w3(32'hbb551520),
	.w4(32'hbc013340),
	.w5(32'hbca7ce94),
	.w6(32'h3bb9e572),
	.w7(32'h3b8fb1a6),
	.w8(32'hbb8806ef),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68a0c1),
	.w1(32'hbae9fb7e),
	.w2(32'hba756056),
	.w3(32'hbb8b1d3d),
	.w4(32'hbb610413),
	.w5(32'hbacbc741),
	.w6(32'hbab4736f),
	.w7(32'hba5d0452),
	.w8(32'h3b055445),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b7bfd),
	.w1(32'h3b5d0d26),
	.w2(32'hba7ef22c),
	.w3(32'h3a0de7c4),
	.w4(32'h3ab6f807),
	.w5(32'hb745193a),
	.w6(32'h3b389315),
	.w7(32'h3ba4ca1f),
	.w8(32'h39108d8a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf8616),
	.w1(32'h3b945377),
	.w2(32'h3bae7e14),
	.w3(32'hbb93fea6),
	.w4(32'hbbc5780b),
	.w5(32'hbc3bff8b),
	.w6(32'h3a163a1c),
	.w7(32'h3c4f072f),
	.w8(32'h3c24eaaf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba250ff),
	.w1(32'h3c959214),
	.w2(32'h3ca4dced),
	.w3(32'hbc49f59c),
	.w4(32'h3ab5168b),
	.w5(32'h3b1720b1),
	.w6(32'h3c84737a),
	.w7(32'h3ca77267),
	.w8(32'h3c8e4c34),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80275d),
	.w1(32'hb9d90839),
	.w2(32'hbbbaa027),
	.w3(32'h3ba2c60f),
	.w4(32'h3bcf599d),
	.w5(32'h3ab79021),
	.w6(32'hb9bc5a96),
	.w7(32'hbc21427d),
	.w8(32'hbb39adda),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ad875),
	.w1(32'hbaa1933d),
	.w2(32'h3af4de78),
	.w3(32'hbb89c228),
	.w4(32'h3c0798ca),
	.w5(32'h3c8ea07c),
	.w6(32'hbc7dfb44),
	.w7(32'hbcaaaa86),
	.w8(32'hbc52f65a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c167f50),
	.w1(32'h3a0cc1a6),
	.w2(32'hbb71f9d5),
	.w3(32'h3c7359b5),
	.w4(32'h3a8211c5),
	.w5(32'hbb47b833),
	.w6(32'h3adaa722),
	.w7(32'hba28c0a0),
	.w8(32'hb98a99ec),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba94e),
	.w1(32'h3b20a97d),
	.w2(32'hb83ff3a0),
	.w3(32'hbb3c63bf),
	.w4(32'h3b02f21b),
	.w5(32'hb81f3fd8),
	.w6(32'h3a4c70fe),
	.w7(32'h393f31b5),
	.w8(32'h3b41e2c1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae39ebe),
	.w1(32'hbbbf53c8),
	.w2(32'hba090364),
	.w3(32'h3b2bef18),
	.w4(32'hbc226ea0),
	.w5(32'hbc070702),
	.w6(32'h3b19751e),
	.w7(32'hbbc0a07c),
	.w8(32'hbb0f3207),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4786d0),
	.w1(32'hbc3263cf),
	.w2(32'hbc1e7608),
	.w3(32'h3b8bc54e),
	.w4(32'h39549f4f),
	.w5(32'h3b45154b),
	.w6(32'hbc7cb0bb),
	.w7(32'hbc552e49),
	.w8(32'hbc1aee70),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc429ca9),
	.w1(32'h3be2b33e),
	.w2(32'hbb900a27),
	.w3(32'hbb49f683),
	.w4(32'h3b2d2bed),
	.w5(32'hbbffa74e),
	.w6(32'h3b8853c3),
	.w7(32'h3b42bdd7),
	.w8(32'h3b1829cf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc424d73),
	.w1(32'h3b74a31c),
	.w2(32'h3bb0b69a),
	.w3(32'hbbad7e30),
	.w4(32'hba125ca4),
	.w5(32'h3abe7323),
	.w6(32'h3b705af4),
	.w7(32'h3bad84fc),
	.w8(32'h3c2c4ae4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1159ba),
	.w1(32'h3b5fe9bc),
	.w2(32'h3c497526),
	.w3(32'h3b978ce1),
	.w4(32'h39117ebd),
	.w5(32'hbc4c78b2),
	.w6(32'h3bfb3e17),
	.w7(32'h3cae9d53),
	.w8(32'h3cea1384),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cad4e),
	.w1(32'hbb255f2b),
	.w2(32'hbb2df186),
	.w3(32'hbc2ec996),
	.w4(32'hbac5de27),
	.w5(32'h3a305e61),
	.w6(32'hbbb90f5f),
	.w7(32'hbbeb3da7),
	.w8(32'h3b232ad1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c376e5b),
	.w1(32'hb917d610),
	.w2(32'hbb946ea4),
	.w3(32'h3c406fd8),
	.w4(32'h3bb4844c),
	.w5(32'hbb200e3e),
	.w6(32'hbbe3f7e4),
	.w7(32'h39008cf3),
	.w8(32'h3bcbd9dd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf341c7),
	.w1(32'hbada99f7),
	.w2(32'hbbac7a98),
	.w3(32'h385b4ba9),
	.w4(32'h3c08fde1),
	.w5(32'hbb5ed008),
	.w6(32'hbb185c8b),
	.w7(32'h3adf1849),
	.w8(32'h3bda57c8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199cd4),
	.w1(32'h3b05e138),
	.w2(32'hba1c5947),
	.w3(32'h3b7e6fb5),
	.w4(32'h3b1b1701),
	.w5(32'hbbc21f50),
	.w6(32'h3b3235c3),
	.w7(32'h38611c70),
	.w8(32'h3b539fa3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14113c),
	.w1(32'hba0cb741),
	.w2(32'h3bd0d5d8),
	.w3(32'hba2ef80f),
	.w4(32'hbba1d374),
	.w5(32'hbb9ebf3a),
	.w6(32'h3c23aea3),
	.w7(32'h3c2cf76d),
	.w8(32'h3c2a29d7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba04141),
	.w1(32'hbb8e5c96),
	.w2(32'hba871c2d),
	.w3(32'hba982c2a),
	.w4(32'hbc4a1f53),
	.w5(32'hbcc9a2c7),
	.w6(32'h3bcc7aa4),
	.w7(32'h3cc2154c),
	.w8(32'h3beea23a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaad9e),
	.w1(32'hbb36e17f),
	.w2(32'hb9a2a6f3),
	.w3(32'hbcae99e8),
	.w4(32'hbc09e996),
	.w5(32'hbbb04f78),
	.w6(32'h3bfb66c6),
	.w7(32'h3bf79e49),
	.w8(32'h3af13e29),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0795b8),
	.w1(32'hb965aafd),
	.w2(32'h3b007517),
	.w3(32'hbc196ef7),
	.w4(32'hbbcd7671),
	.w5(32'hbbfba925),
	.w6(32'h3c492ea8),
	.w7(32'h3c96a93f),
	.w8(32'h3b26c7bd),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb835f20),
	.w1(32'hbbbee7f1),
	.w2(32'h3a8632e8),
	.w3(32'hbc1ba663),
	.w4(32'hbc5a464f),
	.w5(32'hbc369d38),
	.w6(32'h3baeec4a),
	.w7(32'h3b8c4fd6),
	.w8(32'h3c52b649),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc243f9),
	.w1(32'h3baa9e8e),
	.w2(32'h3b213e64),
	.w3(32'hbba63cb7),
	.w4(32'hbc02ba7e),
	.w5(32'hb8cdcf46),
	.w6(32'h3c5a256d),
	.w7(32'h3bd81d29),
	.w8(32'hba338c8e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64c518),
	.w1(32'h3c217c57),
	.w2(32'h3bdd9d68),
	.w3(32'hbc1333be),
	.w4(32'h3a5df6e7),
	.w5(32'hbb19bc00),
	.w6(32'h3b78d651),
	.w7(32'h3c4a6251),
	.w8(32'h3c65a3e2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad037f),
	.w1(32'h3c0cefc6),
	.w2(32'h3c825091),
	.w3(32'hbb28db8d),
	.w4(32'h3be7fef7),
	.w5(32'h3c2241b1),
	.w6(32'h3bcc9f1c),
	.w7(32'h3a97bede),
	.w8(32'h3bf0e058),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6752b2),
	.w1(32'hbc78b4b3),
	.w2(32'hbc00b20a),
	.w3(32'h3bfe9dd4),
	.w4(32'hbc2f4247),
	.w5(32'hbbed84f6),
	.w6(32'h3b8b5aa2),
	.w7(32'h3c174118),
	.w8(32'h3adad5e8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a68b7),
	.w1(32'h3c04faa9),
	.w2(32'h3c252ffa),
	.w3(32'hbc58684e),
	.w4(32'h3ae4d4ac),
	.w5(32'hbc29c03a),
	.w6(32'h3b46448b),
	.w7(32'h3bfd74ca),
	.w8(32'h3c4dfd81),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d13ef),
	.w1(32'h3b2f7eee),
	.w2(32'h3b2a7d90),
	.w3(32'hbbe20eb8),
	.w4(32'hb9a92f41),
	.w5(32'hbb926c32),
	.w6(32'h3c87c91b),
	.w7(32'h3bdec9cd),
	.w8(32'h3c39a0b8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2e503),
	.w1(32'h3be1b501),
	.w2(32'h3ad989dd),
	.w3(32'h3bb05e98),
	.w4(32'h3bff27c6),
	.w5(32'hb9b20fb7),
	.w6(32'h3c0507ab),
	.w7(32'h3c3c1ffd),
	.w8(32'h3ba29a13),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4270f3),
	.w1(32'h3afbc2f1),
	.w2(32'hbb84a315),
	.w3(32'hbc334619),
	.w4(32'hb9c1317a),
	.w5(32'hbad13ac1),
	.w6(32'h3beabbcf),
	.w7(32'h3b60cbf5),
	.w8(32'h3b848469),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f2b7d),
	.w1(32'h3c2b7546),
	.w2(32'h3baa9aee),
	.w3(32'hb883d758),
	.w4(32'hbab2ddfb),
	.w5(32'hbc12889d),
	.w6(32'h3bc9e858),
	.w7(32'h3ae6ea78),
	.w8(32'h3ace9eda),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdee2ae),
	.w1(32'h3bb7b227),
	.w2(32'h3a02b793),
	.w3(32'hbb560cea),
	.w4(32'h3aa1b933),
	.w5(32'h3a13843f),
	.w6(32'h3bb7eb72),
	.w7(32'h3b66c1ca),
	.w8(32'h3b949f68),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79e72e),
	.w1(32'h3c657256),
	.w2(32'h3bfcbf5d),
	.w3(32'h3b0ccc94),
	.w4(32'hbb0fed15),
	.w5(32'hbc2aae97),
	.w6(32'h3ba3ca04),
	.w7(32'h3c9097dd),
	.w8(32'h3cb6857d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75e976),
	.w1(32'hbb554187),
	.w2(32'hbb28846a),
	.w3(32'h3ae45db4),
	.w4(32'h3ad58266),
	.w5(32'h3b0c2518),
	.w6(32'h38c2a1b2),
	.w7(32'h3b5a858e),
	.w8(32'h3b6e7886),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eb157),
	.w1(32'hb9f6fe46),
	.w2(32'hbb1c1ae3),
	.w3(32'h3b276279),
	.w4(32'h3c3d2460),
	.w5(32'h3c03faf9),
	.w6(32'hbbebff16),
	.w7(32'hbc31982b),
	.w8(32'hb959e4e8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbd049),
	.w1(32'h3b87d8ac),
	.w2(32'h3bf8bbfb),
	.w3(32'h3b84c77a),
	.w4(32'h3baa4b08),
	.w5(32'h3c07349e),
	.w6(32'hb9d93222),
	.w7(32'h3b1a752a),
	.w8(32'h3b1da586),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5c4ed),
	.w1(32'h3c243353),
	.w2(32'h3bf7b367),
	.w3(32'h3bce21c0),
	.w4(32'h3bb2553c),
	.w5(32'h3ab3637b),
	.w6(32'h3c342cdd),
	.w7(32'h3c518b6f),
	.w8(32'h3c324bb2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b0bd3),
	.w1(32'h3c2240d8),
	.w2(32'hbb5878a4),
	.w3(32'h3aa94e7b),
	.w4(32'h3a12b7db),
	.w5(32'hbc8a743c),
	.w6(32'h3b05392e),
	.w7(32'h3c65bbd3),
	.w8(32'hbbe624e2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9d454),
	.w1(32'hbaba9337),
	.w2(32'hbb30bcbc),
	.w3(32'hbcb3e883),
	.w4(32'h39fbfd21),
	.w5(32'h3b358348),
	.w6(32'h39c16507),
	.w7(32'h3aca8018),
	.w8(32'hbadadb60),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb985763),
	.w1(32'h3a415f39),
	.w2(32'hbc25208b),
	.w3(32'h3b1e9973),
	.w4(32'hbc14f158),
	.w5(32'hbc96fe83),
	.w6(32'h3b8b03d8),
	.w7(32'h3c3f61a8),
	.w8(32'h3c7213ed),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64bac5),
	.w1(32'h3b9f1db3),
	.w2(32'h3c396b1a),
	.w3(32'hbcb2ec7d),
	.w4(32'hba919fe0),
	.w5(32'hbc29c8fd),
	.w6(32'h3bd1c538),
	.w7(32'h3cf32603),
	.w8(32'h3c3bf0aa),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaee81a),
	.w1(32'h3ca14a6d),
	.w2(32'h3cbf69bd),
	.w3(32'hbc8fc196),
	.w4(32'h3aa7789e),
	.w5(32'h3b105786),
	.w6(32'h3ca8771a),
	.w7(32'h3d0196a1),
	.w8(32'h3c78dc11),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c245189),
	.w1(32'hbbb133a0),
	.w2(32'hbc8470a1),
	.w3(32'hbc116135),
	.w4(32'hbc05afe5),
	.w5(32'h3b8b58eb),
	.w6(32'h3bed9a40),
	.w7(32'h3bd7f55e),
	.w8(32'h3c3e5d12),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c7fe6),
	.w1(32'hb97c52c0),
	.w2(32'h3bc83249),
	.w3(32'h3b8a9617),
	.w4(32'h3c5bd4fe),
	.w5(32'h3bf2b968),
	.w6(32'h3b0d9ef4),
	.w7(32'h3bdf2641),
	.w8(32'h3c0780c1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f411b),
	.w1(32'hbcac56ba),
	.w2(32'hbc8175af),
	.w3(32'h3b93fbec),
	.w4(32'h3bfccb08),
	.w5(32'h3aada723),
	.w6(32'hbcf8dab4),
	.w7(32'hbcbca6a5),
	.w8(32'hbbb7d1d6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b709597),
	.w1(32'h3bb08f9d),
	.w2(32'hbb34f5d6),
	.w3(32'h3c3548d0),
	.w4(32'h3c75b8fa),
	.w5(32'h3c2d2555),
	.w6(32'hbc11d594),
	.w7(32'hbbba9d5b),
	.w8(32'h39c0072d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8b80c),
	.w1(32'hbbe1b12e),
	.w2(32'hbc347845),
	.w3(32'h3c3167a7),
	.w4(32'hbbf4e6fe),
	.w5(32'hbbda4457),
	.w6(32'h3c046f04),
	.w7(32'h3c89d672),
	.w8(32'h3c061efa),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44f082),
	.w1(32'h3bbb8e08),
	.w2(32'hbbe7a4c8),
	.w3(32'h3be96953),
	.w4(32'hba8fe883),
	.w5(32'hbc16a00c),
	.w6(32'h3c5715b6),
	.w7(32'h3c253719),
	.w8(32'hbacb7ca0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4ad81),
	.w1(32'h3bf16b76),
	.w2(32'hb855120a),
	.w3(32'hbc2b590e),
	.w4(32'h3a5788c2),
	.w5(32'hbbaed7a2),
	.w6(32'h3be18260),
	.w7(32'h3b353975),
	.w8(32'h3b742b8f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad0f40),
	.w1(32'h3a3b0c36),
	.w2(32'h3ad2a838),
	.w3(32'hb992e3e1),
	.w4(32'hbad80f3c),
	.w5(32'hbba94390),
	.w6(32'h3beb9315),
	.w7(32'h3bf9d795),
	.w8(32'h3bdf4997),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccab82),
	.w1(32'h3b5d2ab8),
	.w2(32'h3b5c1444),
	.w3(32'hbbc2ed03),
	.w4(32'hbb90b5f6),
	.w5(32'hbbd52542),
	.w6(32'h3b673059),
	.w7(32'h3b45d3b2),
	.w8(32'h3bf1110c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b080eae),
	.w1(32'hbb7aa408),
	.w2(32'h3b0a34c9),
	.w3(32'hbbc97a4e),
	.w4(32'h3c2d17ec),
	.w5(32'h3cba6990),
	.w6(32'hbc083f0d),
	.w7(32'hbc3de41b),
	.w8(32'hbbe44b5d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ab5ac),
	.w1(32'h3aa1942b),
	.w2(32'h39a7bece),
	.w3(32'h3c8854ff),
	.w4(32'h3ae0afc7),
	.w5(32'h3b28543c),
	.w6(32'h3b55f781),
	.w7(32'h3aa06bb7),
	.w8(32'h3b7b2d75),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b012e02),
	.w1(32'hba8ab5d4),
	.w2(32'hbb779082),
	.w3(32'h3aca958d),
	.w4(32'h3c6eb37c),
	.w5(32'h3b4991bc),
	.w6(32'hbc05c2eb),
	.w7(32'hbbd11459),
	.w8(32'h3b59f911),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841f63),
	.w1(32'h3b51078a),
	.w2(32'h3bbd697d),
	.w3(32'h3c0f4d2c),
	.w4(32'h3b828637),
	.w5(32'h3bd4953d),
	.w6(32'h3b8b372f),
	.w7(32'h3bb60ee6),
	.w8(32'h3c09ab83),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3df9d),
	.w1(32'h3c87cbf6),
	.w2(32'h3caff34a),
	.w3(32'h3bf44b63),
	.w4(32'h3c6e25b1),
	.w5(32'h3c971622),
	.w6(32'h3c77730d),
	.w7(32'h3cbc21ce),
	.w8(32'h3c374954),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b7f02),
	.w1(32'h3b505c1f),
	.w2(32'hbb83593e),
	.w3(32'h3c9c1047),
	.w4(32'hba7869ec),
	.w5(32'hbbb96adf),
	.w6(32'h3bdf9af3),
	.w7(32'h3b8257b9),
	.w8(32'h3c78fc00),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be84fcf),
	.w1(32'h3b2293b4),
	.w2(32'h3b93eae4),
	.w3(32'h3b2a6df9),
	.w4(32'h3ba494b5),
	.w5(32'h3ba3a858),
	.w6(32'hbaac9424),
	.w7(32'hb89d8771),
	.w8(32'h3b8ca4a4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf81d3b),
	.w1(32'h3b317302),
	.w2(32'h3a2ebb27),
	.w3(32'h3bdaa242),
	.w4(32'h3ae1e290),
	.w5(32'h3a82836f),
	.w6(32'h3b67c1ca),
	.w7(32'h3b205912),
	.w8(32'h3b45df8f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8585e),
	.w1(32'h3b1cf7fb),
	.w2(32'h3b717ab8),
	.w3(32'h3b1364f8),
	.w4(32'h3c00f2be),
	.w5(32'h3bb70e30),
	.w6(32'h3b887100),
	.w7(32'h3bb262f1),
	.w8(32'h3b25efdd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41e5d0),
	.w1(32'h3c630a30),
	.w2(32'h3c597a67),
	.w3(32'h3b8f6c32),
	.w4(32'h3c7c9db3),
	.w5(32'h3c829022),
	.w6(32'h3c3e39cc),
	.w7(32'h3c368099),
	.w8(32'h3c35b193),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ece05),
	.w1(32'h397f38d5),
	.w2(32'h3a443f03),
	.w3(32'h3c06984d),
	.w4(32'hbad770d6),
	.w5(32'h3b8c048f),
	.w6(32'h3c0d7982),
	.w7(32'hba0e72fc),
	.w8(32'h3bebb7bf),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2ee34),
	.w1(32'hba1fcebf),
	.w2(32'hbb416901),
	.w3(32'h3bb7448c),
	.w4(32'hb9cf5b47),
	.w5(32'hbb4b9646),
	.w6(32'h3c001c87),
	.w7(32'h3bc70f04),
	.w8(32'h3b8ce98f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7a7df),
	.w1(32'h3c076a97),
	.w2(32'h3c0a9033),
	.w3(32'hbac2f529),
	.w4(32'hbaae0821),
	.w5(32'h3b39886d),
	.w6(32'h3c39a3cd),
	.w7(32'h3b5b77bf),
	.w8(32'h3bb079ca),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc3da9),
	.w1(32'hbbdfc8a2),
	.w2(32'hbc56573d),
	.w3(32'h3b79aa23),
	.w4(32'hbc1838be),
	.w5(32'hbc67bf42),
	.w6(32'hbbaf3654),
	.w7(32'hbbdfca9c),
	.w8(32'hbb88cd48),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82be07),
	.w1(32'hba376714),
	.w2(32'h3b22f886),
	.w3(32'hbc4661c2),
	.w4(32'h3a949a59),
	.w5(32'h3b83b8d0),
	.w6(32'hbb15d33d),
	.w7(32'hbb098c77),
	.w8(32'hb906c5fe),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989da5d),
	.w1(32'h3c64c6db),
	.w2(32'h3c891bb1),
	.w3(32'h37e0dcef),
	.w4(32'h3c7f54e6),
	.w5(32'h3c716341),
	.w6(32'h3c616584),
	.w7(32'h3c8aae3e),
	.w8(32'h3ba7c9de),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c181386),
	.w1(32'h3c06cb86),
	.w2(32'hbb2f5a38),
	.w3(32'h3c332b81),
	.w4(32'h3c392838),
	.w5(32'h3b8ec867),
	.w6(32'h3b4ef4a8),
	.w7(32'hbab4180f),
	.w8(32'h3c2ccb8f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfa595),
	.w1(32'hbba147b2),
	.w2(32'hbbfb3d1c),
	.w3(32'h3c5a6efe),
	.w4(32'hbc3f114c),
	.w5(32'hbc3d4c6c),
	.w6(32'h3b329cf8),
	.w7(32'h3b04d750),
	.w8(32'h3b7e131c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e13f36),
	.w1(32'h3b923b81),
	.w2(32'hbbd8817b),
	.w3(32'hbb6b2cae),
	.w4(32'h3affcce2),
	.w5(32'hbb9eb464),
	.w6(32'h3b797a0a),
	.w7(32'hba5a3bf5),
	.w8(32'hbb33ef67),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb022ee),
	.w1(32'h3ba0e56b),
	.w2(32'h3bd30982),
	.w3(32'hbbb8f664),
	.w4(32'h3b5d0f00),
	.w5(32'h3c1f2333),
	.w6(32'h3b64b97e),
	.w7(32'h3b0e8721),
	.w8(32'h3c1c3984),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule