module layer_10_featuremap_302(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4aaba),
	.w1(32'hbba007bd),
	.w2(32'h3bad14ba),
	.w3(32'h3b5a0d2e),
	.w4(32'h3ba49b6f),
	.w5(32'hbb126234),
	.w6(32'hbbb041ad),
	.w7(32'h3b575c0e),
	.w8(32'hbb7e147a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9928b6),
	.w1(32'hba777e09),
	.w2(32'hbb4d5852),
	.w3(32'hbb595235),
	.w4(32'hbb079925),
	.w5(32'hbba97b45),
	.w6(32'hba8408bb),
	.w7(32'hbc01db16),
	.w8(32'h3b33c653),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a848d2d),
	.w1(32'hbb931bd4),
	.w2(32'h39d9f138),
	.w3(32'hbba63f18),
	.w4(32'hbc02b460),
	.w5(32'h3b098a78),
	.w6(32'h3b9e16f0),
	.w7(32'h3b1d040b),
	.w8(32'h3ae83561),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e523cb),
	.w1(32'hba9ddabc),
	.w2(32'hba41b428),
	.w3(32'h3ab19b82),
	.w4(32'hbaad80ea),
	.w5(32'hbbcb38c0),
	.w6(32'h3b54c23b),
	.w7(32'hb853c45a),
	.w8(32'hbc3dd086),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db7c0c),
	.w1(32'hbad128c1),
	.w2(32'h3b527f1b),
	.w3(32'hbba6226e),
	.w4(32'hbb9f0824),
	.w5(32'hbaf8b0eb),
	.w6(32'hbb600b19),
	.w7(32'hbb8d4bd3),
	.w8(32'hbad4af1b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a216c55),
	.w1(32'hbb7c457b),
	.w2(32'h39f49555),
	.w3(32'hbb206730),
	.w4(32'hba8c71ef),
	.w5(32'h386ceaec),
	.w6(32'h3a1efcb2),
	.w7(32'hb88d7e31),
	.w8(32'hbaf838b9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1eccc),
	.w1(32'hbadfb7ca),
	.w2(32'hb94adc0a),
	.w3(32'h3a561a8a),
	.w4(32'hba956de6),
	.w5(32'h3b99ffb8),
	.w6(32'h3bfffb33),
	.w7(32'h3a831fcc),
	.w8(32'h3ab19375),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ec0dd),
	.w1(32'hbba974be),
	.w2(32'h3bdf461d),
	.w3(32'h3b064937),
	.w4(32'hb9a0349c),
	.w5(32'h3b37d8cb),
	.w6(32'hba954e42),
	.w7(32'h3b33d2e0),
	.w8(32'h3b182590),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8291ee),
	.w1(32'h3a8967e4),
	.w2(32'h3b4dd06a),
	.w3(32'h3b057b8f),
	.w4(32'h3b808883),
	.w5(32'h3a0ac1ef),
	.w6(32'hbb261d0f),
	.w7(32'h3b92dba6),
	.w8(32'h38b25290),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06c595),
	.w1(32'hbb7487e6),
	.w2(32'hb98cf851),
	.w3(32'h3a220ce7),
	.w4(32'h3a045dc4),
	.w5(32'hbb50ea52),
	.w6(32'hb92733e2),
	.w7(32'h3a97e4b7),
	.w8(32'hbaf5978f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b0839),
	.w1(32'hbb9377c2),
	.w2(32'hba4e6880),
	.w3(32'hbb299fe3),
	.w4(32'hbb80a23d),
	.w5(32'hbaf37693),
	.w6(32'h3b2408fb),
	.w7(32'hb82bf99d),
	.w8(32'hbb30f1a9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6ac65),
	.w1(32'hbb90984c),
	.w2(32'hbbbd2cf7),
	.w3(32'h3b432f05),
	.w4(32'h3a43017a),
	.w5(32'h3b753c7d),
	.w6(32'h3bd487a4),
	.w7(32'hba0114e6),
	.w8(32'hbb85dd2b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f880),
	.w1(32'hbc144def),
	.w2(32'hbb3521c7),
	.w3(32'hbbaa2570),
	.w4(32'h3bb8d6d9),
	.w5(32'h3b7f4629),
	.w6(32'hbbfd362d),
	.w7(32'h3b1153e0),
	.w8(32'hbb2ea42c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ffd66),
	.w1(32'hbb9bdaa8),
	.w2(32'h3abbf221),
	.w3(32'hbaf62d39),
	.w4(32'hbbea21be),
	.w5(32'hbb98b39d),
	.w6(32'h3ab1caad),
	.w7(32'hbb07b7b5),
	.w8(32'hbb37d34e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0554),
	.w1(32'hbb190f4f),
	.w2(32'hbb12655f),
	.w3(32'hba94df9b),
	.w4(32'hbbaee7c7),
	.w5(32'h3bff4c0f),
	.w6(32'hb99bdf8a),
	.w7(32'hbb42e502),
	.w8(32'h3baeddb1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20e41a),
	.w1(32'h3a8babf7),
	.w2(32'h39276240),
	.w3(32'h3b1dc703),
	.w4(32'hbb77bdec),
	.w5(32'h3ab05c94),
	.w6(32'h3c0c388f),
	.w7(32'hb98ce833),
	.w8(32'hba9e7360),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab46409),
	.w1(32'hbb18e4b9),
	.w2(32'h3a8f28b7),
	.w3(32'h3b8d8d41),
	.w4(32'h3b603213),
	.w5(32'h3a05e975),
	.w6(32'h3b903147),
	.w7(32'hba7b15f8),
	.w8(32'h391f0bf7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26afc8),
	.w1(32'h3a49d9ab),
	.w2(32'hbb2cb706),
	.w3(32'h3af282bc),
	.w4(32'h3acdfb18),
	.w5(32'hbad3e71a),
	.w6(32'hbaf39274),
	.w7(32'hbaa621df),
	.w8(32'hbbad0c32),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e91c0),
	.w1(32'h3b09aae0),
	.w2(32'h3a48bc41),
	.w3(32'hb9d59148),
	.w4(32'hbb6ba30e),
	.w5(32'h3bffb918),
	.w6(32'hbb3c0f01),
	.w7(32'hb83b4504),
	.w8(32'hbb0a14be),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba1fd9),
	.w1(32'hbbef506f),
	.w2(32'hbb3bb228),
	.w3(32'h3b99db80),
	.w4(32'h3c0faa3d),
	.w5(32'h3c241da3),
	.w6(32'h3bc82bcd),
	.w7(32'h3c14c4a8),
	.w8(32'h3ae9ade0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ce58a),
	.w1(32'hbbafd452),
	.w2(32'h3a3eb883),
	.w3(32'hb89c73d5),
	.w4(32'hba39742b),
	.w5(32'h39f25e47),
	.w6(32'hba28a928),
	.w7(32'h3b6ab871),
	.w8(32'h3b44fb4c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa00bb),
	.w1(32'h3938eecb),
	.w2(32'hbb0e1130),
	.w3(32'h39729d79),
	.w4(32'h3a0e594f),
	.w5(32'hbb967bbd),
	.w6(32'h3b211922),
	.w7(32'hb9577eaf),
	.w8(32'h3c0ae444),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf473ed),
	.w1(32'hba513048),
	.w2(32'hbace97e0),
	.w3(32'hb9ac1479),
	.w4(32'h3a8fc1f2),
	.w5(32'h3c0e9313),
	.w6(32'h3c3b57d6),
	.w7(32'h3b75fd62),
	.w8(32'hbbdad277),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4bb7d),
	.w1(32'hbb838ed6),
	.w2(32'h3ad90a39),
	.w3(32'hbbbfaf41),
	.w4(32'hbb67281d),
	.w5(32'h3a9ede4d),
	.w6(32'hbc15b864),
	.w7(32'hbab9a646),
	.w8(32'h388d2171),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb145e8),
	.w1(32'h3c1262b0),
	.w2(32'h3c03a975),
	.w3(32'h3c1cadaa),
	.w4(32'h3b3c4f69),
	.w5(32'hba3a1f61),
	.w6(32'h3be7d2c1),
	.w7(32'hb9696075),
	.w8(32'hbb8483b3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7cc30),
	.w1(32'hbbab0632),
	.w2(32'hbb2a3a78),
	.w3(32'h3b926ac2),
	.w4(32'hba9812cb),
	.w5(32'h3aff6e1e),
	.w6(32'h3bd64d2b),
	.w7(32'h3aa31a84),
	.w8(32'h3b70fee4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b824763),
	.w1(32'h3ae29412),
	.w2(32'h3b47b607),
	.w3(32'hbab0a22c),
	.w4(32'h391785f8),
	.w5(32'h3c1fa4a8),
	.w6(32'h3b67346a),
	.w7(32'h3b1f4dc7),
	.w8(32'h3b83f6cc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c357989),
	.w1(32'h3acaadc1),
	.w2(32'h3b3d352b),
	.w3(32'h3bcba219),
	.w4(32'h3c08f5af),
	.w5(32'h3b7fcdd4),
	.w6(32'hba9ea5a0),
	.w7(32'h3c0cc913),
	.w8(32'h39576382),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a2a3f),
	.w1(32'hbb9527a8),
	.w2(32'hbb535ec0),
	.w3(32'hbaf8ef10),
	.w4(32'hbc2ce9bf),
	.w5(32'hbb8d9067),
	.w6(32'h3b932eb2),
	.w7(32'h39b70ccf),
	.w8(32'hbb805c71),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97bc34),
	.w1(32'hbbffbc1c),
	.w2(32'hbba9b679),
	.w3(32'hba987c0e),
	.w4(32'h3b3559b1),
	.w5(32'hbb9caf1d),
	.w6(32'hbbe5e71a),
	.w7(32'hbaf93c55),
	.w8(32'hbbd284d9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f34e),
	.w1(32'h3bf1c8d1),
	.w2(32'h3b5e224e),
	.w3(32'hbc1d8eb5),
	.w4(32'hbb852166),
	.w5(32'hbb586b8a),
	.w6(32'h3baf943b),
	.w7(32'hb9ea4244),
	.w8(32'h3bdd99c3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233ddb),
	.w1(32'hbbaa11a3),
	.w2(32'hbbd83fae),
	.w3(32'h3c0cddd3),
	.w4(32'h3b0974bb),
	.w5(32'hbbbe3b17),
	.w6(32'h3baecd76),
	.w7(32'hbb4b3326),
	.w8(32'hbae657ab),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3b1d8),
	.w1(32'h3c16a0b7),
	.w2(32'h3b8cf91c),
	.w3(32'hb87b4f76),
	.w4(32'hbac4e228),
	.w5(32'h3ba901fd),
	.w6(32'hb81b36ee),
	.w7(32'h3b9eb328),
	.w8(32'hbabb8d9d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c7e44),
	.w1(32'h3a9f5d92),
	.w2(32'hba7b4e61),
	.w3(32'hbae538fd),
	.w4(32'h3b10013a),
	.w5(32'hbb85ea27),
	.w6(32'hbae67683),
	.w7(32'hbb805418),
	.w8(32'hbbedd77f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa4916),
	.w1(32'h3b9f03b3),
	.w2(32'hba3a9a36),
	.w3(32'h3b40fa7a),
	.w4(32'h3c13d801),
	.w5(32'h3b6a508b),
	.w6(32'hbbd1acac),
	.w7(32'hb9831e48),
	.w8(32'hbb0c02bf),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d0d45),
	.w1(32'h3bd786b9),
	.w2(32'h3bf7a543),
	.w3(32'h38fa1c04),
	.w4(32'hbb800a45),
	.w5(32'hbbcbd9ea),
	.w6(32'hbb98ffc8),
	.w7(32'h3a81abce),
	.w8(32'hbb1e99fe),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b379b),
	.w1(32'h3c881d8f),
	.w2(32'h3ba81154),
	.w3(32'hba232ee0),
	.w4(32'hbae46817),
	.w5(32'hba0b33d5),
	.w6(32'h3b287f0f),
	.w7(32'hbb913f4a),
	.w8(32'h3aa1ea2c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a19d3),
	.w1(32'hbb92a8ab),
	.w2(32'h3b4cdbea),
	.w3(32'hbc0a957d),
	.w4(32'h38d43d43),
	.w5(32'hbba15640),
	.w6(32'hbc446ff2),
	.w7(32'hbae2085a),
	.w8(32'hbba05630),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6f6bb),
	.w1(32'h3c67a844),
	.w2(32'h3c0115c9),
	.w3(32'h3a8b0a2b),
	.w4(32'h3a36da56),
	.w5(32'h3b0ab1bc),
	.w6(32'hbb88707e),
	.w7(32'hbbcd8088),
	.w8(32'hbb62f881),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5a41a),
	.w1(32'hbb834963),
	.w2(32'hbb9ec476),
	.w3(32'h3b345742),
	.w4(32'h3afed739),
	.w5(32'hbb33864a),
	.w6(32'hbb80724b),
	.w7(32'hbb0b5824),
	.w8(32'h3b2d89b6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99673ea),
	.w1(32'h3b833066),
	.w2(32'h3894e647),
	.w3(32'h3bae257c),
	.w4(32'h3b9f8453),
	.w5(32'h3a80be46),
	.w6(32'hba8374bc),
	.w7(32'hb9aeaaea),
	.w8(32'h3afaed0b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c8e9e),
	.w1(32'hbba55c2b),
	.w2(32'hbb039fca),
	.w3(32'h3aa4f0cb),
	.w4(32'hba19f1c3),
	.w5(32'h3c0bb4cd),
	.w6(32'h3bfd426d),
	.w7(32'h3aa8e507),
	.w8(32'h3bdae7e7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eb6cc),
	.w1(32'h3b53423b),
	.w2(32'h3a26a8fa),
	.w3(32'h3bb8783d),
	.w4(32'h3bcd854d),
	.w5(32'h394bb6c7),
	.w6(32'hba1a09e8),
	.w7(32'h3c6d0fe8),
	.w8(32'h391bc062),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69b301),
	.w1(32'h3c0f0109),
	.w2(32'h3b959de0),
	.w3(32'h3b0ca6f2),
	.w4(32'h3b62109c),
	.w5(32'hbaf121cc),
	.w6(32'h3c199f22),
	.w7(32'h3a849b69),
	.w8(32'hbb372722),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01b425),
	.w1(32'hbbe343a6),
	.w2(32'hbbcfaa99),
	.w3(32'h3a0ed205),
	.w4(32'hbb71f7ba),
	.w5(32'hba9111fb),
	.w6(32'h3aaabe5e),
	.w7(32'hbb046d91),
	.w8(32'h3ba55acb),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab67c6e),
	.w1(32'hbac98946),
	.w2(32'hba484606),
	.w3(32'hb94ba04c),
	.w4(32'hbb5714b3),
	.w5(32'hb9a632b1),
	.w6(32'h3c9a810d),
	.w7(32'h3bb7c375),
	.w8(32'h3af4ed3c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a143b42),
	.w1(32'hba981121),
	.w2(32'h3988a6cd),
	.w3(32'hbad4bd84),
	.w4(32'hbb744153),
	.w5(32'h3a5b46ef),
	.w6(32'h3b7c9b34),
	.w7(32'h3a12ed0c),
	.w8(32'h3a541803),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b815b),
	.w1(32'h3bbff8ea),
	.w2(32'h3b1c2b18),
	.w3(32'h3b4825f9),
	.w4(32'h3b671be7),
	.w5(32'h3b00da04),
	.w6(32'hbb3ec0bb),
	.w7(32'h38ff8ad3),
	.w8(32'hba072b7d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8f4e1),
	.w1(32'hbacb266c),
	.w2(32'hba1a4b0b),
	.w3(32'hbbd57591),
	.w4(32'h39c6747d),
	.w5(32'hba36b506),
	.w6(32'hbbaca1ad),
	.w7(32'h3a759fb7),
	.w8(32'h3ba8f2c0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc5b13),
	.w1(32'hbac35440),
	.w2(32'hbaabbb3e),
	.w3(32'h3812e69a),
	.w4(32'h3ab9356d),
	.w5(32'h3b12a1f1),
	.w6(32'h3b660451),
	.w7(32'hba8325d1),
	.w8(32'hbb0ac0bc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea526e),
	.w1(32'h3ae80406),
	.w2(32'h3aa82a09),
	.w3(32'h3bc54a4c),
	.w4(32'h3bd06c83),
	.w5(32'h3aa70958),
	.w6(32'hbb039765),
	.w7(32'hbb212247),
	.w8(32'hbbad2653),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39622e),
	.w1(32'hba6a3f47),
	.w2(32'hbb8c59b7),
	.w3(32'h3afe3b92),
	.w4(32'h3b05f1e0),
	.w5(32'h398cf725),
	.w6(32'hbb30f9d7),
	.w7(32'hbb0714d2),
	.w8(32'hba5b7c9a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc8c0c),
	.w1(32'h3a015439),
	.w2(32'h3b432757),
	.w3(32'h3b0cb181),
	.w4(32'hbb247112),
	.w5(32'hbbbb6c49),
	.w6(32'h3b0abeb7),
	.w7(32'hbbd7d9bc),
	.w8(32'hbbbeac91),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0356b),
	.w1(32'h395c5294),
	.w2(32'hbba61fc6),
	.w3(32'hba067136),
	.w4(32'hbb52872f),
	.w5(32'h3ab51799),
	.w6(32'h3ba4f309),
	.w7(32'hbb539a30),
	.w8(32'hbb03c33d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac23150),
	.w1(32'hb9054a88),
	.w2(32'h3b0bdd4a),
	.w3(32'h3b935041),
	.w4(32'h3bd48460),
	.w5(32'hbb03f485),
	.w6(32'h3b80df9b),
	.w7(32'h3b162391),
	.w8(32'h3aaaf8ac),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cf856),
	.w1(32'hbac3d2fd),
	.w2(32'hbb830c11),
	.w3(32'hb9e00bc4),
	.w4(32'hba661ea5),
	.w5(32'hbab76f93),
	.w6(32'h3b1a5e05),
	.w7(32'h3a97e026),
	.w8(32'h3b0a4a56),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64ff44),
	.w1(32'h3c0e9d99),
	.w2(32'h3b87a605),
	.w3(32'h3c0d8147),
	.w4(32'h3c263117),
	.w5(32'h3535ddde),
	.w6(32'hbb2da96a),
	.w7(32'h3b9e888f),
	.w8(32'h3a321ed2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1d08),
	.w1(32'hbb17a719),
	.w2(32'h3ada3b9d),
	.w3(32'h3ad8e76e),
	.w4(32'hbabc3386),
	.w5(32'hb9e01be4),
	.w6(32'h39a9ba03),
	.w7(32'h39f08374),
	.w8(32'hba0d21ff),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50c0c1),
	.w1(32'hbaf02849),
	.w2(32'hba960b2a),
	.w3(32'h3b310a78),
	.w4(32'h3b46b2d7),
	.w5(32'hbb977667),
	.w6(32'h3aafc757),
	.w7(32'h3a514b8a),
	.w8(32'h3aa2b1b9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0d037),
	.w1(32'h3c4cc79e),
	.w2(32'hba1f3b90),
	.w3(32'hba2c6fdf),
	.w4(32'hbb9c296b),
	.w5(32'hbb335cac),
	.w6(32'h3c435667),
	.w7(32'hbb2044fa),
	.w8(32'hbaed0d11),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfae54),
	.w1(32'h3bd38754),
	.w2(32'h3b26c2ab),
	.w3(32'h3b0f5705),
	.w4(32'h3b83b394),
	.w5(32'h3ab0d1b3),
	.w6(32'hbb8d9688),
	.w7(32'hbb8cd871),
	.w8(32'h3ba8b0ec),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa485fd),
	.w1(32'hbb198c65),
	.w2(32'hba6638bc),
	.w3(32'h3b22d0c8),
	.w4(32'hba369347),
	.w5(32'hbae8ab56),
	.w6(32'h3c9a7550),
	.w7(32'h3b8b1879),
	.w8(32'hbc0eaf3b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be109ad),
	.w1(32'h3c14f35a),
	.w2(32'h3bccd010),
	.w3(32'hb88c298c),
	.w4(32'h3a98d0d9),
	.w5(32'hbb25c47c),
	.w6(32'hb7b8d2c8),
	.w7(32'hba49d342),
	.w8(32'hbb90f9c0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91e2a6),
	.w1(32'h3aab7cf3),
	.w2(32'hbadb28af),
	.w3(32'h3b8ac83d),
	.w4(32'h3b307696),
	.w5(32'hbaa3d54f),
	.w6(32'hbbdbd186),
	.w7(32'hbb74f398),
	.w8(32'hba85779f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3367b5),
	.w1(32'h3b7f9f9d),
	.w2(32'h3b0c7c4b),
	.w3(32'h3a8ec1fc),
	.w4(32'h3aea6027),
	.w5(32'hb934b9db),
	.w6(32'hbb8cb106),
	.w7(32'hb974b9c8),
	.w8(32'hba0938ad),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b565c08),
	.w1(32'h3c0f07fc),
	.w2(32'h3c044d7e),
	.w3(32'h3b8c9863),
	.w4(32'h3b94ee82),
	.w5(32'hbb99636e),
	.w6(32'h3c3a249e),
	.w7(32'h39f96b04),
	.w8(32'hba41d0ed),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa67cda),
	.w1(32'hbb90256f),
	.w2(32'h3a3d2567),
	.w3(32'hbb262c76),
	.w4(32'hbbc8fc57),
	.w5(32'hbbd71fe7),
	.w6(32'h3ba45bb1),
	.w7(32'hba54d86c),
	.w8(32'hbb6c2045),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1371a1),
	.w1(32'h3afbda13),
	.w2(32'hbb3e3e25),
	.w3(32'hbb4b0535),
	.w4(32'hbc0fad8c),
	.w5(32'hbbb98c72),
	.w6(32'hbb171913),
	.w7(32'hbba154d9),
	.w8(32'hbb6b40a7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f8394),
	.w1(32'hbb2b436c),
	.w2(32'h3c3d7dbd),
	.w3(32'h3b4bb9b4),
	.w4(32'h3be6450c),
	.w5(32'hb998aef8),
	.w6(32'hbade1e39),
	.w7(32'h3c249065),
	.w8(32'h3baf2eab),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a859),
	.w1(32'h3bb84f83),
	.w2(32'h3bbbaaa5),
	.w3(32'hbae5109f),
	.w4(32'h3b142f61),
	.w5(32'h3a1d909b),
	.w6(32'hb888b8ef),
	.w7(32'h3b9b720f),
	.w8(32'h39fd473a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cca729),
	.w1(32'h3b3aa58d),
	.w2(32'h3ad49124),
	.w3(32'h380f2ab0),
	.w4(32'h3b7cea9a),
	.w5(32'h3af21010),
	.w6(32'hb7be77b7),
	.w7(32'h3b8245a0),
	.w8(32'hbb6d6f74),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcd75b),
	.w1(32'hbbd8a395),
	.w2(32'h3bc5399b),
	.w3(32'h3adc9f67),
	.w4(32'h37b5c4c9),
	.w5(32'h3bb7334f),
	.w6(32'hbb039ca9),
	.w7(32'hbb8fd793),
	.w8(32'hbbd76c50),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c886f),
	.w1(32'h3bd34af0),
	.w2(32'h3ba9b598),
	.w3(32'h3c0939ab),
	.w4(32'h3ba85b9e),
	.w5(32'h3a603663),
	.w6(32'hbbe02b7e),
	.w7(32'hbb9a068f),
	.w8(32'hba35b1a8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9046),
	.w1(32'h3ba04b78),
	.w2(32'h3af5733a),
	.w3(32'h3b34b679),
	.w4(32'h3b2d2572),
	.w5(32'h3ab217a2),
	.w6(32'hbb92899e),
	.w7(32'hbb47a8ff),
	.w8(32'h3b9fbc4e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e6a3),
	.w1(32'hba976015),
	.w2(32'hba678c80),
	.w3(32'hbad9ee36),
	.w4(32'hbb40ae29),
	.w5(32'h3b272531),
	.w6(32'h3b365ddf),
	.w7(32'h3b182f57),
	.w8(32'hba042bd9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38578bd0),
	.w1(32'hbb35753b),
	.w2(32'h388897ed),
	.w3(32'hba7f1808),
	.w4(32'h3b7bd8e2),
	.w5(32'hbb06ab47),
	.w6(32'hbbdaca5d),
	.w7(32'h3adfbe39),
	.w8(32'h3b9bfceb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53062f),
	.w1(32'hb93be6e2),
	.w2(32'h3b46fe0f),
	.w3(32'h3b07c7ec),
	.w4(32'h3b7f29ef),
	.w5(32'hba1a1866),
	.w6(32'h3c2579b0),
	.w7(32'h3b97c7a3),
	.w8(32'hbabe78bf),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133cb5),
	.w1(32'hba8ca636),
	.w2(32'h3a0b26fb),
	.w3(32'h3b3629e6),
	.w4(32'h38aed0e3),
	.w5(32'h3a8d01e8),
	.w6(32'h3b800d71),
	.w7(32'h3a6e565a),
	.w8(32'hba6b3b22),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895d84),
	.w1(32'hbb0f95c0),
	.w2(32'hba50658f),
	.w3(32'h3ad1f4ab),
	.w4(32'hb9e77ef1),
	.w5(32'hbb4d0e6d),
	.w6(32'h3a8618f9),
	.w7(32'hba7eebff),
	.w8(32'hb9fb0a15),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af11de9),
	.w1(32'h3b60e074),
	.w2(32'h3b54cd84),
	.w3(32'h38894567),
	.w4(32'hbaf214a2),
	.w5(32'h3ba4be50),
	.w6(32'h3ba70ef6),
	.w7(32'hbadd4f77),
	.w8(32'hb83fa4d5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38b96e),
	.w1(32'hbb920002),
	.w2(32'hbb075b5d),
	.w3(32'h3ab2934e),
	.w4(32'h3b8054c6),
	.w5(32'h3bca17e5),
	.w6(32'hbbe1c693),
	.w7(32'h3af1a3d1),
	.w8(32'h3b2c32ab),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c0a30),
	.w1(32'h3bb92921),
	.w2(32'h3b2576fb),
	.w3(32'h3b9060e4),
	.w4(32'h3ac7ac1d),
	.w5(32'hbbb1f029),
	.w6(32'h3b054511),
	.w7(32'h3b7c7c43),
	.w8(32'h3c33cc0a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad67b17),
	.w1(32'hbbbedfb0),
	.w2(32'h3b728022),
	.w3(32'hbaa9edce),
	.w4(32'h3b073e04),
	.w5(32'hbba7ba7e),
	.w6(32'h3c121a17),
	.w7(32'h3bc71a61),
	.w8(32'h3a99d6d0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2d3a5),
	.w1(32'h38f8c068),
	.w2(32'hbb40e731),
	.w3(32'hba3ce501),
	.w4(32'hbc0a6264),
	.w5(32'hbb680394),
	.w6(32'h3aafcf1f),
	.w7(32'hbbbbad46),
	.w8(32'h3c4df508),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba725523),
	.w1(32'hbb7e212a),
	.w2(32'hba3569d0),
	.w3(32'hbbb6c567),
	.w4(32'h3890855d),
	.w5(32'hbbbedb39),
	.w6(32'h3c8823dd),
	.w7(32'h3bfe2c32),
	.w8(32'hbb3b24b8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdf655),
	.w1(32'h3a3edfbc),
	.w2(32'hba23a32a),
	.w3(32'hbb9dc941),
	.w4(32'hbb99506f),
	.w5(32'h3b429878),
	.w6(32'h3c9eb6e6),
	.w7(32'h3c0147ff),
	.w8(32'hb9855154),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d7dd8),
	.w1(32'hbb8f5bc4),
	.w2(32'h3a654546),
	.w3(32'h3990da89),
	.w4(32'hbbb01ca8),
	.w5(32'h3bcc285b),
	.w6(32'h3b68493b),
	.w7(32'hbaaabcd7),
	.w8(32'h3b2ecf98),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e0685),
	.w1(32'hbbaeee2e),
	.w2(32'hbbdc989e),
	.w3(32'h3b82dd27),
	.w4(32'h3b70de87),
	.w5(32'h392a29d8),
	.w6(32'h3c35de56),
	.w7(32'h3bc53861),
	.w8(32'h3b33ddb5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b359edd),
	.w1(32'h3b2a9f1a),
	.w2(32'h3b1355ff),
	.w3(32'h3ae948da),
	.w4(32'h3af7d3d3),
	.w5(32'hbbf1639e),
	.w6(32'h3bbdcf66),
	.w7(32'h3a7385d1),
	.w8(32'hbb0151fe),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86744a),
	.w1(32'hbc464b61),
	.w2(32'hbc008a69),
	.w3(32'hb9664d09),
	.w4(32'hba931dcd),
	.w5(32'h3b58e954),
	.w6(32'hbc448c44),
	.w7(32'hbb965ab0),
	.w8(32'hbc0466c6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae126ae),
	.w1(32'hbb1cf31b),
	.w2(32'hbb7f2ba0),
	.w3(32'hbbdeb6ff),
	.w4(32'h3bf86d83),
	.w5(32'hbb20e31c),
	.w6(32'hbb62ac6d),
	.w7(32'hbb3bd538),
	.w8(32'hbaf59f7b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d4016),
	.w1(32'hbbf021ea),
	.w2(32'hbb8dfc46),
	.w3(32'h3b09df88),
	.w4(32'hbb148704),
	.w5(32'hbab5b366),
	.w6(32'hbbc9113f),
	.w7(32'hbb9295d0),
	.w8(32'h3b32b575),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2bfce),
	.w1(32'h3b87d1c8),
	.w2(32'h3b52085a),
	.w3(32'h394b7346),
	.w4(32'h3afa334a),
	.w5(32'hbac88dc6),
	.w6(32'h3c1e49f5),
	.w7(32'h399ecc5e),
	.w8(32'hbb63ec48),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84803d),
	.w1(32'hbb508436),
	.w2(32'hbb999d7f),
	.w3(32'h3918d0fb),
	.w4(32'hbbc8f5d2),
	.w5(32'h3b940e40),
	.w6(32'hbb44f5e7),
	.w7(32'hbbd417f1),
	.w8(32'h3bb657c9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0166d6),
	.w1(32'hbafa6092),
	.w2(32'h3bbff61d),
	.w3(32'hb9e9ba2f),
	.w4(32'h3bbad7ed),
	.w5(32'hbb794973),
	.w6(32'hbc2786be),
	.w7(32'hba37ec7b),
	.w8(32'h3ac6ac92),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a7826),
	.w1(32'hbc0668bf),
	.w2(32'hbbb3f570),
	.w3(32'hb9b5baa7),
	.w4(32'hba57fb74),
	.w5(32'h3ab62c26),
	.w6(32'hbb7e444f),
	.w7(32'h3ba9166a),
	.w8(32'hba6362c3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d1b9b),
	.w1(32'h398047ea),
	.w2(32'hbbc95bbc),
	.w3(32'h3ba400c3),
	.w4(32'h3b3f7847),
	.w5(32'hbb848054),
	.w6(32'h3abb5150),
	.w7(32'hbb0d1ec2),
	.w8(32'h3a2bbc06),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17c826),
	.w1(32'h3a43a6ab),
	.w2(32'hbb151da6),
	.w3(32'h3a516ea7),
	.w4(32'h3bf90449),
	.w5(32'hbb1fa3ff),
	.w6(32'hbb8fc260),
	.w7(32'hbb463dd2),
	.w8(32'hbb96b9f6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb93b0f),
	.w1(32'h3a08eae6),
	.w2(32'hba08c47f),
	.w3(32'h3af40b2a),
	.w4(32'hba47aa26),
	.w5(32'hbc14ac59),
	.w6(32'h3b0bc5cf),
	.w7(32'hbad713b9),
	.w8(32'h3ad9c26d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba00641),
	.w1(32'h3aec5647),
	.w2(32'hbb55d3f8),
	.w3(32'h3b598291),
	.w4(32'hbb4a4c0a),
	.w5(32'hbc035d0f),
	.w6(32'h3c4c8034),
	.w7(32'hbbb1d95e),
	.w8(32'hbc2d413c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0feb65),
	.w1(32'h39a43ceb),
	.w2(32'hba9c4c58),
	.w3(32'hbc0819b4),
	.w4(32'hbba88712),
	.w5(32'hba026d9e),
	.w6(32'hbbdf2f8f),
	.w7(32'hbace642f),
	.w8(32'hbba0cdc6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6651e7),
	.w1(32'hbc0804e5),
	.w2(32'h3a2da5ec),
	.w3(32'hbafbef85),
	.w4(32'hbc07964b),
	.w5(32'hbb2fad44),
	.w6(32'h3c3e9f68),
	.w7(32'hbb746667),
	.w8(32'hbbef8352),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11e7fe),
	.w1(32'hbc08f514),
	.w2(32'h3c55ccf5),
	.w3(32'hbc102df6),
	.w4(32'hba8ab13b),
	.w5(32'hbb6a80f2),
	.w6(32'h396ff60e),
	.w7(32'hbbe23ddf),
	.w8(32'hbb38ec08),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02aa8d),
	.w1(32'h3bbfee21),
	.w2(32'h39e4b63f),
	.w3(32'hbb9902d5),
	.w4(32'hbb9694d6),
	.w5(32'hbadd6099),
	.w6(32'h3b6d036b),
	.w7(32'hbbb0618f),
	.w8(32'hbb28ca24),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37adb8),
	.w1(32'hbb4acc29),
	.w2(32'hbb5756a6),
	.w3(32'h3a9d5fc7),
	.w4(32'hbb382b7d),
	.w5(32'h3b23fbd8),
	.w6(32'hbbb55045),
	.w7(32'h3b847ed6),
	.w8(32'h3adae438),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3da0a9),
	.w1(32'h3b90869b),
	.w2(32'hba7a1f8c),
	.w3(32'h3b35383e),
	.w4(32'hbb1404ec),
	.w5(32'hbb1e621e),
	.w6(32'h3ace7da2),
	.w7(32'hbb084925),
	.w8(32'hbbed4b24),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e3fb6),
	.w1(32'hbad521cd),
	.w2(32'h3b594a39),
	.w3(32'h3bf9ddf7),
	.w4(32'h3bc3d841),
	.w5(32'hbb119887),
	.w6(32'h3be60046),
	.w7(32'h3ab49be2),
	.w8(32'h3a52d197),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3260a6),
	.w1(32'hbafe1646),
	.w2(32'hba5b8ad0),
	.w3(32'h3b586467),
	.w4(32'hbb6a4202),
	.w5(32'hbb3847ac),
	.w6(32'h3bbee0ad),
	.w7(32'hba934db5),
	.w8(32'hbc2e21a6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc285b28),
	.w1(32'h3ab54fcb),
	.w2(32'hbb04aec3),
	.w3(32'h3b96b65e),
	.w4(32'h3a6d6f4a),
	.w5(32'hba1e5182),
	.w6(32'h3a6a4ee9),
	.w7(32'h39ca42a6),
	.w8(32'hbb574ecc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66170b),
	.w1(32'hba2ead25),
	.w2(32'hbb71a99e),
	.w3(32'hbb11c3ec),
	.w4(32'hbb7dda38),
	.w5(32'h3abb53eb),
	.w6(32'h3974df7e),
	.w7(32'hbb52ff71),
	.w8(32'hbb0d8d50),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eb809),
	.w1(32'hbaf54914),
	.w2(32'h3a90137b),
	.w3(32'h3a26c993),
	.w4(32'hbad80cd5),
	.w5(32'h3a391b81),
	.w6(32'hbbd6acc2),
	.w7(32'hbb10703d),
	.w8(32'h3bcf171b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07472c),
	.w1(32'h3b1de2f8),
	.w2(32'hbb8724c7),
	.w3(32'h3d02d2a0),
	.w4(32'h3c35d4bc),
	.w5(32'hbad5a3bf),
	.w6(32'h3cc4614f),
	.w7(32'h3a1319cc),
	.w8(32'hbaffad10),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07845f),
	.w1(32'hb9e4d2a7),
	.w2(32'h3b20da63),
	.w3(32'hbb8c9cf1),
	.w4(32'hba91d5ed),
	.w5(32'h3c926e1d),
	.w6(32'hba6f547b),
	.w7(32'hba4f50cf),
	.w8(32'hbbe16551),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd95997),
	.w1(32'hbc9283f2),
	.w2(32'h3aca3ca2),
	.w3(32'h3b9f3667),
	.w4(32'h3bef3a61),
	.w5(32'hba2f5fb0),
	.w6(32'h3c2608fc),
	.w7(32'hbb867b68),
	.w8(32'h3a083dd4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74d023),
	.w1(32'hb922fd22),
	.w2(32'h3b6fe2e9),
	.w3(32'hbb5ac64e),
	.w4(32'h3aae3a38),
	.w5(32'hbc3ecdea),
	.w6(32'hb9c840e3),
	.w7(32'hbab80f66),
	.w8(32'h3c0a9c30),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0379b0),
	.w1(32'hbba133e6),
	.w2(32'hbca8436a),
	.w3(32'h3c098420),
	.w4(32'h3a64cb82),
	.w5(32'hbb92dea0),
	.w6(32'h3d1ad5d3),
	.w7(32'hbb47ff6b),
	.w8(32'hba20f876),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52edbc),
	.w1(32'h3b26b219),
	.w2(32'h3aa5cbb4),
	.w3(32'hbbb37d4c),
	.w4(32'hbb8f507d),
	.w5(32'hbbe198ce),
	.w6(32'h37faea14),
	.w7(32'hba76311e),
	.w8(32'hbb2361a0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03d08d),
	.w1(32'hbac895a6),
	.w2(32'h39ec8bfe),
	.w3(32'h3b93273a),
	.w4(32'h3a9e0dd2),
	.w5(32'hb8fdc87b),
	.w6(32'hba6fc579),
	.w7(32'hbb5fd2e4),
	.w8(32'h3bbea05c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a77f0),
	.w1(32'hbb947e44),
	.w2(32'hbb3d80d9),
	.w3(32'h3b41abb6),
	.w4(32'hbb2c7c72),
	.w5(32'h3a9154c6),
	.w6(32'h3ba807df),
	.w7(32'hba437a91),
	.w8(32'hbb26bfca),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18a3ee),
	.w1(32'hbb81fc91),
	.w2(32'hbadb9256),
	.w3(32'h3b117ad0),
	.w4(32'h393631eb),
	.w5(32'h3b93cc5f),
	.w6(32'h3b8ce20c),
	.w7(32'hba9f31b1),
	.w8(32'h3c9ad21e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7af5c1),
	.w1(32'h3cd28b17),
	.w2(32'h3d0a608f),
	.w3(32'h3caf69d3),
	.w4(32'h3c8a7250),
	.w5(32'hbb4f85a8),
	.w6(32'hbad92091),
	.w7(32'h3cff49aa),
	.w8(32'hbac23590),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c6ade),
	.w1(32'h3b8e5bf9),
	.w2(32'hbabf9121),
	.w3(32'hbbb231ff),
	.w4(32'hbb8c5375),
	.w5(32'hbb1d1eda),
	.w6(32'h3b40121b),
	.w7(32'hba023de9),
	.w8(32'h3adee596),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3386e5),
	.w1(32'hba8e9b7b),
	.w2(32'hbb75489b),
	.w3(32'hb943289e),
	.w4(32'h39e48a8c),
	.w5(32'hbc3f31e6),
	.w6(32'hb9fc069c),
	.w7(32'hbc074a3c),
	.w8(32'hbbcd0cea),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae497fe),
	.w1(32'hbafe7219),
	.w2(32'hba4fb5eb),
	.w3(32'hbbff091c),
	.w4(32'hb8ef34fa),
	.w5(32'hbae3ba0d),
	.w6(32'h3b114d38),
	.w7(32'h3b9e024b),
	.w8(32'h3ab2e339),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936a72d),
	.w1(32'hbb07eb6c),
	.w2(32'hbc008dba),
	.w3(32'hbc007dd6),
	.w4(32'hbb9d0934),
	.w5(32'hba8bb860),
	.w6(32'h3be3ddfd),
	.w7(32'hbae245a0),
	.w8(32'hbcb4e45e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cda78),
	.w1(32'hbc827477),
	.w2(32'h3ad7cbe1),
	.w3(32'hbbd4a167),
	.w4(32'h3af30117),
	.w5(32'hbb44cde2),
	.w6(32'hbc591a2f),
	.w7(32'hbb9725b9),
	.w8(32'hba03361e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76252b1),
	.w1(32'hbb3ffa9a),
	.w2(32'hbba134af),
	.w3(32'hb9b08544),
	.w4(32'hba7caf3c),
	.w5(32'h3c59547a),
	.w6(32'h3aa2cf50),
	.w7(32'hbaca67ca),
	.w8(32'hbb4cc0cf),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4016e7),
	.w1(32'hbc32509e),
	.w2(32'hbab36ff8),
	.w3(32'h3bab511f),
	.w4(32'h3894b471),
	.w5(32'h3b70d7aa),
	.w6(32'hbc21ba17),
	.w7(32'hbb94b008),
	.w8(32'h3b7bcae7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e738f),
	.w1(32'hbbf6ab01),
	.w2(32'hbc0bd74d),
	.w3(32'hbb8c75c8),
	.w4(32'hbb8ef11a),
	.w5(32'hbb3afff7),
	.w6(32'hbb349889),
	.w7(32'hbc0436f7),
	.w8(32'h3aca042b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bbd92),
	.w1(32'hbb86fb3d),
	.w2(32'h3ac55fee),
	.w3(32'h3a2afc6a),
	.w4(32'hba6caa64),
	.w5(32'hbb1a57e5),
	.w6(32'h3aaac984),
	.w7(32'hbaf1c999),
	.w8(32'h3b81527d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bd34e),
	.w1(32'hbbb308fd),
	.w2(32'hbba88170),
	.w3(32'hbb4fc97b),
	.w4(32'hbb6e34d6),
	.w5(32'h3a3c3137),
	.w6(32'h3ce1f94b),
	.w7(32'h38d0ac77),
	.w8(32'h3a55d607),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6df261),
	.w1(32'hbb1666f5),
	.w2(32'h3a896c38),
	.w3(32'hbb0128da),
	.w4(32'h3866f04d),
	.w5(32'hbb142330),
	.w6(32'h3ad33e5e),
	.w7(32'hba9d3233),
	.w8(32'hbb5725f6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b5031),
	.w1(32'hbc611f94),
	.w2(32'hbc078f8b),
	.w3(32'hbbf8c204),
	.w4(32'h3ba277f1),
	.w5(32'h3b753dbc),
	.w6(32'h3b848bca),
	.w7(32'h3afed2e0),
	.w8(32'h3a850771),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a3b72),
	.w1(32'hbad29398),
	.w2(32'hb9ff73ba),
	.w3(32'h3b62a913),
	.w4(32'hba8309fe),
	.w5(32'hb9882828),
	.w6(32'h3b8503bd),
	.w7(32'h3a30707f),
	.w8(32'h3a70756d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82da90),
	.w1(32'hba57bb52),
	.w2(32'hbb08beab),
	.w3(32'hbaa6a885),
	.w4(32'hbb3254c1),
	.w5(32'h379b9289),
	.w6(32'h3b7105e5),
	.w7(32'hbb0db726),
	.w8(32'h3b005e13),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e51af),
	.w1(32'hbba605ad),
	.w2(32'hbab33148),
	.w3(32'hbb13f7c9),
	.w4(32'hbbf08775),
	.w5(32'hb9c73d86),
	.w6(32'hbbbc51f4),
	.w7(32'hbb7174d6),
	.w8(32'hba56ceeb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa20bc8),
	.w1(32'hbaef4f5d),
	.w2(32'h3ab0a3dd),
	.w3(32'hbb039e1f),
	.w4(32'hbb654bb3),
	.w5(32'h391d17da),
	.w6(32'hbacfb206),
	.w7(32'hbb0f9565),
	.w8(32'h3b09efec),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31bbf3),
	.w1(32'hbb031e22),
	.w2(32'hbb306895),
	.w3(32'h3ab991a4),
	.w4(32'hbb430215),
	.w5(32'h3aeda871),
	.w6(32'h3b91e64b),
	.w7(32'h38c91ffc),
	.w8(32'h3b655d98),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b36a3),
	.w1(32'h3a3a51ef),
	.w2(32'hba0563f5),
	.w3(32'hbb80cdb0),
	.w4(32'hbbc2bb1f),
	.w5(32'hbb7e1a33),
	.w6(32'h3c41e14b),
	.w7(32'h3add2186),
	.w8(32'hbab56d4b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17e5f1),
	.w1(32'h3c25a2f2),
	.w2(32'hbada4465),
	.w3(32'hbc216896),
	.w4(32'hbb7eb454),
	.w5(32'hba0bbf14),
	.w6(32'h3c47ee03),
	.w7(32'h3af78e66),
	.w8(32'hbb90617c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b361c84),
	.w1(32'h3b5d30b3),
	.w2(32'h3af91f49),
	.w3(32'hbb5cdd77),
	.w4(32'hba7146de),
	.w5(32'h3c7cc320),
	.w6(32'hbc231778),
	.w7(32'hbb86065f),
	.w8(32'hbb2166df),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f42586),
	.w1(32'hbbcd7ab9),
	.w2(32'hbc02c4b2),
	.w3(32'h3ca1395e),
	.w4(32'h3c24bd20),
	.w5(32'h3b922e5f),
	.w6(32'h3b7a3d49),
	.w7(32'hbc0ea6f9),
	.w8(32'hbb18833e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25def3),
	.w1(32'h3b8d0b77),
	.w2(32'h3bf11e0a),
	.w3(32'h3ac7a5fb),
	.w4(32'h3b5e19b6),
	.w5(32'hbb32f1b7),
	.w6(32'hbadde42c),
	.w7(32'h3b846b8c),
	.w8(32'hbb6ff658),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb379c4f),
	.w1(32'hba8def09),
	.w2(32'hbb6d3df3),
	.w3(32'hbaf80386),
	.w4(32'h39b5e7b8),
	.w5(32'h3811fa32),
	.w6(32'h3a7fd1a2),
	.w7(32'hbbcfb35c),
	.w8(32'hbb506862),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb618911),
	.w1(32'h3a59ef3b),
	.w2(32'h3bc6666f),
	.w3(32'hba444098),
	.w4(32'hbb9492f6),
	.w5(32'hbb864712),
	.w6(32'hba453a1b),
	.w7(32'hb9349ca4),
	.w8(32'h3b192477),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2a34b),
	.w1(32'h390781aa),
	.w2(32'hbad5365f),
	.w3(32'hbb47f098),
	.w4(32'h3946eedd),
	.w5(32'hbb00dab7),
	.w6(32'h3a4fdcaa),
	.w7(32'h3a95eae1),
	.w8(32'h3b32b854),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b610373),
	.w1(32'hbb880599),
	.w2(32'hbbc4f170),
	.w3(32'hb9bba0a5),
	.w4(32'hb8de16cb),
	.w5(32'hbbf891c6),
	.w6(32'hb76ab9a5),
	.w7(32'hbb727b99),
	.w8(32'hbca63b74),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc894901),
	.w1(32'hbc02e1bb),
	.w2(32'hbc57901f),
	.w3(32'hbb9d7939),
	.w4(32'hbc27c971),
	.w5(32'hbb849c22),
	.w6(32'hbc522fc1),
	.w7(32'hbc239344),
	.w8(32'hbb16b621),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f244),
	.w1(32'h3a05b6e5),
	.w2(32'hbbc8e2c9),
	.w3(32'hbb920135),
	.w4(32'hbb1ceae6),
	.w5(32'h3a9453f4),
	.w6(32'h3926fc69),
	.w7(32'hbb67592a),
	.w8(32'hbb6a4865),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac61c9f),
	.w1(32'h3a8c09a5),
	.w2(32'h3b8ad90a),
	.w3(32'hbb7d86b2),
	.w4(32'h3a84f4f8),
	.w5(32'h3c7fc612),
	.w6(32'hbbb8084d),
	.w7(32'hb8ce5689),
	.w8(32'hbb9b1308),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea1b8c),
	.w1(32'hbca831cd),
	.w2(32'h3a47b31b),
	.w3(32'hbbbe164b),
	.w4(32'h3b70cf9f),
	.w5(32'h3ad67293),
	.w6(32'h3b188bcf),
	.w7(32'hbc8ab7bf),
	.w8(32'h3c4c35ed),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad993df),
	.w1(32'hbc33776d),
	.w2(32'h3add2c06),
	.w3(32'h3a56ef98),
	.w4(32'h3a991cac),
	.w5(32'hbc34bb26),
	.w6(32'h3b48e0cc),
	.w7(32'hbb59ac51),
	.w8(32'h3be0e113),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15fb81),
	.w1(32'hbc0e022b),
	.w2(32'hbc368b78),
	.w3(32'hbb320169),
	.w4(32'hbba5d51e),
	.w5(32'hba58346e),
	.w6(32'h3cafdb23),
	.w7(32'h3be1d56b),
	.w8(32'hba038f06),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab429a1),
	.w1(32'h3af3cc82),
	.w2(32'h3b192ad1),
	.w3(32'h395dae47),
	.w4(32'hba5bdaf8),
	.w5(32'hb6f84191),
	.w6(32'h39933f6e),
	.w7(32'h3b7e4f49),
	.w8(32'hbbc1829e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaef1ef),
	.w1(32'h398a1c9f),
	.w2(32'hbbabc405),
	.w3(32'hbb48e6aa),
	.w4(32'h39264d5b),
	.w5(32'hbb1961b2),
	.w6(32'hbb6a0172),
	.w7(32'hbb6153b4),
	.w8(32'hbb688edf),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939ca8),
	.w1(32'hbbdb3900),
	.w2(32'hbbd1b367),
	.w3(32'hbbda2dfc),
	.w4(32'hbb8b71ec),
	.w5(32'hbc1518d8),
	.w6(32'hbb9f6115),
	.w7(32'hbbd48b18),
	.w8(32'hbcd3715e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9c2f1),
	.w1(32'h3b6c562a),
	.w2(32'hba5ef135),
	.w3(32'hbb1123e4),
	.w4(32'h3aa109f8),
	.w5(32'hbbb25197),
	.w6(32'hbc36c795),
	.w7(32'hbc0d9ba7),
	.w8(32'h3af4c7be),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa464b3),
	.w1(32'hbc393bf8),
	.w2(32'hbbe704b6),
	.w3(32'hbbc5efc8),
	.w4(32'hbb0b4aba),
	.w5(32'hba458969),
	.w6(32'hbba2648b),
	.w7(32'hbbc19297),
	.w8(32'h3b4c9a77),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3ebcc),
	.w1(32'h3b5f0d21),
	.w2(32'h3a39dd0a),
	.w3(32'h3b0fc4ce),
	.w4(32'h3ad45caf),
	.w5(32'hbc376b15),
	.w6(32'h3b731989),
	.w7(32'h3a0f64da),
	.w8(32'h3b80c445),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16e466),
	.w1(32'h3c516e4e),
	.w2(32'h3c4b2d83),
	.w3(32'hbc66c96b),
	.w4(32'hbc390451),
	.w5(32'h3b92fae5),
	.w6(32'h3926aec2),
	.w7(32'hbb2192ac),
	.w8(32'h3b041e85),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a656d4d),
	.w1(32'h39ea8a48),
	.w2(32'h39f4d240),
	.w3(32'h3bf32d10),
	.w4(32'hbae4e183),
	.w5(32'hbbf66650),
	.w6(32'hbbe37803),
	.w7(32'hb9d5f2eb),
	.w8(32'h37129ef6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7986c),
	.w1(32'hb88e756c),
	.w2(32'hba7ab804),
	.w3(32'hbb50361a),
	.w4(32'hbb1ca516),
	.w5(32'h3c7fbf03),
	.w6(32'h3a351060),
	.w7(32'hba1b0eb7),
	.w8(32'h3bbb2f71),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb21289),
	.w1(32'hbbe8a70a),
	.w2(32'hbbc3ee5f),
	.w3(32'h3bd851aa),
	.w4(32'h3b8c6191),
	.w5(32'h3b0b2da9),
	.w6(32'hbb96fdb9),
	.w7(32'h3c12e560),
	.w8(32'hbaba2322),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3dfb8),
	.w1(32'hbaf08aa1),
	.w2(32'hbaf12519),
	.w3(32'hb956768e),
	.w4(32'hbbefb0bf),
	.w5(32'hba984a60),
	.w6(32'h3c50ef35),
	.w7(32'hb9cf8d3b),
	.w8(32'hbbada089),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983afdb),
	.w1(32'h396c291c),
	.w2(32'h3b0fc563),
	.w3(32'h3b7775e6),
	.w4(32'h3b84ec2b),
	.w5(32'h3a0ed72e),
	.w6(32'hbb335d87),
	.w7(32'h3b016419),
	.w8(32'h3a9b37fc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa55ca2),
	.w1(32'hbb1f5dfe),
	.w2(32'hbbaa7de8),
	.w3(32'hbb9c0259),
	.w4(32'hbb5713ae),
	.w5(32'hbbff4573),
	.w6(32'hbb00781e),
	.w7(32'hbb5c8cc6),
	.w8(32'hbac4e1af),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0ceed),
	.w1(32'h363747d9),
	.w2(32'hbb90aa34),
	.w3(32'h3a19da24),
	.w4(32'h3aa54e05),
	.w5(32'hb98db5ef),
	.w6(32'h3aaf0c9c),
	.w7(32'hba139f53),
	.w8(32'hbbef0574),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567a65),
	.w1(32'hba8d2d40),
	.w2(32'hbb877dda),
	.w3(32'hbb3ea2b7),
	.w4(32'h3a2e8c1b),
	.w5(32'hbc007031),
	.w6(32'hbbea63de),
	.w7(32'hbb882857),
	.w8(32'hbb6ebeb1),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae50b36),
	.w1(32'h3bf1a312),
	.w2(32'h3b886793),
	.w3(32'h3c25d4a1),
	.w4(32'h3bfe086f),
	.w5(32'hbb2ab959),
	.w6(32'h3c91df33),
	.w7(32'h3b80f2a3),
	.w8(32'h3b042636),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba380e69),
	.w1(32'h3b34dc78),
	.w2(32'h3a26401a),
	.w3(32'hba4a361c),
	.w4(32'hbb157274),
	.w5(32'h3a22ac9b),
	.w6(32'h3b2b568a),
	.w7(32'h3b351043),
	.w8(32'h3b9b4555),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b305efc),
	.w1(32'h390f5140),
	.w2(32'h3928166a),
	.w3(32'h3a69e171),
	.w4(32'h3b8cc4b9),
	.w5(32'h3b3f78b0),
	.w6(32'h3b39861f),
	.w7(32'h3b4c396e),
	.w8(32'h3ae4313f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ecbf8),
	.w1(32'hbb9632b7),
	.w2(32'h3a5b36fa),
	.w3(32'h3c07623c),
	.w4(32'h3b174250),
	.w5(32'hbbcfa2dd),
	.w6(32'h3b143267),
	.w7(32'h3bdcf2de),
	.w8(32'h3ae99469),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0970a4),
	.w1(32'h3b58f4d9),
	.w2(32'h3b819645),
	.w3(32'h3af90217),
	.w4(32'hba4a4737),
	.w5(32'hbb532efe),
	.w6(32'h3b06dff8),
	.w7(32'h3b1ec208),
	.w8(32'hbb0aa0ec),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc198b0),
	.w1(32'h39b97673),
	.w2(32'h3ba20de0),
	.w3(32'hbb520a26),
	.w4(32'hbb6b0494),
	.w5(32'hb9c46841),
	.w6(32'hb887709c),
	.w7(32'h3bbd25b0),
	.w8(32'h3a95a63a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a334d46),
	.w1(32'h3b93d653),
	.w2(32'h3b3d5f7e),
	.w3(32'h3b9a2d4c),
	.w4(32'hb8eb35d0),
	.w5(32'hba654c30),
	.w6(32'h3a7bf466),
	.w7(32'hbace31d1),
	.w8(32'hba31fbde),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0e217),
	.w1(32'h3bd387d1),
	.w2(32'h3c026cb8),
	.w3(32'hbbb1220c),
	.w4(32'hbb22fc3b),
	.w5(32'h3aadd8c9),
	.w6(32'hbb1b112f),
	.w7(32'h3b0faf2f),
	.w8(32'h399de7be),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30652e),
	.w1(32'h3b540032),
	.w2(32'h3adeee02),
	.w3(32'hbbdb23e3),
	.w4(32'h39994721),
	.w5(32'hbb1b55df),
	.w6(32'hbb45f619),
	.w7(32'hb89a9c7a),
	.w8(32'hbb127687),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26e284),
	.w1(32'h3a133926),
	.w2(32'hbabb37e2),
	.w3(32'hbbae24cf),
	.w4(32'h3a52f265),
	.w5(32'h3b422518),
	.w6(32'hbb872afd),
	.w7(32'hbb83de1c),
	.w8(32'h3bbe0c14),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71ba68),
	.w1(32'hbbd53f21),
	.w2(32'hbc4d35c7),
	.w3(32'h3cc6fef2),
	.w4(32'h3c9f2014),
	.w5(32'hbaa62b63),
	.w6(32'h3c130c85),
	.w7(32'h3bf32552),
	.w8(32'h3b8645a0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af05686),
	.w1(32'hbb264bde),
	.w2(32'h3b3731a6),
	.w3(32'h3b5ef244),
	.w4(32'h3acd8abc),
	.w5(32'hbbdfc50f),
	.w6(32'h3b9b5055),
	.w7(32'h3b0112c0),
	.w8(32'h3ccc9dc5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e51ff),
	.w1(32'h3d252115),
	.w2(32'h3c398f7f),
	.w3(32'h3d107130),
	.w4(32'h3c5e3b2d),
	.w5(32'hbb680d03),
	.w6(32'h3d6645a7),
	.w7(32'h3cbb3970),
	.w8(32'h3a3d0585),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9340),
	.w1(32'h3c0caa61),
	.w2(32'hbb7b1c61),
	.w3(32'hbbaa1f05),
	.w4(32'hbaa9af15),
	.w5(32'hbbce8c8d),
	.w6(32'h3bcfacba),
	.w7(32'h3a8f9396),
	.w8(32'hbb9cda07),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39ac2e),
	.w1(32'hbbcf239b),
	.w2(32'hbc040a4a),
	.w3(32'hbc2428e5),
	.w4(32'hbc5437ff),
	.w5(32'hbc07b515),
	.w6(32'hbc461f54),
	.w7(32'hbbac4b8d),
	.w8(32'hbbb57fca),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f10f0),
	.w1(32'hbbcc1b1b),
	.w2(32'hbc1b1dbe),
	.w3(32'hbc18ca66),
	.w4(32'hbc28a6b6),
	.w5(32'hbbe12bb2),
	.w6(32'h3a9e948a),
	.w7(32'h3af7e1b9),
	.w8(32'hbbdd156e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fedb9),
	.w1(32'h3992274e),
	.w2(32'h3a811513),
	.w3(32'hbbd0739c),
	.w4(32'hbbdef144),
	.w5(32'hbc2c9113),
	.w6(32'hbc05904a),
	.w7(32'hbb2888ed),
	.w8(32'hbc0cfae0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020504),
	.w1(32'h38c92a2b),
	.w2(32'hbb1b2745),
	.w3(32'h3b8d6b37),
	.w4(32'hba8c9ad4),
	.w5(32'hbb479b60),
	.w6(32'h3c475e6b),
	.w7(32'hbb417231),
	.w8(32'hbb281af5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bf987),
	.w1(32'hba82f26a),
	.w2(32'hbb0fd973),
	.w3(32'hbbf05b1d),
	.w4(32'hbb2812f7),
	.w5(32'hbabbdbca),
	.w6(32'hbb95341c),
	.w7(32'hbba448f2),
	.w8(32'h3b813705),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02c267),
	.w1(32'hbb51f805),
	.w2(32'hbb0363e8),
	.w3(32'hbbc0b72a),
	.w4(32'hbb2bf88b),
	.w5(32'hbba79081),
	.w6(32'hbb95c30c),
	.w7(32'h3bd3c1af),
	.w8(32'hbb750882),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bbc95e),
	.w1(32'hbb393efb),
	.w2(32'hbb64e47a),
	.w3(32'hbb3c8e08),
	.w4(32'h3a99f415),
	.w5(32'hbbc8a179),
	.w6(32'hbae0929c),
	.w7(32'hba8d3058),
	.w8(32'hbbbb574b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc4d73),
	.w1(32'hba893b4a),
	.w2(32'hba10e7f5),
	.w3(32'h3a774835),
	.w4(32'hbac0e637),
	.w5(32'h3c923ed6),
	.w6(32'hba8d2960),
	.w7(32'hba0aa723),
	.w8(32'h3cf696c9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfa151),
	.w1(32'hbbc02990),
	.w2(32'hbc0af5d6),
	.w3(32'h3cb261dc),
	.w4(32'h3c574732),
	.w5(32'hbbb8d9b0),
	.w6(32'h3c107154),
	.w7(32'h3c7d742f),
	.w8(32'hbc370063),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ed1fc),
	.w1(32'hbc1f942a),
	.w2(32'hbbae3b48),
	.w3(32'hbb40d21a),
	.w4(32'hba3b20c3),
	.w5(32'h3bb4f015),
	.w6(32'hbbd8d264),
	.w7(32'hbc3d54b0),
	.w8(32'h3b4de238),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8b611),
	.w1(32'hbbbe3223),
	.w2(32'h3aea9415),
	.w3(32'h3a8a7dd7),
	.w4(32'h3ad1532d),
	.w5(32'hbbcdb9ec),
	.w6(32'hbbddf8e1),
	.w7(32'h3bd834e7),
	.w8(32'h3cd4abfb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ee7e),
	.w1(32'h3b876dbc),
	.w2(32'hbbda3727),
	.w3(32'h3bc101d3),
	.w4(32'h38a74145),
	.w5(32'hba27c0cc),
	.w6(32'h3d07fb1c),
	.w7(32'h3c1f63bb),
	.w8(32'hb8a73880),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8da2e),
	.w1(32'h3916a1dc),
	.w2(32'h3a1f7b8d),
	.w3(32'h3abf4227),
	.w4(32'h39aa2c29),
	.w5(32'hba73c485),
	.w6(32'h3b3202d0),
	.w7(32'h3a4d3123),
	.w8(32'hbb6a5a62),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba234f4),
	.w1(32'h3b57d2ee),
	.w2(32'h3b5d29c6),
	.w3(32'h3bbecb2b),
	.w4(32'h3bf57be4),
	.w5(32'hbc971908),
	.w6(32'h3b240b0d),
	.w7(32'h3b821ed0),
	.w8(32'hbc893dc1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d119e),
	.w1(32'hbc178fe3),
	.w2(32'hba902fde),
	.w3(32'hbc848d9b),
	.w4(32'hbbabd9c6),
	.w5(32'h3b5e3509),
	.w6(32'hbc1bc12e),
	.w7(32'hba640ab8),
	.w8(32'hbad524dd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c137fd9),
	.w1(32'h39ba9791),
	.w2(32'h3c16647e),
	.w3(32'h3942a120),
	.w4(32'hbbbc792c),
	.w5(32'h3b9abba8),
	.w6(32'hbc4de5c3),
	.w7(32'h39694a2e),
	.w8(32'hbac26215),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54177e),
	.w1(32'hbb16bcd9),
	.w2(32'hba458120),
	.w3(32'h39c60aaf),
	.w4(32'h3b7c363f),
	.w5(32'hbb31f01d),
	.w6(32'hbb673519),
	.w7(32'h3b1e7f02),
	.w8(32'hbb78056f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f547b),
	.w1(32'h3bb8983c),
	.w2(32'hb9ac31ee),
	.w3(32'h3b0e2aea),
	.w4(32'hba50fcc9),
	.w5(32'hba8db2be),
	.w6(32'h3b97edd5),
	.w7(32'h3ae3fa52),
	.w8(32'h3b843df0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc950d5),
	.w1(32'h3b87ea08),
	.w2(32'hbad3c90e),
	.w3(32'hbc1c61df),
	.w4(32'hbc32a412),
	.w5(32'hbb3d0338),
	.w6(32'h3c315ae7),
	.w7(32'h3a7ee34f),
	.w8(32'h3a9fb335),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964c05c),
	.w1(32'hbadc4a35),
	.w2(32'h3ae194fb),
	.w3(32'h39f8b6a6),
	.w4(32'h3ab12ba0),
	.w5(32'h39dff060),
	.w6(32'h3872bd2e),
	.w7(32'h3ba0eb83),
	.w8(32'h3afd6686),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84fd4e),
	.w1(32'h3af70b00),
	.w2(32'h3a329e24),
	.w3(32'hbb1b1d17),
	.w4(32'hbb0398c8),
	.w5(32'hba448145),
	.w6(32'h3c0150a1),
	.w7(32'h3999c3e1),
	.w8(32'hbb06b208),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33f17f),
	.w1(32'h3b05b730),
	.w2(32'h3b98c1c1),
	.w3(32'hbb937e39),
	.w4(32'hbacc04e5),
	.w5(32'hbb7ef7df),
	.w6(32'h3b63ce7b),
	.w7(32'h3ae23e5c),
	.w8(32'h3b452397),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a220dd4),
	.w1(32'hbc0a33eb),
	.w2(32'h3b33c517),
	.w3(32'h386d83fe),
	.w4(32'h3b7b0efd),
	.w5(32'hbac85dc3),
	.w6(32'h3cd08b15),
	.w7(32'hbba97da2),
	.w8(32'h3a3c20df),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71b3bf),
	.w1(32'hba9d6e3b),
	.w2(32'h3b6c257f),
	.w3(32'h3a69a005),
	.w4(32'h39f6fddb),
	.w5(32'h3b679203),
	.w6(32'h3b818f2b),
	.w7(32'hbb33bf53),
	.w8(32'hbb9bf68b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a51b8),
	.w1(32'h3aa9cc4d),
	.w2(32'h3ae9bce4),
	.w3(32'hbbb1d51b),
	.w4(32'hbb8d6e47),
	.w5(32'h3b0fd345),
	.w6(32'hbb21dee9),
	.w7(32'hbabed150),
	.w8(32'hba3dca11),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac35c3b),
	.w1(32'hbab4270e),
	.w2(32'h3afa62de),
	.w3(32'h3b637ba0),
	.w4(32'h3a757812),
	.w5(32'h386ac767),
	.w6(32'h3b5f294e),
	.w7(32'h3a8ee92f),
	.w8(32'hbbbc0a7c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6d5ab),
	.w1(32'h3aae909c),
	.w2(32'h3b739761),
	.w3(32'hbb87d5d2),
	.w4(32'hb9f45f6b),
	.w5(32'hbb15669e),
	.w6(32'hbb85b998),
	.w7(32'hb67e6c21),
	.w8(32'hbb089a8b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91cb45),
	.w1(32'h3ba23f2c),
	.w2(32'h3991e8e8),
	.w3(32'hbb9ffcb6),
	.w4(32'hbb4f41f3),
	.w5(32'h3c610270),
	.w6(32'hbab4bada),
	.w7(32'hbb876816),
	.w8(32'hbc8b8c5b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc291bb4),
	.w1(32'hbc5d8f6b),
	.w2(32'h3caa87c1),
	.w3(32'hbcc9f4fd),
	.w4(32'hbc41b995),
	.w5(32'h3a04155b),
	.w6(32'hbc6b3831),
	.w7(32'hbc245401),
	.w8(32'h3b470a4a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a900e4),
	.w1(32'h3b687576),
	.w2(32'h3bc9465b),
	.w3(32'h3bca963e),
	.w4(32'h3baded43),
	.w5(32'h3cd01a91),
	.w6(32'h3c0b3260),
	.w7(32'h3a97d486),
	.w8(32'hbc165fed),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b15e8),
	.w1(32'hbc7b4ce4),
	.w2(32'h3c1a0d45),
	.w3(32'hbb9149d6),
	.w4(32'hb9ee12d7),
	.w5(32'hbb4c160d),
	.w6(32'hbc1d5b03),
	.w7(32'hbc6c8a19),
	.w8(32'h3b6dc7da),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b021883),
	.w1(32'hbb35c9f3),
	.w2(32'hbc0ee449),
	.w3(32'h39203396),
	.w4(32'hbb31f125),
	.w5(32'hbad006c6),
	.w6(32'h3c4007a2),
	.w7(32'hbbab5bfc),
	.w8(32'hbba99c10),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ad2f1),
	.w1(32'h3adc33a5),
	.w2(32'hbb851333),
	.w3(32'hbb66cea6),
	.w4(32'hbaec7524),
	.w5(32'hbc265e5a),
	.w6(32'h3aacace4),
	.w7(32'hbac44242),
	.w8(32'hba23232d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afed561),
	.w1(32'hbb93ee2d),
	.w2(32'h3b931902),
	.w3(32'hbb802c6d),
	.w4(32'hbb1599cb),
	.w5(32'h39787e9e),
	.w6(32'h3ade8837),
	.w7(32'h3930ead8),
	.w8(32'hbb50e386),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18dfc0),
	.w1(32'h3b3093fd),
	.w2(32'h3b4bd5c9),
	.w3(32'h3aefb0d4),
	.w4(32'hb9fe4b8c),
	.w5(32'hb8c4d0a3),
	.w6(32'h3a987d8e),
	.w7(32'h3ab2a59a),
	.w8(32'h3c4ac05b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16af6c),
	.w1(32'h3b82f817),
	.w2(32'hbb92de15),
	.w3(32'h3b0c3eea),
	.w4(32'hbb9470f8),
	.w5(32'h3b1a6759),
	.w6(32'h3c3db0ec),
	.w7(32'hbab92929),
	.w8(32'hba93f64c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8512df),
	.w1(32'h3898af80),
	.w2(32'h3b9f9517),
	.w3(32'hbb941506),
	.w4(32'hbaf9e7bf),
	.w5(32'hbc17e82b),
	.w6(32'hbb1f6f87),
	.w7(32'hbb2ff127),
	.w8(32'h3b7cb2a0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0abe80),
	.w1(32'hbbc6ae62),
	.w2(32'hbc185e90),
	.w3(32'hba55c0b1),
	.w4(32'hbb3a1f02),
	.w5(32'hbb9df196),
	.w6(32'h3af16b85),
	.w7(32'hbc19bf6f),
	.w8(32'hbc17448d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1649fb),
	.w1(32'h3b2ca6f6),
	.w2(32'h3b8716b7),
	.w3(32'hbbd15284),
	.w4(32'h3af1f1cd),
	.w5(32'h3bb99a7a),
	.w6(32'hbbd75af2),
	.w7(32'hba95661d),
	.w8(32'h3bc8710d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6883d),
	.w1(32'hbafe9ad2),
	.w2(32'hbb29cf5d),
	.w3(32'h3ba8b0ef),
	.w4(32'h3b7e232c),
	.w5(32'hb9cf8684),
	.w6(32'h3c14723e),
	.w7(32'h3b231b3c),
	.w8(32'h3b2c8e1d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f9b88),
	.w1(32'hb91edd4d),
	.w2(32'hbb297cbc),
	.w3(32'hbafac5ab),
	.w4(32'hbb1fc80a),
	.w5(32'h3b3ce309),
	.w6(32'h3b8a61db),
	.w7(32'hba5f2dd4),
	.w8(32'hbab534f0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abda7d4),
	.w1(32'h395527aa),
	.w2(32'h3aaa36dd),
	.w3(32'hbb2b8455),
	.w4(32'hb9b10385),
	.w5(32'h3b15a432),
	.w6(32'hb978b17e),
	.w7(32'hbc0cccd8),
	.w8(32'hbbbdbd4b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1cd06),
	.w1(32'h3bd14907),
	.w2(32'h3b8d4a32),
	.w3(32'hbb586a2a),
	.w4(32'hbb953fe6),
	.w5(32'h3b76ef6f),
	.w6(32'h3b1e1d47),
	.w7(32'h39f2a0aa),
	.w8(32'h3c025386),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf72072),
	.w1(32'hbbcf8a41),
	.w2(32'h3b019f05),
	.w3(32'h3c4cc9f0),
	.w4(32'hbb08736e),
	.w5(32'hba1f6f5d),
	.w6(32'h3c6be2fc),
	.w7(32'hbb2dd871),
	.w8(32'hba56ff8b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d30667),
	.w1(32'hba9f26c4),
	.w2(32'hb9c347d3),
	.w3(32'hba9d22d5),
	.w4(32'hba37283e),
	.w5(32'h39d7b98a),
	.w6(32'hbaeacfcf),
	.w7(32'hba8918c8),
	.w8(32'h3a31ea2e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a819dc),
	.w1(32'h39ad11b5),
	.w2(32'hb92cd936),
	.w3(32'h3ad644b4),
	.w4(32'h3a64df1f),
	.w5(32'h39f0f57e),
	.w6(32'h3abbff8d),
	.w7(32'h3aa7ba20),
	.w8(32'hba1d1671),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cf45d),
	.w1(32'hba31ad84),
	.w2(32'h39f8b10f),
	.w3(32'h39078d37),
	.w4(32'h38589448),
	.w5(32'hb62f9b64),
	.w6(32'hbb078124),
	.w7(32'hb9d29fc6),
	.w8(32'hba5761d0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e2316),
	.w1(32'h3991b29f),
	.w2(32'h39d01a36),
	.w3(32'hb9bc88b2),
	.w4(32'h3991fd79),
	.w5(32'h3a1b8acf),
	.w6(32'h3a1952e5),
	.w7(32'hb9a6c6a9),
	.w8(32'h3a2a5c52),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dfce2),
	.w1(32'h399ee615),
	.w2(32'h3a06b95a),
	.w3(32'h39295d5d),
	.w4(32'h3a165605),
	.w5(32'h3aa8046f),
	.w6(32'h396b73a4),
	.w7(32'h3a1a0bf1),
	.w8(32'h3af5773b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf2535),
	.w1(32'h3a62a889),
	.w2(32'h395fcec0),
	.w3(32'h3ab4bef9),
	.w4(32'h39f93776),
	.w5(32'h3a8e7e8a),
	.w6(32'h3ab2b95d),
	.w7(32'h3996e1db),
	.w8(32'hba6e4a7a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979130b),
	.w1(32'hb98c9c8f),
	.w2(32'h39ebcfb6),
	.w3(32'hb92e4cfc),
	.w4(32'hb915331c),
	.w5(32'h39a1d492),
	.w6(32'hba99689d),
	.w7(32'h3861a4e6),
	.w8(32'h390d02c1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ffb3c),
	.w1(32'hb8bbb568),
	.w2(32'hb871d84a),
	.w3(32'h3a1bd13f),
	.w4(32'h38909b84),
	.w5(32'h3a44d395),
	.w6(32'h39e8318e),
	.w7(32'h3923c565),
	.w8(32'h3835ba95),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38d489),
	.w1(32'h3a02cd69),
	.w2(32'h39a42881),
	.w3(32'h38855c15),
	.w4(32'hb94152e3),
	.w5(32'h393fcbce),
	.w6(32'hb9f325ab),
	.w7(32'h39a16ded),
	.w8(32'h39b0cd09),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38815bf0),
	.w1(32'hb9a5fb5c),
	.w2(32'h38cd7832),
	.w3(32'hb8b77bfe),
	.w4(32'hb7c2c219),
	.w5(32'h38d2cca1),
	.w6(32'h39240939),
	.w7(32'h399e5c46),
	.w8(32'hb9890c31),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05f92d),
	.w1(32'hba0eda88),
	.w2(32'h36e34663),
	.w3(32'hba56a49a),
	.w4(32'hb92b34e8),
	.w5(32'hba53b8a3),
	.w6(32'hbab288f2),
	.w7(32'hba2db302),
	.w8(32'hba9f5d6a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba417826),
	.w1(32'hba433657),
	.w2(32'hb8a2ff28),
	.w3(32'hba98305b),
	.w4(32'hba1cd95c),
	.w5(32'h3a444f4a),
	.w6(32'hbabebc48),
	.w7(32'hb9c7f128),
	.w8(32'h39bff84c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ebb38),
	.w1(32'h39dbde4b),
	.w2(32'h39fb4f46),
	.w3(32'h39c82392),
	.w4(32'h3a6d38ea),
	.w5(32'hb976963e),
	.w6(32'hb99c15f2),
	.w7(32'h3a43a1f1),
	.w8(32'hb910eb60),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb894ceae),
	.w1(32'h3a1b3981),
	.w2(32'hb82ce005),
	.w3(32'h39c68739),
	.w4(32'h380f3d74),
	.w5(32'hb974190b),
	.w6(32'h39fbec02),
	.w7(32'h393a86a3),
	.w8(32'hba15bcc1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dc8a90),
	.w1(32'hb9739863),
	.w2(32'hb8d74aca),
	.w3(32'hba3f416c),
	.w4(32'hb94d9fe8),
	.w5(32'h3a41dd06),
	.w6(32'hba68ee5c),
	.w7(32'hba46c371),
	.w8(32'h3a21ed4d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cddb7c),
	.w1(32'h3a08b0b9),
	.w2(32'h39c49871),
	.w3(32'h36c0e273),
	.w4(32'hb9560383),
	.w5(32'hba1002da),
	.w6(32'h3a012966),
	.w7(32'h39f567de),
	.w8(32'h39d6d917),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38021cc5),
	.w1(32'hb9378303),
	.w2(32'h3a01d4d9),
	.w3(32'hba01b2b5),
	.w4(32'hba273591),
	.w5(32'hb8880150),
	.w6(32'hba337e55),
	.w7(32'hb99fe18a),
	.w8(32'hb9c578b3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c7f40),
	.w1(32'h3981dfcf),
	.w2(32'h39ecf32c),
	.w3(32'h37f3c819),
	.w4(32'h39d5b52f),
	.w5(32'hba480c4a),
	.w6(32'h39a8dff0),
	.w7(32'h39457c60),
	.w8(32'hb9a3b492),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bfe73),
	.w1(32'hba8f3b55),
	.w2(32'hba8d9339),
	.w3(32'hba63c66d),
	.w4(32'hba1b49a8),
	.w5(32'h3a05c0d2),
	.w6(32'hb9c65ada),
	.w7(32'hb9f062da),
	.w8(32'hb8e4acce),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9b113),
	.w1(32'hb9c044b0),
	.w2(32'hb96b6008),
	.w3(32'h3a22ab7a),
	.w4(32'h3a00d831),
	.w5(32'h37085a78),
	.w6(32'h3992c3c7),
	.w7(32'h38ca81f2),
	.w8(32'hba0994c7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef4a64),
	.w1(32'hb9ef1bdd),
	.w2(32'hb97a1c89),
	.w3(32'hb88032e9),
	.w4(32'hb9565b03),
	.w5(32'hbaa33c56),
	.w6(32'hb9cb0988),
	.w7(32'hba20ca4d),
	.w8(32'hbb0908bd),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8df43),
	.w1(32'hbb266f48),
	.w2(32'hbaa9305f),
	.w3(32'hbad76866),
	.w4(32'hba9212e8),
	.w5(32'h388bf017),
	.w6(32'hbb8bc527),
	.w7(32'hbb1d4a95),
	.w8(32'h39e1bb38),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981dfa9),
	.w1(32'h39b46665),
	.w2(32'h3951c4c9),
	.w3(32'hb81b7fa7),
	.w4(32'h39a93a99),
	.w5(32'hba159933),
	.w6(32'h39879d84),
	.w7(32'h3a04076d),
	.w8(32'hba7ec1ea),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0597e2),
	.w1(32'hb9b9cf78),
	.w2(32'hb9bee163),
	.w3(32'h3891b88b),
	.w4(32'hba440e4a),
	.w5(32'hb8eaf985),
	.w6(32'hba6bf7b4),
	.w7(32'hba7dd235),
	.w8(32'hb97a87e2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396436b3),
	.w1(32'h3a9fd52a),
	.w2(32'h39e4ad2c),
	.w3(32'h3a1046a3),
	.w4(32'h3645fc2c),
	.w5(32'h39be20b2),
	.w6(32'h3aaa21eb),
	.w7(32'hb755a0c2),
	.w8(32'h3998730b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982b509),
	.w1(32'h392f7849),
	.w2(32'h3913c52e),
	.w3(32'h39d1f5ef),
	.w4(32'hb9868238),
	.w5(32'h3980fdc8),
	.w6(32'h3a8ac79b),
	.w7(32'h38d22f47),
	.w8(32'h3a0adcbd),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d7a79),
	.w1(32'h3a986fa2),
	.w2(32'h3a090f9d),
	.w3(32'h3a4e45e9),
	.w4(32'h3a4bf722),
	.w5(32'h3a24efc4),
	.w6(32'h3ac0c7b2),
	.w7(32'h3a176a51),
	.w8(32'hb9047df5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be86cf),
	.w1(32'h39ac2538),
	.w2(32'h3a8a52e9),
	.w3(32'h3987ad64),
	.w4(32'hb9499151),
	.w5(32'hba1f8a59),
	.w6(32'h3a03bb77),
	.w7(32'h397e199e),
	.w8(32'hb92125eb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f66813),
	.w1(32'hb98a446b),
	.w2(32'h39185509),
	.w3(32'hba27fca2),
	.w4(32'hb9814e89),
	.w5(32'hb9555e5c),
	.w6(32'h3a23a0a8),
	.w7(32'h3a169b6b),
	.w8(32'h399620a0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38760955),
	.w1(32'h390127aa),
	.w2(32'h39c35708),
	.w3(32'h393c72a4),
	.w4(32'hb932df35),
	.w5(32'hb9284264),
	.w6(32'hba351c02),
	.w7(32'hb9de141f),
	.w8(32'hb9d965b2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule