module layer_10_featuremap_135(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeed25b),
	.w1(32'hba8aa190),
	.w2(32'h3981ab17),
	.w3(32'hbada2daa),
	.w4(32'h3b0be70c),
	.w5(32'h3b4ae528),
	.w6(32'hbbc73c7e),
	.w7(32'hbbca1e10),
	.w8(32'hbc106724),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba50b1d),
	.w1(32'h3adaf879),
	.w2(32'h3b71f176),
	.w3(32'hbb2cdd32),
	.w4(32'h3789567a),
	.w5(32'h3a62c3f1),
	.w6(32'h3a3f03bd),
	.w7(32'h3ae61603),
	.w8(32'hb9a021e9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16be86),
	.w1(32'h3a96b7a3),
	.w2(32'h3b357590),
	.w3(32'hba7cb5ae),
	.w4(32'hb9b69707),
	.w5(32'hbaa8141f),
	.w6(32'hbab15468),
	.w7(32'hba3188e8),
	.w8(32'hbb4a2afe),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad4ea4),
	.w1(32'hbb8a2a89),
	.w2(32'hbb88961a),
	.w3(32'hbb41d58e),
	.w4(32'hbb32a8ef),
	.w5(32'hbb2f2c55),
	.w6(32'h3ada1b6d),
	.w7(32'h3b28c7ab),
	.w8(32'h3abbc272),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b70bd),
	.w1(32'hbb92427f),
	.w2(32'hbb3ae09c),
	.w3(32'hbb8a9182),
	.w4(32'hbb8430bd),
	.w5(32'hbb6cd231),
	.w6(32'hbb5a1260),
	.w7(32'hbaf80e32),
	.w8(32'hb875f1b0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91fcc0),
	.w1(32'hbad79708),
	.w2(32'hbae6b580),
	.w3(32'hba0bcf57),
	.w4(32'hbacfe62e),
	.w5(32'hbabe7790),
	.w6(32'hba996ce6),
	.w7(32'hba08978f),
	.w8(32'h38fc6d76),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11a09a),
	.w1(32'h39851759),
	.w2(32'h3b402116),
	.w3(32'hba59a0e7),
	.w4(32'hba924d62),
	.w5(32'h397d90b9),
	.w6(32'hb9ec2860),
	.w7(32'hb95b484b),
	.w8(32'hbae4c29b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba207155),
	.w1(32'hbb60640e),
	.w2(32'hbb96f027),
	.w3(32'hbabf989d),
	.w4(32'hbb407d89),
	.w5(32'hbb47e3b0),
	.w6(32'hbb2c2b50),
	.w7(32'hbb41a19b),
	.w8(32'hbaffc7f4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cd44b),
	.w1(32'hb923802f),
	.w2(32'h3a027203),
	.w3(32'hbb01a1fd),
	.w4(32'hba4e1d63),
	.w5(32'hb8f8530c),
	.w6(32'h392fe139),
	.w7(32'hb9a956f7),
	.w8(32'hba474ca3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a78852),
	.w1(32'h3bceb44d),
	.w2(32'h3be0f17f),
	.w3(32'hb81b0566),
	.w4(32'h3b9dd1b6),
	.w5(32'h3b86be35),
	.w6(32'h3bde3010),
	.w7(32'h3be4ed65),
	.w8(32'h3b2c0270),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18db95),
	.w1(32'h3b590bb2),
	.w2(32'h3b38f5ac),
	.w3(32'h3ada87be),
	.w4(32'hba80fbd8),
	.w5(32'hbab02c10),
	.w6(32'h3a302401),
	.w7(32'hba83aa9c),
	.w8(32'hb7f9e28d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dea06),
	.w1(32'hbb40a349),
	.w2(32'hbbd11bde),
	.w3(32'hba8c41a1),
	.w4(32'hbad2ff8b),
	.w5(32'hbb632483),
	.w6(32'hbb222ddc),
	.w7(32'hbb47bb91),
	.w8(32'hbb30f0b8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63eb2f),
	.w1(32'hbaa96a18),
	.w2(32'hba9b324e),
	.w3(32'hbb404e4a),
	.w4(32'hba79f194),
	.w5(32'hba17ae94),
	.w6(32'hba9547a0),
	.w7(32'hba97e431),
	.w8(32'hb950085f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36a2d3),
	.w1(32'hba427536),
	.w2(32'hbb52835b),
	.w3(32'h3a0468ed),
	.w4(32'h3a300c54),
	.w5(32'hbad7577e),
	.w6(32'h39b087fe),
	.w7(32'hbb070890),
	.w8(32'h39f0c66d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacc165),
	.w1(32'hbaf822b3),
	.w2(32'hbba3686a),
	.w3(32'h39b84fda),
	.w4(32'hbb83c187),
	.w5(32'hbba4cd7a),
	.w6(32'h3b309a3b),
	.w7(32'h3b113a3b),
	.w8(32'h3a40c566),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0e780),
	.w1(32'h3a148c6a),
	.w2(32'h3b08d708),
	.w3(32'hbb60cad7),
	.w4(32'h39dfb5a8),
	.w5(32'h3a7884af),
	.w6(32'h3a14aacb),
	.w7(32'h3ab6de23),
	.w8(32'h3a67b913),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380912af),
	.w1(32'hba170e96),
	.w2(32'h3990f51a),
	.w3(32'hb9435e40),
	.w4(32'h3621972a),
	.w5(32'hba8838ef),
	.w6(32'h3799e4dd),
	.w7(32'hba41a4dc),
	.w8(32'hbab3f503),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac09f84),
	.w1(32'h3b9906b7),
	.w2(32'h3bb0a918),
	.w3(32'hb83be7f5),
	.w4(32'h3ae6fa5f),
	.w5(32'h3b25c2f8),
	.w6(32'h3b78eba6),
	.w7(32'h3b676f2a),
	.w8(32'hb89e9ea5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7d6db),
	.w1(32'h38ad1986),
	.w2(32'h39c19220),
	.w3(32'hba1fcf71),
	.w4(32'hbac7c558),
	.w5(32'hb88a182a),
	.w6(32'hb9f56c8b),
	.w7(32'hba1bf854),
	.w8(32'hbb11c2e4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fbada),
	.w1(32'hb9f2df47),
	.w2(32'h3a05028f),
	.w3(32'hba91f332),
	.w4(32'hba4b08d1),
	.w5(32'h389c2056),
	.w6(32'hb9d569a8),
	.w7(32'h39e748eb),
	.w8(32'h38adda17),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921775e),
	.w1(32'hbabcd861),
	.w2(32'hbae5416a),
	.w3(32'hb95d5db1),
	.w4(32'hba80abf9),
	.w5(32'hbac02f5d),
	.w6(32'hba67de79),
	.w7(32'hbab50ffa),
	.w8(32'hba05e576),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88afba),
	.w1(32'hbb264f54),
	.w2(32'hbb8118e2),
	.w3(32'hba56366e),
	.w4(32'h3ac1cebe),
	.w5(32'h3abe763c),
	.w6(32'hbbb066d8),
	.w7(32'hbbdcec9c),
	.w8(32'hbbdf2f9e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21cdc9),
	.w1(32'h3a8b3c50),
	.w2(32'h3b219a5d),
	.w3(32'h39d96894),
	.w4(32'h3b683ea4),
	.w5(32'h3b8f2579),
	.w6(32'h3b2211d7),
	.w7(32'h3b4e02ec),
	.w8(32'h3b775931),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3862c905),
	.w1(32'hbb528e39),
	.w2(32'hbb823f75),
	.w3(32'h3b32ae3a),
	.w4(32'hbb3a7c71),
	.w5(32'hbb6e73a7),
	.w6(32'hbb1b912f),
	.w7(32'hbb65899b),
	.w8(32'hbb3c3586),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea38c),
	.w1(32'h3aac5581),
	.w2(32'h3b48a63e),
	.w3(32'hbb4d2735),
	.w4(32'hb97ff1b4),
	.w5(32'h3a787650),
	.w6(32'h3ad4cb2c),
	.w7(32'h3b71e078),
	.w8(32'h3a86d780),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3951d1d1),
	.w1(32'h3b44489c),
	.w2(32'h3a8fc3d4),
	.w3(32'hb9f8e854),
	.w4(32'h3b00f5a6),
	.w5(32'h39d92975),
	.w6(32'h3ada5dbf),
	.w7(32'h3a5871c4),
	.w8(32'h39ed6891),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9d72f),
	.w1(32'hba1b741a),
	.w2(32'h383e28b9),
	.w3(32'hb963ca82),
	.w4(32'hba688f77),
	.w5(32'hb96814d7),
	.w6(32'hba107bcf),
	.w7(32'hb91d65dc),
	.w8(32'h39232fbd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba479411),
	.w1(32'hbabf6603),
	.w2(32'hbb12bf33),
	.w3(32'hba47904a),
	.w4(32'h3a4dab1e),
	.w5(32'hba364c5e),
	.w6(32'h3addee78),
	.w7(32'h3b1a0009),
	.w8(32'hba2e8106),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6f494),
	.w1(32'hbab54831),
	.w2(32'h3a6ca13f),
	.w3(32'hbacc0857),
	.w4(32'hbb16dab9),
	.w5(32'hba863664),
	.w6(32'hbb85f21e),
	.w7(32'hbb521cb6),
	.w8(32'hbb2287c7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8b969),
	.w1(32'hba38a765),
	.w2(32'hbaae9ee5),
	.w3(32'h3a09f50c),
	.w4(32'hb89f1d57),
	.w5(32'hba78925a),
	.w6(32'hba8ff561),
	.w7(32'hba38f985),
	.w8(32'hba325df0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac70e6),
	.w1(32'hba8bbe3f),
	.w2(32'hba89a534),
	.w3(32'hb9547c33),
	.w4(32'hba4c3a07),
	.w5(32'hba74c75a),
	.w6(32'hba3c6715),
	.w7(32'hba771971),
	.w8(32'hba0e530e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17ea01),
	.w1(32'hba2746ec),
	.w2(32'hba3c43cf),
	.w3(32'hb9b6bae7),
	.w4(32'hba26fceb),
	.w5(32'hba446437),
	.w6(32'hb91c74b7),
	.w7(32'hba3aa0c9),
	.w8(32'hb9e51b73),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b30f83),
	.w1(32'hba948529),
	.w2(32'h3a9ae006),
	.w3(32'h39525acb),
	.w4(32'hbb1acc67),
	.w5(32'h3ad6dd33),
	.w6(32'hba223596),
	.w7(32'h3a6ad8f0),
	.w8(32'hb9f29e31),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b18e1),
	.w1(32'h3987a141),
	.w2(32'h3b0d92b6),
	.w3(32'h3accc20b),
	.w4(32'hb93c794a),
	.w5(32'h3b205b85),
	.w6(32'hba1dab5d),
	.w7(32'h3a156aeb),
	.w8(32'hb91e3e53),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b8b7c),
	.w1(32'h3b7c5b65),
	.w2(32'h3b6dbd5a),
	.w3(32'h3b2be64e),
	.w4(32'h3b0b463c),
	.w5(32'h3b088ccc),
	.w6(32'h3b77e100),
	.w7(32'h3b8db777),
	.w8(32'hb9f2009e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab40ec5),
	.w1(32'hba06f391),
	.w2(32'hb8fbcdfc),
	.w3(32'h3a02c9c7),
	.w4(32'hba36e068),
	.w5(32'hb99ba370),
	.w6(32'h39f84005),
	.w7(32'h39ba170d),
	.w8(32'h39e78f62),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a826e30),
	.w1(32'h3b20249a),
	.w2(32'h3b56c347),
	.w3(32'h3ab25bc8),
	.w4(32'h3a916c6e),
	.w5(32'hb71edc7c),
	.w6(32'h3b4ce7c6),
	.w7(32'h3b26544c),
	.w8(32'h39a993ce),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9325c7),
	.w1(32'h3a6b0eb8),
	.w2(32'h3b2fc4e3),
	.w3(32'hbaa93fe3),
	.w4(32'hb8fa3ce5),
	.w5(32'h399d86f4),
	.w6(32'hb9423721),
	.w7(32'hba0fa685),
	.w8(32'hbb2768e1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd6c7d),
	.w1(32'hbb8e8a87),
	.w2(32'hbb82b0c1),
	.w3(32'hbb0ece5a),
	.w4(32'hbb575192),
	.w5(32'hbb30f185),
	.w6(32'hbb906af1),
	.w7(32'hbb60e0cb),
	.w8(32'hbaf121a2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134ee9),
	.w1(32'hb91c81d8),
	.w2(32'hb902aae5),
	.w3(32'hbb140753),
	.w4(32'hba1b7fa3),
	.w5(32'hb9daa383),
	.w6(32'hb9c43482),
	.w7(32'hba903b96),
	.w8(32'hbb046139),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16b61a),
	.w1(32'hbac0114e),
	.w2(32'hbb2c5391),
	.w3(32'hb9187df9),
	.w4(32'hb97dc9fa),
	.w5(32'hbad0d04f),
	.w6(32'hbac638d7),
	.w7(32'hbb0c0f12),
	.w8(32'hba554435),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0646e9),
	.w1(32'h3b247177),
	.w2(32'h3b3143e0),
	.w3(32'hbad2db04),
	.w4(32'hbab1c5bb),
	.w5(32'hba7e1270),
	.w6(32'h3b29a399),
	.w7(32'h3b302bd1),
	.w8(32'h39d389b0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac89e84),
	.w1(32'hb8b31eef),
	.w2(32'hb9b72d44),
	.w3(32'hb99e7e09),
	.w4(32'h366bc326),
	.w5(32'h3959d60d),
	.w6(32'h39bc1df0),
	.w7(32'hb8ab17fe),
	.w8(32'h38938af2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f8e52),
	.w1(32'h3bcb3f1d),
	.w2(32'h3c0def88),
	.w3(32'h3ad88528),
	.w4(32'h3b525659),
	.w5(32'h3b9ec09e),
	.w6(32'h3bb4e535),
	.w7(32'h3ba4b1e0),
	.w8(32'h3b105149),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40ed34),
	.w1(32'h3b071659),
	.w2(32'h3b1ed87c),
	.w3(32'h39887ffd),
	.w4(32'h3a24d9a8),
	.w5(32'hb9e2dc02),
	.w6(32'h3b0c5f8d),
	.w7(32'h3a8c32fb),
	.w8(32'h39506d92),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae55315),
	.w1(32'h39aae8bb),
	.w2(32'hba37c457),
	.w3(32'hb93a6330),
	.w4(32'hba65c0e3),
	.w5(32'hbad212b2),
	.w6(32'hb99fb4cf),
	.w7(32'hba44804f),
	.w8(32'hbb24bc1b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95b074),
	.w1(32'hbafae720),
	.w2(32'hbb8fdea4),
	.w3(32'hbae7eace),
	.w4(32'hbafb3fae),
	.w5(32'hb9611105),
	.w6(32'h3a870872),
	.w7(32'hbaa8ac69),
	.w8(32'hbaf44c61),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f9e31),
	.w1(32'h3adf6074),
	.w2(32'h3b50b992),
	.w3(32'hbae03ae0),
	.w4(32'h39f534b6),
	.w5(32'h3ac80b21),
	.w6(32'hbab64ab0),
	.w7(32'hb8c8c428),
	.w8(32'h39dc6f45),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a999e22),
	.w1(32'h3a0758e7),
	.w2(32'h3a1cbb15),
	.w3(32'h3a5ee328),
	.w4(32'h3a0c4fd2),
	.w5(32'h3a62f489),
	.w6(32'h398bd09a),
	.w7(32'h3879878c),
	.w8(32'h3a516c8e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e62009),
	.w1(32'hbb400999),
	.w2(32'hbb42f933),
	.w3(32'h3949e25b),
	.w4(32'hbb1b878a),
	.w5(32'hbb21118d),
	.w6(32'hbb3c1bb3),
	.w7(32'hbb3b1d1e),
	.w8(32'hbacf9bea),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8121a2),
	.w1(32'h3a788c9b),
	.w2(32'h3b052f11),
	.w3(32'hbb63cd2e),
	.w4(32'h3697b417),
	.w5(32'h3a952ada),
	.w6(32'h37c55960),
	.w7(32'h39e52353),
	.w8(32'hbab057b1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeced6f),
	.w1(32'hba4212c2),
	.w2(32'hb94d3d00),
	.w3(32'hbaecf34a),
	.w4(32'hbb14a4d8),
	.w5(32'hbafacd99),
	.w6(32'h399b70de),
	.w7(32'h3b0c7764),
	.w8(32'hbb6ea606),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84bac9),
	.w1(32'hb8b0d6be),
	.w2(32'h3b697542),
	.w3(32'hbb533b07),
	.w4(32'hba80600a),
	.w5(32'h3a83a3ed),
	.w6(32'hb9f48db9),
	.w7(32'h3afe4c59),
	.w8(32'h3a71545b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2937e),
	.w1(32'hbb4c98ce),
	.w2(32'hbaeeef2b),
	.w3(32'hba8c80c3),
	.w4(32'hbac2cee8),
	.w5(32'hbb2f11ab),
	.w6(32'hbaa8171b),
	.w7(32'hb9995662),
	.w8(32'h3b3d0ff3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8532a2),
	.w1(32'h3b446fc8),
	.w2(32'h3bac55b4),
	.w3(32'h3b0ab974),
	.w4(32'h3b27ccdb),
	.w5(32'h3b56d858),
	.w6(32'h3b01d7c0),
	.w7(32'h3b6419fe),
	.w8(32'h3b49dbeb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854357),
	.w1(32'hbb027c7d),
	.w2(32'hbb030b7f),
	.w3(32'h3b3a3e8a),
	.w4(32'hbadb2b1a),
	.w5(32'hbae7ad78),
	.w6(32'hbab44388),
	.w7(32'hbb2b808e),
	.w8(32'hba789f06),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16cc28),
	.w1(32'h3b429426),
	.w2(32'h3b2c833d),
	.w3(32'hbab797d2),
	.w4(32'h3a6c6026),
	.w5(32'hb9448887),
	.w6(32'h3b0abda9),
	.w7(32'h3a60c69b),
	.w8(32'h3a2693ce),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390563d7),
	.w1(32'hbb138adc),
	.w2(32'hbb3dfebe),
	.w3(32'hbafaa309),
	.w4(32'hbac4d721),
	.w5(32'hba97fa51),
	.w6(32'hbb5e67fb),
	.w7(32'hbb06d6a5),
	.w8(32'hbb39dc39),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94b04c),
	.w1(32'h3934551a),
	.w2(32'h3b217588),
	.w3(32'hbb1453b6),
	.w4(32'hba81f5d1),
	.w5(32'h39b57ba2),
	.w6(32'h39eb3bef),
	.w7(32'h3a292c73),
	.w8(32'hbb292c96),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05674f),
	.w1(32'hbb476fc1),
	.w2(32'hbb5cb098),
	.w3(32'hbb020b9f),
	.w4(32'hbb21b52f),
	.w5(32'hbb31f70e),
	.w6(32'hbb1110ad),
	.w7(32'hbb322484),
	.w8(32'hbb05cb05),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3470ea),
	.w1(32'h3a91c59b),
	.w2(32'h3b03b06c),
	.w3(32'hbb1d106a),
	.w4(32'h3a933aef),
	.w5(32'h3a8b4f3d),
	.w6(32'h3a642dbb),
	.w7(32'h39614ab3),
	.w8(32'hbaf0a4d5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39602641),
	.w1(32'hbaf9519f),
	.w2(32'hbb21fb2e),
	.w3(32'h3979d323),
	.w4(32'hbac20931),
	.w5(32'hbb12f237),
	.w6(32'hbb000923),
	.w7(32'hbb3ccd15),
	.w8(32'hbb1e6874),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb215caa),
	.w1(32'hb98516e1),
	.w2(32'hba8a68aa),
	.w3(32'hbaf75f9b),
	.w4(32'hba345c1d),
	.w5(32'hb917bb1f),
	.w6(32'h39f01b33),
	.w7(32'hbaff40cf),
	.w8(32'hbb352d4e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64bccf),
	.w1(32'h3b8f7f8b),
	.w2(32'h3baea17d),
	.w3(32'h3b085342),
	.w4(32'h3b1547d8),
	.w5(32'h3b2ff164),
	.w6(32'h3b86aeb8),
	.w7(32'h3b970350),
	.w8(32'h3a8dc76a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6c13a),
	.w1(32'h39c1bc73),
	.w2(32'h3af829c9),
	.w3(32'h370b3e61),
	.w4(32'hbb017cee),
	.w5(32'h39f17c57),
	.w6(32'h39606412),
	.w7(32'h3ab35b3e),
	.w8(32'hb9f8485d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946adfa),
	.w1(32'hba825674),
	.w2(32'hbb2195a7),
	.w3(32'hba91b15a),
	.w4(32'h398c8da7),
	.w5(32'hb8e24b39),
	.w6(32'hba9f99a8),
	.w7(32'hba9fc35b),
	.w8(32'hba1c58b5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab286c4),
	.w1(32'hbb79557c),
	.w2(32'hbb83f0c6),
	.w3(32'h392dd65f),
	.w4(32'hbb07452e),
	.w5(32'hbab46ac8),
	.w6(32'hbb60b248),
	.w7(32'hbb4837a0),
	.w8(32'hbad59acf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96cb61),
	.w1(32'h3ad9f81c),
	.w2(32'h3aedf660),
	.w3(32'hbb174d3c),
	.w4(32'h3adee6f1),
	.w5(32'h3a9291e4),
	.w6(32'h3a6a2994),
	.w7(32'h3a670b27),
	.w8(32'h3ac6b09c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a122cbf),
	.w1(32'hbad5fd0e),
	.w2(32'h3a22c258),
	.w3(32'h3a14eabb),
	.w4(32'hbad23f91),
	.w5(32'hb9994006),
	.w6(32'hba9547b5),
	.w7(32'h390f9059),
	.w8(32'h398cae36),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd9463),
	.w1(32'h3a5271b9),
	.w2(32'hb8791f48),
	.w3(32'hb9a8f229),
	.w4(32'h3a9a3a92),
	.w5(32'hb9724676),
	.w6(32'h3aa09892),
	.w7(32'h3ab48951),
	.w8(32'hb9358b87),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9117d7),
	.w1(32'h3b46c40b),
	.w2(32'h3b817ee6),
	.w3(32'hba64936c),
	.w4(32'h39468c02),
	.w5(32'h3a6435c3),
	.w6(32'h3b27918f),
	.w7(32'h3b2491bd),
	.w8(32'hb9d5edb6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81cdff),
	.w1(32'hbb2bf6da),
	.w2(32'hbae72089),
	.w3(32'hba5f2369),
	.w4(32'hbb165e67),
	.w5(32'hbac53f45),
	.w6(32'hbb025f17),
	.w7(32'hbadb9d8d),
	.w8(32'hba845617),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba996122),
	.w1(32'hbb216f2e),
	.w2(32'hbb12c2ab),
	.w3(32'hba9fb6f1),
	.w4(32'hbb0ec87d),
	.w5(32'hbb10a1b6),
	.w6(32'hbaddb3ef),
	.w7(32'hbaf63527),
	.w8(32'hbabd0b33),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163f63),
	.w1(32'hba633a78),
	.w2(32'hba6ec4f4),
	.w3(32'hbb048850),
	.w4(32'hba1e2cc7),
	.w5(32'hba220959),
	.w6(32'h383d1599),
	.w7(32'hb946b922),
	.w8(32'h391837c1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98960a4),
	.w1(32'h3abcec2e),
	.w2(32'h3b372acd),
	.w3(32'hba0f497c),
	.w4(32'hbacdf9c4),
	.w5(32'hb9c59445),
	.w6(32'h39892a6d),
	.w7(32'h3a2f141c),
	.w8(32'hbae09580),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a97303),
	.w1(32'hbba966c3),
	.w2(32'hbc084b06),
	.w3(32'hbac6b675),
	.w4(32'hbb6e5051),
	.w5(32'hbac3030a),
	.w6(32'hbb2eb1aa),
	.w7(32'hbb37e3c1),
	.w8(32'hbac3aa95),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5330a4),
	.w1(32'hbafd4648),
	.w2(32'hbb5044a3),
	.w3(32'hb98f1c4c),
	.w4(32'hba7e3fc0),
	.w5(32'hbb06809d),
	.w6(32'hba91dac3),
	.w7(32'hbb081007),
	.w8(32'hb9deb034),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08957a),
	.w1(32'hba86367b),
	.w2(32'h392d9846),
	.w3(32'hbaac1a6a),
	.w4(32'hbade354c),
	.w5(32'hba67583e),
	.w6(32'hbb2074ab),
	.w7(32'hbae2c233),
	.w8(32'hbb1f56fc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c9e480),
	.w1(32'h3b4ae2e6),
	.w2(32'h3b2f28b1),
	.w3(32'h397c53f6),
	.w4(32'h3b43019f),
	.w5(32'h3bb33f29),
	.w6(32'h3af92a71),
	.w7(32'h3b4f640b),
	.w8(32'h3b9e88e0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b888e01),
	.w1(32'hbad47ff0),
	.w2(32'hbad222bf),
	.w3(32'h3baf2336),
	.w4(32'hbabffe92),
	.w5(32'hbaac5475),
	.w6(32'hbabd34a9),
	.w7(32'hbadbf2e6),
	.w8(32'hb9f918c5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ae03c),
	.w1(32'hbaaf76b8),
	.w2(32'hba439798),
	.w3(32'hb9ca0101),
	.w4(32'hba50947c),
	.w5(32'hbad22bb1),
	.w6(32'hba881f8d),
	.w7(32'hbaa71449),
	.w8(32'hba33db56),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55cf3e),
	.w1(32'h3a9638a6),
	.w2(32'h3b6c599d),
	.w3(32'hba899f91),
	.w4(32'hb9496e58),
	.w5(32'hba728b51),
	.w6(32'h3a948bb7),
	.w7(32'h3ad1213b),
	.w8(32'h39eade64),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8a6ac),
	.w1(32'h38ccc9f6),
	.w2(32'h3accb49b),
	.w3(32'hb9b4c434),
	.w4(32'hbacd2e39),
	.w5(32'hbaaffca2),
	.w6(32'hb98823e4),
	.w7(32'h3a837b03),
	.w8(32'h37fb31cf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90acad4),
	.w1(32'hb91e2d4e),
	.w2(32'h3b0d9ce0),
	.w3(32'hbaefaa81),
	.w4(32'h38b41052),
	.w5(32'h39ee29e6),
	.w6(32'hbaf57651),
	.w7(32'hba529975),
	.w8(32'hbaef1c62),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390845db),
	.w1(32'h3ace957e),
	.w2(32'h3aa764eb),
	.w3(32'hba1e23bd),
	.w4(32'hba406347),
	.w5(32'hbac05279),
	.w6(32'hba9bbd85),
	.w7(32'hbb00cf30),
	.w8(32'h3a07672f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98a333),
	.w1(32'hb939da3d),
	.w2(32'hb90437f1),
	.w3(32'h3b07fd36),
	.w4(32'hba2d4db0),
	.w5(32'hbaf7cace),
	.w6(32'hb9dec77a),
	.w7(32'hba9eb4c5),
	.w8(32'hba8ab176),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9cfe4),
	.w1(32'h3b0366b1),
	.w2(32'h37f85350),
	.w3(32'hbb1c9df3),
	.w4(32'h3aa77006),
	.w5(32'h3b15c3c9),
	.w6(32'h3a94183b),
	.w7(32'hb9d13a14),
	.w8(32'h3a031aca),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6af51),
	.w1(32'hba6a9d8d),
	.w2(32'hba8a10c4),
	.w3(32'h3b2b663a),
	.w4(32'hba210b95),
	.w5(32'hba8099ee),
	.w6(32'hba2ba5f7),
	.w7(32'hba77e390),
	.w8(32'hba09d90f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803926),
	.w1(32'h3b7dfa82),
	.w2(32'h3bea38d5),
	.w3(32'hba5023cc),
	.w4(32'h3b339303),
	.w5(32'h3b807f5f),
	.w6(32'h3b2eefe4),
	.w7(32'h3baadc05),
	.w8(32'h3b760f57),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bc759),
	.w1(32'hbac33aca),
	.w2(32'hbac9b251),
	.w3(32'h3b2d09f1),
	.w4(32'hba984a3d),
	.w5(32'hba5bb0de),
	.w6(32'hba9e50d0),
	.w7(32'hba89b7ef),
	.w8(32'hb7d06a5a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba961fbd),
	.w1(32'hbaabcb16),
	.w2(32'hbab474f5),
	.w3(32'hba903fa5),
	.w4(32'hba337583),
	.w5(32'hba6f9b2c),
	.w6(32'hbaa4c407),
	.w7(32'hbab6c0ff),
	.w8(32'hba9b8d0f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae4558),
	.w1(32'h3b5f93e8),
	.w2(32'h3ba43fce),
	.w3(32'hba5829cd),
	.w4(32'h3afcb6c7),
	.w5(32'h3b0e60aa),
	.w6(32'h3b722853),
	.w7(32'h3b7c75ae),
	.w8(32'h3b09832a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad443d1),
	.w1(32'h3b329a2c),
	.w2(32'h3bb0a13c),
	.w3(32'h39da9008),
	.w4(32'h3a7ed9de),
	.w5(32'h3b1a87ec),
	.w6(32'h3b29fde6),
	.w7(32'h3b826d2f),
	.w8(32'h3ac962fc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64c553),
	.w1(32'hba0534e5),
	.w2(32'h3a444457),
	.w3(32'h3acc36ae),
	.w4(32'hb6570d8e),
	.w5(32'h39f06c72),
	.w6(32'hba60103e),
	.w7(32'h38cd6574),
	.w8(32'h3ab5b083),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7abda18),
	.w1(32'h3aaa6f18),
	.w2(32'h3b395aec),
	.w3(32'h38c823b3),
	.w4(32'h39c13a37),
	.w5(32'h396d73ec),
	.w6(32'hb99d08e8),
	.w7(32'hb9606b6a),
	.w8(32'hbb159b7e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c30336),
	.w1(32'hbaf7cc5d),
	.w2(32'hbae1365c),
	.w3(32'hba58b2cb),
	.w4(32'h3b43692a),
	.w5(32'h3b961f64),
	.w6(32'hbb4c7908),
	.w7(32'hbb8e2613),
	.w8(32'hbae3f1c9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b210041),
	.w1(32'h39b7c9de),
	.w2(32'h3aba79bc),
	.w3(32'h3b931303),
	.w4(32'h3b12cbda),
	.w5(32'h3b12b75d),
	.w6(32'h3a594113),
	.w7(32'h3adafbb8),
	.w8(32'h3afc73cb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e1669),
	.w1(32'hba250ece),
	.w2(32'h3a8c2ae1),
	.w3(32'h3b4e1f14),
	.w4(32'h3a0ef358),
	.w5(32'h3b170e3d),
	.w6(32'hba8be47e),
	.w7(32'hb9fc8fe1),
	.w8(32'h3a58a31d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f3fbe),
	.w1(32'h393955e3),
	.w2(32'h3a9850a2),
	.w3(32'hbaf412ee),
	.w4(32'hbac09a2a),
	.w5(32'hba23937e),
	.w6(32'h3a71c3ae),
	.w7(32'h3aa29f13),
	.w8(32'hb9caeb9d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b5722),
	.w1(32'h3b945bb0),
	.w2(32'h3bd8bac6),
	.w3(32'hbac92dc8),
	.w4(32'h3b3cc45c),
	.w5(32'h3b56264e),
	.w6(32'h3b979c78),
	.w7(32'h3bc7d6da),
	.w8(32'h3b61a67f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920b45),
	.w1(32'hbb297edf),
	.w2(32'h39fd6770),
	.w3(32'h3b569d8d),
	.w4(32'hbba5fc3c),
	.w5(32'hbad4fc17),
	.w6(32'hb9d92ec7),
	.w7(32'hba31d15e),
	.w8(32'hbb6b292d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4dbd3),
	.w1(32'hbb90e1f0),
	.w2(32'hbadd66c4),
	.w3(32'hbb68e9e4),
	.w4(32'h3a118fb3),
	.w5(32'h3b66b942),
	.w6(32'hbb906977),
	.w7(32'hbaf71a37),
	.w8(32'h39c0408e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ea1cb),
	.w1(32'hbb4daffc),
	.w2(32'hbba289d0),
	.w3(32'h3b5b74c8),
	.w4(32'hbb0b6814),
	.w5(32'hbb637483),
	.w6(32'hbb254065),
	.w7(32'hbb8c7122),
	.w8(32'hba91ef8d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2529cf),
	.w1(32'hbb31d955),
	.w2(32'h364970c7),
	.w3(32'hbabf0e98),
	.w4(32'hbb2e752b),
	.w5(32'hba03c52d),
	.w6(32'hbb356754),
	.w7(32'hbae7115c),
	.w8(32'h3a8c108e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86bbc8),
	.w1(32'hbb0033db),
	.w2(32'hbb2d8683),
	.w3(32'hba750ea6),
	.w4(32'hba4ca584),
	.w5(32'hbae06c07),
	.w6(32'hba078c4b),
	.w7(32'hbaed4f7f),
	.w8(32'hba249c3d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5e893),
	.w1(32'hba37e268),
	.w2(32'hb9c2d6a2),
	.w3(32'hba5b7e03),
	.w4(32'hba9917fb),
	.w5(32'hba0f7cc2),
	.w6(32'hb9941eaf),
	.w7(32'hb97e626e),
	.w8(32'hb96c19d5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5850d),
	.w1(32'h3aa0af4c),
	.w2(32'h3b545f95),
	.w3(32'hba174e02),
	.w4(32'hbac2558f),
	.w5(32'hbab6514a),
	.w6(32'hba57ef5b),
	.w7(32'h3935e4a3),
	.w8(32'hbb01a460),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2a90c),
	.w1(32'hbabf8b91),
	.w2(32'hbacebd7f),
	.w3(32'hbac57bec),
	.w4(32'hb9f132bf),
	.w5(32'hba90dbe7),
	.w6(32'hba73bec1),
	.w7(32'hba97f6d4),
	.w8(32'hb9e5ac0b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5d667),
	.w1(32'hbaebb6cb),
	.w2(32'hbb08ad4e),
	.w3(32'hbae1d5b7),
	.w4(32'hba0769d5),
	.w5(32'hba64367b),
	.w6(32'hbb027084),
	.w7(32'hba8e9e7e),
	.w8(32'h3a650858),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf02d49),
	.w1(32'hbabc67d3),
	.w2(32'h39c134b3),
	.w3(32'hbb13d475),
	.w4(32'hbaeb1d18),
	.w5(32'hbaaa46e7),
	.w6(32'hba8956a9),
	.w7(32'h3996e0bc),
	.w8(32'h3aab2e56),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0bbe),
	.w1(32'hbad33838),
	.w2(32'hbae4584d),
	.w3(32'h39d5d55d),
	.w4(32'hba8729e2),
	.w5(32'hbaf2c7cf),
	.w6(32'hbaac1244),
	.w7(32'hba5530ab),
	.w8(32'hba784cab),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1677b7),
	.w1(32'hbb6dd6b3),
	.w2(32'hbb7bfa6f),
	.w3(32'hbaf69ad8),
	.w4(32'hbb1b3da1),
	.w5(32'hbaf1cbd2),
	.w6(32'hbb09f099),
	.w7(32'hbaa128de),
	.w8(32'hbaec1493),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a8527),
	.w1(32'hbaf78484),
	.w2(32'hbabd9261),
	.w3(32'h3ae1da7a),
	.w4(32'hbb3e2ee4),
	.w5(32'hbb5d415b),
	.w6(32'hba8bc0e0),
	.w7(32'hba82bbfa),
	.w8(32'hbac431bb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6fe29),
	.w1(32'hb9cba0ca),
	.w2(32'hb9ec41cd),
	.w3(32'hbad82d66),
	.w4(32'hbb3ae422),
	.w5(32'hbb232e3d),
	.w6(32'hb9c38a28),
	.w7(32'hba0334f0),
	.w8(32'hbb869057),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cda80),
	.w1(32'hba6e2388),
	.w2(32'hbb03126e),
	.w3(32'hbb6ca1fa),
	.w4(32'hbaa63f3b),
	.w5(32'hba859b29),
	.w6(32'hba18d28b),
	.w7(32'hba86547f),
	.w8(32'h3803be5a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9361de2),
	.w1(32'hbb055cc1),
	.w2(32'hbb5a5a57),
	.w3(32'hb98151a8),
	.w4(32'hba6774bd),
	.w5(32'hbb0dde20),
	.w6(32'hbabbb93b),
	.w7(32'hbb20fe83),
	.w8(32'hba2b9823),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16623b),
	.w1(32'hbb1266ab),
	.w2(32'hbb40128d),
	.w3(32'hbac1a98f),
	.w4(32'hbafc9ff5),
	.w5(32'hbb1a6b18),
	.w6(32'hbb06bfb9),
	.w7(32'hbb304a07),
	.w8(32'hbad6aa9b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd136),
	.w1(32'hbb27e9aa),
	.w2(32'hbb65f1fd),
	.w3(32'hbae98e70),
	.w4(32'hbb0ecfbf),
	.w5(32'hbb4031df),
	.w6(32'hbb192a1b),
	.w7(32'hbb3c8900),
	.w8(32'hbae27fe7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26ed2a),
	.w1(32'hbaf65a49),
	.w2(32'hbb75cd6c),
	.w3(32'hbaf97fcb),
	.w4(32'hb87880b6),
	.w5(32'hbadfe4c8),
	.w6(32'hbb21273d),
	.w7(32'hbb190631),
	.w8(32'hbb227863),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82e687),
	.w1(32'hb89c7e44),
	.w2(32'hba55b190),
	.w3(32'hba3244b6),
	.w4(32'hbad66853),
	.w5(32'hbb3311c9),
	.w6(32'hba72a4c0),
	.w7(32'hbac93f57),
	.w8(32'hbb970f68),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb59249),
	.w1(32'h399cee2c),
	.w2(32'h3a952e5f),
	.w3(32'hbb604f24),
	.w4(32'h38deeead),
	.w5(32'h386d42ef),
	.w6(32'h3a9068e5),
	.w7(32'h3b14c3ce),
	.w8(32'h3b214a00),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a6d71),
	.w1(32'hba008aa1),
	.w2(32'h3a82a5fe),
	.w3(32'h3aa6daf3),
	.w4(32'hb9a5da7b),
	.w5(32'h3a7227cc),
	.w6(32'h38b558ec),
	.w7(32'h3ac07992),
	.w8(32'h3a8be2f0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20ae41),
	.w1(32'hbb5dbbfd),
	.w2(32'hbb865990),
	.w3(32'h3a3eb241),
	.w4(32'hbb2f562d),
	.w5(32'hbb5f0844),
	.w6(32'hbb41dcb6),
	.w7(32'hbb5f47f6),
	.w8(32'hbb3434d3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb637f92),
	.w1(32'hbb438f26),
	.w2(32'hbba0f4fd),
	.w3(32'hbb3a9b60),
	.w4(32'h3afcb054),
	.w5(32'h3a1b9559),
	.w6(32'hbbd11b4c),
	.w7(32'hbbc545db),
	.w8(32'hbb9a4f5a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf96485),
	.w1(32'h3a062383),
	.w2(32'h3b1eaed3),
	.w3(32'hb99f6a52),
	.w4(32'h3968d8cc),
	.w5(32'h3ad58a47),
	.w6(32'hb92032eb),
	.w7(32'h3a86ed9d),
	.w8(32'h3b0000b8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a50da),
	.w1(32'hbaa44d11),
	.w2(32'hbabed641),
	.w3(32'h3b021ed7),
	.w4(32'hba8618dc),
	.w5(32'hbaa020f8),
	.w6(32'hba83a3a9),
	.w7(32'hbaa54acf),
	.w8(32'hb9fedc9b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba609db1),
	.w1(32'hb7bcb2d8),
	.w2(32'hb7807310),
	.w3(32'hba23177b),
	.w4(32'h384da006),
	.w5(32'h37d59e5a),
	.w6(32'hb7e9a0b2),
	.w7(32'h38044130),
	.w8(32'h37f331e7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38f8f7),
	.w1(32'hb8ce4495),
	.w2(32'h398542f9),
	.w3(32'hb958d436),
	.w4(32'hb9a71fc1),
	.w5(32'hb916528c),
	.w6(32'hb7474679),
	.w7(32'hb984afef),
	.w8(32'hb95e97d2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a475d5),
	.w1(32'h399aea57),
	.w2(32'h3a0850da),
	.w3(32'hb91a3cc6),
	.w4(32'h393e166a),
	.w5(32'h390e52e1),
	.w6(32'h3981cfab),
	.w7(32'h39ec34f0),
	.w8(32'h39cc867d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb860dd0c),
	.w1(32'hb8640d68),
	.w2(32'hb746883e),
	.w3(32'hb887608f),
	.w4(32'hb7fc75ff),
	.w5(32'h375cdf61),
	.w6(32'hb812ba79),
	.w7(32'hb743ea73),
	.w8(32'h38051d6b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37838927),
	.w1(32'h395ffcf1),
	.w2(32'h39774957),
	.w3(32'h39449500),
	.w4(32'h38f64c4d),
	.w5(32'h393a54e0),
	.w6(32'h38cecbfb),
	.w7(32'hb7f2922a),
	.w8(32'h37c729e4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70d9f96),
	.w1(32'hb7479703),
	.w2(32'hb828b3d6),
	.w3(32'h371e5f20),
	.w4(32'h378c0739),
	.w5(32'hb7474b5c),
	.w6(32'hb80bb670),
	.w7(32'hb74cfd12),
	.w8(32'hb79a9a48),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94712e5),
	.w1(32'h39592db8),
	.w2(32'h39c35e57),
	.w3(32'hb8603aa8),
	.w4(32'h3988c3fc),
	.w5(32'h39ba2d32),
	.w6(32'h3618afdd),
	.w7(32'h398fe2b7),
	.w8(32'h39cd6bb4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a2b136),
	.w1(32'h392f8b67),
	.w2(32'h3838cc2a),
	.w3(32'h3883a0ef),
	.w4(32'h39274f30),
	.w5(32'hb861be5a),
	.w6(32'hb75e6d5f),
	.w7(32'h38a6f4c7),
	.w8(32'hb7f6bbec),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f3fc7),
	.w1(32'hb94dabd2),
	.w2(32'h393f56c4),
	.w3(32'hb983ff6f),
	.w4(32'hb8a18ce9),
	.w5(32'h39c4d3b3),
	.w6(32'h390be751),
	.w7(32'h3906d028),
	.w8(32'h39ff149b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3693f27c),
	.w1(32'h369ec90a),
	.w2(32'hb843a606),
	.w3(32'h388e08e3),
	.w4(32'h382b3620),
	.w5(32'hb87d3977),
	.w6(32'hb88c65d7),
	.w7(32'hb80f6dcf),
	.w8(32'hb8901388),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90620bd),
	.w1(32'hb94ce164),
	.w2(32'h38e4e749),
	.w3(32'hb9914149),
	.w4(32'h3875f617),
	.w5(32'h382b06e3),
	.w6(32'hb922f158),
	.w7(32'hb77951d4),
	.w8(32'h3979c985),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1548c5),
	.w1(32'hba0c3d7e),
	.w2(32'hb9982153),
	.w3(32'hb9c31407),
	.w4(32'hb9b9c3d6),
	.w5(32'hb71dc0b6),
	.w6(32'hb9302e6b),
	.w7(32'hb923fc6e),
	.w8(32'h38109634),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38efa46f),
	.w1(32'hb92da1d2),
	.w2(32'hb99478d5),
	.w3(32'h3938d101),
	.w4(32'hb8c6637e),
	.w5(32'hb9bfa352),
	.w6(32'hb885721e),
	.w7(32'hb95f5710),
	.w8(32'hb9d9009e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39861f1d),
	.w1(32'h392ffc20),
	.w2(32'h39b583d1),
	.w3(32'h39a0d824),
	.w4(32'h39006407),
	.w5(32'h38f55d29),
	.w6(32'h39a697c4),
	.w7(32'h38eb5dc9),
	.w8(32'h39ba0141),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384b5ae3),
	.w1(32'h3787f2ae),
	.w2(32'h3698f376),
	.w3(32'h38499b2d),
	.w4(32'h3882b995),
	.w5(32'h3840aef7),
	.w6(32'h38a4552d),
	.w7(32'h38d25715),
	.w8(32'h38eefc1f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98306a1),
	.w1(32'h399e998d),
	.w2(32'h3939806b),
	.w3(32'h3768def8),
	.w4(32'h39e26836),
	.w5(32'h3720bbca),
	.w6(32'hb8703835),
	.w7(32'h39de7b1e),
	.w8(32'hb57ed2d5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93bab5f),
	.w1(32'hb8db7870),
	.w2(32'hb9711ad4),
	.w3(32'hb7b7b8d2),
	.w4(32'hb751a7ea),
	.w5(32'hb9a4e9e4),
	.w6(32'h38ce7a12),
	.w7(32'h38ad19c9),
	.w8(32'hb819cf33),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8013aa3),
	.w1(32'hb7a484c1),
	.w2(32'h368a259f),
	.w3(32'hb623e768),
	.w4(32'hb7daa2de),
	.w5(32'hb760c164),
	.w6(32'hb80d50ab),
	.w7(32'hb7d6bec2),
	.w8(32'hb7b68914),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ce3359),
	.w1(32'h3729f979),
	.w2(32'hb40917de),
	.w3(32'hb6e2976a),
	.w4(32'h362cdb19),
	.w5(32'hb5fa1f7b),
	.w6(32'h35b8c1f1),
	.w7(32'h37486ddb),
	.w8(32'h37336182),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8127a31),
	.w1(32'hb7971b07),
	.w2(32'hb71513b6),
	.w3(32'hb60bc4d0),
	.w4(32'hb55111f3),
	.w5(32'h384a9928),
	.w6(32'h34bbccaf),
	.w7(32'h37ee2999),
	.w8(32'h382868a0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971993f),
	.w1(32'hb9950608),
	.w2(32'hb9431ef6),
	.w3(32'hb96bebad),
	.w4(32'hb93d647c),
	.w5(32'hb901b1fc),
	.w6(32'hb9ac8e37),
	.w7(32'hb96308ee),
	.w8(32'hb97aa79e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a62ed),
	.w1(32'hb91a27fd),
	.w2(32'hb8452cd6),
	.w3(32'hb93ea118),
	.w4(32'hb8756dcc),
	.w5(32'h38adf4e9),
	.w6(32'hb912d1fe),
	.w7(32'hb7405557),
	.w8(32'h3910d504),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3733eec9),
	.w1(32'h37a26a93),
	.w2(32'h37afe049),
	.w3(32'h375640a3),
	.w4(32'h3793c6c4),
	.w5(32'h37eb1ce7),
	.w6(32'h380a7705),
	.w7(32'h37d27e1e),
	.w8(32'h38042900),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38407c5d),
	.w1(32'h384cb067),
	.w2(32'h3802d0b0),
	.w3(32'h38a509f1),
	.w4(32'h388b0aa1),
	.w5(32'h37275ea9),
	.w6(32'h398f80a8),
	.w7(32'h399ea8ae),
	.w8(32'h39b04eee),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ac6c5),
	.w1(32'hb996f992),
	.w2(32'h398731db),
	.w3(32'hba2f5cab),
	.w4(32'h3a065c43),
	.w5(32'h3a4bd509),
	.w6(32'hb9436900),
	.w7(32'h3a396a72),
	.w8(32'h3a7a01d2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962471b),
	.w1(32'h396635fe),
	.w2(32'h390e62b8),
	.w3(32'h39c3000a),
	.w4(32'h39a28613),
	.w5(32'h39e9c4e2),
	.w6(32'h3a001f72),
	.w7(32'h39e024a9),
	.w8(32'h394ea58e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f9e7a),
	.w1(32'h38a60e5a),
	.w2(32'hb9817c47),
	.w3(32'hb91fd71c),
	.w4(32'h3a02f893),
	.w5(32'h38752170),
	.w6(32'hb8719736),
	.w7(32'h39d9ab54),
	.w8(32'h39a0b80d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f14214),
	.w1(32'hba088084),
	.w2(32'hb9708e67),
	.w3(32'hb9d65306),
	.w4(32'hb9b729cc),
	.w5(32'hb9536839),
	.w6(32'hb9ff5345),
	.w7(32'hb9062b4c),
	.w8(32'h39dd0298),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82a80b),
	.w1(32'h39c669f4),
	.w2(32'h39b36644),
	.w3(32'hba88d884),
	.w4(32'hb9912276),
	.w5(32'h39d66ac2),
	.w6(32'hbaade1a2),
	.w7(32'hb79fb809),
	.w8(32'h3aa86fdb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab33cb2),
	.w1(32'h3a56855a),
	.w2(32'h3984c34a),
	.w3(32'h3a8918f0),
	.w4(32'h39ed8369),
	.w5(32'h38420618),
	.w6(32'h3a02615d),
	.w7(32'h39ddc964),
	.w8(32'h38aa53fb),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a82857),
	.w1(32'hb91e9fc6),
	.w2(32'hb9c21ffa),
	.w3(32'hb900e1ad),
	.w4(32'hb97eda92),
	.w5(32'hba03e825),
	.w6(32'hb9289b6d),
	.w7(32'hb9b32a1a),
	.w8(32'hba330b9e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935dd25),
	.w1(32'hb9859042),
	.w2(32'hb9a60f65),
	.w3(32'h37507557),
	.w4(32'hb8a5ab47),
	.w5(32'hb917ab58),
	.w6(32'hb80f1e42),
	.w7(32'hb9576d8d),
	.w8(32'hb9959fce),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89649f7),
	.w1(32'hb8b4be3f),
	.w2(32'hb766b925),
	.w3(32'hb87d07f9),
	.w4(32'hb783402c),
	.w5(32'h382303b3),
	.w6(32'hb7141924),
	.w7(32'h37a2b403),
	.w8(32'h385dc419),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fa0672),
	.w1(32'h33dc1e59),
	.w2(32'h371ab300),
	.w3(32'hb6627f52),
	.w4(32'h361e7895),
	.w5(32'h3710fc03),
	.w6(32'h36965844),
	.w7(32'hb6804319),
	.w8(32'h372ca741),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882e866),
	.w1(32'h38fac179),
	.w2(32'h399324b1),
	.w3(32'h388eb510),
	.w4(32'h3842b5eb),
	.w5(32'h393cebb5),
	.w6(32'h398b07d5),
	.w7(32'h397c575b),
	.w8(32'h39bf4f89),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8beed64),
	.w1(32'hb8c08a9d),
	.w2(32'hb8be1261),
	.w3(32'hb8e9401b),
	.w4(32'hb912db66),
	.w5(32'hb89d40b1),
	.w6(32'hb8ded812),
	.w7(32'hb91c64d7),
	.w8(32'hb916825b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c31a2),
	.w1(32'h3991b49f),
	.w2(32'h38bc9c32),
	.w3(32'h39a965d0),
	.w4(32'h39a0f0e2),
	.w5(32'hb8b17d26),
	.w6(32'h3986f462),
	.w7(32'h38bd2a5c),
	.w8(32'h38f10bad),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f2add),
	.w1(32'hb99ccdf3),
	.w2(32'hb9b35cb7),
	.w3(32'h38c40766),
	.w4(32'hb97d2d7a),
	.w5(32'hb9abdc64),
	.w6(32'h388620d9),
	.w7(32'hb9ad2650),
	.w8(32'hb9b556f4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e985af),
	.w1(32'h38f2d3f1),
	.w2(32'h39204253),
	.w3(32'hb89671dc),
	.w4(32'h38d8c317),
	.w5(32'h397dc753),
	.w6(32'hb8815150),
	.w7(32'h39012630),
	.w8(32'h395d1ef0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f3d02),
	.w1(32'hb8d17bd4),
	.w2(32'hb902fdd7),
	.w3(32'hb8d27314),
	.w4(32'hb91428bd),
	.w5(32'hb94d7fd8),
	.w6(32'hb9842b76),
	.w7(32'hb9a31c3e),
	.w8(32'hb919e327),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9b877),
	.w1(32'hb8a5614c),
	.w2(32'h3908001c),
	.w3(32'hb9917d53),
	.w4(32'hb8fdcb31),
	.w5(32'h38f52637),
	.w6(32'hb9233529),
	.w7(32'hb80ae943),
	.w8(32'hb80ddcfb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a368191),
	.w1(32'h39f8f449),
	.w2(32'h39bf0087),
	.w3(32'h3a4920dd),
	.w4(32'h39aaf2c5),
	.w5(32'hb8031c07),
	.w6(32'h399c390d),
	.w7(32'hb90efffd),
	.w8(32'hb8fc8e93),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a113c10),
	.w1(32'h3a953da1),
	.w2(32'hb61e6944),
	.w3(32'h3a64800c),
	.w4(32'h395bb28e),
	.w5(32'hb9eeecb4),
	.w6(32'h3a9147a6),
	.w7(32'h3a10beb0),
	.w8(32'hb8eeaa27),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ab1d2),
	.w1(32'hba4e63e2),
	.w2(32'hb9664893),
	.w3(32'hba248883),
	.w4(32'hba1ce7b7),
	.w5(32'hb8ca3503),
	.w6(32'hba6adb94),
	.w7(32'hba7c000d),
	.w8(32'hba4f0f1f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba523be4),
	.w1(32'hba0e8b2e),
	.w2(32'hba40e974),
	.w3(32'hb9462658),
	.w4(32'hb9df70ac),
	.w5(32'hba66cbbc),
	.w6(32'h38f9f820),
	.w7(32'hb9336027),
	.w8(32'hba0670a0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f2378),
	.w1(32'hb840292b),
	.w2(32'hb90428a1),
	.w3(32'hb89aa332),
	.w4(32'h387041c1),
	.w5(32'hb79ec7f4),
	.w6(32'hb8bc4d0d),
	.w7(32'h37c21927),
	.w8(32'hb81c3766),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9270be7),
	.w1(32'h394d8228),
	.w2(32'h375e4727),
	.w3(32'h37a4547d),
	.w4(32'h39c30c40),
	.w5(32'hb91aafc9),
	.w6(32'h39ca644a),
	.w7(32'hb8247565),
	.w8(32'hb73a7c57),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3874bb33),
	.w1(32'h393025b4),
	.w2(32'h39ff7e8f),
	.w3(32'h389222db),
	.w4(32'h39783ef4),
	.w5(32'h3a1b5e55),
	.w6(32'h39494027),
	.w7(32'h395172ff),
	.w8(32'h39e2cfa3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a010fa7),
	.w1(32'h39648ad2),
	.w2(32'hb8c10aba),
	.w3(32'h39a7007c),
	.w4(32'hb91f6ebf),
	.w5(32'h393872ae),
	.w6(32'h39a582f0),
	.w7(32'h395fee8c),
	.w8(32'h3a39e824),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dcb9b2),
	.w1(32'hba222833),
	.w2(32'hb9e3a34f),
	.w3(32'hb9af56fa),
	.w4(32'hba708bec),
	.w5(32'hba644f06),
	.w6(32'hba254ead),
	.w7(32'hba9dcbdf),
	.w8(32'hba63e3ac),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad6003),
	.w1(32'h39ea5a70),
	.w2(32'hb8fd839f),
	.w3(32'h39c59be4),
	.w4(32'h39287bd3),
	.w5(32'hb9699ba2),
	.w6(32'h3a197757),
	.w7(32'h391b1d17),
	.w8(32'hb90480af),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77116ab),
	.w1(32'hb65d3379),
	.w2(32'h3540b64f),
	.w3(32'hb7879416),
	.w4(32'hb59385d5),
	.w5(32'h3567f808),
	.w6(32'hb72b7601),
	.w7(32'h3677e45b),
	.w8(32'h3702c2a7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a73c71),
	.w1(32'hb86a3e5d),
	.w2(32'hb8852740),
	.w3(32'hb6b10b69),
	.w4(32'h367a2eaf),
	.w5(32'h3708baa5),
	.w6(32'hb8ba796a),
	.w7(32'hb77ce234),
	.w8(32'hb8462e06),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5483d),
	.w1(32'hb902a313),
	.w2(32'hb8dc94dc),
	.w3(32'h380e7581),
	.w4(32'h3733e6be),
	.w5(32'hb802391f),
	.w6(32'h38469934),
	.w7(32'hb8125e44),
	.w8(32'hb8d02933),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7af4c91),
	.w1(32'h37d62058),
	.w2(32'h38d5ece5),
	.w3(32'h36496da0),
	.w4(32'h3939f6d8),
	.w5(32'h39975c4f),
	.w6(32'h388ed3ad),
	.w7(32'h38f85e7e),
	.w8(32'h399c1fd3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb785fcd9),
	.w1(32'h3703982f),
	.w2(32'hb675e2ae),
	.w3(32'hb74c206c),
	.w4(32'h37034a1d),
	.w5(32'h3610797f),
	.w6(32'h36895acd),
	.w7(32'h34a2aa73),
	.w8(32'h35941e5e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375ba3d7),
	.w1(32'h37878b28),
	.w2(32'h38327a36),
	.w3(32'hb8aaabcd),
	.w4(32'hb8e02fc1),
	.w5(32'hb7f2cef6),
	.w6(32'hb91ba610),
	.w7(32'hb888edc6),
	.w8(32'h385106dc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85bc62a),
	.w1(32'h38a486e4),
	.w2(32'h37e202d9),
	.w3(32'h37830312),
	.w4(32'h38d04874),
	.w5(32'h35279316),
	.w6(32'h36bda102),
	.w7(32'h3890c4f5),
	.w8(32'h387d6d72),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba043fbc),
	.w1(32'hba0f0b9c),
	.w2(32'hb9b1bcfd),
	.w3(32'hba04ba95),
	.w4(32'hb9ba660f),
	.w5(32'hb89517df),
	.w6(32'hb9ea8e9a),
	.w7(32'hb997b289),
	.w8(32'hb860302e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a47964),
	.w1(32'hb8a533af),
	.w2(32'hb8fa2cda),
	.w3(32'h3920521c),
	.w4(32'hb8792ae3),
	.w5(32'hb900c78b),
	.w6(32'hb7f736ae),
	.w7(32'hb5cca0c6),
	.w8(32'hb891a878),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a4ca3),
	.w1(32'hb920d741),
	.w2(32'hb91c7ee3),
	.w3(32'hb8d8502f),
	.w4(32'hb8acc30e),
	.w5(32'hb920b855),
	.w6(32'hb952b59c),
	.w7(32'hb976053e),
	.w8(32'hb9a1b924),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba030fea),
	.w1(32'hb9b63d77),
	.w2(32'h3a545de2),
	.w3(32'hba6f191d),
	.w4(32'hba223b9d),
	.w5(32'h3a27265f),
	.w6(32'hb9b34d87),
	.w7(32'h39ac2697),
	.w8(32'h3ab98da9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac9a17),
	.w1(32'h3a129e70),
	.w2(32'hba00dbe7),
	.w3(32'h3a4387b4),
	.w4(32'h39af09e9),
	.w5(32'hb995a07c),
	.w6(32'h39f29df6),
	.w7(32'h3905bf22),
	.w8(32'h38c1f7d5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983c28d),
	.w1(32'hb863cc4a),
	.w2(32'h38400198),
	.w3(32'hb8e97ce7),
	.w4(32'hb9653a5d),
	.w5(32'h378bbc1a),
	.w6(32'hb99d4f45),
	.w7(32'hb9c73f7e),
	.w8(32'hb93b21fb),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380c8bd2),
	.w1(32'h38012e99),
	.w2(32'h36dec379),
	.w3(32'h3786cb46),
	.w4(32'h37abb97b),
	.w5(32'h374f4080),
	.w6(32'h371eb42b),
	.w7(32'h36d41022),
	.w8(32'h37098ea5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e677f1),
	.w1(32'h38e8b5d8),
	.w2(32'h381e9827),
	.w3(32'hb930624d),
	.w4(32'hb90bac9b),
	.w5(32'h3847c2b0),
	.w6(32'hb962d38f),
	.w7(32'h38fc143b),
	.w8(32'h399f4f5f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807d71c),
	.w1(32'hb7953086),
	.w2(32'h3683cdcf),
	.w3(32'hb7bd6caf),
	.w4(32'hb72a7652),
	.w5(32'h36d69103),
	.w6(32'h37c3014c),
	.w7(32'h37fe858f),
	.w8(32'h372967d8),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9810543),
	.w1(32'hb9489fa0),
	.w2(32'hb92348f3),
	.w3(32'hb915ca8d),
	.w4(32'hb94d4901),
	.w5(32'hb87a9997),
	.w6(32'hb8a34848),
	.w7(32'h3772f649),
	.w8(32'h3834ec2a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8962684),
	.w1(32'hb825708e),
	.w2(32'h38c738a8),
	.w3(32'h382b2302),
	.w4(32'hb936a425),
	.w5(32'hb88c6868),
	.w6(32'h38d910e1),
	.w7(32'hb9f07e89),
	.w8(32'hba08a9ec),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3935688f),
	.w1(32'h395d5f74),
	.w2(32'h379a1868),
	.w3(32'h3974e234),
	.w4(32'h3942ac59),
	.w5(32'hb7d97cbd),
	.w6(32'hb4217eb0),
	.w7(32'h392c8d50),
	.w8(32'h389874e3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39276e61),
	.w1(32'h377b636c),
	.w2(32'hb991793d),
	.w3(32'h3947356e),
	.w4(32'h38c35ab3),
	.w5(32'hb9986e46),
	.w6(32'h390577a0),
	.w7(32'h36f9a642),
	.w8(32'hb9991b7c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10c99e),
	.w1(32'hb9f7879d),
	.w2(32'h39896628),
	.w3(32'hba0cf757),
	.w4(32'hb94dc9ca),
	.w5(32'h399a6aa8),
	.w6(32'hb98b74d3),
	.w7(32'h3951e8e5),
	.w8(32'h39d7e7c4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98196fd),
	.w1(32'hb7cacadc),
	.w2(32'hb894ef79),
	.w3(32'hb9366d66),
	.w4(32'hb830d547),
	.w5(32'hb94ccd3c),
	.w6(32'hb91e92bb),
	.w7(32'hb993ca2c),
	.w8(32'hb9cf8303),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37303335),
	.w1(32'h36a7fed5),
	.w2(32'hb5c08914),
	.w3(32'h37209b3c),
	.w4(32'hb63b3ab0),
	.w5(32'hb71ec555),
	.w6(32'h3728d7ee),
	.w7(32'hb5f4468a),
	.w8(32'hb6899a36),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36697ec0),
	.w1(32'h391ff875),
	.w2(32'h395906b9),
	.w3(32'hb88393bd),
	.w4(32'h391bcc23),
	.w5(32'h397602fb),
	.w6(32'h380876ad),
	.w7(32'h38dca7bd),
	.w8(32'h39885809),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ef17e2),
	.w1(32'h378e376b),
	.w2(32'h37b55697),
	.w3(32'hb6213f6e),
	.w4(32'h36bd010b),
	.w5(32'h36fd82d6),
	.w6(32'h37304b1b),
	.w7(32'h37a5d3c9),
	.w8(32'h378a1afe),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9603907),
	.w1(32'hb8d1e667),
	.w2(32'hb84a2415),
	.w3(32'hb8cf88d9),
	.w4(32'hb5c37418),
	.w5(32'h38bf305d),
	.w6(32'hb8a1a228),
	.w7(32'hb6c0e629),
	.w8(32'h38c6cf61),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987c0ea),
	.w1(32'h39906c0d),
	.w2(32'hb8219859),
	.w3(32'h3a2bb936),
	.w4(32'h3a0ca61c),
	.w5(32'h38a2a8e7),
	.w6(32'h3a2da998),
	.w7(32'h3a0a55aa),
	.w8(32'h37c8f078),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980c786),
	.w1(32'hb9810d05),
	.w2(32'hb973a565),
	.w3(32'hb8993cac),
	.w4(32'hb902e730),
	.w5(32'hb8c83891),
	.w6(32'hb8e10c87),
	.w7(32'hb93bbc38),
	.w8(32'hb9176028),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d578b2),
	.w1(32'hb93ee153),
	.w2(32'hb9b326f4),
	.w3(32'hb87805c2),
	.w4(32'hb91535a2),
	.w5(32'hb98091ca),
	.w6(32'hb94ce88d),
	.w7(32'hb985084f),
	.w8(32'hb9bc0517),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9068259),
	.w1(32'hb5a9264c),
	.w2(32'hb974fb2f),
	.w3(32'h37616323),
	.w4(32'h38656419),
	.w5(32'hb8c3eb06),
	.w6(32'hb916689c),
	.w7(32'hb906e0c9),
	.w8(32'hb8dcff01),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37220903),
	.w1(32'hb849864f),
	.w2(32'h396a6147),
	.w3(32'hb90e41b4),
	.w4(32'hb828941a),
	.w5(32'h371c2d05),
	.w6(32'hb8420cc3),
	.w7(32'h36d720c9),
	.w8(32'h392bb551),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e023b3),
	.w1(32'h38ed3d20),
	.w2(32'hb999ee6d),
	.w3(32'h3a5cf48e),
	.w4(32'h39962f3c),
	.w5(32'hb99c08e8),
	.w6(32'h3a7ea7ae),
	.w7(32'h3986a62b),
	.w8(32'hb9a8eb31),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ada05),
	.w1(32'hb8071f66),
	.w2(32'hb5854d0f),
	.w3(32'hb830836c),
	.w4(32'hb816898b),
	.w5(32'h36b27e4d),
	.w6(32'hb83d7306),
	.w7(32'hb85ccb43),
	.w8(32'hb7a4986d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79044dd),
	.w1(32'hb53a24ba),
	.w2(32'hb6747ce1),
	.w3(32'hb73167d5),
	.w4(32'h36d7d55e),
	.w5(32'h36ba1460),
	.w6(32'hb6375bce),
	.w7(32'hb6a9d514),
	.w8(32'h35b45b88),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e389f3),
	.w1(32'hb873d187),
	.w2(32'h379f6e3a),
	.w3(32'h396ee73a),
	.w4(32'hb8e14fcf),
	.w5(32'h38bf5b90),
	.w6(32'h38d34fb2),
	.w7(32'hb91eafb8),
	.w8(32'h346883c8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941c641),
	.w1(32'h3944325b),
	.w2(32'h39b255b4),
	.w3(32'h39860ff0),
	.w4(32'h396e2592),
	.w5(32'h39277f5a),
	.w6(32'h3a06c236),
	.w7(32'h3987ba5a),
	.w8(32'h3997cb66),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de2275),
	.w1(32'h3a355e2b),
	.w2(32'h3a243f87),
	.w3(32'h3a34ee91),
	.w4(32'h3a46dcd8),
	.w5(32'h39e81924),
	.w6(32'h3a22295d),
	.w7(32'h3a319833),
	.w8(32'h399e74b0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99afa89),
	.w1(32'hb91d0946),
	.w2(32'h380733fe),
	.w3(32'hb99402b1),
	.w4(32'hb8d528c2),
	.w5(32'h39aca2b4),
	.w6(32'hb80a06bf),
	.w7(32'hb67bca78),
	.w8(32'h38dc022d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c8a758),
	.w1(32'h37c2d603),
	.w2(32'h38949436),
	.w3(32'hb7f50386),
	.w4(32'h37e91a76),
	.w5(32'h389f4232),
	.w6(32'h36676278),
	.w7(32'h38892bb6),
	.w8(32'h389ce76f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb829cf3b),
	.w1(32'h387fc7ec),
	.w2(32'h3931db1d),
	.w3(32'h37ace190),
	.w4(32'h37dbf72a),
	.w5(32'h38f294e9),
	.w6(32'h391f4ed2),
	.w7(32'h385e5c89),
	.w8(32'h3871e46e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9849bdc),
	.w1(32'hb9b55d3b),
	.w2(32'hba02e75f),
	.w3(32'hb7df5297),
	.w4(32'hb9d74e9a),
	.w5(32'hb9c46b56),
	.w6(32'hb667152f),
	.w7(32'hb9027c3e),
	.w8(32'hb9104da9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea7ce8),
	.w1(32'hb9372321),
	.w2(32'h397f13b7),
	.w3(32'hb96c83e9),
	.w4(32'h388a5c72),
	.w5(32'h39db2277),
	.w6(32'h39828e6f),
	.w7(32'h39502bbd),
	.w8(32'h39fe6756),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb930afdb),
	.w1(32'hb949bc0b),
	.w2(32'hb8368440),
	.w3(32'hb93698ea),
	.w4(32'hb98edbbd),
	.w5(32'h3881c7b3),
	.w6(32'hb8b3f608),
	.w7(32'hb896ecc8),
	.w8(32'h38a69c7e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8922f2a),
	.w1(32'hb920e1ac),
	.w2(32'hb99f6379),
	.w3(32'h3903b4b3),
	.w4(32'hb7166eaa),
	.w5(32'hb90e0f6c),
	.w6(32'hb89585af),
	.w7(32'hb92cc039),
	.w8(32'hb9605dad),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ca0a6),
	.w1(32'h397c4093),
	.w2(32'h38711a34),
	.w3(32'h3972971c),
	.w4(32'h39ad254b),
	.w5(32'h393f9382),
	.w6(32'h38c84fcc),
	.w7(32'h39784058),
	.w8(32'h39cac7a7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b14a90),
	.w1(32'hb6ed6ce6),
	.w2(32'hb6f00379),
	.w3(32'hb72027d0),
	.w4(32'hb6bfeca8),
	.w5(32'hb6b42a05),
	.w6(32'h361d75e1),
	.w7(32'hb6a0cd5f),
	.w8(32'hb6f3103b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3651023f),
	.w1(32'h35c04b13),
	.w2(32'hb6b769bf),
	.w3(32'h3633dd78),
	.w4(32'hb677b227),
	.w5(32'hb6bb9880),
	.w6(32'h36869f23),
	.w7(32'h36516801),
	.w8(32'hb61d6687),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e10a5d),
	.w1(32'h3841c1b0),
	.w2(32'h38ab7cfa),
	.w3(32'hb855f9f7),
	.w4(32'hb583aa68),
	.w5(32'h388b448a),
	.w6(32'hb7750c0c),
	.w7(32'h37c7ae59),
	.w8(32'h38b45b48),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37297872),
	.w1(32'h35f90972),
	.w2(32'hb783abea),
	.w3(32'hb64ff4b6),
	.w4(32'hb6c54085),
	.w5(32'hb6c9b313),
	.w6(32'hb7206c7e),
	.w7(32'hb78dbad8),
	.w8(32'hb607495f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8afd1a6),
	.w1(32'hb91739e0),
	.w2(32'hb8fe12dc),
	.w3(32'hb868ca31),
	.w4(32'hb95dd0a2),
	.w5(32'hb8e6637b),
	.w6(32'hb81555e1),
	.w7(32'hb928ae1d),
	.w8(32'hb93bc0b8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb874e703),
	.w1(32'h396f260b),
	.w2(32'h3a6b1b9c),
	.w3(32'h3a0cb5b9),
	.w4(32'h3a4897b9),
	.w5(32'h3a2fb9c9),
	.w6(32'h3a8cbe2a),
	.w7(32'h3a39fa98),
	.w8(32'h3a5e27ae),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392bd00b),
	.w1(32'h38db97b1),
	.w2(32'h38bf1840),
	.w3(32'h399a3e7f),
	.w4(32'h39706b2b),
	.w5(32'h38dab639),
	.w6(32'h3991b2e1),
	.w7(32'h39455e84),
	.w8(32'h391d800c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370bbf46),
	.w1(32'h37221033),
	.w2(32'hb6f09536),
	.w3(32'hb704687a),
	.w4(32'h36dd1d6d),
	.w5(32'hb796e19d),
	.w6(32'hb796e567),
	.w7(32'h35d41727),
	.w8(32'hb69d0b8b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960aca2),
	.w1(32'h389f390b),
	.w2(32'h39b6cffd),
	.w3(32'h394d26f2),
	.w4(32'hb900fc6d),
	.w5(32'h39a8129d),
	.w6(32'h39b6a765),
	.w7(32'h37ea8f5e),
	.w8(32'h39d021ec),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b2e03b),
	.w1(32'h384a2676),
	.w2(32'hb73435af),
	.w3(32'h386db445),
	.w4(32'h38e9f759),
	.w5(32'h37a43296),
	.w6(32'h3952315a),
	.w7(32'h3977b015),
	.w8(32'h386f5533),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366b6a4b),
	.w1(32'h36c6bf75),
	.w2(32'h36b94d50),
	.w3(32'h36378e8f),
	.w4(32'h369f22d7),
	.w5(32'h364d62c2),
	.w6(32'h36139421),
	.w7(32'h368aea8a),
	.w8(32'h36f44013),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f5d74),
	.w1(32'hb8f8d82e),
	.w2(32'hb90e717f),
	.w3(32'h373c8586),
	.w4(32'hb8fb1eb3),
	.w5(32'h37a0c1ee),
	.w6(32'h3885a7c9),
	.w7(32'hb93f29ff),
	.w8(32'hb86f054f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9823563),
	.w1(32'hb9520fa7),
	.w2(32'hb90b60cc),
	.w3(32'hb990b0e6),
	.w4(32'hb97d3773),
	.w5(32'hb8cdb208),
	.w6(32'hb948f5a4),
	.w7(32'hb8be7339),
	.w8(32'h381e7df2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f5df3f),
	.w1(32'h38b239fd),
	.w2(32'hb86995bd),
	.w3(32'h38dcd21e),
	.w4(32'hb8a94881),
	.w5(32'hb7e70fd0),
	.w6(32'hb66971af),
	.w7(32'hb93c8847),
	.w8(32'hb8bafd21),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36acc584),
	.w1(32'h3638d114),
	.w2(32'h36b9ebbf),
	.w3(32'h35fcb01e),
	.w4(32'hb5ee292b),
	.w5(32'h364042c3),
	.w6(32'h37020706),
	.w7(32'hb6527e78),
	.w8(32'h36e144d8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e57818),
	.w1(32'hb7bde2bb),
	.w2(32'hb7276ca9),
	.w3(32'hb6db94e6),
	.w4(32'hb6bf6cdf),
	.w5(32'h36c246b1),
	.w6(32'h35e25803),
	.w7(32'hb72cf453),
	.w8(32'h369dcdd3),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934a45a),
	.w1(32'hb9730e02),
	.w2(32'hb99bc937),
	.w3(32'hb806bc08),
	.w4(32'hb8805706),
	.w5(32'hb9033ad4),
	.w6(32'hb9003785),
	.w7(32'hb9000ca8),
	.w8(32'hb93d61eb),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cd1337),
	.w1(32'h394380ea),
	.w2(32'h392d8e9d),
	.w3(32'h38f61414),
	.w4(32'h3928114e),
	.w5(32'h393bf31e),
	.w6(32'h396e2de9),
	.w7(32'h3901dae4),
	.w8(32'h399e3629),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c94115),
	.w1(32'h391b8536),
	.w2(32'h38ac0b3e),
	.w3(32'h3841a8fc),
	.w4(32'h37da71ce),
	.w5(32'h3927318c),
	.w6(32'h38c9de13),
	.w7(32'h374491c4),
	.w8(32'h3911fd08),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a0f09),
	.w1(32'h39cbf269),
	.w2(32'h39a4581a),
	.w3(32'h39760c42),
	.w4(32'h39e65727),
	.w5(32'h39819fca),
	.w6(32'h39f62000),
	.w7(32'h39887319),
	.w8(32'h3909c912),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b9d1c),
	.w1(32'hb8dd41ee),
	.w2(32'hb946fe5d),
	.w3(32'hb7f301ca),
	.w4(32'hb8155703),
	.w5(32'hb8f51a39),
	.w6(32'hb8884a03),
	.w7(32'hb8a6038a),
	.w8(32'hb9402858),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb734c65d),
	.w1(32'h381cfd47),
	.w2(32'h37fc2a39),
	.w3(32'hb6f26e02),
	.w4(32'h37ac384e),
	.w5(32'h380bec2a),
	.w6(32'hb5b40765),
	.w7(32'h36a60975),
	.w8(32'h383a82ea),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37874674),
	.w1(32'h37e952c3),
	.w2(32'h376e23a7),
	.w3(32'h38033014),
	.w4(32'h379a365c),
	.w5(32'h37a8b02d),
	.w6(32'h38031211),
	.w7(32'h3813f642),
	.w8(32'h37693f15),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3575835d),
	.w1(32'h363ff3a8),
	.w2(32'h36092e45),
	.w3(32'h376d21fd),
	.w4(32'h3735c686),
	.w5(32'hb6f835e7),
	.w6(32'h37c8ab39),
	.w7(32'h373a2414),
	.w8(32'hb7a0fe86),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce83eb),
	.w1(32'h3980304c),
	.w2(32'h39cd3b0c),
	.w3(32'h3844ad3b),
	.w4(32'h398296c5),
	.w5(32'h39f8a4de),
	.w6(32'h3838a9fc),
	.w7(32'h39a47088),
	.w8(32'h3a0675c1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1db5d),
	.w1(32'h38e2715f),
	.w2(32'h384694bb),
	.w3(32'h398b56c8),
	.w4(32'hb702cbe7),
	.w5(32'h392f77ab),
	.w6(32'h3979f618),
	.w7(32'h39873213),
	.w8(32'h39a59e68),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a20463),
	.w1(32'hb883a282),
	.w2(32'hb9508579),
	.w3(32'h37886ada),
	.w4(32'hb93bdfa3),
	.w5(32'hba0f15b3),
	.w6(32'hb9219394),
	.w7(32'hb99ca134),
	.w8(32'hb9fedd29),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ec180),
	.w1(32'hb9a60ed1),
	.w2(32'hb97d62b4),
	.w3(32'hb954e190),
	.w4(32'hb989c134),
	.w5(32'hb966fa37),
	.w6(32'hb9582214),
	.w7(32'hb98df49a),
	.w8(32'hb984a2dc),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b8fc59),
	.w1(32'h37d16b19),
	.w2(32'h37c48afc),
	.w3(32'hb79e4bd6),
	.w4(32'hb804e253),
	.w5(32'h38d67de5),
	.w6(32'hb87e9319),
	.w7(32'h36754c69),
	.w8(32'h3912a1ee),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e5d02d),
	.w1(32'hb818d910),
	.w2(32'h38a1a28f),
	.w3(32'hb8624d10),
	.w4(32'hb7c00185),
	.w5(32'h38cc4647),
	.w6(32'hb8923555),
	.w7(32'hb81a691d),
	.w8(32'h38ab6c83),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782cfc8),
	.w1(32'hb76c2ebb),
	.w2(32'hb8754f64),
	.w3(32'h36d1c8c9),
	.w4(32'h363db82d),
	.w5(32'hb892226e),
	.w6(32'h3711b0a2),
	.w7(32'hb74bcb72),
	.w8(32'hb8a859e2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980a066),
	.w1(32'h390550ec),
	.w2(32'h38f0cf9d),
	.w3(32'hb9343dbe),
	.w4(32'h39c35b33),
	.w5(32'h39b18b91),
	.w6(32'hb8930a55),
	.w7(32'h39304beb),
	.w8(32'h39e633b9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3840f5d7),
	.w1(32'h38d1b803),
	.w2(32'h390a55d3),
	.w3(32'h388b9118),
	.w4(32'h38fd8a16),
	.w5(32'h39442ed9),
	.w6(32'h389cd6fd),
	.w7(32'h38f6e96f),
	.w8(32'h394bb179),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3766a598),
	.w1(32'h37933630),
	.w2(32'hb9024019),
	.w3(32'h39abbcbb),
	.w4(32'hb67c6f3d),
	.w5(32'hb8ab3e75),
	.w6(32'h38d12292),
	.w7(32'hb933a390),
	.w8(32'hb922390f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule