module layer_6_featuremap_74(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7568e4),
	.w1(32'hb98e622b),
	.w2(32'h3b2630e1),
	.w3(32'hbbaa07a8),
	.w4(32'hbb359986),
	.w5(32'hbb1198e1),
	.w6(32'hba8c6181),
	.w7(32'h375ccb65),
	.w8(32'h3a6388f3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba053524),
	.w1(32'h3ab70b47),
	.w2(32'h39343fa3),
	.w3(32'h3a29d184),
	.w4(32'hba7dde98),
	.w5(32'h3b391ab2),
	.w6(32'h3b1bc7ad),
	.w7(32'h3b00cef5),
	.w8(32'h3b668057),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11fad6),
	.w1(32'h3c234f51),
	.w2(32'hbc04ec52),
	.w3(32'h3c27a859),
	.w4(32'hbc78a54e),
	.w5(32'hbbe35171),
	.w6(32'h3c8cb927),
	.w7(32'hbc2e5ce4),
	.w8(32'hbbf67096),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7c051),
	.w1(32'hb97e9b54),
	.w2(32'hbae93db0),
	.w3(32'hbb39bae0),
	.w4(32'h3906966f),
	.w5(32'hba127c5d),
	.w6(32'hbb4af6e5),
	.w7(32'h3a7bc420),
	.w8(32'h3aeffe97),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d7b75),
	.w1(32'hba1fcb98),
	.w2(32'hbc1a0efc),
	.w3(32'h3ccbf063),
	.w4(32'hbcd58919),
	.w5(32'h3c9f39b5),
	.w6(32'h3c462e97),
	.w7(32'hbcf5561e),
	.w8(32'h3c6d54e1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12cf55),
	.w1(32'hbaee52eb),
	.w2(32'hbb5b558f),
	.w3(32'hbb5f1931),
	.w4(32'hbb9416bd),
	.w5(32'h3afd80f4),
	.w6(32'hbb26e4f3),
	.w7(32'hbba1b64f),
	.w8(32'hb8150a00),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b1960),
	.w1(32'hbb8d72cf),
	.w2(32'hbada2c3b),
	.w3(32'hbbd1017e),
	.w4(32'h3b685f2a),
	.w5(32'hbb204bb1),
	.w6(32'hbbed2ddf),
	.w7(32'h3bb1370e),
	.w8(32'hba6fd5e3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af46829),
	.w1(32'h3b02d7d3),
	.w2(32'hbd4908e6),
	.w3(32'hbc75f512),
	.w4(32'h3af7f697),
	.w5(32'h3bf6a134),
	.w6(32'hbc915a2c),
	.w7(32'hbcc93147),
	.w8(32'h3c09f1fd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d28811b),
	.w1(32'h3babd9d7),
	.w2(32'hba8f92b2),
	.w3(32'hbb4b65a3),
	.w4(32'hbbc5bd6d),
	.w5(32'hbb4243c9),
	.w6(32'h3c4191f0),
	.w7(32'hbbdd0595),
	.w8(32'hbc283260),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc434b78),
	.w1(32'hbb00ec40),
	.w2(32'h3a6eb4c6),
	.w3(32'hbb5b4a91),
	.w4(32'hbb7f0ae1),
	.w5(32'hba5dd55a),
	.w6(32'hba10e01e),
	.w7(32'hbaec2ffa),
	.w8(32'h3b0a3b57),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a981edc),
	.w1(32'hbd0028c2),
	.w2(32'hbcd22249),
	.w3(32'hbc9b761e),
	.w4(32'hbd37e5be),
	.w5(32'hbcf3a4bc),
	.w6(32'hbd0eff93),
	.w7(32'hbd39d481),
	.w8(32'hbd2cb50b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa5804),
	.w1(32'h3b99e7ac),
	.w2(32'h3bf5f375),
	.w3(32'h3b780592),
	.w4(32'h3aa81fac),
	.w5(32'h3b1156e5),
	.w6(32'h3af7e5b2),
	.w7(32'hbb4201e2),
	.w8(32'hbb0403ae),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b2726),
	.w1(32'hbbd42e1d),
	.w2(32'h3ac28f0b),
	.w3(32'hbbc70eb5),
	.w4(32'h3b9f9861),
	.w5(32'h3af35e7c),
	.w6(32'hbb8b34ac),
	.w7(32'h3bdee7bd),
	.w8(32'h3b6fcb03),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a286c93),
	.w1(32'hbb9d5c0b),
	.w2(32'h3c45748f),
	.w3(32'hbb3e39f1),
	.w4(32'h3b437e7a),
	.w5(32'h395bdded),
	.w6(32'hbba18167),
	.w7(32'h3b868f77),
	.w8(32'h3a3e4896),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfba95),
	.w1(32'h37a9a671),
	.w2(32'h3bb06798),
	.w3(32'hbaab0d3b),
	.w4(32'h3b3bbe1a),
	.w5(32'hba9ef2d5),
	.w6(32'hbb872190),
	.w7(32'h3b5b598e),
	.w8(32'h3afc2af2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be143e2),
	.w1(32'hbb69d974),
	.w2(32'h38860875),
	.w3(32'hbbb60ee2),
	.w4(32'h3b4182ba),
	.w5(32'hbaaf423d),
	.w6(32'hbb9a8e76),
	.w7(32'h3a2c610f),
	.w8(32'hbb288908),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5db58),
	.w1(32'hbbacc6ab),
	.w2(32'h3ca89cd2),
	.w3(32'h3ad52787),
	.w4(32'h3c5dec27),
	.w5(32'hba203064),
	.w6(32'h3bfae84f),
	.w7(32'h3cc580c1),
	.w8(32'h3c4f0b69),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad24738),
	.w1(32'hbbd0a5b8),
	.w2(32'hbb442046),
	.w3(32'hbbf6f476),
	.w4(32'hbaf5c596),
	.w5(32'hbbf57637),
	.w6(32'hbbc005a7),
	.w7(32'h3a2be3c0),
	.w8(32'hbb77d117),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b7d4),
	.w1(32'hba42ad1d),
	.w2(32'h398747f1),
	.w3(32'h39837b7e),
	.w4(32'hb93c7cd4),
	.w5(32'h39a3e3d2),
	.w6(32'hb8a714ee),
	.w7(32'hb94f08e2),
	.w8(32'h3a85c409),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd18e2),
	.w1(32'hbc33b7ed),
	.w2(32'h3ce7b779),
	.w3(32'h3c80ec98),
	.w4(32'h3b60e486),
	.w5(32'h3bad9ff0),
	.w6(32'h3c44483b),
	.w7(32'h3c31bde6),
	.w8(32'h3c640861),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be052),
	.w1(32'h3a301d8e),
	.w2(32'hbb2f4c3b),
	.w3(32'hba0d5082),
	.w4(32'hbb6cc89a),
	.w5(32'hbb3ec072),
	.w6(32'hba3f590e),
	.w7(32'hbaf51467),
	.w8(32'hbb4b34f6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c0398e),
	.w1(32'hbaf7d1e0),
	.w2(32'h3a576f69),
	.w3(32'h3c06a195),
	.w4(32'hbc08e910),
	.w5(32'h3b66f3a7),
	.w6(32'h3b16f80a),
	.w7(32'hbb90f2c5),
	.w8(32'h3b96c368),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa27fbf),
	.w1(32'h3cdbe033),
	.w2(32'hbc83a44e),
	.w3(32'hbab64bcd),
	.w4(32'hbc05934e),
	.w5(32'h3becacad),
	.w6(32'h3c97420e),
	.w7(32'hbcb401bb),
	.w8(32'h3c8cadd3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4489ab),
	.w1(32'hbc9505a4),
	.w2(32'h3ce5e6c9),
	.w3(32'hbccbd2c3),
	.w4(32'h3d0ee25c),
	.w5(32'hbc0da169),
	.w6(32'hbd30091a),
	.w7(32'h3cde24c0),
	.w8(32'h3ba20dad),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc429410),
	.w1(32'h3c2300af),
	.w2(32'h3badb010),
	.w3(32'hbc92c26e),
	.w4(32'h3c20a9f3),
	.w5(32'hbbdc3064),
	.w6(32'hbbcdae93),
	.w7(32'h3c381194),
	.w8(32'hbbb49599),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade2a9d),
	.w1(32'h3cf7d024),
	.w2(32'h3c7a0819),
	.w3(32'h3c8fb834),
	.w4(32'hbc387df3),
	.w5(32'h3a90de75),
	.w6(32'h3d034123),
	.w7(32'h3b9b3783),
	.w8(32'h3c59ac2b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a1f1),
	.w1(32'hbb06c8fe),
	.w2(32'hbbc5860b),
	.w3(32'hba96938c),
	.w4(32'h3b3daae7),
	.w5(32'hbafa55a1),
	.w6(32'h3a8c14dd),
	.w7(32'h3a3c22f8),
	.w8(32'h3b2fd381),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb212e4b),
	.w1(32'hbaaa5c9a),
	.w2(32'h3b4908e7),
	.w3(32'hba8a2850),
	.w4(32'h3b998f3a),
	.w5(32'hba146b5a),
	.w6(32'hbb34af99),
	.w7(32'h3bbb422b),
	.w8(32'h3a3ba62f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bcaf0),
	.w1(32'h3a45bf21),
	.w2(32'h3ab981a8),
	.w3(32'h3b33de70),
	.w4(32'h3b025b14),
	.w5(32'hbbbb5207),
	.w6(32'h39248d98),
	.w7(32'h391b1a6b),
	.w8(32'hbbc5c245),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f1ec0),
	.w1(32'hbbfa91d5),
	.w2(32'hbc8c65d4),
	.w3(32'hbc30e2f4),
	.w4(32'hbbeb93aa),
	.w5(32'hbc9f1fcb),
	.w6(32'hbcb0eae6),
	.w7(32'h3be5dc8c),
	.w8(32'hbc894f5b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58fc0b),
	.w1(32'h3bb987fc),
	.w2(32'hbc056097),
	.w3(32'h3d103226),
	.w4(32'hbbfb9d04),
	.w5(32'h39b7f640),
	.w6(32'h3c83fb0d),
	.w7(32'hbc8a278a),
	.w8(32'h3bd53dbb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44beac),
	.w1(32'h3a9c8f1f),
	.w2(32'h3b9b7493),
	.w3(32'h3a9ebad3),
	.w4(32'hbb7a49d4),
	.w5(32'hbb12806d),
	.w6(32'h3a04866e),
	.w7(32'h3c0c2131),
	.w8(32'hbc38c821),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf9ffc),
	.w1(32'h3bc4b0a1),
	.w2(32'hbb4f062a),
	.w3(32'hbd43be49),
	.w4(32'h3c42b8d2),
	.w5(32'h3ca1bf78),
	.w6(32'hbcbdcda7),
	.w7(32'h3c94cbc6),
	.w8(32'h3c9fb8bc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1600d2),
	.w1(32'h3c2f21de),
	.w2(32'hbc59f38c),
	.w3(32'h3c84e30a),
	.w4(32'hbc8bc71d),
	.w5(32'h3b429be7),
	.w6(32'h3cd5edcc),
	.w7(32'hbcf743bb),
	.w8(32'h3c2df118),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac6911),
	.w1(32'h3bbca5dc),
	.w2(32'hbb7dd621),
	.w3(32'h3bc9edaa),
	.w4(32'hbb59bf3a),
	.w5(32'h392dbe2b),
	.w6(32'h3bfdd6f1),
	.w7(32'hbbad579c),
	.w8(32'h3a93187f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393896d9),
	.w1(32'h3bc3d96a),
	.w2(32'h3b159f21),
	.w3(32'h3b2cb2fe),
	.w4(32'hbb44219f),
	.w5(32'hbad2a227),
	.w6(32'h3adcd72d),
	.w7(32'hbb9c7241),
	.w8(32'hbbceed18),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ed1f1),
	.w1(32'hba347633),
	.w2(32'h3b8ce501),
	.w3(32'hba74d7bc),
	.w4(32'hbae3f26b),
	.w5(32'h3b97da04),
	.w6(32'h39f5298d),
	.w7(32'hbb6f60bd),
	.w8(32'h3b1432cd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c85f),
	.w1(32'h3aae3cb8),
	.w2(32'h3b8b42ba),
	.w3(32'h3b8784cb),
	.w4(32'h3980dc4c),
	.w5(32'hbb1c5a23),
	.w6(32'h3b02ba7d),
	.w7(32'h39f57889),
	.w8(32'hbaff50ce),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02dd7b),
	.w1(32'hbc086fb5),
	.w2(32'h3c23ab76),
	.w3(32'h3954cb0a),
	.w4(32'h3aaeb154),
	.w5(32'h3bbefb9c),
	.w6(32'h3b9cba18),
	.w7(32'hba1c0f79),
	.w8(32'hbc19a313),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a88a4),
	.w1(32'hbd82a875),
	.w2(32'h3d90bcca),
	.w3(32'hbd0502bf),
	.w4(32'h3d2f6bf9),
	.w5(32'hbcdba653),
	.w6(32'hbd83ac9e),
	.w7(32'h3db6e5d6),
	.w8(32'hbd4c1e33),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd27105f),
	.w1(32'h3c9a1990),
	.w2(32'hbccec7ce),
	.w3(32'h3c6ce981),
	.w4(32'h3b0f02dc),
	.w5(32'hba8dfc54),
	.w6(32'h3c7266e4),
	.w7(32'hbc450fe0),
	.w8(32'h3c62d078),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba33f04),
	.w1(32'hba4de303),
	.w2(32'hbaea79f6),
	.w3(32'hbaf06aa7),
	.w4(32'hba5c8e47),
	.w5(32'hbb8507dc),
	.w6(32'hbb525eed),
	.w7(32'hb9ee44e3),
	.w8(32'hbb2e21e6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39095066),
	.w1(32'h3c239ee3),
	.w2(32'hbb9a1886),
	.w3(32'hba2f0a6b),
	.w4(32'hbbb68e68),
	.w5(32'hb9d81ab5),
	.w6(32'h3be46401),
	.w7(32'hbbcceb20),
	.w8(32'h3b08baba),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0834a5),
	.w1(32'hbad11b41),
	.w2(32'hb9dac8ec),
	.w3(32'hbc44a7b3),
	.w4(32'hbc197d71),
	.w5(32'hbb6d1ad4),
	.w6(32'hbc32f7f1),
	.w7(32'hbc53e1b2),
	.w8(32'hbb644f28),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b400d89),
	.w1(32'hbb41b7b7),
	.w2(32'hbb80b6c4),
	.w3(32'hbb34c000),
	.w4(32'hbad4e108),
	.w5(32'hbaee1fd8),
	.w6(32'hbb218331),
	.w7(32'hbb0c010a),
	.w8(32'hbaa22cb1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15052d),
	.w1(32'hbccf44df),
	.w2(32'hbcc5a9fb),
	.w3(32'hbcae8633),
	.w4(32'hbcd127e7),
	.w5(32'hbc197016),
	.w6(32'hbd105715),
	.w7(32'hbd254711),
	.w8(32'hbcb2dc22),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaab0c1),
	.w1(32'hbab6482d),
	.w2(32'h3c1c922c),
	.w3(32'hbb6d3d3c),
	.w4(32'h3bdb4621),
	.w5(32'hbc51acd4),
	.w6(32'hbbaea218),
	.w7(32'h3baa01bb),
	.w8(32'hbc091d84),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba107867),
	.w1(32'h3bf55d51),
	.w2(32'h3d865f30),
	.w3(32'h3ca423fc),
	.w4(32'h3ca1ff3d),
	.w5(32'h3bf3b7e7),
	.w6(32'h3d2c855f),
	.w7(32'h3d918d92),
	.w8(32'h3d055818),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ce384),
	.w1(32'h3b2031c9),
	.w2(32'hbb6fce52),
	.w3(32'h3aaa317b),
	.w4(32'h39f0fd8e),
	.w5(32'h3bc36da7),
	.w6(32'h3b02a926),
	.w7(32'hba06bc6a),
	.w8(32'h3b3bc544),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7526ce),
	.w1(32'hbb6d68a5),
	.w2(32'hbcbd9666),
	.w3(32'hbc0b02fa),
	.w4(32'hbc728b9f),
	.w5(32'h3c553637),
	.w6(32'h3b89a06f),
	.w7(32'hbc9b9ec6),
	.w8(32'h3cac7941),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca5467),
	.w1(32'h3a11dbc5),
	.w2(32'hbb9fbbdf),
	.w3(32'h39f7f445),
	.w4(32'hbabbb6dc),
	.w5(32'hb9b06663),
	.w6(32'hba888caa),
	.w7(32'hbb11c9c2),
	.w8(32'hb9a3104c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f227c),
	.w1(32'hbaff7415),
	.w2(32'hbb3d5116),
	.w3(32'h3ad3cd5c),
	.w4(32'hbb04d54d),
	.w5(32'hbbb8155a),
	.w6(32'hba0e752e),
	.w7(32'hbb5cea8a),
	.w8(32'hbb4d287a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7f304),
	.w1(32'h37d9e2b7),
	.w2(32'hbb487f9e),
	.w3(32'hbb963319),
	.w4(32'h3bbaad19),
	.w5(32'hbb55a503),
	.w6(32'hbba724b8),
	.w7(32'h3b4ff00d),
	.w8(32'hbb776fc5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cf12f),
	.w1(32'h3b885e65),
	.w2(32'h3998d1ad),
	.w3(32'h3b868fa0),
	.w4(32'h3b9e29ca),
	.w5(32'hbbdb7366),
	.w6(32'h3b31b442),
	.w7(32'h3b6fe902),
	.w8(32'hbc3dd7b0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14e2ad),
	.w1(32'h3b445a38),
	.w2(32'h3a6ec052),
	.w3(32'h3ae74b6f),
	.w4(32'hba3dd8dd),
	.w5(32'h39c4b381),
	.w6(32'h3a5024eb),
	.w7(32'h3ba20d0f),
	.w8(32'h3b4d233e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51f16c),
	.w1(32'h3cfac471),
	.w2(32'h3ce6d68a),
	.w3(32'h3c12173b),
	.w4(32'h3cb72e3a),
	.w5(32'h3c9c5349),
	.w6(32'h3d04fb38),
	.w7(32'h3d14d7cc),
	.w8(32'h3d1595c5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c465e36),
	.w1(32'hbaf6d4a0),
	.w2(32'h39cb8352),
	.w3(32'hbbf59479),
	.w4(32'hbb7f95e2),
	.w5(32'hbbb49328),
	.w6(32'h3a9e2f5a),
	.w7(32'h3b9a020e),
	.w8(32'h3b32908e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19556e),
	.w1(32'hba2a7f6e),
	.w2(32'hbc255556),
	.w3(32'h3c24358a),
	.w4(32'h3c3c1586),
	.w5(32'h3bfe45a4),
	.w6(32'hbbe8b196),
	.w7(32'hbc066641),
	.w8(32'h3ba9ca79),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19fb0d),
	.w1(32'h39cf406d),
	.w2(32'h3a77f1f4),
	.w3(32'h39051da1),
	.w4(32'hbab2ca08),
	.w5(32'h389112b1),
	.w6(32'hbabd3fe0),
	.w7(32'hba9be75b),
	.w8(32'hbb098252),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b034ca6),
	.w1(32'h3cb33985),
	.w2(32'h3c901690),
	.w3(32'hbc9fec1d),
	.w4(32'h3c0653b1),
	.w5(32'h3baf91c3),
	.w6(32'hbbab92af),
	.w7(32'h3c9c5a6f),
	.w8(32'h3ce0ea6a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadd1ee),
	.w1(32'hbb6e452c),
	.w2(32'hbbf501e1),
	.w3(32'h3b84b14d),
	.w4(32'hb9c2d15c),
	.w5(32'hba977443),
	.w6(32'h3b87c1a3),
	.w7(32'hb9c9cefe),
	.w8(32'hbb9a4529),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43be49),
	.w1(32'hbd2b5433),
	.w2(32'hbdb22551),
	.w3(32'hbd8325ba),
	.w4(32'hbda91dd3),
	.w5(32'hbd53a2e8),
	.w6(32'hbdc22c35),
	.w7(32'hbe11dfd0),
	.w8(32'hbdbbf08e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2fd8ab),
	.w1(32'hbc92da37),
	.w2(32'h3c0ec4af),
	.w3(32'h3c36b605),
	.w4(32'h3c7d5f92),
	.w5(32'h3bf822c9),
	.w6(32'hbcd0ca02),
	.w7(32'hbc099fae),
	.w8(32'hbbf8a985),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0d1b),
	.w1(32'h3bcf9797),
	.w2(32'h3b9f8f1d),
	.w3(32'h3b88fff8),
	.w4(32'hbaff1eff),
	.w5(32'hbbabb58d),
	.w6(32'h3c275b85),
	.w7(32'h3bc3ea6d),
	.w8(32'hbadb1e0d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule