module layer_10_featuremap_463(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h355a205e),
	.w1(32'h34142a07),
	.w2(32'hb4217be9),
	.w3(32'h350a0cb7),
	.w4(32'hb4d087ea),
	.w5(32'hb5087ee6),
	.w6(32'hb3858560),
	.w7(32'hb582903d),
	.w8(32'hb53be5a7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb804ab28),
	.w1(32'hb48e7956),
	.w2(32'hb87e0dbc),
	.w3(32'hb8a04bdf),
	.w4(32'hb8839a81),
	.w5(32'hb8bdc8ba),
	.w6(32'hb8cd5030),
	.w7(32'hb87944b4),
	.w8(32'hb88d2c2e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35085594),
	.w1(32'hb395a26a),
	.w2(32'hb4695da9),
	.w3(32'hb453d585),
	.w4(32'hb5293a4c),
	.w5(32'hb5590956),
	.w6(32'hb516cbba),
	.w7(32'hb5a45aa6),
	.w8(32'hb5753273),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37858263),
	.w1(32'h37ddd66a),
	.w2(32'h38270d10),
	.w3(32'h37ee93cd),
	.w4(32'h37efed6f),
	.w5(32'h37fef75e),
	.w6(32'h37ce4099),
	.w7(32'h3818ec8f),
	.w8(32'h381c5230),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70356ae),
	.w1(32'hb7222cbc),
	.w2(32'hb74b3ec6),
	.w3(32'hb6dff532),
	.w4(32'hb731d5ff),
	.w5(32'hb743ceb1),
	.w6(32'hb729811e),
	.w7(32'hb714c4e3),
	.w8(32'hb6f47382),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35642f2b),
	.w1(32'h34be7ffd),
	.w2(32'h34b4c47e),
	.w3(32'h349d4515),
	.w4(32'h337b39a5),
	.w5(32'hb45c1299),
	.w6(32'hb4b49d24),
	.w7(32'hb53faf32),
	.w8(32'hb47a3239),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e59945),
	.w1(32'hb9101142),
	.w2(32'hb9807a8a),
	.w3(32'h39541393),
	.w4(32'hb821d526),
	.w5(32'hb932fb73),
	.w6(32'h396a37b8),
	.w7(32'h388627d4),
	.w8(32'hb949d8ad),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd9e90),
	.w1(32'hb9b92fa8),
	.w2(32'hb9a1257f),
	.w3(32'hb9bc1476),
	.w4(32'hb9383ea5),
	.w5(32'hb9573c9d),
	.w6(32'h352b6b32),
	.w7(32'hb8a3d677),
	.w8(32'hb844c553),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3543b945),
	.w1(32'h3801db0b),
	.w2(32'h37ae8984),
	.w3(32'h353153ed),
	.w4(32'h37bdcf9e),
	.w5(32'h37bd9965),
	.w6(32'hb72b966d),
	.w7(32'hb58e9539),
	.w8(32'h37b99a8e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a20063),
	.w1(32'hb923695d),
	.w2(32'hb925a948),
	.w3(32'hb95bc208),
	.w4(32'hb78caa65),
	.w5(32'hb84837fa),
	.w6(32'h38ed2b54),
	.w7(32'h39243e49),
	.w8(32'hb8824668),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ef485),
	.w1(32'hb8a2f227),
	.w2(32'hb81c0970),
	.w3(32'hb76d0a57),
	.w4(32'hb7beddef),
	.w5(32'hb6685e27),
	.w6(32'hb8190170),
	.w7(32'hb846f5d4),
	.w8(32'hb7761605),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7272859),
	.w1(32'hb9189f6e),
	.w2(32'hb91b1e05),
	.w3(32'h38e46325),
	.w4(32'hb84447f6),
	.w5(32'hb8dc9801),
	.w6(32'h39467f04),
	.w7(32'h3931a01d),
	.w8(32'hb830f934),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fc4e2),
	.w1(32'hb94d881b),
	.w2(32'hb9362501),
	.w3(32'hb88c501e),
	.w4(32'h36f46cf8),
	.w5(32'hb7f6c900),
	.w6(32'h39085801),
	.w7(32'h38c7059e),
	.w8(32'hb89ad142),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df080a),
	.w1(32'hb967ca76),
	.w2(32'hb981e33f),
	.w3(32'hb90fa6a5),
	.w4(32'hb94dba4a),
	.w5(32'hb9414eb9),
	.w6(32'hb84a0e2d),
	.w7(32'hb8ddb668),
	.w8(32'hb934f241),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c73f2c),
	.w1(32'h3839f644),
	.w2(32'h38a3fc2b),
	.w3(32'hb6b4bfa9),
	.w4(32'h388cb939),
	.w5(32'h3898d0cd),
	.w6(32'h38399373),
	.w7(32'h38e81c18),
	.w8(32'h38eef371),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6dc1d),
	.w1(32'hb95fb550),
	.w2(32'hb9588733),
	.w3(32'hb9b94cb6),
	.w4(32'hb979c342),
	.w5(32'hb95249ae),
	.w6(32'hb913af50),
	.w7(32'hb8b1b287),
	.w8(32'hb95e0025),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75a2b6d),
	.w1(32'hb83dfbc5),
	.w2(32'hb7f1a792),
	.w3(32'hb7f596d5),
	.w4(32'hb8b73dd2),
	.w5(32'hb863bf06),
	.w6(32'hb45c447a),
	.w7(32'hb78e85a3),
	.w8(32'h367c6a8e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b6d6f),
	.w1(32'hb948f6f2),
	.w2(32'hb97640c3),
	.w3(32'hb8a90f82),
	.w4(32'hb8a49cc4),
	.w5(32'hb8374d57),
	.w6(32'h391a6470),
	.w7(32'h38c447dd),
	.w8(32'hb897da39),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e3f0a3),
	.w1(32'hb892a038),
	.w2(32'hb8b36235),
	.w3(32'h36b65bea),
	.w4(32'h38675d62),
	.w5(32'h37f48a3c),
	.w6(32'h39044d5c),
	.w7(32'h38cd8908),
	.w8(32'h339c7236),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3690e53c),
	.w1(32'h36255f54),
	.w2(32'h35db2705),
	.w3(32'h3648b1cf),
	.w4(32'h35bb85de),
	.w5(32'h3599caa8),
	.w6(32'hb5a04cad),
	.w7(32'h36001d70),
	.w8(32'h33cd3df4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368473e7),
	.w1(32'h363bfc8b),
	.w2(32'h35d10bdf),
	.w3(32'h360785ca),
	.w4(32'hb4321504),
	.w5(32'hb5d86912),
	.w6(32'h3421c662),
	.w7(32'hb60e5c13),
	.w8(32'hb5e81c29),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb699d5b9),
	.w1(32'h37b4156b),
	.w2(32'hb78390ae),
	.w3(32'hb8024ed9),
	.w4(32'h37362c75),
	.w5(32'hb7a7beee),
	.w6(32'hb7f95a2a),
	.w7(32'h381772ee),
	.w8(32'h37fef5dd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba214622),
	.w1(32'hb9dde64b),
	.w2(32'hb8faa56d),
	.w3(32'hb909a8a4),
	.w4(32'hb8076add),
	.w5(32'h37df47fa),
	.w6(32'h3934a7a1),
	.w7(32'h39cf0107),
	.w8(32'h3830c7e2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c55bc),
	.w1(32'hb906b361),
	.w2(32'hb84c9153),
	.w3(32'hb8c22f9b),
	.w4(32'h383a08ce),
	.w5(32'h38e538cb),
	.w6(32'h38e22e73),
	.w7(32'h393f4e0e),
	.w8(32'h38ef1415),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e49718),
	.w1(32'h38d382b6),
	.w2(32'h38a92175),
	.w3(32'hb8aba675),
	.w4(32'h38caba17),
	.w5(32'h38adff05),
	.w6(32'hb8852532),
	.w7(32'h38e4c157),
	.w8(32'h387521b6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888d2fe),
	.w1(32'hb80a2d2f),
	.w2(32'h36d05303),
	.w3(32'hb82721d4),
	.w4(32'h36a3810b),
	.w5(32'h37af9824),
	.w6(32'h36bd2c46),
	.w7(32'h37dbc0eb),
	.w8(32'h3739abca),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f32927),
	.w1(32'h36b41374),
	.w2(32'h36804bbf),
	.w3(32'h35e35e7f),
	.w4(32'hb5bb686f),
	.w5(32'hb6836057),
	.w6(32'hb7007dac),
	.w7(32'hb73804cd),
	.w8(32'hb714e7e4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6890ca6),
	.w1(32'h371dce94),
	.w2(32'h3883da89),
	.w3(32'hb96d8766),
	.w4(32'h3901a443),
	.w5(32'h3934ca8f),
	.w6(32'h392b76d7),
	.w7(32'h38d20a58),
	.w8(32'h3995efaa),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be80fb),
	.w1(32'hb8a5aa35),
	.w2(32'hb84ebc07),
	.w3(32'hb8c6bbd1),
	.w4(32'hb8ada35c),
	.w5(32'hb8253051),
	.w6(32'hb8c7459e),
	.w7(32'hb8441401),
	.w8(32'h375756ff),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ad139),
	.w1(32'h380d7147),
	.w2(32'h391da174),
	.w3(32'hb50d33ba),
	.w4(32'h392f0544),
	.w5(32'h39563ab8),
	.w6(32'h397ed2bc),
	.w7(32'h395b46db),
	.w8(32'h398e206f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6022714),
	.w1(32'hb6871d23),
	.w2(32'hb5ea197a),
	.w3(32'hb64de65c),
	.w4(32'hb7187218),
	.w5(32'hb61519af),
	.w6(32'h36165cdc),
	.w7(32'h34ab10ee),
	.w8(32'h35e83142),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb801fb2a),
	.w1(32'hb80894d2),
	.w2(32'hb7f0786c),
	.w3(32'hb7b85a0b),
	.w4(32'hb8048430),
	.w5(32'hb7962ca5),
	.w6(32'hb7a2b4d0),
	.w7(32'hb65e0a9b),
	.w8(32'hb609c9c4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec14ab),
	.w1(32'hb8f4ee6b),
	.w2(32'hb8f33bc7),
	.w3(32'hb77049ab),
	.w4(32'hb7ce7d7b),
	.w5(32'hb7fc2a10),
	.w6(32'h388c2b40),
	.w7(32'h382eef09),
	.w8(32'hb84e7df9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36528280),
	.w1(32'hb6d67a79),
	.w2(32'hb81e8576),
	.w3(32'hb7a68a5e),
	.w4(32'hb763d945),
	.w5(32'hb8167265),
	.w6(32'hb80dadd8),
	.w7(32'hb775ae1b),
	.w8(32'hb808c1be),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35baf1c3),
	.w1(32'hb68f42cc),
	.w2(32'hb7580b30),
	.w3(32'hb6f13741),
	.w4(32'hb78edb3c),
	.w5(32'hb6e1cb14),
	.w6(32'h37bafc65),
	.w7(32'h3706a372),
	.w8(32'hb70579ca),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ab9e8),
	.w1(32'hb8b64e4f),
	.w2(32'hb8da1dbc),
	.w3(32'h3908f52c),
	.w4(32'hb7849490),
	.w5(32'hb823d94a),
	.w6(32'h38e2994b),
	.w7(32'h38600043),
	.w8(32'hb8443c30),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941530b),
	.w1(32'hb9a68d39),
	.w2(32'hb9523c81),
	.w3(32'hb8ce3640),
	.w4(32'hb963bb54),
	.w5(32'hb945654b),
	.w6(32'h38b5e028),
	.w7(32'h39823e6f),
	.w8(32'hb72c1797),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38972a37),
	.w1(32'h397a71c0),
	.w2(32'h392aa8ac),
	.w3(32'hb940ee89),
	.w4(32'h3905161c),
	.w5(32'h39025f51),
	.w6(32'hb7f52f92),
	.w7(32'h39c3ad28),
	.w8(32'h39f08ebe),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8323709),
	.w1(32'h39486a23),
	.w2(32'h38ab1f36),
	.w3(32'hb7d6b527),
	.w4(32'h39b3bdd2),
	.w5(32'h399a2d27),
	.w6(32'h39140930),
	.w7(32'h39a21900),
	.w8(32'h39f60ad1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4c2ce),
	.w1(32'h389b4aad),
	.w2(32'h38b1f5d5),
	.w3(32'h380583c1),
	.w4(32'h38b16e6d),
	.w5(32'h3893e5ab),
	.w6(32'h37bd8c4d),
	.w7(32'h38d70760),
	.w8(32'h38a1a59d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375e9be2),
	.w1(32'h36aed1d6),
	.w2(32'h35d431aa),
	.w3(32'hb68d801e),
	.w4(32'hb6ce8212),
	.w5(32'hb692466f),
	.w6(32'h36876a47),
	.w7(32'h35f17475),
	.w8(32'h35bd9f50),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376e71bc),
	.w1(32'h378fa02c),
	.w2(32'h374199db),
	.w3(32'h374df8cc),
	.w4(32'h37036778),
	.w5(32'h36d0052b),
	.w6(32'h36a861f6),
	.w7(32'hb57039ce),
	.w8(32'hb3d609bb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8afa815),
	.w1(32'hb8c32199),
	.w2(32'hb855c109),
	.w3(32'hb8d1a1b6),
	.w4(32'hb8b75947),
	.w5(32'h36a9e2f2),
	.w6(32'hb870620c),
	.w7(32'hb8810ab0),
	.w8(32'hb86bc733),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb4722),
	.w1(32'hb9aa44e4),
	.w2(32'hb91f01ed),
	.w3(32'hb996ab4b),
	.w4(32'h372c0f90),
	.w5(32'h387c35dd),
	.w6(32'h38d3ab60),
	.w7(32'h39208b25),
	.w8(32'h38b135df),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d77bf),
	.w1(32'hb8659f9f),
	.w2(32'h38044da9),
	.w3(32'hb883e0da),
	.w4(32'h38cb6a84),
	.w5(32'h39073ead),
	.w6(32'h3870dfc3),
	.w7(32'h39256cfb),
	.w8(32'h39164e2d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94904a7),
	.w1(32'hb8071453),
	.w2(32'h37d0c8de),
	.w3(32'h37dc91d5),
	.w4(32'h3923857e),
	.w5(32'h393a767f),
	.w6(32'h38cb0c94),
	.w7(32'h394b57dc),
	.w8(32'h38de9645),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bf705),
	.w1(32'hb6dc4762),
	.w2(32'h375c86dd),
	.w3(32'hb7bf01c8),
	.w4(32'h38bfb744),
	.w5(32'h38d06c32),
	.w6(32'h3916600c),
	.w7(32'h3928213b),
	.w8(32'h391417ad),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a93358),
	.w1(32'hb97f13b2),
	.w2(32'hb9287957),
	.w3(32'hb7e2d6a1),
	.w4(32'h375a2719),
	.w5(32'h38c2260e),
	.w6(32'h39ba8f20),
	.w7(32'h398e5e20),
	.w8(32'h3847ab90),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f8dd88),
	.w1(32'h36923f88),
	.w2(32'h3768191a),
	.w3(32'hb750e1a9),
	.w4(32'h3726aedd),
	.w5(32'h3782a7bf),
	.w6(32'hb7abfac0),
	.w7(32'h373f53b7),
	.w8(32'h3786f56d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ae6b0),
	.w1(32'h38680d6d),
	.w2(32'h3862fbd9),
	.w3(32'h384d0e73),
	.w4(32'h38b59bd2),
	.w5(32'h38ce979f),
	.w6(32'h37b773c9),
	.w7(32'h384c7013),
	.w8(32'h38aada31),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f55011),
	.w1(32'hb7942990),
	.w2(32'hb7260fc8),
	.w3(32'hb69e98f2),
	.w4(32'h380148a2),
	.w5(32'h38184968),
	.w6(32'h37824714),
	.w7(32'h3862ae9f),
	.w8(32'h38612e1f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e0996),
	.w1(32'hb8df61cb),
	.w2(32'hb8884361),
	.w3(32'hb81798c2),
	.w4(32'hb7815a7d),
	.w5(32'hb84d2166),
	.w6(32'h37e22ccc),
	.w7(32'h37deeeee),
	.w8(32'hb8e12c28),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a0459a),
	.w1(32'hb878627b),
	.w2(32'hb853221b),
	.w3(32'hb885955d),
	.w4(32'hb807725a),
	.w5(32'hb82d8ea3),
	.w6(32'hb7941f57),
	.w7(32'hb74ff54e),
	.w8(32'hb809347f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9734184),
	.w1(32'hb939409e),
	.w2(32'hb97e8c11),
	.w3(32'hb8daff38),
	.w4(32'hb85b5d71),
	.w5(32'hb89bfcad),
	.w6(32'h3956a623),
	.w7(32'h3902a7a3),
	.w8(32'hb873f387),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8461ea3),
	.w1(32'hb7dee55d),
	.w2(32'hb861f56d),
	.w3(32'hb7866659),
	.w4(32'h37e03aee),
	.w5(32'hb7a2d268),
	.w6(32'hb7210ca9),
	.w7(32'hb6a83860),
	.w8(32'hb7c39090),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6055a7f),
	.w1(32'h36b2e817),
	.w2(32'h36ad17a3),
	.w3(32'hb6630736),
	.w4(32'h36b77829),
	.w5(32'h360d7250),
	.w6(32'h36cd5a19),
	.w7(32'h36c929f2),
	.w8(32'hb548ce1f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35bbbe51),
	.w1(32'h363827e8),
	.w2(32'h362b49d2),
	.w3(32'h34916626),
	.w4(32'h351a31e9),
	.w5(32'h34d3496d),
	.w6(32'hb629900c),
	.w7(32'hb5f762c7),
	.w8(32'hb595c881),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3765e1bf),
	.w1(32'h37bff253),
	.w2(32'h37b17aea),
	.w3(32'h36244435),
	.w4(32'h37364278),
	.w5(32'h37a2b59c),
	.w6(32'h372d651e),
	.w7(32'h3793dc57),
	.w8(32'h37ac409d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7996692),
	.w1(32'hb72ecaef),
	.w2(32'hb726c49b),
	.w3(32'hb70e4960),
	.w4(32'h35a61fc6),
	.w5(32'h37a12713),
	.w6(32'h3651751f),
	.w7(32'h37d0988c),
	.w8(32'h37bbbacf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f8aa5d),
	.w1(32'hb83f98a4),
	.w2(32'hb79ed1ed),
	.w3(32'hb763b58d),
	.w4(32'hb811283e),
	.w5(32'hb78521d3),
	.w6(32'h37bbe5d1),
	.w7(32'h3653334d),
	.w8(32'h3787602b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a022e),
	.w1(32'hb89f1831),
	.w2(32'hb895ceca),
	.w3(32'hb892dd88),
	.w4(32'h370b96a4),
	.w5(32'hb8028231),
	.w6(32'h37d23c1c),
	.w7(32'h37e71ac5),
	.w8(32'hb80ea21c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d7bd6),
	.w1(32'hb9651e4e),
	.w2(32'hb96e6c89),
	.w3(32'hb9407853),
	.w4(32'hb8ca5cbb),
	.w5(32'hb9390326),
	.w6(32'hb8183e25),
	.w7(32'hb85004ac),
	.w8(32'hb9184de2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3697ca0d),
	.w1(32'h364b1600),
	.w2(32'h35d8201f),
	.w3(32'h360e7c70),
	.w4(32'h3555082f),
	.w5(32'hb54f74e3),
	.w6(32'h34b65041),
	.w7(32'hb5baa0fa),
	.w8(32'hb46dcec7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363631ef),
	.w1(32'h365333a9),
	.w2(32'h36620503),
	.w3(32'h35439220),
	.w4(32'h361605b5),
	.w5(32'h35b35c2f),
	.w6(32'h35143441),
	.w7(32'h351513a7),
	.w8(32'h34b9f5ca),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7817127),
	.w1(32'hb77359b9),
	.w2(32'hb7389abd),
	.w3(32'hb77dc804),
	.w4(32'hb6d4af6f),
	.w5(32'hb69048ce),
	.w6(32'hb75ac369),
	.w7(32'hb5c24879),
	.w8(32'hb5df1b55),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ae7ea7),
	.w1(32'h363c4283),
	.w2(32'hb5167611),
	.w3(32'h3592748d),
	.w4(32'hb583527d),
	.w5(32'hb667b713),
	.w6(32'hb5ad723a),
	.w7(32'hb6473177),
	.w8(32'hb67fa820),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95124cb),
	.w1(32'hb9a4755b),
	.w2(32'hb9ed9d81),
	.w3(32'hb9e87a8e),
	.w4(32'hb9ba0d5a),
	.w5(32'hb9a601e5),
	.w6(32'h382d2ae2),
	.w7(32'hb9178f0c),
	.w8(32'hb94edf4a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bc85a),
	.w1(32'hb984a6b7),
	.w2(32'hb9976120),
	.w3(32'h36e5fc8a),
	.w4(32'hb824f831),
	.w5(32'hb8fa4a4d),
	.w6(32'hb8a56ddc),
	.w7(32'hb8ae6974),
	.w8(32'hb99023ed),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985e28e),
	.w1(32'hb91e7c7d),
	.w2(32'hb98a4409),
	.w3(32'hb8bdaff4),
	.w4(32'h377c842a),
	.w5(32'hb91d11b7),
	.w6(32'hb8229cc2),
	.w7(32'h3840a02c),
	.w8(32'hb91afd56),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c56e3c),
	.w1(32'hbbb81ff6),
	.w2(32'hbbf43525),
	.w3(32'hb86e37d7),
	.w4(32'hbbce46d7),
	.w5(32'hbbcbdc7d),
	.w6(32'hb62746e0),
	.w7(32'hbba3c1de),
	.w8(32'hbbb98769),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf20053),
	.w1(32'hbc06b07e),
	.w2(32'hbb87c4d3),
	.w3(32'hbb930be5),
	.w4(32'hbbe9b770),
	.w5(32'hbb79284a),
	.w6(32'hbbab3de9),
	.w7(32'hbc02febc),
	.w8(32'hbc0ab71c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcefe79),
	.w1(32'hbbe5f6c9),
	.w2(32'hbc0f21e3),
	.w3(32'hbbce250c),
	.w4(32'hbc15e197),
	.w5(32'hbbb3fce4),
	.w6(32'hbbd7b5a5),
	.w7(32'hbbd116eb),
	.w8(32'hbbe61a9f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b6f04),
	.w1(32'hbbb90773),
	.w2(32'hba229bbc),
	.w3(32'hbc3207c3),
	.w4(32'hbc05d879),
	.w5(32'hbb26c6c2),
	.w6(32'hbc57682d),
	.w7(32'hbba53d2a),
	.w8(32'hbb9a14a3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7499a),
	.w1(32'h3b4ed995),
	.w2(32'hbbc30b1b),
	.w3(32'h3a7fec85),
	.w4(32'h3a5ee6ed),
	.w5(32'hbbe71ebd),
	.w6(32'hbb30c1ed),
	.w7(32'hba97fb14),
	.w8(32'hbb399d54),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205e52),
	.w1(32'hb984c716),
	.w2(32'hbba2287f),
	.w3(32'hbb18aefd),
	.w4(32'hbbbb3ac0),
	.w5(32'hbbb92ae0),
	.w6(32'hbb4fbe93),
	.w7(32'hbb2ac897),
	.w8(32'hbbe38f66),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad82dbc),
	.w1(32'h3b5cca4e),
	.w2(32'h3ae30e08),
	.w3(32'hbb3ffd71),
	.w4(32'hbb42fe0d),
	.w5(32'hba6ba081),
	.w6(32'hbb28f2c6),
	.w7(32'hbbf3dd29),
	.w8(32'hbc268f8f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989e7dc),
	.w1(32'hb9003c6c),
	.w2(32'h3bcc0ca1),
	.w3(32'hbb8479bf),
	.w4(32'h3bd14072),
	.w5(32'h3bdc2858),
	.w6(32'hbc045113),
	.w7(32'h3bb7ae1b),
	.w8(32'h3bc3fd1f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a9516),
	.w1(32'h3b1337a5),
	.w2(32'h3b86a71d),
	.w3(32'h3b78ecd5),
	.w4(32'h3bb33b38),
	.w5(32'h3ac7b07a),
	.w6(32'h3b82380f),
	.w7(32'h3b1fb6cf),
	.w8(32'hbb834a00),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24c304),
	.w1(32'h3b8c229e),
	.w2(32'h398fcab6),
	.w3(32'h3ba96a13),
	.w4(32'h3b22beeb),
	.w5(32'h3a385992),
	.w6(32'h39c4f67b),
	.w7(32'h3b3a4c4f),
	.w8(32'h3ad063ec),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f5e35),
	.w1(32'hbb9f3c3b),
	.w2(32'hbc1e037a),
	.w3(32'h3b9b7775),
	.w4(32'hbb81c5b8),
	.w5(32'h3aa656e8),
	.w6(32'h3a178b28),
	.w7(32'hbbc65aab),
	.w8(32'hba468861),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55ebbc),
	.w1(32'h3a4ca056),
	.w2(32'hbb53d005),
	.w3(32'hbbc5fa54),
	.w4(32'h3b82819e),
	.w5(32'hbb224aba),
	.w6(32'hbb21c1d9),
	.w7(32'h3bf8e2b2),
	.w8(32'h3c420ab8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6af519),
	.w1(32'hbc02c4b1),
	.w2(32'hbbb0392d),
	.w3(32'h3b352078),
	.w4(32'hbbaa90ef),
	.w5(32'hbb263c90),
	.w6(32'h3c1da797),
	.w7(32'hbb9d4bfa),
	.w8(32'hb96feb36),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83ed5c),
	.w1(32'hbb3aee16),
	.w2(32'hb9f10fb9),
	.w3(32'hbacc66de),
	.w4(32'hbaa24ab6),
	.w5(32'hbadebd97),
	.w6(32'hba7adca3),
	.w7(32'h3a8b66f0),
	.w8(32'hb92cdf09),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a546acf),
	.w1(32'h3b2034d7),
	.w2(32'h38023edf),
	.w3(32'hba6a8102),
	.w4(32'h39b10ab7),
	.w5(32'h3b420aa6),
	.w6(32'h3b50557c),
	.w7(32'h3b818d36),
	.w8(32'h3bfdcc2c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33728f),
	.w1(32'hbc2685c7),
	.w2(32'hbc1b8c26),
	.w3(32'h3b7f308f),
	.w4(32'hbc328fce),
	.w5(32'hbbbb095c),
	.w6(32'h3b90ea9b),
	.w7(32'hbc3ddf7a),
	.w8(32'hbc3e209b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd74ccc),
	.w1(32'hbb444732),
	.w2(32'hb877c4e2),
	.w3(32'hbbb6079b),
	.w4(32'hbc272d56),
	.w5(32'hbba2c844),
	.w6(32'hbbfc66fa),
	.w7(32'hbaeb5196),
	.w8(32'hbc080dad),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb245b1e),
	.w1(32'hbb116d3b),
	.w2(32'h3ae73294),
	.w3(32'hbba30801),
	.w4(32'hbc416a7b),
	.w5(32'hba28b99c),
	.w6(32'hbb88296a),
	.w7(32'hbb4eee73),
	.w8(32'hbbf24b24),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa68252),
	.w1(32'h3b072523),
	.w2(32'hb93b6c74),
	.w3(32'hbaca5b9f),
	.w4(32'hb9a1405a),
	.w5(32'hb952b663),
	.w6(32'hbb6f8077),
	.w7(32'h3b78e780),
	.w8(32'h3b180f23),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfefe7f),
	.w1(32'hbbc67be9),
	.w2(32'hbb990c96),
	.w3(32'h3ab08c24),
	.w4(32'h3ad04545),
	.w5(32'h3adc483e),
	.w6(32'hba5b6b31),
	.w7(32'hbb9571b9),
	.w8(32'h3b070ded),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb539f15),
	.w1(32'hba1eaa86),
	.w2(32'hbb74f401),
	.w3(32'h3b8d441a),
	.w4(32'hbb5c366a),
	.w5(32'hbc1220c3),
	.w6(32'h3a852137),
	.w7(32'hbb3fc7aa),
	.w8(32'hbb5d3f1e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b014e),
	.w1(32'hbc388454),
	.w2(32'hbb27f907),
	.w3(32'hbb43f588),
	.w4(32'hbb902a60),
	.w5(32'h3ae2aadb),
	.w6(32'hbabe87ff),
	.w7(32'hbc01c5a6),
	.w8(32'h39d7911d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae84ec2),
	.w1(32'h3b39b2c6),
	.w2(32'hbc034562),
	.w3(32'hbab55640),
	.w4(32'hbc0aae45),
	.w5(32'hbc0a3354),
	.w6(32'hbb825587),
	.w7(32'hbc27f591),
	.w8(32'hbb97837d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba659ac),
	.w1(32'h3bdf759c),
	.w2(32'hba9011ae),
	.w3(32'hbc0a7b5d),
	.w4(32'h3bad26d2),
	.w5(32'h3bb246da),
	.w6(32'hbc0ed92c),
	.w7(32'h3c2817fd),
	.w8(32'h3c46f7c4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8454),
	.w1(32'h3b63f1a2),
	.w2(32'hba402515),
	.w3(32'hb8f0cc41),
	.w4(32'h3bb5268a),
	.w5(32'h3aa9030f),
	.w6(32'h3c09558f),
	.w7(32'h3a61c373),
	.w8(32'h3acc24df),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5411c1),
	.w1(32'hbc24befa),
	.w2(32'hbbf1c25e),
	.w3(32'h3a6ba08c),
	.w4(32'hbb9c8cab),
	.w5(32'h39e899f5),
	.w6(32'h39c840a9),
	.w7(32'hbc0716e9),
	.w8(32'hbbda0f71),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba91a7b),
	.w1(32'h3b55002e),
	.w2(32'h3adea9ea),
	.w3(32'hbbe03a0a),
	.w4(32'h3ad7f47a),
	.w5(32'h3b82e048),
	.w6(32'hbbda2217),
	.w7(32'h3b94d856),
	.w8(32'hbb7548c6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7cbeb),
	.w1(32'h3b187330),
	.w2(32'hb90dcfce),
	.w3(32'hbbcda902),
	.w4(32'hbb85c7c2),
	.w5(32'hbb2e891e),
	.w6(32'hbb5fac2e),
	.w7(32'hbbe53de6),
	.w8(32'hbbffbd8a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82167a),
	.w1(32'hbb6973d6),
	.w2(32'hba9a454a),
	.w3(32'hbabe097c),
	.w4(32'hb8b2cb74),
	.w5(32'h3b095fa6),
	.w6(32'hbbf931a1),
	.w7(32'h3b2cb87c),
	.w8(32'h3adf480b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc237fe3),
	.w1(32'h3b009bd1),
	.w2(32'h3bbc55b0),
	.w3(32'hbb8614d7),
	.w4(32'h3ba25f6a),
	.w5(32'h3c384cbb),
	.w6(32'hba090125),
	.w7(32'hbb83c560),
	.w8(32'hba03df35),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b259),
	.w1(32'hbba54379),
	.w2(32'hbc22fb2c),
	.w3(32'hbb5b5d96),
	.w4(32'hbc040511),
	.w5(32'hbc1ff989),
	.w6(32'hbc46116d),
	.w7(32'hbba9a3a1),
	.w8(32'hbba71bc3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fb7ea),
	.w1(32'hbb977ef9),
	.w2(32'hbbb26298),
	.w3(32'hbc3a9b88),
	.w4(32'hbb72cfba),
	.w5(32'hbb9145fa),
	.w6(32'hbbbcb1bc),
	.w7(32'hbbddb5ea),
	.w8(32'hbb286955),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2373df),
	.w1(32'hbaa15340),
	.w2(32'h3b13c038),
	.w3(32'hbb92f322),
	.w4(32'hbb1e80ff),
	.w5(32'h3b9db797),
	.w6(32'hbaf0a447),
	.w7(32'hbaaf3cd4),
	.w8(32'hbb059d0a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab170a1),
	.w1(32'h3ba2720e),
	.w2(32'hbad774c4),
	.w3(32'hbb16a3ab),
	.w4(32'h3a90e7e4),
	.w5(32'hb90c4f5c),
	.w6(32'hb90dcc98),
	.w7(32'h3aa5a41a),
	.w8(32'hbb05f9ad),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74d446),
	.w1(32'h3afd6298),
	.w2(32'hbbbbb2b5),
	.w3(32'hbb88c2a9),
	.w4(32'hba4f0046),
	.w5(32'hbbbc9a97),
	.w6(32'hbb4385a2),
	.w7(32'hba8ec558),
	.w8(32'hbbf5e38a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa23d3),
	.w1(32'hbaee0389),
	.w2(32'hbaccbf10),
	.w3(32'h3b8e092c),
	.w4(32'h3b0e6432),
	.w5(32'h3b945c12),
	.w6(32'hbb13b077),
	.w7(32'h3a7d201c),
	.w8(32'h3ad5db63),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae85b1e),
	.w1(32'hbb8d9ec3),
	.w2(32'hbb4facec),
	.w3(32'h3b742ec9),
	.w4(32'hbade67e0),
	.w5(32'h39b9943e),
	.w6(32'h3bead5de),
	.w7(32'hbab1fab6),
	.w8(32'hbabb1645),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67d704),
	.w1(32'h3a011bb6),
	.w2(32'h3acf0772),
	.w3(32'h3ae3c8b5),
	.w4(32'hba3810d1),
	.w5(32'hb9ab402a),
	.w6(32'h3922b66e),
	.w7(32'h3a845970),
	.w8(32'hbad78c20),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1470c),
	.w1(32'hbb2e1ff0),
	.w2(32'hbb591efa),
	.w3(32'h3aa9bd29),
	.w4(32'hba8f03a3),
	.w5(32'hbbe5f76f),
	.w6(32'h3b1596f1),
	.w7(32'hbc0fbbed),
	.w8(32'hbc1c1144),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4732c),
	.w1(32'hbb3f341c),
	.w2(32'hbba46511),
	.w3(32'hbc79ecc1),
	.w4(32'hbbb439f4),
	.w5(32'hbb0dddb6),
	.w6(32'hbc2efc83),
	.w7(32'hbae3a4b4),
	.w8(32'hbb47c3fa),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbadd0a),
	.w1(32'h3bffbd77),
	.w2(32'h3b4dcede),
	.w3(32'hbba3d320),
	.w4(32'h3b1f0129),
	.w5(32'h3bd63523),
	.w6(32'h3a3a35a7),
	.w7(32'h3a2351e7),
	.w8(32'h3b913417),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccc797),
	.w1(32'h3ba8e3dc),
	.w2(32'hbb7f793d),
	.w3(32'hbb47b97c),
	.w4(32'hbb139705),
	.w5(32'hbc4b258e),
	.w6(32'h3b62a969),
	.w7(32'hbbcbdd1d),
	.w8(32'hbc2ba46f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12769f),
	.w1(32'h3b0d1fd6),
	.w2(32'h3ae76719),
	.w3(32'hbc279ed3),
	.w4(32'hba5da5e5),
	.w5(32'h3ba82274),
	.w6(32'hbbb35335),
	.w7(32'h3a73f15a),
	.w8(32'h3a2751a9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fdb18),
	.w1(32'h3a0dc840),
	.w2(32'hbb8608a2),
	.w3(32'h3a592e8f),
	.w4(32'hbb491025),
	.w5(32'hbb2c5937),
	.w6(32'h3aceb07b),
	.w7(32'h3a766f17),
	.w8(32'hbb509633),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0b300),
	.w1(32'h3a884946),
	.w2(32'hbb83bbb2),
	.w3(32'h3b044e4e),
	.w4(32'hbbd55588),
	.w5(32'hbc2bbbbf),
	.w6(32'h3b82977e),
	.w7(32'hbb556096),
	.w8(32'hbac6a087),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b198692),
	.w1(32'h3c007a16),
	.w2(32'hba82cc36),
	.w3(32'h3b424049),
	.w4(32'h3b7381fd),
	.w5(32'hbc40dfe4),
	.w6(32'h3672ddb8),
	.w7(32'h3bf0d956),
	.w8(32'hbb0a6665),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b013601),
	.w1(32'hbb1ed297),
	.w2(32'h3b21fe1c),
	.w3(32'hba995492),
	.w4(32'hbaaf6ec3),
	.w5(32'h3ac62cd1),
	.w6(32'h3b0183dc),
	.w7(32'hbb1ee850),
	.w8(32'hbb494949),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a212e),
	.w1(32'hbae3c3f5),
	.w2(32'h3aacae2f),
	.w3(32'hbb2bf782),
	.w4(32'hbb9af3be),
	.w5(32'h3a3871ad),
	.w6(32'hb9e194e4),
	.w7(32'hbb37a250),
	.w8(32'hbb3195ad),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b772ab8),
	.w1(32'h3babed33),
	.w2(32'hba085a5c),
	.w3(32'h3b0de6b0),
	.w4(32'h3b35adf6),
	.w5(32'hb9900597),
	.w6(32'hba9475a4),
	.w7(32'h3a173a6f),
	.w8(32'h391294b7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9553cca),
	.w1(32'h3a8d479e),
	.w2(32'hbba959fc),
	.w3(32'hbb1e8781),
	.w4(32'h3b038f21),
	.w5(32'hbb00f2c3),
	.w6(32'hb8a92a51),
	.w7(32'h3b35589d),
	.w8(32'hbb9904bb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b928654),
	.w1(32'hbb801fa8),
	.w2(32'hbb7f284d),
	.w3(32'h3bb483c6),
	.w4(32'hbb1cd72a),
	.w5(32'hbb69b19e),
	.w6(32'h3b256837),
	.w7(32'hbbce83f0),
	.w8(32'hbc20d164),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7a194),
	.w1(32'hbc1c0471),
	.w2(32'h3aba9c64),
	.w3(32'h3aae4092),
	.w4(32'hbb6ad15d),
	.w5(32'h3c05df09),
	.w6(32'h3bc8faa1),
	.w7(32'hbb708824),
	.w8(32'h3c0f4a01),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea2fac),
	.w1(32'h3b0eab3f),
	.w2(32'hbc1ca862),
	.w3(32'h3b9a7e14),
	.w4(32'hbb92a98a),
	.w5(32'hbc00344f),
	.w6(32'h3b69d1bb),
	.w7(32'hbc00d2ce),
	.w8(32'hbc1f6008),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53df91),
	.w1(32'hbbdfc40f),
	.w2(32'hbad812a5),
	.w3(32'hbc05e69e),
	.w4(32'hbbe04a83),
	.w5(32'hbadc64b0),
	.w6(32'hbbeb8733),
	.w7(32'hbbe96f50),
	.w8(32'hbba16e8c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb938b38),
	.w1(32'h3ba41121),
	.w2(32'hbaff6008),
	.w3(32'hbc03521f),
	.w4(32'h38cca1d5),
	.w5(32'hbaafc3fd),
	.w6(32'hbbeb0237),
	.w7(32'h3a4d0bd9),
	.w8(32'hbb8f6d87),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb952a1a),
	.w1(32'h39a357ea),
	.w2(32'hbbffdc08),
	.w3(32'hbc14acfb),
	.w4(32'h3a25aef8),
	.w5(32'h3a9a2d3c),
	.w6(32'hba8c92e8),
	.w7(32'h3aa9f614),
	.w8(32'hbb61426b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a227f),
	.w1(32'h3ba8cabf),
	.w2(32'hbb12b51c),
	.w3(32'hbc3527ad),
	.w4(32'hbb05a0fa),
	.w5(32'hbb920871),
	.w6(32'hbbcfc79b),
	.w7(32'hbb0c9b4a),
	.w8(32'hbb9507eb),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98458f7),
	.w1(32'hbb23e81d),
	.w2(32'hbb80cd6b),
	.w3(32'hbaae1b6a),
	.w4(32'hbbc44117),
	.w5(32'hbc3fc779),
	.w6(32'h3af2e0ff),
	.w7(32'hbb162fd0),
	.w8(32'hbc001f6b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb481e4e),
	.w1(32'hbba0ec16),
	.w2(32'hbb7c9dcf),
	.w3(32'hbbef3a3b),
	.w4(32'hbbbb0eeb),
	.w5(32'hbb06351a),
	.w6(32'hbc0ac1de),
	.w7(32'hbbad086f),
	.w8(32'hbb829d6e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcadd96),
	.w1(32'hbb06b43f),
	.w2(32'hbb574b58),
	.w3(32'hbb494258),
	.w4(32'hbad05537),
	.w5(32'hbb889e41),
	.w6(32'hbb9fe94e),
	.w7(32'hbb2e869e),
	.w8(32'hb9c7bd3e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f550e),
	.w1(32'hbbb8df01),
	.w2(32'hbbde99ca),
	.w3(32'hbbf30e4a),
	.w4(32'hbbf4fb08),
	.w5(32'hbbdc53ed),
	.w6(32'hb8c9aafd),
	.w7(32'hbb88218c),
	.w8(32'hbc117c59),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1c600),
	.w1(32'hb7de3e6c),
	.w2(32'hbb938775),
	.w3(32'hbb98241a),
	.w4(32'h3b4b9dd6),
	.w5(32'hbb8be1ad),
	.w6(32'hbb704d4e),
	.w7(32'h3a8e5a07),
	.w8(32'hbb88347c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30cd87),
	.w1(32'h3b0c0468),
	.w2(32'h3adf9977),
	.w3(32'hbb5f8b02),
	.w4(32'hba3b3183),
	.w5(32'h3b893c6e),
	.w6(32'hbb2e8d8c),
	.w7(32'h3bafbc88),
	.w8(32'h3b9f2507),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca8295),
	.w1(32'hbacc151b),
	.w2(32'hbb867f1f),
	.w3(32'h3b6347d6),
	.w4(32'h3b2b5531),
	.w5(32'h3a92e77d),
	.w6(32'hbb4ded87),
	.w7(32'hba08727d),
	.w8(32'h3af41b00),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b073),
	.w1(32'h39581ff0),
	.w2(32'h3a05c915),
	.w3(32'hbbb8bd54),
	.w4(32'hbc19e21a),
	.w5(32'hbc23b2da),
	.w6(32'h3b55c1d8),
	.w7(32'hbb733abd),
	.w8(32'hbbc9918f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf223c),
	.w1(32'h3b432c5d),
	.w2(32'h3ade33ba),
	.w3(32'h3adfbe6b),
	.w4(32'h3afd6247),
	.w5(32'h3b840a8d),
	.w6(32'hbac68786),
	.w7(32'hba57c715),
	.w8(32'h3a9e9a91),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93d1f5),
	.w1(32'h3b180560),
	.w2(32'hbaf9c39f),
	.w3(32'h3b7f6196),
	.w4(32'h3ba32ffe),
	.w5(32'hbb3d24ee),
	.w6(32'hbae283df),
	.w7(32'hbb700487),
	.w8(32'hbac45ea7),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae16462),
	.w1(32'h3b876081),
	.w2(32'hbc0ff2fb),
	.w3(32'hba89a4e2),
	.w4(32'hbb629479),
	.w5(32'hbc5f033a),
	.w6(32'hbb8bc203),
	.w7(32'hbb19f486),
	.w8(32'hbc290cfc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6ddf9),
	.w1(32'hbc2664f0),
	.w2(32'hbc118751),
	.w3(32'hbb0f7088),
	.w4(32'hbbcc662b),
	.w5(32'hbb5686ce),
	.w6(32'hbba5319e),
	.w7(32'hbac6903a),
	.w8(32'h3ac9eb52),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16dcd),
	.w1(32'h39bcde53),
	.w2(32'hbb8548ad),
	.w3(32'hbb46bc2e),
	.w4(32'h3af85a1a),
	.w5(32'hb8d016c5),
	.w6(32'hbb1bf898),
	.w7(32'hbb05b69d),
	.w8(32'hbb6534d8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaacaa7),
	.w1(32'hbae60eb6),
	.w2(32'hb9f514e7),
	.w3(32'hba121d0c),
	.w4(32'h3bbc1672),
	.w5(32'h3b871739),
	.w6(32'hbbd7954a),
	.w7(32'h3b8b45aa),
	.w8(32'h3c21d0f9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cabf2),
	.w1(32'hbb130bf3),
	.w2(32'h3a39cb79),
	.w3(32'h3b9c51bd),
	.w4(32'hbaeb51c2),
	.w5(32'hbb62ee53),
	.w6(32'h3c0fa7fd),
	.w7(32'h3b2f2f5d),
	.w8(32'hbbbb972b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c173a5e),
	.w1(32'hbc09928a),
	.w2(32'hbc3d60fd),
	.w3(32'h3be71006),
	.w4(32'hbc30a006),
	.w5(32'hbc62f33a),
	.w6(32'h3bcd7779),
	.w7(32'hbc208d35),
	.w8(32'hbc5506c2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8d7a7),
	.w1(32'hbb7763cb),
	.w2(32'hbb959bd1),
	.w3(32'hbc1f0ec4),
	.w4(32'hbbe8a947),
	.w5(32'h39dbfd6a),
	.w6(32'hbc267377),
	.w7(32'hbbe91d6f),
	.w8(32'hbc0faae9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6750d7),
	.w1(32'hbbb1442e),
	.w2(32'hbbbf9af1),
	.w3(32'hbc3718ea),
	.w4(32'hbad41342),
	.w5(32'hbbc37afb),
	.w6(32'hbbf097b3),
	.w7(32'hbaa1deba),
	.w8(32'hbb7b2d2b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb51075),
	.w1(32'hbb562381),
	.w2(32'hbab6f32f),
	.w3(32'hbbadeec7),
	.w4(32'h3a31b59c),
	.w5(32'h3b303122),
	.w6(32'hbb34f59a),
	.w7(32'h39b3dc9f),
	.w8(32'h3b1412c8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51da90),
	.w1(32'hbaf00a85),
	.w2(32'hba506fcb),
	.w3(32'h3b9442e6),
	.w4(32'h3b980f7c),
	.w5(32'hbb40b841),
	.w6(32'h3a4efe43),
	.w7(32'hb91a4a40),
	.w8(32'h3b89e1aa),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c8d5c),
	.w1(32'h3aafcc39),
	.w2(32'hbb028f16),
	.w3(32'hbb84b3ba),
	.w4(32'hb9caa2dc),
	.w5(32'h3bc46dbc),
	.w6(32'h3b7cb2b8),
	.w7(32'hbaf5151c),
	.w8(32'h3b371e90),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0224e),
	.w1(32'hbab258a4),
	.w2(32'hba99798c),
	.w3(32'h39cdb9b6),
	.w4(32'hbbd1ce66),
	.w5(32'hbbd8ebb4),
	.w6(32'hba053d29),
	.w7(32'h3b0b3b22),
	.w8(32'hbc2da8f0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e5b6d),
	.w1(32'h3b0d06ad),
	.w2(32'h38382a1c),
	.w3(32'h3b4cc3a3),
	.w4(32'hbb37b44f),
	.w5(32'hbacca1da),
	.w6(32'hbbd91938),
	.w7(32'hb9328e60),
	.w8(32'h3a3461f9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30c74b),
	.w1(32'h3ae9acb5),
	.w2(32'hbb90ce70),
	.w3(32'h3b11d562),
	.w4(32'h3aff9795),
	.w5(32'hbc1e0a46),
	.w6(32'h3aae11e7),
	.w7(32'h3bc7ce5f),
	.w8(32'hbbb8c472),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0719c2),
	.w1(32'hbb40306c),
	.w2(32'hbc08a376),
	.w3(32'hbc035ba2),
	.w4(32'hbb7d4d0f),
	.w5(32'hbc158ef7),
	.w6(32'hbbd53338),
	.w7(32'hbb3d6025),
	.w8(32'hbaf24cc6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376001),
	.w1(32'h3b5f4d5c),
	.w2(32'h3bb42dc3),
	.w3(32'hbb71691c),
	.w4(32'h3b8184a6),
	.w5(32'h3b811c54),
	.w6(32'hb9c84883),
	.w7(32'h3bb059e1),
	.w8(32'h3b910432),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52d16d),
	.w1(32'hbb3bb6f0),
	.w2(32'h3b6565a8),
	.w3(32'h3b7b91c7),
	.w4(32'hbc0fcbc2),
	.w5(32'hbb0c4449),
	.w6(32'h3bbb2cc9),
	.w7(32'hbb607d41),
	.w8(32'hba5265e5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b968c8d),
	.w1(32'h3c54652e),
	.w2(32'h3c557788),
	.w3(32'hbb9d5b0b),
	.w4(32'h3b993a15),
	.w5(32'hbba3460a),
	.w6(32'hbb9d681e),
	.w7(32'h3bcd010b),
	.w8(32'h3b55e02f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c035c97),
	.w1(32'h3c119c89),
	.w2(32'hba22b607),
	.w3(32'h3ad8e320),
	.w4(32'h3b99d521),
	.w5(32'hbbcc9199),
	.w6(32'h3b263594),
	.w7(32'hbbd1c230),
	.w8(32'hbc1477e3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bbdf6),
	.w1(32'hbc3dedf7),
	.w2(32'hbb975a1b),
	.w3(32'hbb302d2f),
	.w4(32'hbc49eb2e),
	.w5(32'hbb6fc295),
	.w6(32'hbbcb908d),
	.w7(32'hbc168b0f),
	.w8(32'hbb1f7d3c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b67b6),
	.w1(32'hbb9df9e7),
	.w2(32'hbb9ed853),
	.w3(32'hbb13ce76),
	.w4(32'hbb0fc039),
	.w5(32'hbb4664d2),
	.w6(32'hb9eefa7c),
	.w7(32'hbbc3fe63),
	.w8(32'hbbfde267),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb261f5),
	.w1(32'hbb9b0408),
	.w2(32'hbbff0fc4),
	.w3(32'hbc2c8c07),
	.w4(32'hbbf1d031),
	.w5(32'hbbe799a3),
	.w6(32'hbb66a4a8),
	.w7(32'hba61a620),
	.w8(32'h39070257),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbab1dd),
	.w1(32'h3a627668),
	.w2(32'hbb7a7ce5),
	.w3(32'h3b6e8b8b),
	.w4(32'hba3b27b1),
	.w5(32'hbbb26fa5),
	.w6(32'h3b97df58),
	.w7(32'hbbe2d39e),
	.w8(32'hbbf3cf69),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf8572),
	.w1(32'hbbc6959e),
	.w2(32'hbc1a1aa4),
	.w3(32'hba628123),
	.w4(32'hbbb0e247),
	.w5(32'hbc721961),
	.w6(32'hbbfb29e0),
	.w7(32'hbbcc5432),
	.w8(32'hbc566934),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07dcb1),
	.w1(32'hbb53ed0f),
	.w2(32'hbc01dde0),
	.w3(32'hbbd1ed2d),
	.w4(32'hbac9d728),
	.w5(32'hbb7a7198),
	.w6(32'hbae5f8a2),
	.w7(32'h3a75069f),
	.w8(32'hba037882),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc206a9c),
	.w1(32'hba074b1a),
	.w2(32'hbb247969),
	.w3(32'hbb62903f),
	.w4(32'hbb75fcb1),
	.w5(32'hbac961cd),
	.w6(32'hbb8cc3e6),
	.w7(32'h39f1a3e5),
	.w8(32'h3a7c1142),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bef97),
	.w1(32'hbb95fa66),
	.w2(32'hbbb295c2),
	.w3(32'hbb20557b),
	.w4(32'h3b93c9ac),
	.w5(32'hb9a5a37f),
	.w6(32'hbb1922d0),
	.w7(32'h3b1fc196),
	.w8(32'h3b8c9f5b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc05792),
	.w1(32'hba89d0ea),
	.w2(32'hbb9dbb53),
	.w3(32'hba107713),
	.w4(32'hbb4de30d),
	.w5(32'hbb645bfa),
	.w6(32'h3b6f53ab),
	.w7(32'hbae2e77f),
	.w8(32'h3a19802e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fcecd),
	.w1(32'hbb878d4a),
	.w2(32'hbb05bb5e),
	.w3(32'h39a1a580),
	.w4(32'hbba0d8a6),
	.w5(32'h3b2884b2),
	.w6(32'h3afca701),
	.w7(32'hbbdbbcae),
	.w8(32'hbb8a4084),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba702a23),
	.w1(32'hbc35088c),
	.w2(32'hbba1d519),
	.w3(32'hbaab8f0b),
	.w4(32'hbc179620),
	.w5(32'hbc385dbd),
	.w6(32'hbb8fee23),
	.w7(32'hbbada93b),
	.w8(32'hbbebc5ed),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3838d0b0),
	.w1(32'h3a969db9),
	.w2(32'h3b613398),
	.w3(32'hb8be52c7),
	.w4(32'hbb61803f),
	.w5(32'hba27b16c),
	.w6(32'hba65c0de),
	.w7(32'h3a0ad625),
	.w8(32'hbb85defc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cd130),
	.w1(32'h38b46015),
	.w2(32'h3a44a37e),
	.w3(32'hbba0c9d7),
	.w4(32'hbbd41b68),
	.w5(32'h3aa619fa),
	.w6(32'h3a0e6bdd),
	.w7(32'hbb3c003f),
	.w8(32'h399af8b5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b994ac3),
	.w1(32'hbb03336b),
	.w2(32'hbb34d54b),
	.w3(32'hb9e36edb),
	.w4(32'hbb00480e),
	.w5(32'hbb358a72),
	.w6(32'hb9a2a034),
	.w7(32'hbb7fb82d),
	.w8(32'hbc042d50),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b77ff),
	.w1(32'hbbb26f5a),
	.w2(32'hb95d1aa8),
	.w3(32'hbbd3138d),
	.w4(32'hbb6fa948),
	.w5(32'hba3939ff),
	.w6(32'hbb5f087a),
	.w7(32'hbbb0addd),
	.w8(32'hbbe234f6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2faf3),
	.w1(32'h3ae9ad48),
	.w2(32'hbb6a85f5),
	.w3(32'hbb0f51f3),
	.w4(32'h3ac17be5),
	.w5(32'hbb761eef),
	.w6(32'hbb1b9974),
	.w7(32'h3b70f4c8),
	.w8(32'hba8808af),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e5868),
	.w1(32'h3a8f908a),
	.w2(32'h3c00b5b6),
	.w3(32'hbc101250),
	.w4(32'hbb41be95),
	.w5(32'h3c32efd9),
	.w6(32'hb919bde3),
	.w7(32'h3bbe982a),
	.w8(32'h3c578d21),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fcf97),
	.w1(32'hbc01bcfc),
	.w2(32'hbc05b897),
	.w3(32'h3b4b2eda),
	.w4(32'hbbf162f3),
	.w5(32'hbc0079f2),
	.w6(32'h3ace13f9),
	.w7(32'hbc0286d0),
	.w8(32'hbbd91663),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d9f46),
	.w1(32'hbbb86f08),
	.w2(32'hbc1d951c),
	.w3(32'hbbff4816),
	.w4(32'hbba8aa5d),
	.w5(32'hbc5ad25c),
	.w6(32'hbbc0736c),
	.w7(32'hbb43e5ba),
	.w8(32'hbbdc7e6c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc501e1d),
	.w1(32'h3b807da7),
	.w2(32'hb7577a4b),
	.w3(32'hbc0ed201),
	.w4(32'hbb35181d),
	.w5(32'hbb1eb674),
	.w6(32'hbbda6d60),
	.w7(32'h3a1ab510),
	.w8(32'h39b157e8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1304c),
	.w1(32'hbb8ab7e4),
	.w2(32'hbae5e1eb),
	.w3(32'h3b1e8d6f),
	.w4(32'hbc2e7dbd),
	.w5(32'hbb70cd66),
	.w6(32'h38bc0268),
	.w7(32'hbbe3794d),
	.w8(32'hbbbeb411),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b054687),
	.w1(32'h3c182cc8),
	.w2(32'h3b2af3c9),
	.w3(32'h3ac11570),
	.w4(32'h3ba99881),
	.w5(32'hbacb6e5d),
	.w6(32'h3b31efb7),
	.w7(32'h3bdb909b),
	.w8(32'h39e58bc8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc57e8),
	.w1(32'hba8da0a6),
	.w2(32'h3b43fc5d),
	.w3(32'h3b15f73c),
	.w4(32'h3b153663),
	.w5(32'hbb555843),
	.w6(32'hbb2bbb06),
	.w7(32'hbad16f57),
	.w8(32'hba8bce71),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7ac45),
	.w1(32'h3a9f17b4),
	.w2(32'h3b82a5a9),
	.w3(32'h3b3da4a8),
	.w4(32'h3b477344),
	.w5(32'h3b9df740),
	.w6(32'h3bb95f0e),
	.w7(32'h3a84e3e0),
	.w8(32'h3b7f48a8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeda462),
	.w1(32'h3af677b7),
	.w2(32'hbc16c68a),
	.w3(32'h3aa7fec9),
	.w4(32'hbb6a9bb0),
	.w5(32'hbc04f0e6),
	.w6(32'hba02c8b2),
	.w7(32'h38e9fd8d),
	.w8(32'hbb838e33),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1efeb9),
	.w1(32'hbac722d1),
	.w2(32'hbae039b9),
	.w3(32'hbc091449),
	.w4(32'h3b76a24f),
	.w5(32'h3a49cabe),
	.w6(32'hbbb1dd4b),
	.w7(32'h3a057e9e),
	.w8(32'h3b445ad0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb168193),
	.w1(32'h3bb19834),
	.w2(32'h3bd6300d),
	.w3(32'h3b1e7b4a),
	.w4(32'h3bad39ee),
	.w5(32'h3b8f8ef1),
	.w6(32'h3b59ac2b),
	.w7(32'h3bab7e4a),
	.w8(32'h3b9d05df),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab63ceb),
	.w1(32'hbb715adc),
	.w2(32'h3a1897a6),
	.w3(32'h3b6ba9db),
	.w4(32'hbbdd0226),
	.w5(32'h3a9235a2),
	.w6(32'hbadb5c66),
	.w7(32'hbbcbee21),
	.w8(32'hbb57408c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a840a76),
	.w1(32'h3af66f3d),
	.w2(32'hbab31685),
	.w3(32'hbaa3dadd),
	.w4(32'hbb02894d),
	.w5(32'hbb8994ac),
	.w6(32'hbb7650fe),
	.w7(32'h3b2b716f),
	.w8(32'hbb3bd01b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03185a),
	.w1(32'h3982d3b8),
	.w2(32'h3ac54529),
	.w3(32'hba9d343b),
	.w4(32'hbb5b1844),
	.w5(32'hbaa7863b),
	.w6(32'hbade6497),
	.w7(32'hb9db897e),
	.w8(32'h3ba1b9b7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19cb8d),
	.w1(32'hbb195e58),
	.w2(32'hbbfc192c),
	.w3(32'hbb046766),
	.w4(32'hbbb8f2d0),
	.w5(32'hbbd3e589),
	.w6(32'h3bade31c),
	.w7(32'hbba4e2ce),
	.w8(32'hbc010320),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01a214),
	.w1(32'hbb8fec1d),
	.w2(32'hbba60594),
	.w3(32'hbc16c322),
	.w4(32'hbbaa53fe),
	.w5(32'hbb8933c8),
	.w6(32'hbc0035ee),
	.w7(32'hbb7d04af),
	.w8(32'hbb6d68f6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b7796),
	.w1(32'hba1816b5),
	.w2(32'hba8ffae5),
	.w3(32'hbc031d23),
	.w4(32'hbc384841),
	.w5(32'hbb573cc6),
	.w6(32'hbb8896e7),
	.w7(32'hbc2963cd),
	.w8(32'hbbee0f26),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfd06e),
	.w1(32'h3b892d6a),
	.w2(32'hb9ec1c94),
	.w3(32'hbbbaf126),
	.w4(32'hbb373b4a),
	.w5(32'hbb022004),
	.w6(32'hbc315289),
	.w7(32'hb95e8241),
	.w8(32'h3ad86f6b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf5ccf),
	.w1(32'hbc03b250),
	.w2(32'hbb72edc3),
	.w3(32'hbbc4c50b),
	.w4(32'hbc103e33),
	.w5(32'h39f3a924),
	.w6(32'hbb8647eb),
	.w7(32'hbba7cd28),
	.w8(32'hba45efa0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf8020),
	.w1(32'h3b32ac70),
	.w2(32'h3b1302c9),
	.w3(32'hbb312896),
	.w4(32'h3ba9b179),
	.w5(32'h3b4af381),
	.w6(32'h3a842a2f),
	.w7(32'h3b46f7ac),
	.w8(32'h37f01b8a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dcc9c),
	.w1(32'hbb582712),
	.w2(32'h3a860d6a),
	.w3(32'hbb314b04),
	.w4(32'h3ab6acaa),
	.w5(32'h3baa52e7),
	.w6(32'h399ecf67),
	.w7(32'h3a038c50),
	.w8(32'h3bc0a2ef),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2f7a2),
	.w1(32'h3b0509e5),
	.w2(32'hb96964fa),
	.w3(32'h3a4a6382),
	.w4(32'hba09e9e6),
	.w5(32'hbb856c1b),
	.w6(32'h3b59192e),
	.w7(32'h3b3c5a46),
	.w8(32'h3b6840a0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0b8f3),
	.w1(32'h3a108d4a),
	.w2(32'h3a7f3557),
	.w3(32'hba95c8fc),
	.w4(32'hb9c8853f),
	.w5(32'hba68c50f),
	.w6(32'h3a595b01),
	.w7(32'h3b8bbdea),
	.w8(32'h3af70ba9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72565d),
	.w1(32'hbaef2170),
	.w2(32'hbbf385e2),
	.w3(32'h3b041787),
	.w4(32'h3a23e4d6),
	.w5(32'hbc5653ee),
	.w6(32'h3ba51bfa),
	.w7(32'h3c14e107),
	.w8(32'h3b4c7303),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae45aa9),
	.w1(32'h3a6967dd),
	.w2(32'h3aea24d0),
	.w3(32'h3bbf3006),
	.w4(32'hbb5523af),
	.w5(32'hbb297b68),
	.w6(32'h3befcafe),
	.w7(32'hbb976aa6),
	.w8(32'hbabe4830),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd0938),
	.w1(32'h3b9142b0),
	.w2(32'h3aad3730),
	.w3(32'h3a2340f0),
	.w4(32'h3b658c65),
	.w5(32'h3bafdb3b),
	.w6(32'hbb3b645e),
	.w7(32'h3b1fc3c7),
	.w8(32'hbb80c25a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28efe4),
	.w1(32'h3b1b0edc),
	.w2(32'h3a7f0ec8),
	.w3(32'hbba3fb36),
	.w4(32'h3b01d090),
	.w5(32'h3b8d812e),
	.w6(32'hbbb1c5bc),
	.w7(32'h3ab6dd22),
	.w8(32'h3a5bec31),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a841162),
	.w1(32'h393b543d),
	.w2(32'h3b3d0e85),
	.w3(32'hbb51cf02),
	.w4(32'hbbbeec7c),
	.w5(32'hbb7e21c3),
	.w6(32'h3a191fb3),
	.w7(32'h3a8e5d36),
	.w8(32'hbb655449),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b807002),
	.w1(32'h3be4c633),
	.w2(32'hbb89b07e),
	.w3(32'hbb18fb7c),
	.w4(32'h3b67bd18),
	.w5(32'h3c0abb0e),
	.w6(32'hbb80c73a),
	.w7(32'hb99c0e01),
	.w8(32'h3b42a520),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb176584),
	.w1(32'h3b030c3e),
	.w2(32'hb8bd6222),
	.w3(32'h3c6a183e),
	.w4(32'hbb0b13ce),
	.w5(32'h3c057aab),
	.w6(32'h3c848b21),
	.w7(32'h3ae33db8),
	.w8(32'h3b92d03b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca8953),
	.w1(32'hbac13e4b),
	.w2(32'h3b28cd34),
	.w3(32'hbaee742f),
	.w4(32'h3a327505),
	.w5(32'h38328bf4),
	.w6(32'h3a6c2a68),
	.w7(32'h3b187c92),
	.w8(32'hba8fb41c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc8ec9),
	.w1(32'h3c3d739d),
	.w2(32'h3b7ced8c),
	.w3(32'h3aec5d96),
	.w4(32'h3bddabba),
	.w5(32'h3c554f78),
	.w6(32'h3aebf686),
	.w7(32'hbc64f75d),
	.w8(32'hbc145304),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4949bd),
	.w1(32'hbbc3a3d8),
	.w2(32'hbb9343cd),
	.w3(32'h3b7ab481),
	.w4(32'h3af7d3c4),
	.w5(32'h3ba5a5f1),
	.w6(32'h39841488),
	.w7(32'h39c3224a),
	.w8(32'h3bac1f35),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a9586),
	.w1(32'hbbe644b3),
	.w2(32'h3aaed189),
	.w3(32'h3ac931df),
	.w4(32'hbb627f93),
	.w5(32'h3a6dd93a),
	.w6(32'h3b4e921b),
	.w7(32'h3b3bab69),
	.w8(32'h3ac182b6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d0180),
	.w1(32'hbc1ce5ef),
	.w2(32'h38ac1b63),
	.w3(32'h3a62eff9),
	.w4(32'h3b400783),
	.w5(32'h3bcb9dac),
	.w6(32'hbb5f1208),
	.w7(32'hbbe48ce0),
	.w8(32'h3ad3b1e7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44587e),
	.w1(32'hbb04f697),
	.w2(32'h3abeda3d),
	.w3(32'h3b2dc1d9),
	.w4(32'h389f1cce),
	.w5(32'hbbd5bd96),
	.w6(32'h3a4131ed),
	.w7(32'h3b4b51af),
	.w8(32'h3ba44ba2),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21a25b),
	.w1(32'hbbc02bc6),
	.w2(32'h3ba094dd),
	.w3(32'h3ba782ad),
	.w4(32'hbbaf377e),
	.w5(32'hb9e4c44b),
	.w6(32'h3b1627f7),
	.w7(32'hba9f8be4),
	.w8(32'hbb914026),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397075aa),
	.w1(32'h39f0d07b),
	.w2(32'h3b557e1d),
	.w3(32'hb9c15225),
	.w4(32'h3b71a740),
	.w5(32'hbba11e49),
	.w6(32'hbb693980),
	.w7(32'h3c4d60cc),
	.w8(32'h3c08ec96),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05ea57),
	.w1(32'h3b699faf),
	.w2(32'h3be2069b),
	.w3(32'h3c04e14c),
	.w4(32'hb94d6ce3),
	.w5(32'hba326318),
	.w6(32'h3bb34185),
	.w7(32'hba6cabf4),
	.w8(32'h3ad1037e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9e57),
	.w1(32'hba9b84d9),
	.w2(32'hbb07c12e),
	.w3(32'h3b83d1b0),
	.w4(32'hbb2bfe72),
	.w5(32'hbadc82c0),
	.w6(32'h3a966d49),
	.w7(32'hbb33e68d),
	.w8(32'hbb0e7d69),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe6b70),
	.w1(32'hba33ac3b),
	.w2(32'h3bbe49cd),
	.w3(32'h3ab430e8),
	.w4(32'hba5cd968),
	.w5(32'h3beab8cd),
	.w6(32'h3b79a004),
	.w7(32'h3ab81d0b),
	.w8(32'hbb48f02a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2002b1),
	.w1(32'h3bf4d6a8),
	.w2(32'h3ac44387),
	.w3(32'h3b86bb30),
	.w4(32'h37c153ae),
	.w5(32'h3cbe77a4),
	.w6(32'hbaa4cc4a),
	.w7(32'hbb2bad82),
	.w8(32'hbb18cec5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e5a33),
	.w1(32'hbc31bd22),
	.w2(32'hbbd43e0a),
	.w3(32'h3ba55e37),
	.w4(32'h3b16a3d2),
	.w5(32'hbb6f4552),
	.w6(32'h3b9c01c3),
	.w7(32'hba332bab),
	.w8(32'hb9abc502),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40becf),
	.w1(32'hba74e4d9),
	.w2(32'h3c33c8b0),
	.w3(32'h3a065b02),
	.w4(32'hbb9c8b5c),
	.w5(32'hbb4a05c9),
	.w6(32'hbad06af6),
	.w7(32'h39ab9bc0),
	.w8(32'h3b8de95d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfadf36),
	.w1(32'h3a34b4b8),
	.w2(32'h3bf41471),
	.w3(32'hbb9b6b9e),
	.w4(32'hbb7aeeb0),
	.w5(32'hbafd3f0f),
	.w6(32'hbb8a698a),
	.w7(32'h3b476ffe),
	.w8(32'h3ad6ae7a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5c061),
	.w1(32'hb9882729),
	.w2(32'hb9daad0c),
	.w3(32'hba876e2a),
	.w4(32'hbb0957c2),
	.w5(32'hba5109f9),
	.w6(32'hba7b8dc2),
	.w7(32'hba85caf6),
	.w8(32'h39c8f724),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948f44),
	.w1(32'hba89fc5f),
	.w2(32'h3b857cd5),
	.w3(32'h3b877191),
	.w4(32'h3c37d713),
	.w5(32'h3af30f5b),
	.w6(32'hbb922540),
	.w7(32'hba1fb30c),
	.w8(32'h3bf5a324),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae47982),
	.w1(32'hbb434372),
	.w2(32'hbac67a6d),
	.w3(32'h3909eef3),
	.w4(32'hbbe0dcd3),
	.w5(32'hb9802c5d),
	.w6(32'h3b0fdc9d),
	.w7(32'hbb981a56),
	.w8(32'hbbfd7d84),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2e7de),
	.w1(32'hbb8f3648),
	.w2(32'hbb9c0323),
	.w3(32'h3a841b37),
	.w4(32'hbb00a655),
	.w5(32'h3bbeac41),
	.w6(32'hbb770ba0),
	.w7(32'h3b2d580e),
	.w8(32'h3a03c145),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9251b0),
	.w1(32'h3bb4d9a3),
	.w2(32'hba91ab9c),
	.w3(32'h3b829c19),
	.w4(32'hbab5b3c2),
	.w5(32'h3c34d857),
	.w6(32'hbadf5688),
	.w7(32'h3af9ac75),
	.w8(32'hbae31c09),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b723bd),
	.w1(32'hbb30c956),
	.w2(32'h3b36f776),
	.w3(32'h3b4fda8b),
	.w4(32'hbba5cf63),
	.w5(32'hbb495b96),
	.w6(32'h3bb58cae),
	.w7(32'h3ba403f6),
	.w8(32'h3b7b1690),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bfe10),
	.w1(32'hbb03785d),
	.w2(32'hbb307132),
	.w3(32'h3a7791b1),
	.w4(32'hbc26a0c4),
	.w5(32'h38b9b769),
	.w6(32'hbac15d71),
	.w7(32'hbb87db9c),
	.w8(32'hbc16b10f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18aaa2),
	.w1(32'hbb3c21df),
	.w2(32'hbc0d4907),
	.w3(32'h3b1cc232),
	.w4(32'h3a8d1335),
	.w5(32'hba35f670),
	.w6(32'hbbbc1c1f),
	.w7(32'hba9f47af),
	.w8(32'hbbf89c19),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51ea7b),
	.w1(32'h3afed667),
	.w2(32'h3b4a78be),
	.w3(32'hbbc22840),
	.w4(32'h39a85e29),
	.w5(32'hba9b093a),
	.w6(32'hbb7fad17),
	.w7(32'h3b1e7bf7),
	.w8(32'hbb1e38a8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acadd27),
	.w1(32'h3a50d4eb),
	.w2(32'h3bb59a94),
	.w3(32'hbadff470),
	.w4(32'hba13f9ef),
	.w5(32'h3c05bfc1),
	.w6(32'h3b3faada),
	.w7(32'hbbba8737),
	.w8(32'h3bb2cf45),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6272c8),
	.w1(32'h3aa2455c),
	.w2(32'h3bbfb670),
	.w3(32'hbb1765db),
	.w4(32'h3bab7f2b),
	.w5(32'h3ae76d9e),
	.w6(32'h38875f94),
	.w7(32'hba29ce8b),
	.w8(32'h38bcede3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa02ec0),
	.w1(32'h3c48a073),
	.w2(32'h3a4f9d2e),
	.w3(32'h3c0364d8),
	.w4(32'h3c5f4f96),
	.w5(32'h3c812107),
	.w6(32'hbb6e0d47),
	.w7(32'hbc1fd24d),
	.w8(32'hbadfb895),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cd7ea),
	.w1(32'hbb12705b),
	.w2(32'h3b71447a),
	.w3(32'h3b513040),
	.w4(32'hbb92d320),
	.w5(32'hbb953cc7),
	.w6(32'h3bbfba47),
	.w7(32'h3b296ccf),
	.w8(32'h3aa61f05),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b990a25),
	.w1(32'h3bb20bea),
	.w2(32'hbb886920),
	.w3(32'hb9b77822),
	.w4(32'h3b323e0d),
	.w5(32'h3ca3ddb5),
	.w6(32'hbafed31a),
	.w7(32'hbba53c8f),
	.w8(32'h36592665),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1a51d),
	.w1(32'hbb5a4f4b),
	.w2(32'hbc14c4dd),
	.w3(32'h3bc0f539),
	.w4(32'hb9b35532),
	.w5(32'hbba6f3e5),
	.w6(32'h3be4bb0b),
	.w7(32'hbb7e4ab5),
	.w8(32'hbc21259d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb64a24),
	.w1(32'hba95b9ff),
	.w2(32'hbbad7f53),
	.w3(32'hbbb09e1e),
	.w4(32'h3b26cb6c),
	.w5(32'h3bd34290),
	.w6(32'hbb055c1a),
	.w7(32'hbb900aec),
	.w8(32'hb9f40e38),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb603534),
	.w1(32'h38abb453),
	.w2(32'hbbc245ad),
	.w3(32'hbac69cf6),
	.w4(32'hbae9cb6e),
	.w5(32'h3c391893),
	.w6(32'hba2b03e5),
	.w7(32'hbafa1445),
	.w8(32'hb8f3d691),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63c514),
	.w1(32'hbb7cf534),
	.w2(32'hbb8d26df),
	.w3(32'h3a2a9c38),
	.w4(32'hbaf63e06),
	.w5(32'hbb03fb60),
	.w6(32'h3beb58b8),
	.w7(32'hba9956a1),
	.w8(32'h39b240aa),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29555c),
	.w1(32'hbaae5233),
	.w2(32'h3b853538),
	.w3(32'h3af536ed),
	.w4(32'hbb1fc130),
	.w5(32'hbb9849f0),
	.w6(32'h3b6eb2f6),
	.w7(32'h3aa25337),
	.w8(32'h3b06e72c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8960fe),
	.w1(32'h3aebff20),
	.w2(32'hbb8478d2),
	.w3(32'h3b96fbd2),
	.w4(32'h3aa0f3f9),
	.w5(32'h3c51c128),
	.w6(32'hbb5ced0d),
	.w7(32'h3af3fbcf),
	.w8(32'hbaf3665d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80c5e),
	.w1(32'h3bb1e046),
	.w2(32'hbaf7c61d),
	.w3(32'hbb029d60),
	.w4(32'h3c25980f),
	.w5(32'h3cc84f94),
	.w6(32'h3a815cc5),
	.w7(32'hbbdf2bdb),
	.w8(32'hba220014),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34c543),
	.w1(32'hbb84207d),
	.w2(32'hbc38087f),
	.w3(32'h3c313a75),
	.w4(32'h3b3548a1),
	.w5(32'h3cbe5cb6),
	.w6(32'h3c35eebc),
	.w7(32'h3a2f6f7f),
	.w8(32'h3ad61f14),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4c11),
	.w1(32'hbb245843),
	.w2(32'hbb479344),
	.w3(32'hbb348cb0),
	.w4(32'h3b9c4b69),
	.w5(32'h3c0427f5),
	.w6(32'h3b22115f),
	.w7(32'h3bbcad98),
	.w8(32'hbacc7af6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be9767),
	.w1(32'hbb871a33),
	.w2(32'hbbc821d9),
	.w3(32'h393b16b6),
	.w4(32'h3b4b080e),
	.w5(32'hbb22186d),
	.w6(32'hbb993b29),
	.w7(32'hbb826c41),
	.w8(32'hbab355cb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5aead),
	.w1(32'hbb9b8740),
	.w2(32'hbb7525d8),
	.w3(32'h3a4e2959),
	.w4(32'hbadf702d),
	.w5(32'hbba32187),
	.w6(32'h3bc16cd4),
	.w7(32'h3b66c740),
	.w8(32'hbbab14d8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba96aab),
	.w1(32'hbb723dca),
	.w2(32'h3b0853fb),
	.w3(32'hbba40447),
	.w4(32'hbbef0435),
	.w5(32'hbbc3861f),
	.w6(32'h3a9f05c7),
	.w7(32'hba7a0420),
	.w8(32'hb9d3e5e0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba14fe1),
	.w1(32'hbb2d746b),
	.w2(32'h3b9cc39e),
	.w3(32'hbb21ad95),
	.w4(32'hbbc90c30),
	.w5(32'hbb239c33),
	.w6(32'hbbd01994),
	.w7(32'h3b90c392),
	.w8(32'h3aeab74a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcccc65),
	.w1(32'h3b63e565),
	.w2(32'h3a69e2bf),
	.w3(32'hb90568c7),
	.w4(32'h3be26b1a),
	.w5(32'h3b53c35e),
	.w6(32'h3bc04a07),
	.w7(32'h3c02571a),
	.w8(32'h3bf8cbc0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ca671),
	.w1(32'h3b783f8f),
	.w2(32'hbb8fc2dc),
	.w3(32'hba0778af),
	.w4(32'h3b0e37ab),
	.w5(32'h3c0ce9f1),
	.w6(32'h3b8a8a3d),
	.w7(32'h3b4021c9),
	.w8(32'hbb0eb6bd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b057abf),
	.w1(32'hbaa2c042),
	.w2(32'hba0f517f),
	.w3(32'hbb63bf9a),
	.w4(32'hbbdb8557),
	.w5(32'hbb1e50bd),
	.w6(32'h3ab9096f),
	.w7(32'hb9fa562d),
	.w8(32'h3aa76bc2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8385e7),
	.w1(32'hbb3de529),
	.w2(32'h3b73d80f),
	.w3(32'hbbc80d88),
	.w4(32'hbb06a34f),
	.w5(32'hba9c79f9),
	.w6(32'h3b381fff),
	.w7(32'h3b001490),
	.w8(32'h3b1b3621),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03e4a8),
	.w1(32'hbbb2553c),
	.w2(32'hbb102886),
	.w3(32'h3af96b42),
	.w4(32'hbb843d51),
	.w5(32'hbad2891d),
	.w6(32'h3b0a37cf),
	.w7(32'hbad8fedc),
	.w8(32'hbb04d38a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1959),
	.w1(32'hbb9ca488),
	.w2(32'h3ae1df54),
	.w3(32'hbbb22ed1),
	.w4(32'hbbdc6f25),
	.w5(32'hbb1f5cc6),
	.w6(32'h39f85105),
	.w7(32'hbb29828f),
	.w8(32'hbb137d6c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782dcd9),
	.w1(32'hbb8a5962),
	.w2(32'hbb7f0f71),
	.w3(32'hbb06bfcd),
	.w4(32'h3ba90349),
	.w5(32'hbb315022),
	.w6(32'hbbe3c4e0),
	.w7(32'h3c0c3937),
	.w8(32'h3b3ab14f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1a10),
	.w1(32'hbae8ab1d),
	.w2(32'h3ab60815),
	.w3(32'hb9e2ec51),
	.w4(32'hbb4d13c9),
	.w5(32'hbbbf7e88),
	.w6(32'hbb00497f),
	.w7(32'hba38bfa8),
	.w8(32'hbbcb9daa),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f33d0),
	.w1(32'hbb15cbb9),
	.w2(32'hbc084868),
	.w3(32'hbb236b0a),
	.w4(32'hbaac09d3),
	.w5(32'h3b4e7e8a),
	.w6(32'hbb0547e6),
	.w7(32'h39850ecb),
	.w8(32'hbb678036),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9506636),
	.w1(32'h3ba9075e),
	.w2(32'hbbbc351a),
	.w3(32'h3bbbb43b),
	.w4(32'hbaa4b807),
	.w5(32'h3c8faf08),
	.w6(32'h3b811cb4),
	.w7(32'hbb402b2d),
	.w8(32'hbad3e4ed),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97f0e0),
	.w1(32'h3b2ffe33),
	.w2(32'h3af26fd9),
	.w3(32'h3b418abb),
	.w4(32'h3aab2944),
	.w5(32'hbb43ff6e),
	.w6(32'h3c27c49f),
	.w7(32'hba906c05),
	.w8(32'hbb52e9d1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b4ffc),
	.w1(32'hbbbc3d81),
	.w2(32'hbc0de1a9),
	.w3(32'hbb41f557),
	.w4(32'hbc54f95d),
	.w5(32'hbc4c687a),
	.w6(32'hbaa5ea66),
	.w7(32'hbb1a9213),
	.w8(32'hbbcc88da),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3368e7),
	.w1(32'hbb428570),
	.w2(32'hbaf0bb9d),
	.w3(32'hbc57d772),
	.w4(32'hba3ecf98),
	.w5(32'hbb060403),
	.w6(32'hbbe4623a),
	.w7(32'h3a59e90a),
	.w8(32'hbb3b75fe),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule