module layer_10_featuremap_501(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff3943),
	.w1(32'h3a19966d),
	.w2(32'h3ad9b9cb),
	.w3(32'h39a8ca6d),
	.w4(32'hbaaec09d),
	.w5(32'hbaa2f1cd),
	.w6(32'hb989ddd5),
	.w7(32'hbae731b1),
	.w8(32'hbb075ea1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb0a55),
	.w1(32'hba165dd7),
	.w2(32'h3ac3b626),
	.w3(32'h3a899ace),
	.w4(32'h3a747e5d),
	.w5(32'h3aafdb21),
	.w6(32'h3ae72e06),
	.w7(32'hba877602),
	.w8(32'hba0b4bab),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd63a8),
	.w1(32'h3afa8e38),
	.w2(32'h398a295a),
	.w3(32'hbb1012a1),
	.w4(32'h3b8b2fb7),
	.w5(32'h3b040589),
	.w6(32'hbb1dc2e9),
	.w7(32'h3ab70b34),
	.w8(32'h3ae9b99d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07399c),
	.w1(32'hbb3cc208),
	.w2(32'hbafc3d46),
	.w3(32'hb92682a8),
	.w4(32'hbb56071b),
	.w5(32'hbb76e741),
	.w6(32'h3b229b79),
	.w7(32'hbb4d675d),
	.w8(32'hbb508ec4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba566d83),
	.w1(32'hba0d93d2),
	.w2(32'hb91725fc),
	.w3(32'hbb1fccea),
	.w4(32'hb9bbe2fc),
	.w5(32'hba3c9cf7),
	.w6(32'hb926437c),
	.w7(32'hbaa48cfe),
	.w8(32'h399d2e46),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad11d34),
	.w1(32'hba43eded),
	.w2(32'hba7fec8d),
	.w3(32'hb9e9d36e),
	.w4(32'hbb2937a3),
	.w5(32'h3b07e409),
	.w6(32'hba39851b),
	.w7(32'h3abbab5d),
	.w8(32'h3b1ef6bb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b251b8b),
	.w1(32'h3aaa5026),
	.w2(32'h39f63fa3),
	.w3(32'h3aba0078),
	.w4(32'h3b890f61),
	.w5(32'hb97be09d),
	.w6(32'h3b119b9d),
	.w7(32'h3acba04f),
	.w8(32'hbb1ec1e2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba36f84),
	.w1(32'hbbb5d447),
	.w2(32'hbc0bc017),
	.w3(32'hbc15f8f3),
	.w4(32'hbb5ee90b),
	.w5(32'hbb72a182),
	.w6(32'hbc2f8817),
	.w7(32'hbc035d24),
	.w8(32'hbb82eb4e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bce05),
	.w1(32'hbb09c6ce),
	.w2(32'h3aa4aa6c),
	.w3(32'h3a8cd6b0),
	.w4(32'hba8e45bb),
	.w5(32'h3ac8fd61),
	.w6(32'h3ae026ac),
	.w7(32'hbaceceb7),
	.w8(32'h3ae48166),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e8415),
	.w1(32'hba498f67),
	.w2(32'h3b8d9cd8),
	.w3(32'hbae9f0c8),
	.w4(32'hbb0de2bd),
	.w5(32'h3a89de4c),
	.w6(32'h3ad8c5b7),
	.w7(32'hba750579),
	.w8(32'hbb53cdf7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3a917),
	.w1(32'hba9478fb),
	.w2(32'hbb16ce55),
	.w3(32'hbae7a95f),
	.w4(32'hba4863a5),
	.w5(32'hbb14a57e),
	.w6(32'h396ec53e),
	.w7(32'hbb1715d5),
	.w8(32'hbaef2970),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a4ac),
	.w1(32'h3aad8dc0),
	.w2(32'hbb6eeb6a),
	.w3(32'hbaa64d24),
	.w4(32'h3b1575e9),
	.w5(32'h39940b30),
	.w6(32'h3a968db9),
	.w7(32'h3b9f3dc8),
	.w8(32'h3a5a037b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8cdcb),
	.w1(32'h3adc98b1),
	.w2(32'h3b8f96f0),
	.w3(32'hb9dfdd25),
	.w4(32'hb94d344d),
	.w5(32'hb8a66f11),
	.w6(32'h38ad67a6),
	.w7(32'h3a492a68),
	.w8(32'hbb8b6473),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bc02e),
	.w1(32'h3b408728),
	.w2(32'h3aa42687),
	.w3(32'hba7bc4a8),
	.w4(32'h399ef9bd),
	.w5(32'hba3b14a3),
	.w6(32'hb9e2d06f),
	.w7(32'h390a1d5b),
	.w8(32'hb96d6894),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7b0ef),
	.w1(32'hbb0b5231),
	.w2(32'hbabc9722),
	.w3(32'h39f7a43d),
	.w4(32'hbaedc8db),
	.w5(32'h3a7504b6),
	.w6(32'h392edc9c),
	.w7(32'h398de2f7),
	.w8(32'hba95cd4a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3557d),
	.w1(32'h3b40a06e),
	.w2(32'h3a5dbd94),
	.w3(32'hbaf51acc),
	.w4(32'h39b95257),
	.w5(32'hbab76418),
	.w6(32'hbb1b1edc),
	.w7(32'hb9b7d388),
	.w8(32'hbb7f7d4e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51a913),
	.w1(32'hbb29ec8e),
	.w2(32'hba79452f),
	.w3(32'h3a561cbe),
	.w4(32'h39a45fa3),
	.w5(32'hbaa11b4b),
	.w6(32'hba0dd1fe),
	.w7(32'h39f0eb28),
	.w8(32'hba9066d2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f72b0),
	.w1(32'hbb97df37),
	.w2(32'hbbf63c2b),
	.w3(32'hbc1c015a),
	.w4(32'hbbc1f242),
	.w5(32'hbbf655ea),
	.w6(32'hbc0d6006),
	.w7(32'hbc118d1d),
	.w8(32'hbbcb167d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f5c13),
	.w1(32'hbb0cc325),
	.w2(32'hbb15996d),
	.w3(32'hbb02b4da),
	.w4(32'hbb1d681c),
	.w5(32'hbaab72fe),
	.w6(32'hba6590e7),
	.w7(32'hbac618aa),
	.w8(32'hbae1aaa1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1d7bf),
	.w1(32'hbb7512a6),
	.w2(32'hbb889cf5),
	.w3(32'hbafe0dcf),
	.w4(32'hbb0748f7),
	.w5(32'hbbed5417),
	.w6(32'hb99b37a1),
	.w7(32'hb7f12fcc),
	.w8(32'hbbb97bae),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5fb20),
	.w1(32'hba19b07b),
	.w2(32'hb9d072c5),
	.w3(32'hbba65769),
	.w4(32'hbaf2c86c),
	.w5(32'h3b101403),
	.w6(32'hbb808c13),
	.w7(32'hbac08298),
	.w8(32'h3ab51f91),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab70343),
	.w1(32'hbab9cfff),
	.w2(32'hbabaa074),
	.w3(32'h3ac85b3a),
	.w4(32'hbadd40ec),
	.w5(32'h39aec1dd),
	.w6(32'h3acd8494),
	.w7(32'hbaa4f7ca),
	.w8(32'hb97741c4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdafd37),
	.w1(32'hbc17eba2),
	.w2(32'hbc1e0348),
	.w3(32'hbc026007),
	.w4(32'hbc0806d8),
	.w5(32'hbb9b2310),
	.w6(32'hbc535627),
	.w7(32'hbba4afe1),
	.w8(32'hbbb8c0fb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0072f),
	.w1(32'h3815f872),
	.w2(32'h3b15897c),
	.w3(32'h39f603fc),
	.w4(32'hbae3d97b),
	.w5(32'hb909c454),
	.w6(32'h3b2eff26),
	.w7(32'hba7b8f62),
	.w8(32'hbaddff11),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb789a28),
	.w1(32'hba84d6ca),
	.w2(32'h3b3f4aa7),
	.w3(32'hbabc8693),
	.w4(32'h3b2a98bb),
	.w5(32'h3b4ac8a6),
	.w6(32'h3aebe68e),
	.w7(32'h3b0dd360),
	.w8(32'h3aa27245),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb194891),
	.w1(32'hba963c81),
	.w2(32'hba5080ce),
	.w3(32'hbb53c34b),
	.w4(32'h396089d2),
	.w5(32'h39e09abe),
	.w6(32'hbb035158),
	.w7(32'h38421be9),
	.w8(32'hbaf89017),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90a4b2),
	.w1(32'h3b4750eb),
	.w2(32'h3a049e1e),
	.w3(32'h3ac65b91),
	.w4(32'hba369c50),
	.w5(32'h3940f302),
	.w6(32'hbac07ffb),
	.w7(32'hba4bce8e),
	.w8(32'hba186f47),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83ad34),
	.w1(32'hbb06c442),
	.w2(32'h3b1a1f0a),
	.w3(32'h38e550f8),
	.w4(32'h3b3dc09e),
	.w5(32'h3ae866ff),
	.w6(32'h3b7f9cff),
	.w7(32'h3b5019f8),
	.w8(32'h3ac04f9f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5072a8d),
	.w1(32'hbb2eb49d),
	.w2(32'hba4260d8),
	.w3(32'hba961960),
	.w4(32'hb9ff8347),
	.w5(32'h3a044aae),
	.w6(32'h3a453437),
	.w7(32'hba54db51),
	.w8(32'hb81a5132),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f003fc),
	.w1(32'h3bbdc328),
	.w2(32'h3c032ba1),
	.w3(32'h3ad9a71a),
	.w4(32'h3b7578d3),
	.w5(32'h3bd21c77),
	.w6(32'h3bbb6eb4),
	.w7(32'h3bb8beba),
	.w8(32'h3b9bc18b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b7fb7),
	.w1(32'hbbb31c6b),
	.w2(32'hbb6df6b2),
	.w3(32'h3aebe685),
	.w4(32'hbb9c270e),
	.w5(32'hbb6e7e63),
	.w6(32'h3a2530ec),
	.w7(32'hbb4a5edf),
	.w8(32'hbb05cccb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7da811),
	.w1(32'h3a95457a),
	.w2(32'hba43b2da),
	.w3(32'hba57f224),
	.w4(32'h3b270635),
	.w5(32'hb6e1d3e7),
	.w6(32'hbad09078),
	.w7(32'h3a70b526),
	.w8(32'h38bf79be),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e1527),
	.w1(32'hbad07e53),
	.w2(32'hba17dca8),
	.w3(32'hba11dae8),
	.w4(32'hba2e4a61),
	.w5(32'hb9eda323),
	.w6(32'h3a484857),
	.w7(32'hbafd644e),
	.w8(32'hbacfca67),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eca73),
	.w1(32'h3a83c99b),
	.w2(32'h3b8ffd7a),
	.w3(32'hbb0c4812),
	.w4(32'h3b208ebe),
	.w5(32'h3afef6fb),
	.w6(32'h3a84b062),
	.w7(32'h3a7041f6),
	.w8(32'hbb090275),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca32ec),
	.w1(32'hb9cde6f5),
	.w2(32'h3894db37),
	.w3(32'hba35d2cf),
	.w4(32'hb8d0291f),
	.w5(32'h39d6bc0d),
	.w6(32'h3971e3b5),
	.w7(32'hbb3a08ad),
	.w8(32'hbb22097f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab41321),
	.w1(32'hbaa46213),
	.w2(32'hba3192f3),
	.w3(32'hbb135616),
	.w4(32'h391099a5),
	.w5(32'hba2c7f6c),
	.w6(32'hbb56c7dc),
	.w7(32'hbb140352),
	.w8(32'hbb402e24),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01ba00),
	.w1(32'h3b654629),
	.w2(32'h3b0c77aa),
	.w3(32'hbbb37966),
	.w4(32'h3b0534ce),
	.w5(32'h3c12a8dd),
	.w6(32'hbbb4313c),
	.w7(32'h3b8c512e),
	.w8(32'h3b84fdb9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57b232),
	.w1(32'hbb78f2d9),
	.w2(32'h3b12508c),
	.w3(32'h3ba319ac),
	.w4(32'h3c0791fb),
	.w5(32'h3bcfc045),
	.w6(32'h3bd1c1b2),
	.w7(32'h3bcd9322),
	.w8(32'h3ba936f3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ef92f),
	.w1(32'h3b11096d),
	.w2(32'h3b9ceed0),
	.w3(32'h3bed1682),
	.w4(32'h3bc12873),
	.w5(32'h3bf85005),
	.w6(32'h3c3c3cc2),
	.w7(32'h3b99c936),
	.w8(32'h3bd488a8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa41c6a),
	.w1(32'hbaadad7d),
	.w2(32'hb9d5d2e7),
	.w3(32'h3a8d097a),
	.w4(32'h3b170b9a),
	.w5(32'h3b194e77),
	.w6(32'h3aff98fd),
	.w7(32'h3b010351),
	.w8(32'hba04e6dd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d8cfe),
	.w1(32'hba36fa44),
	.w2(32'hbb038ae1),
	.w3(32'h3a67d3ce),
	.w4(32'hbb67347b),
	.w5(32'h399694a7),
	.w6(32'h37a671ea),
	.w7(32'hbaeccb5e),
	.w8(32'hbb44f4a1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb022ae1),
	.w1(32'hb8aeaf67),
	.w2(32'hb94900ba),
	.w3(32'hbaee63e1),
	.w4(32'hba0af3a8),
	.w5(32'h3abee7ab),
	.w6(32'hbb24ace6),
	.w7(32'hbacca9a7),
	.w8(32'hba8f330b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba545967),
	.w1(32'h3b2d9a15),
	.w2(32'h3b3d105a),
	.w3(32'hbac0c2ea),
	.w4(32'h3b33df2d),
	.w5(32'h3aa431b0),
	.w6(32'hbabe256a),
	.w7(32'h3af1ae46),
	.w8(32'h3a13ccd6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61f338),
	.w1(32'h3b106772),
	.w2(32'h3abdad48),
	.w3(32'hbb2ed958),
	.w4(32'hbaa184c8),
	.w5(32'hbb79ff18),
	.w6(32'hbac635dc),
	.w7(32'hbb0d54f3),
	.w8(32'hbbc16724),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18536e),
	.w1(32'hbaa13cb6),
	.w2(32'h3b5f1b2d),
	.w3(32'hb9cb4454),
	.w4(32'h3a76ff55),
	.w5(32'h3b4d86c5),
	.w6(32'h3b1b021c),
	.w7(32'h3b06f591),
	.w8(32'h3a9c076e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ae7d9),
	.w1(32'h3ae101cc),
	.w2(32'h3b6bcec2),
	.w3(32'hbb01cbab),
	.w4(32'h393a8376),
	.w5(32'h3b473002),
	.w6(32'h3ae5034b),
	.w7(32'h39c97b8b),
	.w8(32'h3a0b3d12),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac34cf3),
	.w1(32'hbb1acdc8),
	.w2(32'hba7d3cf8),
	.w3(32'h3a13a7ae),
	.w4(32'hbabbdbbb),
	.w5(32'h3ac3eafd),
	.w6(32'hba81a132),
	.w7(32'hbb2d5872),
	.w8(32'h39d2b1e7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9958c3),
	.w1(32'hbbc6af5f),
	.w2(32'hbc302e7a),
	.w3(32'hbba174d4),
	.w4(32'hbbf2f8f9),
	.w5(32'hbc2253ff),
	.w6(32'hbc08ba2b),
	.w7(32'hbc2f31df),
	.w8(32'hbc26f0db),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8194fd),
	.w1(32'h3b25dc73),
	.w2(32'h3ad83177),
	.w3(32'hbb0e2cbd),
	.w4(32'h3a6a0ef0),
	.w5(32'h3aa6ca46),
	.w6(32'hbb0b1b19),
	.w7(32'h3a3c6db7),
	.w8(32'h3ab14f15),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6d732),
	.w1(32'h3add264e),
	.w2(32'hb9181664),
	.w3(32'hba3f47bb),
	.w4(32'h3aebbc8e),
	.w5(32'h3af34607),
	.w6(32'hbaf6148c),
	.w7(32'h3a6324c6),
	.w8(32'h399a2feb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1a243),
	.w1(32'hbb171bdb),
	.w2(32'hbb5f377b),
	.w3(32'h3a95dd8f),
	.w4(32'hbb321862),
	.w5(32'hbb2e36bb),
	.w6(32'h39a9ca20),
	.w7(32'hbb08c5d2),
	.w8(32'hba8a67dc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe38690),
	.w1(32'hbb092b67),
	.w2(32'hbad9a9ff),
	.w3(32'hbb2295f2),
	.w4(32'hbab30d10),
	.w5(32'hbadd5766),
	.w6(32'hba9f318a),
	.w7(32'hbb4c8570),
	.w8(32'hbb887476),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e937f),
	.w1(32'h3b5f6c9b),
	.w2(32'h3ade1218),
	.w3(32'hbb5b94c0),
	.w4(32'h3ae6617a),
	.w5(32'h3b243a08),
	.w6(32'hbb6fc8b8),
	.w7(32'h3a75c68d),
	.w8(32'h3b6f1952),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a082b),
	.w1(32'h3a5d84f8),
	.w2(32'hbabdcf70),
	.w3(32'hbb81c59c),
	.w4(32'hbb87d791),
	.w5(32'hbb10b48f),
	.w6(32'hbb544652),
	.w7(32'hbb80ecac),
	.w8(32'hb9d25391),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe9c62),
	.w1(32'hbb34b798),
	.w2(32'hba8a781a),
	.w3(32'h39b9080b),
	.w4(32'h3b49e62c),
	.w5(32'h3b4c8e61),
	.w6(32'h3a9fb55a),
	.w7(32'h3a9a1220),
	.w8(32'hb9de879c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86604c),
	.w1(32'h3a81fa04),
	.w2(32'h3b96e422),
	.w3(32'h3967d9a9),
	.w4(32'h3aec60f2),
	.w5(32'h3babcd9d),
	.w6(32'h38895f11),
	.w7(32'h3a866014),
	.w8(32'h3b19f619),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0deeec),
	.w1(32'h3a87ef31),
	.w2(32'h3a797db5),
	.w3(32'hbaad5ad9),
	.w4(32'hba2a0b87),
	.w5(32'h3a2fda56),
	.w6(32'hb9634acd),
	.w7(32'hb9de4696),
	.w8(32'h3afdae89),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a75e6d),
	.w1(32'hba293749),
	.w2(32'hbb1cf0e5),
	.w3(32'hb88ea0d7),
	.w4(32'hba85b704),
	.w5(32'hba8ed129),
	.w6(32'h3b0d779c),
	.w7(32'hbb0a98b7),
	.w8(32'hb9bfeed9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7da5a5),
	.w1(32'h3ab98f7c),
	.w2(32'hbaa31ecd),
	.w3(32'h3a28dd80),
	.w4(32'h3add03d9),
	.w5(32'h3a6fffc5),
	.w6(32'h3999281c),
	.w7(32'h3a51bcaf),
	.w8(32'hba8a12b5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0d3c),
	.w1(32'hbb4a0b78),
	.w2(32'hbab40f21),
	.w3(32'h39d46872),
	.w4(32'hba910ba8),
	.w5(32'hbb7fcead),
	.w6(32'hbaa6626e),
	.w7(32'hbb7a9bef),
	.w8(32'hb9a33dcd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabed632),
	.w1(32'hbb30a55f),
	.w2(32'hbb6f5149),
	.w3(32'hbb42876f),
	.w4(32'hbb254709),
	.w5(32'h39480632),
	.w6(32'hbaec4e5c),
	.w7(32'hbb986f1e),
	.w8(32'hbb61b662),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb696379),
	.w1(32'hbb860071),
	.w2(32'hbb26fe1f),
	.w3(32'hbbabee8d),
	.w4(32'hbb529dd8),
	.w5(32'hbb24fa04),
	.w6(32'hbb8cb01d),
	.w7(32'hbb206419),
	.w8(32'hbae6a0f4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae04de5),
	.w1(32'hba977575),
	.w2(32'hba27b94b),
	.w3(32'hbabf88f3),
	.w4(32'hba8c5369),
	.w5(32'hbad97eca),
	.w6(32'hba0cfdc9),
	.w7(32'hbaeac046),
	.w8(32'hbaa92cd0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba956875),
	.w1(32'h3a93e7ae),
	.w2(32'hba18fe5f),
	.w3(32'hbaea39f9),
	.w4(32'hba019339),
	.w5(32'h3a58e822),
	.w6(32'h39e5cc7b),
	.w7(32'h3ad42bc4),
	.w8(32'h3b340f4b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb867875b),
	.w1(32'h3b9c605b),
	.w2(32'h3b908598),
	.w3(32'h3ac84b36),
	.w4(32'h3ba921e8),
	.w5(32'h3b2caad8),
	.w6(32'h3a8f6383),
	.w7(32'h3bbe1bf1),
	.w8(32'h3b95611c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74763b),
	.w1(32'h3b5a5567),
	.w2(32'h3b73c11d),
	.w3(32'h3b668caa),
	.w4(32'h3ae93bf0),
	.w5(32'h3b0b9266),
	.w6(32'h3b80bf7f),
	.w7(32'h394761d8),
	.w8(32'hba115a91),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9562fb),
	.w1(32'hba2fc444),
	.w2(32'hbb008316),
	.w3(32'h39e5d666),
	.w4(32'hbafe2567),
	.w5(32'hbb251c4c),
	.w6(32'hbad07e37),
	.w7(32'h397d4fcb),
	.w8(32'hb97533ab),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba393da3),
	.w1(32'h3b850c40),
	.w2(32'h3bfb8a04),
	.w3(32'h3935a9c9),
	.w4(32'h3b83338f),
	.w5(32'h3bd5cdc8),
	.w6(32'hba669428),
	.w7(32'hbb250b71),
	.w8(32'hbb6f8c69),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40bc27),
	.w1(32'hbc10fc24),
	.w2(32'hbbf845d9),
	.w3(32'hbb811cff),
	.w4(32'hbb475bcb),
	.w5(32'hbb4e5de0),
	.w6(32'hbb5bbdc1),
	.w7(32'hbc16ce73),
	.w8(32'hbb969e41),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a15da),
	.w1(32'h3c079bd1),
	.w2(32'h3bf2962f),
	.w3(32'h3a2c9e04),
	.w4(32'h3c120f10),
	.w5(32'h3c3ad02e),
	.w6(32'h3ba3eb27),
	.w7(32'h3bc54d00),
	.w8(32'h3bc6f3f5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9a87f),
	.w1(32'hbb10652a),
	.w2(32'hbae14b8c),
	.w3(32'h3b3a645e),
	.w4(32'hbb1f917e),
	.w5(32'hbaaba181),
	.w6(32'h3b06503f),
	.w7(32'hbb561355),
	.w8(32'hbaeb9270),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015e72),
	.w1(32'hbb1ef997),
	.w2(32'hbb409d8b),
	.w3(32'hbaaa56fa),
	.w4(32'hbb223e4c),
	.w5(32'hbb481a69),
	.w6(32'hbb0a7bd6),
	.w7(32'h38e150bc),
	.w8(32'h3b038bf7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e84df7),
	.w1(32'h3a93790c),
	.w2(32'h3a3665a1),
	.w3(32'h3a9aa9e2),
	.w4(32'h3b43d82d),
	.w5(32'h3b1831d7),
	.w6(32'h3bceafea),
	.w7(32'h3aba3df5),
	.w8(32'h3b3da4b1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe079f4),
	.w1(32'hbb52d9f2),
	.w2(32'hbb6bb575),
	.w3(32'hbbcc8a40),
	.w4(32'hbb1e1aa5),
	.w5(32'hbab6ff66),
	.w6(32'hbbcfd2a1),
	.w7(32'hba824981),
	.w8(32'h38e6c456),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a8797),
	.w1(32'hbb314260),
	.w2(32'hbb7d08d1),
	.w3(32'h3a7ceff8),
	.w4(32'hba34095d),
	.w5(32'hba79254c),
	.w6(32'h3ae26c3c),
	.w7(32'hb92d9726),
	.w8(32'h3a3925ae),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833fb9),
	.w1(32'hbabd004e),
	.w2(32'hbb900a9f),
	.w3(32'hbaf773b3),
	.w4(32'hbb216ec1),
	.w5(32'hbb0aa37f),
	.w6(32'hbb402145),
	.w7(32'hba1c987d),
	.w8(32'h3a733b61),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b080424),
	.w1(32'h39ff10ca),
	.w2(32'hbbcc156c),
	.w3(32'hba3e20a7),
	.w4(32'hbb1cbcaf),
	.w5(32'hbba5eb3e),
	.w6(32'hbb817f04),
	.w7(32'hbb8cf2dc),
	.w8(32'hbb618d21),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6112c6),
	.w1(32'hba9e47b3),
	.w2(32'hbb06d5db),
	.w3(32'h3b7b64e3),
	.w4(32'h3a88d181),
	.w5(32'hbb112213),
	.w6(32'h3b9b758e),
	.w7(32'h3939ffce),
	.w8(32'hbb497745),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7441e7),
	.w1(32'hbb061760),
	.w2(32'hbada7c3a),
	.w3(32'hbbb7e983),
	.w4(32'hbb20a307),
	.w5(32'hbb6f8457),
	.w6(32'hbbc02acd),
	.w7(32'hbb89601c),
	.w8(32'hbb9633d8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb6715),
	.w1(32'h3ae3b69c),
	.w2(32'h39d34b64),
	.w3(32'hbb003872),
	.w4(32'h3b343c7f),
	.w5(32'h3a81e9b4),
	.w6(32'hba75c1b1),
	.w7(32'h3b6043fc),
	.w8(32'h3a1208c1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa19a3c),
	.w1(32'h3c60a569),
	.w2(32'h3c3ba86d),
	.w3(32'h3a9b6168),
	.w4(32'h3c63bd82),
	.w5(32'h3c2135a3),
	.w6(32'h3a8ac972),
	.w7(32'h3c351684),
	.w8(32'h3c05143d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c498c53),
	.w1(32'h3b028eb4),
	.w2(32'hbacc9b24),
	.w3(32'h3c4353f3),
	.w4(32'h3b860c5f),
	.w5(32'h3a4ac8e9),
	.w6(32'h3c0c94dc),
	.w7(32'h3b5fa342),
	.w8(32'h3a7d3aa9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21d602),
	.w1(32'h3af82c60),
	.w2(32'hba076749),
	.w3(32'hb7deb390),
	.w4(32'hbac148ea),
	.w5(32'hbba50459),
	.w6(32'h39829112),
	.w7(32'hbb7be32e),
	.w8(32'hbbd1b7ef),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa535b5),
	.w1(32'h3a42ff8f),
	.w2(32'hbadfc093),
	.w3(32'hbb35bc16),
	.w4(32'hbb337a9a),
	.w5(32'hbaf5ffb6),
	.w6(32'hbb775504),
	.w7(32'hbb40a6b6),
	.w8(32'hbb718eb1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c0c94),
	.w1(32'hbb1f5324),
	.w2(32'hbb4357d2),
	.w3(32'hbafa21d2),
	.w4(32'hbb11317b),
	.w5(32'hbb1c2619),
	.w6(32'hbb7d6f97),
	.w7(32'hbb37697c),
	.w8(32'hbb130438),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917cc2),
	.w1(32'hbafb5d4c),
	.w2(32'hb98a6a88),
	.w3(32'hbb285ab6),
	.w4(32'hbb0d7df8),
	.w5(32'h39b420e6),
	.w6(32'hbb1e67d1),
	.w7(32'hb84e1ac9),
	.w8(32'h3aa056fa),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5feb95),
	.w1(32'hba82f002),
	.w2(32'h3b054beb),
	.w3(32'h3a30cb69),
	.w4(32'h3a803659),
	.w5(32'h3a714e40),
	.w6(32'h3b98132d),
	.w7(32'hbb2ebbae),
	.w8(32'hbb0380cc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83353a),
	.w1(32'h3a8df4d4),
	.w2(32'h3a889fde),
	.w3(32'h3a31c91a),
	.w4(32'h3a503ed8),
	.w5(32'hba3444ef),
	.w6(32'hbabf92f9),
	.w7(32'h3a965dad),
	.w8(32'hbaf4b5a2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8b46),
	.w1(32'hba2dc4ab),
	.w2(32'h39f082af),
	.w3(32'hbb4b6502),
	.w4(32'hbb6d6fca),
	.w5(32'hbb0f3d7b),
	.w6(32'hbb8259f7),
	.w7(32'hbb482ff4),
	.w8(32'hbb31c0c9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9644d0),
	.w1(32'hbbaa614c),
	.w2(32'hbbb577d0),
	.w3(32'hbc2a494b),
	.w4(32'hbbf1b0c7),
	.w5(32'hbbcf6b17),
	.w6(32'hbc6c706a),
	.w7(32'hbbe61aec),
	.w8(32'hbbe41416),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7f942),
	.w1(32'h3b8dcae9),
	.w2(32'h3a570b54),
	.w3(32'h3b2e1843),
	.w4(32'h3bc65ac9),
	.w5(32'h3a828374),
	.w6(32'h3adcaef1),
	.w7(32'h3b74f846),
	.w8(32'h37b63cd4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb022),
	.w1(32'h3b114777),
	.w2(32'h3adfc157),
	.w3(32'hbbcea1f9),
	.w4(32'h3afcbe01),
	.w5(32'h3b8ac01f),
	.w6(32'hbb7b21d8),
	.w7(32'h3b96a2b6),
	.w8(32'h3b14e516),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950211c),
	.w1(32'h3b8ca44d),
	.w2(32'h3bd248f0),
	.w3(32'h3a863e56),
	.w4(32'h3b5ad282),
	.w5(32'h3ba39cb4),
	.w6(32'h3af2d7bc),
	.w7(32'h3a81f14e),
	.w8(32'h3b1881cb),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bf49c),
	.w1(32'hbb0f41ea),
	.w2(32'hbb255360),
	.w3(32'hbb8deeb8),
	.w4(32'hbb869c84),
	.w5(32'hbb09c15d),
	.w6(32'hbb295347),
	.w7(32'hbbd3885e),
	.w8(32'hbbaf48d8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e5e76),
	.w1(32'h3afb8166),
	.w2(32'h3b3cc92a),
	.w3(32'hb8d4f981),
	.w4(32'hbac7e707),
	.w5(32'hba07185f),
	.w6(32'h3aa4048b),
	.w7(32'hbaa95b08),
	.w8(32'hbb10d39a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a59ea),
	.w1(32'hbbd5d67e),
	.w2(32'hbb48f62a),
	.w3(32'h39d7377c),
	.w4(32'hbbb16117),
	.w5(32'h3a8fe4f2),
	.w6(32'hba95e2fe),
	.w7(32'hbb17f739),
	.w8(32'h3a1d8b0e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfa752),
	.w1(32'hbae74b36),
	.w2(32'hbb436361),
	.w3(32'hba976dc6),
	.w4(32'hbb36adf5),
	.w5(32'hbb4d4f67),
	.w6(32'hb9b61f5d),
	.w7(32'hbaa1b739),
	.w8(32'hbb7f5649),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfda5b),
	.w1(32'hbad15060),
	.w2(32'h3a99d0d0),
	.w3(32'hbbb3754b),
	.w4(32'hbb662708),
	.w5(32'hbae2d9c9),
	.w6(32'hbba4bb72),
	.w7(32'hbb4f8700),
	.w8(32'hbb6f69ec),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba517e6d),
	.w1(32'h3bf02c53),
	.w2(32'h3c0993ea),
	.w3(32'h3b6ac6b7),
	.w4(32'h3c1c27c6),
	.w5(32'h3c6e0c0a),
	.w6(32'h3b753ee6),
	.w7(32'h3bf12aec),
	.w8(32'h3c1796de),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b5ce6),
	.w1(32'hbc1a0ef4),
	.w2(32'hbc311427),
	.w3(32'hbbd632bb),
	.w4(32'hbc3e5afc),
	.w5(32'hbbce30bf),
	.w6(32'hbb59e95e),
	.w7(32'hbc123016),
	.w8(32'hbb8b16f6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcc6ef),
	.w1(32'h3a4e825c),
	.w2(32'h3b2cac7f),
	.w3(32'h3adf708f),
	.w4(32'h3b989e76),
	.w5(32'h3ba9ca90),
	.w6(32'hb9cd96c0),
	.w7(32'h3b0c8187),
	.w8(32'h3ba2244c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7f2fc),
	.w1(32'h3b999a99),
	.w2(32'h3c1d20f2),
	.w3(32'hbaa5364d),
	.w4(32'h3b8a08b0),
	.w5(32'h3bfc195b),
	.w6(32'h3941b696),
	.w7(32'h3b97d821),
	.w8(32'h3b92ea19),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965f3e9),
	.w1(32'hbb11adaf),
	.w2(32'hbbf1b17e),
	.w3(32'h3ac2b0e9),
	.w4(32'hbab00b52),
	.w5(32'hbb3c9a3b),
	.w6(32'h3ac12598),
	.w7(32'h392c8f93),
	.w8(32'hbb4d0dbf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac97ed),
	.w1(32'h3aff6fcd),
	.w2(32'h3b3ad2ba),
	.w3(32'h3a8a11bd),
	.w4(32'h3aab22b0),
	.w5(32'h3a2c7528),
	.w6(32'h3a6506a1),
	.w7(32'h3aadb9a6),
	.w8(32'hba1c270b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb2801),
	.w1(32'h3b936a22),
	.w2(32'hbb49161a),
	.w3(32'hbc078e79),
	.w4(32'hbbc09b40),
	.w5(32'hbba6e177),
	.w6(32'hbc471372),
	.w7(32'hbbadc725),
	.w8(32'hba780fa0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b9a0),
	.w1(32'h3b15b51d),
	.w2(32'h3b1e8cc8),
	.w3(32'h3b867edb),
	.w4(32'h3b5c87df),
	.w5(32'h3aa209c2),
	.w6(32'h3b4bdc17),
	.w7(32'h3b0b05f3),
	.w8(32'h399ff5ee),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefb4ee),
	.w1(32'hbb83773e),
	.w2(32'hbb69ebe6),
	.w3(32'hbb65978c),
	.w4(32'hbb17e1a2),
	.w5(32'hbb64cde4),
	.w6(32'hbb90f2a4),
	.w7(32'hbb075499),
	.w8(32'hbb042ccc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9246),
	.w1(32'hbabb7ec4),
	.w2(32'hbbbc26c2),
	.w3(32'hbb144843),
	.w4(32'hbada03f9),
	.w5(32'hbb8b3d4e),
	.w6(32'h3939307e),
	.w7(32'h39abcfd2),
	.w8(32'hbb6599a8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb645d14),
	.w1(32'h3c5832b3),
	.w2(32'h3c534b1b),
	.w3(32'hbb665e38),
	.w4(32'h3ba05cb0),
	.w5(32'h3ba50b32),
	.w6(32'hbb36d77e),
	.w7(32'h3b433213),
	.w8(32'h3b04504c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb6438),
	.w1(32'h3a1290ac),
	.w2(32'h3b13d458),
	.w3(32'h3c04099e),
	.w4(32'hbb2d76c2),
	.w5(32'hba53f37c),
	.w6(32'h3c19c7c8),
	.w7(32'hbb680a57),
	.w8(32'hbb4f8cf2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5c079),
	.w1(32'hbacbbffc),
	.w2(32'h3ab4c18f),
	.w3(32'hbb7ef463),
	.w4(32'h3b3e7f95),
	.w5(32'h3adec328),
	.w6(32'hbae04502),
	.w7(32'h3beb2725),
	.w8(32'h3c0e9692),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b196f),
	.w1(32'hbb07e8c8),
	.w2(32'hb9d91dd3),
	.w3(32'h3b60918c),
	.w4(32'hbac94b10),
	.w5(32'hbac48a3a),
	.w6(32'h3c423d22),
	.w7(32'hba47416a),
	.w8(32'hbab0d1c5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab82d86),
	.w1(32'h3be5c8e1),
	.w2(32'h3c324719),
	.w3(32'hbba329f4),
	.w4(32'h3c25ed3a),
	.w5(32'h3c867f11),
	.w6(32'hba8ccb5e),
	.w7(32'h3c41b9f7),
	.w8(32'h3c49e99d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bddd5),
	.w1(32'hbbb12a1a),
	.w2(32'hbbcb526a),
	.w3(32'h3be6b4bd),
	.w4(32'hbc0209e3),
	.w5(32'hbbf55c37),
	.w6(32'h3b898766),
	.w7(32'hbbcced69),
	.w8(32'hbb8e6494),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dfbf8),
	.w1(32'h3c0b144e),
	.w2(32'h3c2a48fc),
	.w3(32'hbb275575),
	.w4(32'h3c04553a),
	.w5(32'h3c27a642),
	.w6(32'h3afef0d6),
	.w7(32'h3c04c656),
	.w8(32'h3c0c8305),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf68a00),
	.w1(32'h3a46f0c8),
	.w2(32'hbb5369f6),
	.w3(32'h3c1686bd),
	.w4(32'hb9058785),
	.w5(32'hbb5bfcfb),
	.w6(32'h3c1f3728),
	.w7(32'hbaca4e38),
	.w8(32'hbb9a22d8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f806d),
	.w1(32'h3ac7b03a),
	.w2(32'h3ac8fbc9),
	.w3(32'hbb9d0393),
	.w4(32'h3b12285d),
	.w5(32'h3b870289),
	.w6(32'hbbc53c0a),
	.w7(32'h3b4b7c8e),
	.w8(32'h3b7558c9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17e926),
	.w1(32'h3a10d23c),
	.w2(32'hb9930961),
	.w3(32'h39aea59b),
	.w4(32'h3af7f788),
	.w5(32'hba7efc80),
	.w6(32'h3b006e9a),
	.w7(32'h3b148f28),
	.w8(32'h3a89a121),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8422f9),
	.w1(32'hbaa47112),
	.w2(32'hba853cf7),
	.w3(32'h3b4a097a),
	.w4(32'h36fecf3a),
	.w5(32'h3a26d4ec),
	.w6(32'h3bb3edcf),
	.w7(32'h3b04860c),
	.w8(32'h3a573796),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11e216),
	.w1(32'h3ab00a4a),
	.w2(32'hb9648b17),
	.w3(32'hb9001f7b),
	.w4(32'h3aaf4e83),
	.w5(32'hbaac0acb),
	.w6(32'h3a818127),
	.w7(32'h3ae9d38a),
	.w8(32'hb9f4e713),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9859a5),
	.w1(32'h3b820d6c),
	.w2(32'h3aaf90bd),
	.w3(32'hbb8b2c3a),
	.w4(32'h3b731923),
	.w5(32'h3ae23882),
	.w6(32'hbaddce97),
	.w7(32'h3b11a739),
	.w8(32'h3ae9d1b7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87e37c),
	.w1(32'h3b80018f),
	.w2(32'hbb7db94b),
	.w3(32'hb825f2f1),
	.w4(32'hbb159743),
	.w5(32'hbba13219),
	.w6(32'hba2674c8),
	.w7(32'hbb9b302c),
	.w8(32'hbb810ac1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6be46),
	.w1(32'h3a0e9122),
	.w2(32'h3ade08bb),
	.w3(32'hba126e1b),
	.w4(32'h3a759bd9),
	.w5(32'h3a93858e),
	.w6(32'h3af1f65e),
	.w7(32'hba95589b),
	.w8(32'hbb29d627),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391be31a),
	.w1(32'hbac3858d),
	.w2(32'h3a991590),
	.w3(32'hbaf85e58),
	.w4(32'hbb403c1d),
	.w5(32'h3ad170b1),
	.w6(32'hbafb1e25),
	.w7(32'hb9f08ede),
	.w8(32'h3ada646e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf317a9),
	.w1(32'h3a9b0850),
	.w2(32'hbb030823),
	.w3(32'hbaf2e616),
	.w4(32'hba38ae6b),
	.w5(32'hbb374b8d),
	.w6(32'hba2d5411),
	.w7(32'h3abd68dc),
	.w8(32'h3afdadd6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0482a7),
	.w1(32'h3aa41e78),
	.w2(32'h3adadc97),
	.w3(32'h3b029c75),
	.w4(32'hb948f7fa),
	.w5(32'hb94f2585),
	.w6(32'h3bd3ac10),
	.w7(32'hb8d73a2a),
	.w8(32'h3a303c92),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39134872),
	.w1(32'hbbcefd0b),
	.w2(32'hbba09523),
	.w3(32'h3a13d74a),
	.w4(32'hbb98b69d),
	.w5(32'hbb918d07),
	.w6(32'h3aaf3358),
	.w7(32'hbb865156),
	.w8(32'hbb5d5b30),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaff27b),
	.w1(32'h3b75ceda),
	.w2(32'h3b293036),
	.w3(32'hbbde32e6),
	.w4(32'h3b84a380),
	.w5(32'h3b388135),
	.w6(32'hbbfabb40),
	.w7(32'h3ae3bb4e),
	.w8(32'hbb1785a9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97459b),
	.w1(32'h3b88a424),
	.w2(32'h3b98aadd),
	.w3(32'h39615ef9),
	.w4(32'hbab0d158),
	.w5(32'h39dd7cfd),
	.w6(32'hb7bf2a13),
	.w7(32'hbaf9ff59),
	.w8(32'hba05fe26),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1a8ba),
	.w1(32'hb905e4e9),
	.w2(32'h3a418428),
	.w3(32'h3b2b3f8c),
	.w4(32'hba737f69),
	.w5(32'hb8fb6b3e),
	.w6(32'h3ab03fa4),
	.w7(32'hb98cc17b),
	.w8(32'h397d4ff0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a629f9a),
	.w1(32'h38a93ae2),
	.w2(32'hbb8affda),
	.w3(32'hb93bc9f8),
	.w4(32'hba907fc2),
	.w5(32'hbbae691a),
	.w6(32'h3a7c31a8),
	.w7(32'hbab4aec7),
	.w8(32'hbb7d397a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4890c8),
	.w1(32'hbb3e4b2a),
	.w2(32'hbabe7e06),
	.w3(32'hbb21bdac),
	.w4(32'hbb83a9c5),
	.w5(32'hbb5665dd),
	.w6(32'h3a323f97),
	.w7(32'hbb0a9346),
	.w8(32'hba091c45),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f5ffb),
	.w1(32'h3a8c550e),
	.w2(32'h3b3fc70a),
	.w3(32'hbb5f504c),
	.w4(32'hbb331506),
	.w5(32'hb8b31e03),
	.w6(32'h39dc0ddb),
	.w7(32'hbb00b22f),
	.w8(32'hbaa468f4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b259fa4),
	.w1(32'h3b3852f5),
	.w2(32'h3bb20888),
	.w3(32'h3af0d33f),
	.w4(32'h3b6a1aed),
	.w5(32'h3bf43805),
	.w6(32'h3b03c723),
	.w7(32'h3b57bf1f),
	.w8(32'h3b7c4e44),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75ae1f),
	.w1(32'hbb764532),
	.w2(32'hbb9cf4a8),
	.w3(32'hba3e29e0),
	.w4(32'hbb2a1eb1),
	.w5(32'h3a34174a),
	.w6(32'hbb240b0b),
	.w7(32'h39e94e96),
	.w8(32'h3b1b4277),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3160b6),
	.w1(32'hba3bb918),
	.w2(32'hbafe472e),
	.w3(32'h3bbad230),
	.w4(32'h3b1b17b4),
	.w5(32'h3aabdf00),
	.w6(32'h3bc99b83),
	.w7(32'h384fb092),
	.w8(32'hbaebe032),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb73e50),
	.w1(32'hbad17d11),
	.w2(32'h3ae5962d),
	.w3(32'hbb3d650a),
	.w4(32'h39b42aca),
	.w5(32'h3b3a138a),
	.w6(32'hbb6b3948),
	.w7(32'h37cdf1ff),
	.w8(32'h3b04b55e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2a764),
	.w1(32'hba22b64c),
	.w2(32'hbbd8fbaa),
	.w3(32'hbb00ddc6),
	.w4(32'hbbb5cf7c),
	.w5(32'hbc169c03),
	.w6(32'hbb6bfaca),
	.w7(32'hbbd1117d),
	.w8(32'hbc08be8b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb57ce7),
	.w1(32'hbb04511a),
	.w2(32'hbb3983f1),
	.w3(32'hbbb94fc1),
	.w4(32'hbb05d74e),
	.w5(32'hbaef81b3),
	.w6(32'hbb8a79b1),
	.w7(32'hba81d40f),
	.w8(32'hb9fde52d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf42731),
	.w1(32'h3b966a41),
	.w2(32'h3b8d6d39),
	.w3(32'hbb4a1b66),
	.w4(32'h3b63ad8c),
	.w5(32'h3b752c21),
	.w6(32'hba7acbc0),
	.w7(32'h3b813b1f),
	.w8(32'h3b13d73f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0ab60),
	.w1(32'hba9536de),
	.w2(32'hbb695aa7),
	.w3(32'h39b84381),
	.w4(32'hbb332841),
	.w5(32'hbbc1b69d),
	.w6(32'h38726872),
	.w7(32'hbb91b2a1),
	.w8(32'hbbdc9ac4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe329d7),
	.w1(32'h3b83a1a2),
	.w2(32'h3b8e5cd1),
	.w3(32'hbb5da002),
	.w4(32'h3b929679),
	.w5(32'h3b279b37),
	.w6(32'hbacd367b),
	.w7(32'h3b1ad536),
	.w8(32'hb9a9ae4c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba183b60),
	.w1(32'hbb9de147),
	.w2(32'hbbc6465b),
	.w3(32'hbb0a9027),
	.w4(32'hbb9de86e),
	.w5(32'hbb8c2b30),
	.w6(32'hbb808757),
	.w7(32'hbba4fec3),
	.w8(32'hbb282684),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39f280),
	.w1(32'hba8317ea),
	.w2(32'hbb716d19),
	.w3(32'hbb13bf12),
	.w4(32'h3a290d86),
	.w5(32'hbaebf072),
	.w6(32'hba9e0c86),
	.w7(32'hb9916a2c),
	.w8(32'hbb3c1a17),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acd5ec),
	.w1(32'h3a2b9d42),
	.w2(32'hb97815cd),
	.w3(32'h3a9e6073),
	.w4(32'h3b3db088),
	.w5(32'h3af6d1a5),
	.w6(32'h399e4bdd),
	.w7(32'h3bb3f0f5),
	.w8(32'h3bca7972),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918881c),
	.w1(32'h3abfcf90),
	.w2(32'h3b0b4963),
	.w3(32'h3b3f01ca),
	.w4(32'h3b4dd07e),
	.w5(32'h3b67b734),
	.w6(32'h3be4da70),
	.w7(32'h3b6ac685),
	.w8(32'h3bab9f0b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf66016),
	.w1(32'hbb757506),
	.w2(32'hbb75df6b),
	.w3(32'hb961a214),
	.w4(32'hbb7748bc),
	.w5(32'hbb159570),
	.w6(32'hb8bd263b),
	.w7(32'hbb923481),
	.w8(32'hbb576913),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab457f2),
	.w1(32'hbb6e3598),
	.w2(32'hbbd2af28),
	.w3(32'h3a35f0c6),
	.w4(32'hbbbd609d),
	.w5(32'hbc031229),
	.w6(32'h3b0400c5),
	.w7(32'hbbded41c),
	.w8(32'hbc00f675),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc026f3),
	.w1(32'hbbfa430e),
	.w2(32'hbbcaea1b),
	.w3(32'hbb9e4f2d),
	.w4(32'hbbfde08d),
	.w5(32'hbba6405b),
	.w6(32'hbb7520ef),
	.w7(32'hbbda2982),
	.w8(32'hbba3d5b3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839441),
	.w1(32'h395a4f6d),
	.w2(32'hb93da536),
	.w3(32'hbbe10023),
	.w4(32'hbb0b4712),
	.w5(32'hb7fb402d),
	.w6(32'hbbbe206e),
	.w7(32'hbb274736),
	.w8(32'hbb3403a2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f387b),
	.w1(32'h3a903bec),
	.w2(32'h3b47aa83),
	.w3(32'hba9d145a),
	.w4(32'hbb29a223),
	.w5(32'h3b43efb8),
	.w6(32'hbacac93e),
	.w7(32'hba323824),
	.w8(32'hba0a31cb),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b1d3d),
	.w1(32'hbbc40368),
	.w2(32'hbc208eee),
	.w3(32'h3a04b20a),
	.w4(32'hbbbc1abc),
	.w5(32'hbbd4b5f9),
	.w6(32'hbae3dfcb),
	.w7(32'hbbfeb797),
	.w8(32'hbc0332b5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f75e),
	.w1(32'hbb102eef),
	.w2(32'h398bb766),
	.w3(32'hbb8ce0c3),
	.w4(32'hb9587490),
	.w5(32'h3a0a5307),
	.w6(32'hbb4b305d),
	.w7(32'hbab85b7f),
	.w8(32'h381f618e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62f4df),
	.w1(32'h39e18366),
	.w2(32'h39e7b3b4),
	.w3(32'hbb7b57d4),
	.w4(32'h3a0e2a18),
	.w5(32'h3a61deb4),
	.w6(32'hbb1fc56f),
	.w7(32'h3b102038),
	.w8(32'h3a983f7e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83b5a3),
	.w1(32'hbc17574a),
	.w2(32'hbbfc082b),
	.w3(32'h3be9707f),
	.w4(32'hbc1dd54f),
	.w5(32'hbbfe5164),
	.w6(32'h3c0b3806),
	.w7(32'hbc0c51a2),
	.w8(32'hbc0e5c31),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbaaa6),
	.w1(32'h3b8f16bc),
	.w2(32'h3aa1cc87),
	.w3(32'hbbdefe04),
	.w4(32'h3a8840f6),
	.w5(32'h39c95266),
	.w6(32'hbbe302e7),
	.w7(32'h39c738f1),
	.w8(32'h39f493a3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70932a),
	.w1(32'hbb8b8d00),
	.w2(32'hba35330b),
	.w3(32'hba230c9e),
	.w4(32'h3aa2a41f),
	.w5(32'h3acd69ed),
	.w6(32'h3a233017),
	.w7(32'h3ad5be8e),
	.w8(32'h3b54f9d8),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba583c),
	.w1(32'h3b6bf22f),
	.w2(32'h3b9aee33),
	.w3(32'h3b13f7d0),
	.w4(32'h3bddacf4),
	.w5(32'h3bd9c0d7),
	.w6(32'h3bb32b20),
	.w7(32'h3bc5722b),
	.w8(32'h3bd729c4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967de5d),
	.w1(32'hbbe965d7),
	.w2(32'hbbb31a54),
	.w3(32'h394e74b9),
	.w4(32'hbbcd0c30),
	.w5(32'hbb89b527),
	.w6(32'hba1531eb),
	.w7(32'hbb7a5027),
	.w8(32'hbad1d8ce),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d767d),
	.w1(32'h3b11ac84),
	.w2(32'hbac63906),
	.w3(32'hbb44f258),
	.w4(32'h3b5326d6),
	.w5(32'hbad69658),
	.w6(32'hbaa79410),
	.w7(32'h3accd6b8),
	.w8(32'hba004478),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fb47d),
	.w1(32'hbb0043fd),
	.w2(32'hbb45a293),
	.w3(32'hbb88fb18),
	.w4(32'hbb432004),
	.w5(32'hbb3bbf3a),
	.w6(32'hbb323aba),
	.w7(32'hbbb677bc),
	.w8(32'hbbbba69a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7e3e2),
	.w1(32'h3bb36ee1),
	.w2(32'h3b674fe1),
	.w3(32'h3b822e2d),
	.w4(32'h3abc6177),
	.w5(32'h3b0307ab),
	.w6(32'h37007f29),
	.w7(32'h3ae696dd),
	.w8(32'h3a9eaa67),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac37fb4),
	.w1(32'hb9a7ebae),
	.w2(32'hbac156bb),
	.w3(32'h3b09adef),
	.w4(32'hbae56ff3),
	.w5(32'hbb9526d6),
	.w6(32'hb7bfef02),
	.w7(32'hbbb245dd),
	.w8(32'hbc18ba94),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb496fb5),
	.w1(32'h3b03ff0f),
	.w2(32'h3ad57a44),
	.w3(32'hbb6ee6f3),
	.w4(32'h3b5945ac),
	.w5(32'h39b2d4dd),
	.w6(32'hbc0014d9),
	.w7(32'h3b87efc4),
	.w8(32'h3b587176),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa2e4f),
	.w1(32'h3b0a9c3f),
	.w2(32'h3b06a92f),
	.w3(32'h3be78dad),
	.w4(32'h3b97933f),
	.w5(32'h3b8b8f94),
	.w6(32'h3c0c8bec),
	.w7(32'h3b309f42),
	.w8(32'h3a994697),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadb21c),
	.w1(32'h3c0707fa),
	.w2(32'h3b9d5ccb),
	.w3(32'h3930a9a3),
	.w4(32'h3c22e078),
	.w5(32'h3bab41a7),
	.w6(32'hb9ab2534),
	.w7(32'h3c1044e7),
	.w8(32'h3bb7977f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba31977),
	.w1(32'hba13ff63),
	.w2(32'hbaa66e38),
	.w3(32'h3bb86810),
	.w4(32'hbb275d8a),
	.w5(32'h398492a7),
	.w6(32'h3bc3758d),
	.w7(32'hba693c31),
	.w8(32'h39e3c3aa),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e86c2),
	.w1(32'h3b3cf779),
	.w2(32'h3b0589bb),
	.w3(32'hbaebf6c7),
	.w4(32'h3b0bd6d4),
	.w5(32'h3a1b1160),
	.w6(32'hb949b0bb),
	.w7(32'h3a3fdfd7),
	.w8(32'h3996623e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33b736),
	.w1(32'hbad99750),
	.w2(32'hbb847b00),
	.w3(32'h39d4b45c),
	.w4(32'hbba9c472),
	.w5(32'hbb8ed886),
	.w6(32'hbb80bca1),
	.w7(32'hbc228893),
	.w8(32'hbc08b2d6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa85e77),
	.w1(32'h3a2281ed),
	.w2(32'h3b1f3a49),
	.w3(32'hba4b83c3),
	.w4(32'h39f605ce),
	.w5(32'h3b226b3e),
	.w6(32'hbb16de96),
	.w7(32'h3acc61d2),
	.w8(32'h3b58fc24),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba911d33),
	.w1(32'h3b9779fe),
	.w2(32'h3bcf777e),
	.w3(32'hba58ce78),
	.w4(32'h3ba598a1),
	.w5(32'h3b4dd520),
	.w6(32'h3b1744d8),
	.w7(32'h3b331dee),
	.w8(32'h39c60810),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b555d40),
	.w1(32'hb988ad4f),
	.w2(32'hb8d79f0f),
	.w3(32'h3b913050),
	.w4(32'hba2ea6d6),
	.w5(32'hba163d89),
	.w6(32'h3bb2b01a),
	.w7(32'hb98aeb84),
	.w8(32'h3907ea98),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab564e4),
	.w1(32'hbb88ba8e),
	.w2(32'hbb6a5898),
	.w3(32'h3b151dea),
	.w4(32'hbb9fa607),
	.w5(32'hbb894f20),
	.w6(32'h3b8ace7f),
	.w7(32'hbb9a9567),
	.w8(32'hbba8483b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ba3b5),
	.w1(32'hbbb19eab),
	.w2(32'hbb9de558),
	.w3(32'hbb6052ae),
	.w4(32'hbb49a488),
	.w5(32'hbaac947f),
	.w6(32'hbb8c4dc5),
	.w7(32'hbb1c1447),
	.w8(32'hbae0ea7a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb457a82),
	.w1(32'hbb9339d3),
	.w2(32'hbb9fe9a3),
	.w3(32'hbbb96fec),
	.w4(32'hbbd7d0b2),
	.w5(32'hbbb90185),
	.w6(32'hbbde4b76),
	.w7(32'hbba7c55c),
	.w8(32'hbba1e5e4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803bcc),
	.w1(32'h3aa3940c),
	.w2(32'hbaae3223),
	.w3(32'hbb433555),
	.w4(32'hba77d471),
	.w5(32'hbb1beee0),
	.w6(32'h395c7c1a),
	.w7(32'hba3c6871),
	.w8(32'hbad0986d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a85d2c),
	.w1(32'hbbb73cc1),
	.w2(32'hbaa71455),
	.w3(32'hbb3e2113),
	.w4(32'hbbc3df30),
	.w5(32'hba8d945a),
	.w6(32'hbb0c9c32),
	.w7(32'hbb336484),
	.w8(32'hba6ccdba),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939c359),
	.w1(32'hbb039175),
	.w2(32'hbb82984c),
	.w3(32'h3ad8fa66),
	.w4(32'h3a8d15ea),
	.w5(32'hba878f3b),
	.w6(32'h3aa4726a),
	.w7(32'h3a89d047),
	.w8(32'h3a913a4f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f44f6),
	.w1(32'hbb9572e3),
	.w2(32'hbb9914e9),
	.w3(32'hbbc2b8fc),
	.w4(32'hbb74cda5),
	.w5(32'hbb6e6985),
	.w6(32'hbb39a3df),
	.w7(32'hbb0dae5e),
	.w8(32'hbb848a66),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8fe14),
	.w1(32'hbbaf9644),
	.w2(32'hbba46282),
	.w3(32'hbb85173a),
	.w4(32'hbb94b50c),
	.w5(32'hbba054c7),
	.w6(32'hbb89dcd8),
	.w7(32'hbba296f3),
	.w8(32'hbba93d66),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b70c4),
	.w1(32'h39dac739),
	.w2(32'h39e77ea1),
	.w3(32'hba2c12ab),
	.w4(32'h3ace8af2),
	.w5(32'h3b990e69),
	.w6(32'hbb02c4b4),
	.w7(32'h3a9fc833),
	.w8(32'h3ac83edd),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ef14c),
	.w1(32'h3a847492),
	.w2(32'h38cd86ae),
	.w3(32'h3b14d418),
	.w4(32'h3aa7c083),
	.w5(32'hba16fed9),
	.w6(32'hbab8fb66),
	.w7(32'hba577729),
	.w8(32'hbb74ec80),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b817ca4),
	.w1(32'hbb3a2d01),
	.w2(32'hbb82680f),
	.w3(32'h3afb3f44),
	.w4(32'hbae6cc94),
	.w5(32'hbb835fc2),
	.w6(32'hbb2eb84c),
	.w7(32'hbb5200d0),
	.w8(32'hbb84ac86),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd48740),
	.w1(32'h397075da),
	.w2(32'h3b217bd4),
	.w3(32'hbbf3d86d),
	.w4(32'h3afc12c3),
	.w5(32'h3b6ec733),
	.w6(32'hbbd8cdf2),
	.w7(32'hb894fd33),
	.w8(32'h3a05918a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41395d),
	.w1(32'h3b603cb7),
	.w2(32'h3b885e02),
	.w3(32'h3babcd29),
	.w4(32'h3b45d58d),
	.w5(32'h3ba4605c),
	.w6(32'h3bd457c1),
	.w7(32'h3b72d58d),
	.w8(32'h3b91169c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66faac),
	.w1(32'h3b50fb02),
	.w2(32'h3b1ba1b3),
	.w3(32'h3ab81471),
	.w4(32'h3b43b273),
	.w5(32'h3b1ecf87),
	.w6(32'h3a5bc93f),
	.w7(32'h3b5c1b5b),
	.w8(32'h3ac65c04),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23eaa8),
	.w1(32'hba2fb4a4),
	.w2(32'hbb8af349),
	.w3(32'hba7c19c1),
	.w4(32'hbab8fc90),
	.w5(32'hbb3c59b6),
	.w6(32'hba5f73b4),
	.w7(32'hba41686b),
	.w8(32'hbb571bc0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa402ee),
	.w1(32'hbaa8b966),
	.w2(32'hbb8aa4a1),
	.w3(32'hbba66358),
	.w4(32'hbb142876),
	.w5(32'hbb9f71fb),
	.w6(32'hbba85504),
	.w7(32'hba58b5bc),
	.w8(32'hbbfa09ea),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa4a0),
	.w1(32'hbac260a1),
	.w2(32'h3b948036),
	.w3(32'h3b035a14),
	.w4(32'h3b8dc946),
	.w5(32'h3bcf6d92),
	.w6(32'h3b73cc60),
	.w7(32'h3b9d8a92),
	.w8(32'h3bbf9beb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7748),
	.w1(32'h3bda2114),
	.w2(32'h3bb4c9c5),
	.w3(32'hbaad9fbe),
	.w4(32'h3bf9ed4b),
	.w5(32'h3c0cde1f),
	.w6(32'h3b132bd5),
	.w7(32'h3c03038d),
	.w8(32'h3c06c016),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5898db),
	.w1(32'hbba30db9),
	.w2(32'hbbc2eb5a),
	.w3(32'h3ba3b7b5),
	.w4(32'hbba6dca1),
	.w5(32'hbbcb31ad),
	.w6(32'h3bcd709c),
	.w7(32'hbb901bdb),
	.w8(32'hbb6c151d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63b4aa),
	.w1(32'h3aaf9b82),
	.w2(32'h3a7770d6),
	.w3(32'hbb412df7),
	.w4(32'hb7a18ce7),
	.w5(32'hba9f318d),
	.w6(32'hb9f4b0cc),
	.w7(32'hba051d83),
	.w8(32'hba944cb4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e045e),
	.w1(32'h3c25f9b4),
	.w2(32'h3bbf5b3a),
	.w3(32'hbb3fee2e),
	.w4(32'h3c1c08c4),
	.w5(32'h3b9f82b2),
	.w6(32'hbb751316),
	.w7(32'h3c212852),
	.w8(32'h3bc14252),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c128a6a),
	.w1(32'hbaa03cff),
	.w2(32'h3a4cddb2),
	.w3(32'h3c0bd365),
	.w4(32'hbb5ef311),
	.w5(32'h3b09f102),
	.w6(32'h3c18b388),
	.w7(32'hbabba50a),
	.w8(32'hbaa87e7e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2bc49),
	.w1(32'h39670d93),
	.w2(32'h3b03519b),
	.w3(32'hbb326f3c),
	.w4(32'hb9ff93ae),
	.w5(32'hbb55725d),
	.w6(32'hbb758e09),
	.w7(32'hba99f13f),
	.w8(32'hbb3a015e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b919236),
	.w1(32'h3c051129),
	.w2(32'h3c4fd0ae),
	.w3(32'h3aa8c142),
	.w4(32'h3c42405c),
	.w5(32'h3c571c9f),
	.w6(32'h3b9e65a9),
	.w7(32'h3c2e714e),
	.w8(32'h3c158ae6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829c85),
	.w1(32'hbb905672),
	.w2(32'hbb27704c),
	.w3(32'h3bff3b04),
	.w4(32'hbb4cf355),
	.w5(32'hbb40d569),
	.w6(32'h3bd2c77b),
	.w7(32'hbb31d508),
	.w8(32'hbb020c27),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d1035),
	.w1(32'h3ba2e35a),
	.w2(32'hba0de7b8),
	.w3(32'h3a53183d),
	.w4(32'hbb0a7e5c),
	.w5(32'hbc08f2e1),
	.w6(32'h3b612c89),
	.w7(32'hbb4f9962),
	.w8(32'hbc40ed0a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6f21b),
	.w1(32'hba652740),
	.w2(32'h3ad797d7),
	.w3(32'hbc1d4238),
	.w4(32'hbb292f99),
	.w5(32'hbacf902c),
	.w6(32'hbb8ce239),
	.w7(32'hbb31ea0b),
	.w8(32'h3ad1ebcd),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f8250),
	.w1(32'hbae70650),
	.w2(32'h3991833e),
	.w3(32'hbb98e607),
	.w4(32'h3a0f052b),
	.w5(32'h3b9cd0f6),
	.w6(32'hbb36a93f),
	.w7(32'hbb31579f),
	.w8(32'hbbc923f0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f1aae),
	.w1(32'h3b5bce1d),
	.w2(32'h3c6edb9f),
	.w3(32'h3aa02e92),
	.w4(32'hbaf8d29f),
	.w5(32'h3cc8da6c),
	.w6(32'hbb47a3a0),
	.w7(32'hbbfda4a3),
	.w8(32'h3c357409),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ec73e),
	.w1(32'hbb3ad289),
	.w2(32'h3b5ef402),
	.w3(32'h3c3f1d46),
	.w4(32'hbb9a8054),
	.w5(32'hbb1c36a4),
	.w6(32'h3c39b1c8),
	.w7(32'hbaaca685),
	.w8(32'hb9c6fc08),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa88f0),
	.w1(32'hbb900ebb),
	.w2(32'hbb43326c),
	.w3(32'hbb137e11),
	.w4(32'h3b5e78f9),
	.w5(32'h3bafe8bf),
	.w6(32'h3b638389),
	.w7(32'hbc1e28dc),
	.w8(32'hbb1cc5d7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34f5d3),
	.w1(32'hbac51d5a),
	.w2(32'hbae1c598),
	.w3(32'h3c2030da),
	.w4(32'h3bdcd4bc),
	.w5(32'h3c08f75d),
	.w6(32'h395f3aac),
	.w7(32'h3a2f7ae1),
	.w8(32'h39aae5ab),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7b2c0),
	.w1(32'hbb831c4f),
	.w2(32'h3b1404b1),
	.w3(32'hbab6615b),
	.w4(32'hbb03904b),
	.w5(32'hbaa86ee2),
	.w6(32'h3b943d94),
	.w7(32'hba406984),
	.w8(32'hba7ae148),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba475ca1),
	.w1(32'h3aad4161),
	.w2(32'h38477df7),
	.w3(32'hb98b7865),
	.w4(32'h3acb8e8f),
	.w5(32'h3c571c02),
	.w6(32'h386741a0),
	.w7(32'h3b148f77),
	.w8(32'hb9d11ed1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cab49),
	.w1(32'hba8f9c86),
	.w2(32'h3a9727fc),
	.w3(32'h3bb10827),
	.w4(32'h3b5ed76d),
	.w5(32'h3b855407),
	.w6(32'h3a2639da),
	.w7(32'h3b861089),
	.w8(32'h3ba00d47),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac8c7e),
	.w1(32'hbadeb918),
	.w2(32'h3b355895),
	.w3(32'hbb2624a8),
	.w4(32'hbc04ff97),
	.w5(32'h3975a673),
	.w6(32'h3b49d850),
	.w7(32'hbc184336),
	.w8(32'hbbc1b978),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0551fa),
	.w1(32'h3bb814f6),
	.w2(32'h3bc12910),
	.w3(32'hbb405a13),
	.w4(32'h3a978b17),
	.w5(32'hbbb68f51),
	.w6(32'h3a69bdc4),
	.w7(32'h3bb6cd6e),
	.w8(32'hbac1efff),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b895386),
	.w1(32'h3a9367e1),
	.w2(32'hbba12651),
	.w3(32'h3b4dc106),
	.w4(32'h3aeda125),
	.w5(32'h3aa9d1ca),
	.w6(32'h3a49c884),
	.w7(32'h39c621ff),
	.w8(32'hba8eff79),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94973d),
	.w1(32'hbabb4143),
	.w2(32'hbbb9d688),
	.w3(32'hbb768f0c),
	.w4(32'hbabc8dbc),
	.w5(32'hbbc5f4f8),
	.w6(32'hbb149d4e),
	.w7(32'hba4119d9),
	.w8(32'hbb8a16e5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa13f2),
	.w1(32'hba027e0a),
	.w2(32'h3b861399),
	.w3(32'hbae2af11),
	.w4(32'hbb1c1adb),
	.w5(32'hba4b9281),
	.w6(32'hba8948a5),
	.w7(32'h38b13f2d),
	.w8(32'h3b9dbc40),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c7b70),
	.w1(32'h3b1bbc9a),
	.w2(32'h3bca9ed6),
	.w3(32'hbc2c7c60),
	.w4(32'hbb516802),
	.w5(32'h3ca3ce2a),
	.w6(32'hbc34e135),
	.w7(32'hbc647a3f),
	.w8(32'hbb13e52a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c88c54),
	.w1(32'h3b455e6d),
	.w2(32'h3c5db7da),
	.w3(32'h3bbbe9ee),
	.w4(32'hba574737),
	.w5(32'h3bb3522c),
	.w6(32'h3bc0b9ba),
	.w7(32'hbad50a23),
	.w8(32'h3ba7781a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83fa81),
	.w1(32'hbadbece8),
	.w2(32'hbb81ada3),
	.w3(32'h38b38a01),
	.w4(32'h38f2b7a8),
	.w5(32'h3b176b36),
	.w6(32'hbbbcb95d),
	.w7(32'h3ad3dc34),
	.w8(32'hba633875),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acebf9d),
	.w1(32'h3bc697cc),
	.w2(32'h3b0474e5),
	.w3(32'h3b39a56a),
	.w4(32'h3b903a14),
	.w5(32'h3ac80ec5),
	.w6(32'hba864353),
	.w7(32'hbb1cc980),
	.w8(32'hbaad1bdd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54e99d),
	.w1(32'hbb6571c3),
	.w2(32'hbb9673da),
	.w3(32'h3ab944e7),
	.w4(32'hbb378fb3),
	.w5(32'hbb692a9b),
	.w6(32'h3b4466e3),
	.w7(32'hbbf34e0d),
	.w8(32'hbbfcf8d5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99e231),
	.w1(32'hba2c4623),
	.w2(32'h3af6aa2b),
	.w3(32'hbb8feed5),
	.w4(32'h3b81d57e),
	.w5(32'h3be88889),
	.w6(32'hbb222386),
	.w7(32'h3ba071a2),
	.w8(32'h3afc862a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf47ac),
	.w1(32'hbbe4e4dd),
	.w2(32'hbc9a87f8),
	.w3(32'hbc0ae626),
	.w4(32'hbae9b5a8),
	.w5(32'hbbf170eb),
	.w6(32'hbc029e20),
	.w7(32'hbb49c44a),
	.w8(32'hbbd4bef9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc809383),
	.w1(32'hba4c9bee),
	.w2(32'hbb686501),
	.w3(32'hbc7a4f19),
	.w4(32'hbb863098),
	.w5(32'hbba32fa0),
	.w6(32'hbc2f682c),
	.w7(32'hbb9bf075),
	.w8(32'hbaf3e3da),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39824e39),
	.w1(32'hba952421),
	.w2(32'hb9ba9bec),
	.w3(32'h3b3f80ab),
	.w4(32'h3a300adf),
	.w5(32'h3991373a),
	.w6(32'hbb205126),
	.w7(32'h3c1bc1d3),
	.w8(32'h3c0222f9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb669a0),
	.w1(32'hba3bf269),
	.w2(32'h3a3ee451),
	.w3(32'hbb59e367),
	.w4(32'h3b841ecb),
	.w5(32'hbba8c661),
	.w6(32'h3b45a09f),
	.w7(32'h3c27e130),
	.w8(32'h3bc352fb),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb975d22),
	.w1(32'hba9435d0),
	.w2(32'hbabb1d89),
	.w3(32'hbc039590),
	.w4(32'h3b53634a),
	.w5(32'h3be80735),
	.w6(32'hbb5ca614),
	.w7(32'hbbfb72c6),
	.w8(32'hbac3833a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba735a6d),
	.w1(32'hb9a0b879),
	.w2(32'h3b5e6377),
	.w3(32'h3b0dd829),
	.w4(32'hbb84ae2e),
	.w5(32'hba225c36),
	.w6(32'hbaa00362),
	.w7(32'hbb88ab19),
	.w8(32'hbb342f65),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93a6a0),
	.w1(32'hbb6f68ed),
	.w2(32'h3ac05fbb),
	.w3(32'hbbf2c3bb),
	.w4(32'hbc133688),
	.w5(32'hbb967274),
	.w6(32'hbba07b60),
	.w7(32'hbc135faa),
	.w8(32'hbc3a97e7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedb3af),
	.w1(32'hbbae0c66),
	.w2(32'h3acc3d5b),
	.w3(32'hbb068170),
	.w4(32'hbc1bea93),
	.w5(32'hbbaabb39),
	.w6(32'hbb5b08b1),
	.w7(32'h3b0a5343),
	.w8(32'hbbfb2642),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4311d),
	.w1(32'hbab268e0),
	.w2(32'h39fec55b),
	.w3(32'h3a272370),
	.w4(32'hbbee4eda),
	.w5(32'hbba9171e),
	.w6(32'hbb6d4bc1),
	.w7(32'hbbc23f3b),
	.w8(32'hbc2a916e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77d868),
	.w1(32'hbb2b7c48),
	.w2(32'hb9baa91f),
	.w3(32'h3c13aade),
	.w4(32'hbc0f64f9),
	.w5(32'hbab62e8e),
	.w6(32'h3b97e10c),
	.w7(32'hbbeb1151),
	.w8(32'hbc18e9c5),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbac7b),
	.w1(32'hbb9a1dfb),
	.w2(32'hba1b5a25),
	.w3(32'h3a683014),
	.w4(32'hbb756eef),
	.w5(32'hbb267a3a),
	.w6(32'h3bede254),
	.w7(32'hb953beec),
	.w8(32'hbab14cee),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9d6d0),
	.w1(32'hbb645ffa),
	.w2(32'hbaab097f),
	.w3(32'hbb9e7df4),
	.w4(32'hbb9722ba),
	.w5(32'h3a7f2603),
	.w6(32'h3b7a6c40),
	.w7(32'hbb7f598f),
	.w8(32'hbb54b6cf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2c2ff),
	.w1(32'h3b546ce4),
	.w2(32'hbad22410),
	.w3(32'hbc4dfcf3),
	.w4(32'hbb84bd59),
	.w5(32'hbbbd28a5),
	.w6(32'hbc1fd522),
	.w7(32'hbc40c0ca),
	.w8(32'hbc01937a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b581950),
	.w1(32'h3b0d6bfb),
	.w2(32'hbb6d0bb2),
	.w3(32'hbb64c3e6),
	.w4(32'hb9e7b6cf),
	.w5(32'h3c4f584b),
	.w6(32'hbb8b31a6),
	.w7(32'hbbad7d22),
	.w8(32'hba8717b2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26e621),
	.w1(32'hbb84770a),
	.w2(32'hbb8a5ef1),
	.w3(32'h3b42bc3e),
	.w4(32'hbb53503d),
	.w5(32'hbbcfaa05),
	.w6(32'h3b9f899d),
	.w7(32'hbb33cdb1),
	.w8(32'hbb8076d0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cd729),
	.w1(32'hbb0323da),
	.w2(32'hbb0a7d71),
	.w3(32'hbb295d9a),
	.w4(32'hbb130b60),
	.w5(32'hbb147259),
	.w6(32'hbb835471),
	.w7(32'hba808fd3),
	.w8(32'hbb203fe9),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72affd),
	.w1(32'h3a439d7c),
	.w2(32'hb96109fb),
	.w3(32'h39404eac),
	.w4(32'h3a95b695),
	.w5(32'hbb53b731),
	.w6(32'hba9d6f8c),
	.w7(32'h3b04d1f4),
	.w8(32'h3b78b0b2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233455),
	.w1(32'h3b29c1c0),
	.w2(32'h3bda80d7),
	.w3(32'hbb762d7a),
	.w4(32'hba48aaba),
	.w5(32'h3c720f7b),
	.w6(32'hbb86b969),
	.w7(32'hbbd8d440),
	.w8(32'h3b859c3a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901cf7),
	.w1(32'hbbba4e75),
	.w2(32'h3b31cf45),
	.w3(32'hba7bcf76),
	.w4(32'hbc34422e),
	.w5(32'hb994ed59),
	.w6(32'h3b8cc17a),
	.w7(32'hbb064321),
	.w8(32'hbb8e0ef1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6b3b5),
	.w1(32'hbb25338a),
	.w2(32'h3b789621),
	.w3(32'hba4adece),
	.w4(32'hba6f7b90),
	.w5(32'h3bfd36ab),
	.w6(32'hbafe4b7f),
	.w7(32'hbb8fdd45),
	.w8(32'h3a309a83),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01999c),
	.w1(32'h3be6a301),
	.w2(32'h3baf4337),
	.w3(32'h3a659b78),
	.w4(32'h3b1eb23e),
	.w5(32'h3b3e3e36),
	.w6(32'h3a18ce84),
	.w7(32'hb86205e5),
	.w8(32'hb9a3abc1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42db31),
	.w1(32'hbafba2e0),
	.w2(32'h3bb44ba0),
	.w3(32'h3bb29e71),
	.w4(32'hbae406f3),
	.w5(32'h3bd01abb),
	.w6(32'h39fabe50),
	.w7(32'hbae1bd6d),
	.w8(32'hbb49f800),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a0974e),
	.w1(32'hb75eab51),
	.w2(32'h3b747463),
	.w3(32'hbb5d104b),
	.w4(32'hbc09b9e8),
	.w5(32'hbb3b68f9),
	.w6(32'hbbc6e0d1),
	.w7(32'hbba72729),
	.w8(32'hbb620e28),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5678f2),
	.w1(32'hbb882496),
	.w2(32'h3bf257cf),
	.w3(32'hba8f67d8),
	.w4(32'hbbdfb7fc),
	.w5(32'hbc0aef73),
	.w6(32'hbb0a2bfe),
	.w7(32'hbb5168c7),
	.w8(32'hbc0b7933),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b444ac7),
	.w1(32'h3b0caa48),
	.w2(32'h3aafdcd3),
	.w3(32'h3a3b7420),
	.w4(32'h3a96e575),
	.w5(32'hbbb92d5a),
	.w6(32'h3ae4c0b3),
	.w7(32'h3b8e04d1),
	.w8(32'hbb10dd93),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37e7b3),
	.w1(32'h3b3b1a22),
	.w2(32'h3bf21dd7),
	.w3(32'hbb5bccf4),
	.w4(32'h3aa0d4d4),
	.w5(32'h3bdb6b5e),
	.w6(32'hb6522ee8),
	.w7(32'hbb29e475),
	.w8(32'h3b220b4e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c120dd9),
	.w1(32'hbb16b98a),
	.w2(32'h3ae88473),
	.w3(32'h3c15774a),
	.w4(32'hba04db4c),
	.w5(32'h3b7125d4),
	.w6(32'h3bb7635a),
	.w7(32'hbb9009e2),
	.w8(32'h3b8a2488),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5dcd2),
	.w1(32'hbba3d202),
	.w2(32'hba0339d8),
	.w3(32'h3b4f07a9),
	.w4(32'h3ace5e44),
	.w5(32'hb8f33022),
	.w6(32'h3bd3c1d5),
	.w7(32'h3c2d60f4),
	.w8(32'h3ae2667e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad9900),
	.w1(32'hbc05512c),
	.w2(32'hbbe861eb),
	.w3(32'hbba8dc01),
	.w4(32'hbbc55321),
	.w5(32'hbb196f18),
	.w6(32'hbb5b925b),
	.w7(32'hbb882445),
	.w8(32'hbbc22e1d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb578387),
	.w1(32'h3abb6da0),
	.w2(32'h3be9908d),
	.w3(32'hba7dc969),
	.w4(32'hbb2d2929),
	.w5(32'h3bca31e3),
	.w6(32'h39aa8a1f),
	.w7(32'hbb858ff9),
	.w8(32'hba01ac5e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7666d7),
	.w1(32'hba9a7943),
	.w2(32'hba72b432),
	.w3(32'h3b0b0ce9),
	.w4(32'h3b470125),
	.w5(32'hbb5dd0d4),
	.w6(32'hbab92f28),
	.w7(32'h3a9e5c4c),
	.w8(32'hb9e4266f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2ffab),
	.w1(32'h3b0e70ce),
	.w2(32'h3b24ffb4),
	.w3(32'h3b994753),
	.w4(32'hba1780cc),
	.w5(32'hbb9e61e7),
	.w6(32'hba383282),
	.w7(32'hbba9156b),
	.w8(32'hbb08b21e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdfbb5),
	.w1(32'hb9c99684),
	.w2(32'hb9328476),
	.w3(32'hbab6e888),
	.w4(32'hbb8d8876),
	.w5(32'hbc39549e),
	.w6(32'hbace5e4a),
	.w7(32'hbab19660),
	.w8(32'hbbcf0749),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7585f1),
	.w1(32'hba66a1eb),
	.w2(32'hbb89ad32),
	.w3(32'hbafe159e),
	.w4(32'h39918a65),
	.w5(32'hbbf2e15d),
	.w6(32'hbb92dd7c),
	.w7(32'h3bedb71c),
	.w8(32'hbb4a9b09),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7612a0),
	.w1(32'hbb989e6e),
	.w2(32'h3bd4e780),
	.w3(32'hbbf43987),
	.w4(32'hbb7db820),
	.w5(32'h3c08c027),
	.w6(32'hbaa842c3),
	.w7(32'hbafa1e46),
	.w8(32'hbb462a43),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff61c4),
	.w1(32'hbb8086ee),
	.w2(32'hbb7c7125),
	.w3(32'h379c5a9f),
	.w4(32'hbc011f1c),
	.w5(32'hbc11b610),
	.w6(32'hba3f5cc3),
	.w7(32'hbc89255e),
	.w8(32'hbc2c2e83),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58079d),
	.w1(32'hbb63f966),
	.w2(32'hba6699f1),
	.w3(32'hbb2da545),
	.w4(32'h39c9cab8),
	.w5(32'hbb0e86ac),
	.w6(32'hba832af6),
	.w7(32'hbabc7405),
	.w8(32'hbb470550),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4b946),
	.w1(32'h3a7e0dfe),
	.w2(32'h3bca2665),
	.w3(32'hbb8bdfc2),
	.w4(32'hbb6f83d5),
	.w5(32'h3abe4eed),
	.w6(32'hbbd666a4),
	.w7(32'hbb776984),
	.w8(32'hb7aca66f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule