module layer_8_featuremap_153(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34229f),
	.w1(32'h3b6a0ec1),
	.w2(32'h3bb6048a),
	.w3(32'hba728644),
	.w4(32'h3bacd637),
	.w5(32'h3b8c2884),
	.w6(32'h39910ad1),
	.w7(32'h3ac4f452),
	.w8(32'hbb3f76b9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dd4c7),
	.w1(32'hbbcf9731),
	.w2(32'h3c4486ed),
	.w3(32'hbb0c7133),
	.w4(32'h3c4e6332),
	.w5(32'h3bdb703c),
	.w6(32'hbb841d7f),
	.w7(32'h3c3826a9),
	.w8(32'h3b5392f7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdb764),
	.w1(32'h3b82b2a4),
	.w2(32'h3bb8786c),
	.w3(32'h3aa8f23b),
	.w4(32'hba78fd3d),
	.w5(32'hbba65c01),
	.w6(32'h3a897d66),
	.w7(32'h3b0a8931),
	.w8(32'hbbb1bdda),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dfd0c),
	.w1(32'h3a6aa134),
	.w2(32'hbc0538a0),
	.w3(32'hbc0a3550),
	.w4(32'h39971a60),
	.w5(32'hbc157e1e),
	.w6(32'hbbb421eb),
	.w7(32'hbb6a2640),
	.w8(32'hbbf18bc2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f0199),
	.w1(32'hbc0240df),
	.w2(32'h3b456a09),
	.w3(32'hbc127b60),
	.w4(32'h3b09a381),
	.w5(32'hb9d126fa),
	.w6(32'hbc2efcfc),
	.w7(32'h3b074693),
	.w8(32'hbaed32bd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1b937),
	.w1(32'h3a82c5f2),
	.w2(32'hbc009878),
	.w3(32'hba26f1b2),
	.w4(32'hb9a5b074),
	.w5(32'hbc1a6b27),
	.w6(32'h3b4fd23b),
	.w7(32'h3989e53d),
	.w8(32'hbc1a4c37),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeefa55),
	.w1(32'hba480355),
	.w2(32'hbc75b304),
	.w3(32'hbb80cc44),
	.w4(32'hb8f40791),
	.w5(32'hbbe19e7c),
	.w6(32'hbbe94114),
	.w7(32'hbbc10cb2),
	.w8(32'hbc2312f1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33074c),
	.w1(32'hbb04343d),
	.w2(32'h3c1f1cf3),
	.w3(32'hbc175fa1),
	.w4(32'h3c98a784),
	.w5(32'h3ba1b974),
	.w6(32'hbc0b0040),
	.w7(32'h3c26d2c8),
	.w8(32'h3b2b7eca),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772e6c8),
	.w1(32'h3914162d),
	.w2(32'h3a9a232b),
	.w3(32'h3ad7e575),
	.w4(32'h3b8418a3),
	.w5(32'h3b3e2aa7),
	.w6(32'hbb119b1e),
	.w7(32'h3b2560fd),
	.w8(32'h3ad325d8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad6834),
	.w1(32'hbb5ee248),
	.w2(32'h3b375b38),
	.w3(32'hbb91ea72),
	.w4(32'h3c6155df),
	.w5(32'h39dd88e2),
	.w6(32'hbb73c60b),
	.w7(32'h3c64c7ae),
	.w8(32'hbc2669bf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d40f8),
	.w1(32'hbbda94c2),
	.w2(32'hb9d3af50),
	.w3(32'hbc2554e8),
	.w4(32'hbaa1cd0f),
	.w5(32'hbb47cc42),
	.w6(32'hbc969d57),
	.w7(32'h3b787d03),
	.w8(32'hba19bf07),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6c8c7),
	.w1(32'hbab664c7),
	.w2(32'h3c09f7e7),
	.w3(32'hbc121164),
	.w4(32'h3c3a0ef4),
	.w5(32'hbbeb3440),
	.w6(32'hbaf86faa),
	.w7(32'h3c091720),
	.w8(32'hbbbfbf5e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6be9ec),
	.w1(32'hbb70f772),
	.w2(32'hbc09e52b),
	.w3(32'h3b4cb8a8),
	.w4(32'hbb8f4934),
	.w5(32'hbbc81986),
	.w6(32'hbb2adef6),
	.w7(32'hba2910f3),
	.w8(32'h3bc8440e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb774ea3),
	.w1(32'h3a46dba9),
	.w2(32'hbc462839),
	.w3(32'hbb185f49),
	.w4(32'hbab69bc6),
	.w5(32'hba2cb2b7),
	.w6(32'hbad688fc),
	.w7(32'hbb96379d),
	.w8(32'hbbd21d8b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852448),
	.w1(32'hb908bc0a),
	.w2(32'hbb9ce735),
	.w3(32'h3a659fde),
	.w4(32'hbb815686),
	.w5(32'hbbbe1d06),
	.w6(32'h3b978a66),
	.w7(32'hbba90ee3),
	.w8(32'hbc12d704),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf83ca),
	.w1(32'hb9062615),
	.w2(32'hbb178096),
	.w3(32'hbb994076),
	.w4(32'h3b29b2fe),
	.w5(32'h3b24f072),
	.w6(32'hbb2865b4),
	.w7(32'hbc762698),
	.w8(32'hbc81e6a4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b35c8),
	.w1(32'hbc56bb55),
	.w2(32'h3b4cc789),
	.w3(32'h392eb15f),
	.w4(32'h3c1887d3),
	.w5(32'hbcb31deb),
	.w6(32'hbc080d4f),
	.w7(32'h3c02bff9),
	.w8(32'h3c0a0063),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e987),
	.w1(32'hbc7d4b0a),
	.w2(32'hbc229556),
	.w3(32'hbbc2f29f),
	.w4(32'hbbfdc783),
	.w5(32'h3b7b4005),
	.w6(32'hbbee78e9),
	.w7(32'hbcba330f),
	.w8(32'hbbf7d3c7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41a935),
	.w1(32'h3bd544e8),
	.w2(32'hbcc068a9),
	.w3(32'hb886e15e),
	.w4(32'h3cad4ecc),
	.w5(32'hbc3f1b16),
	.w6(32'hbc978dca),
	.w7(32'hbb99f57c),
	.w8(32'h3d1912dd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad2414),
	.w1(32'h3c0cc9e2),
	.w2(32'hba89ea40),
	.w3(32'h3c1efb00),
	.w4(32'hbb8ecfba),
	.w5(32'hbca12870),
	.w6(32'hbc6b9d3f),
	.w7(32'hbba32a31),
	.w8(32'h3d318e4f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4b784),
	.w1(32'h3c08999d),
	.w2(32'hbc0bbabb),
	.w3(32'h3a72b44e),
	.w4(32'h3b34c8c9),
	.w5(32'h3cb8616f),
	.w6(32'hbc66cd75),
	.w7(32'hbc82f149),
	.w8(32'h3c2e1aa1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1aed31),
	.w1(32'hba74f447),
	.w2(32'hbceff666),
	.w3(32'hbc49c882),
	.w4(32'hbc56864f),
	.w5(32'h3c2759b3),
	.w6(32'h3ce36e41),
	.w7(32'h3ccb3495),
	.w8(32'hbc9c97ac),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7d4fa7),
	.w1(32'h3ac9efa2),
	.w2(32'h3cd1addf),
	.w3(32'hbc350805),
	.w4(32'hba84347e),
	.w5(32'h3c376de4),
	.w6(32'h3c1d969d),
	.w7(32'hb98921a2),
	.w8(32'hbc437c78),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8a843),
	.w1(32'hbc6149ae),
	.w2(32'h3c92e902),
	.w3(32'h3ab35fd9),
	.w4(32'hba93e958),
	.w5(32'h3bbde8b4),
	.w6(32'hbba0d224),
	.w7(32'h3c46b9af),
	.w8(32'hbbc67d4e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85894c),
	.w1(32'hbb9af11e),
	.w2(32'h3bbdab9f),
	.w3(32'hbc069f6c),
	.w4(32'h3b94ec08),
	.w5(32'h3beba4e3),
	.w6(32'h3903e66a),
	.w7(32'hbabaada7),
	.w8(32'h3b5a3c39),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fd0ce),
	.w1(32'hbb6fd466),
	.w2(32'h3c6443e7),
	.w3(32'h3b05d561),
	.w4(32'h3c3391fd),
	.w5(32'hbbd221fe),
	.w6(32'h3a87c054),
	.w7(32'hbbba35cf),
	.w8(32'hba70d9b0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a2beb),
	.w1(32'hbcb90419),
	.w2(32'hbcbd62b8),
	.w3(32'h3c7ac385),
	.w4(32'h3ba76793),
	.w5(32'hbc2f73ee),
	.w6(32'hbb9c0791),
	.w7(32'h3cb73926),
	.w8(32'hbb5a53fe),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff8ea3),
	.w1(32'h3caca1d3),
	.w2(32'h3c3cab0c),
	.w3(32'h3cde56d9),
	.w4(32'h3cd94e0e),
	.w5(32'hbbec1fd6),
	.w6(32'h3b22d28b),
	.w7(32'h3d04a5f7),
	.w8(32'h3ad18064),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf30c66),
	.w1(32'hbc89f5f0),
	.w2(32'h3c39f446),
	.w3(32'hbc46575c),
	.w4(32'hbbf43a56),
	.w5(32'hbc4ea64b),
	.w6(32'hbcc8ccce),
	.w7(32'h3c216d0e),
	.w8(32'h3c9a5263),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1931cb),
	.w1(32'h3c519b7b),
	.w2(32'h3cd0b757),
	.w3(32'h3cde3f59),
	.w4(32'hbac6f3cc),
	.w5(32'h3c6bf770),
	.w6(32'hbcf1db00),
	.w7(32'hbc8eeee5),
	.w8(32'hbc0b96ae),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc016137),
	.w1(32'hbb9aba45),
	.w2(32'h3ba0d87e),
	.w3(32'hbc0e631c),
	.w4(32'h3bfdda99),
	.w5(32'h3b019f39),
	.w6(32'h3c9f770c),
	.w7(32'h3c044e50),
	.w8(32'h3b894c1c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a1a5b),
	.w1(32'h3be3a97d),
	.w2(32'h3c4a0a98),
	.w3(32'h3bb78270),
	.w4(32'hbbe2833a),
	.w5(32'hba095e92),
	.w6(32'h3bb4cb75),
	.w7(32'hbc1b8b7a),
	.w8(32'hbc6bd830),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a625d),
	.w1(32'hb82c2322),
	.w2(32'hbc8c14fd),
	.w3(32'h3b29a1ea),
	.w4(32'h3bf393bc),
	.w5(32'h3ca9922b),
	.w6(32'hbc7ee277),
	.w7(32'hbc83e573),
	.w8(32'h3d0584e3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc630739),
	.w1(32'h3c44ff18),
	.w2(32'h3b2a1e7f),
	.w3(32'hbc556cb1),
	.w4(32'h3b190fc8),
	.w5(32'h3c863766),
	.w6(32'h3d1c8473),
	.w7(32'hbc1e7010),
	.w8(32'h3c44ca4a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce199a0),
	.w1(32'hbb3453be),
	.w2(32'h3bb72918),
	.w3(32'hbbd750db),
	.w4(32'hbb06330f),
	.w5(32'h3b577494),
	.w6(32'h3cb3012c),
	.w7(32'hba623d88),
	.w8(32'h3ba41aff),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba991710),
	.w1(32'hb90fe5c5),
	.w2(32'h3c819eb7),
	.w3(32'h3aeccc8e),
	.w4(32'hbbe2c410),
	.w5(32'hbc34b38e),
	.w6(32'h3b85224f),
	.w7(32'h3c3533a8),
	.w8(32'hbc70dbb3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac1b96),
	.w1(32'h3c2cecc9),
	.w2(32'h3c13e3e2),
	.w3(32'hbb56056e),
	.w4(32'hbcacf4a7),
	.w5(32'h3a9d1611),
	.w6(32'hbc976310),
	.w7(32'h3b2e0b46),
	.w8(32'hbb809d0c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd940c7),
	.w1(32'h3bc94987),
	.w2(32'hbc1bea6f),
	.w3(32'hbbc249ac),
	.w4(32'hbb05f02d),
	.w5(32'hbbf5640b),
	.w6(32'hbcc8a5c3),
	.w7(32'h3af0579f),
	.w8(32'hbc0a3f12),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88824d),
	.w1(32'hbb4ee025),
	.w2(32'h3c9fd1ba),
	.w3(32'h3c3237e1),
	.w4(32'h3b87c1a3),
	.w5(32'hbd0ad2c6),
	.w6(32'h3c42ce13),
	.w7(32'h39ad59d7),
	.w8(32'h3d4a5a67),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeb0ea),
	.w1(32'h3c94c7c9),
	.w2(32'hbb9cc433),
	.w3(32'hbc8aba78),
	.w4(32'hbbe7a63c),
	.w5(32'h398fa414),
	.w6(32'hbd3b7aa2),
	.w7(32'hbc5ebdb0),
	.w8(32'hbb73ec4e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc525bc5),
	.w1(32'hbb2d29da),
	.w2(32'hbb44e94b),
	.w3(32'h3b142998),
	.w4(32'h3979d174),
	.w5(32'hbb28e568),
	.w6(32'h3ab08eeb),
	.w7(32'h3bbdd7ab),
	.w8(32'h3a76634f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf12364),
	.w1(32'hbc186da3),
	.w2(32'h3cb95368),
	.w3(32'h3b8723c1),
	.w4(32'hbb62dc73),
	.w5(32'h3c147bbb),
	.w6(32'hbc371e13),
	.w7(32'hbc12315c),
	.w8(32'hbd227899),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe34b7),
	.w1(32'h3c3ab1d9),
	.w2(32'h3bd7c4be),
	.w3(32'h3c5102bd),
	.w4(32'h3b2e9fa9),
	.w5(32'h3ba2e80d),
	.w6(32'h3c0f97be),
	.w7(32'hbc681634),
	.w8(32'h3ce43a8a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b3ab2),
	.w1(32'h3bebb7ec),
	.w2(32'hbc0cf18a),
	.w3(32'hbc159997),
	.w4(32'h3a0e0f42),
	.w5(32'hbbf6f684),
	.w6(32'h3c9efeb4),
	.w7(32'h3b19a250),
	.w8(32'h3b8745ab),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aeb43),
	.w1(32'h3a9f2550),
	.w2(32'h3c21ed6e),
	.w3(32'hbb20626f),
	.w4(32'hbacb027f),
	.w5(32'hbd057464),
	.w6(32'hbbc33e33),
	.w7(32'h3ca341e4),
	.w8(32'hbc8f7f68),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac01b80),
	.w1(32'hbcd269ef),
	.w2(32'h3ca23295),
	.w3(32'h3ab48e52),
	.w4(32'hbc328b43),
	.w5(32'hbb972397),
	.w6(32'hbc2aaa46),
	.w7(32'h3bfdab18),
	.w8(32'hbcc757f8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bb152),
	.w1(32'hbb369153),
	.w2(32'hbc903d38),
	.w3(32'h3b3e67a3),
	.w4(32'hbca542bf),
	.w5(32'hbcabd001),
	.w6(32'hbc2ae571),
	.w7(32'hbb84c28e),
	.w8(32'h3cc444aa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee74a0),
	.w1(32'h3c23cca5),
	.w2(32'hba453a33),
	.w3(32'hb9b5d338),
	.w4(32'hbb466d6c),
	.w5(32'hbbeb94f5),
	.w6(32'hbb987136),
	.w7(32'hbbb0ba98),
	.w8(32'hbbbca526),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d119ca7),
	.w1(32'hbc5bb991),
	.w2(32'hbb48a130),
	.w3(32'hbc10fbdd),
	.w4(32'hba20887c),
	.w5(32'hbc3c8dcf),
	.w6(32'h3c091c4e),
	.w7(32'h3c17cd57),
	.w8(32'hbc4de64a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48a01b),
	.w1(32'h3bd89cfe),
	.w2(32'hbc893b9d),
	.w3(32'hbc732f51),
	.w4(32'hbcf54d67),
	.w5(32'hbd425477),
	.w6(32'hbca391c8),
	.w7(32'h3c569b9a),
	.w8(32'hbbd7b6a3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95c916),
	.w1(32'hbc985215),
	.w2(32'h3d2ada05),
	.w3(32'hbd5b5d25),
	.w4(32'hbc20868c),
	.w5(32'hb9e9a1bb),
	.w6(32'hbd830414),
	.w7(32'hbcb0b1b1),
	.w8(32'hbd353015),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83149f),
	.w1(32'hbc59344d),
	.w2(32'hbcb0fd31),
	.w3(32'hbb260bb1),
	.w4(32'h3b54b515),
	.w5(32'h3c4e2e65),
	.w6(32'h3c083094),
	.w7(32'hbc154445),
	.w8(32'hbbb48b16),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1598b7),
	.w1(32'hbb596485),
	.w2(32'hbbbe2f16),
	.w3(32'h3b9a6c27),
	.w4(32'h3c8e1430),
	.w5(32'h3be4a712),
	.w6(32'h3d27ce91),
	.w7(32'hba1a93bc),
	.w8(32'hbb247253),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c472372),
	.w1(32'h3c2c87af),
	.w2(32'hbc1fdedb),
	.w3(32'hbbd37a01),
	.w4(32'hb9a33a21),
	.w5(32'hbbda2ee5),
	.w6(32'hbbd916ce),
	.w7(32'h3967d733),
	.w8(32'hba3285d4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebc434),
	.w1(32'hba0a9afa),
	.w2(32'hbb9dd589),
	.w3(32'hbb1f6b57),
	.w4(32'hbc17d16f),
	.w5(32'hbc8ce34f),
	.w6(32'hbba6e518),
	.w7(32'h3b47c8b2),
	.w8(32'h3d0ca5de),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b88c7),
	.w1(32'h3c2274db),
	.w2(32'hbced2fa1),
	.w3(32'hbbdd5c98),
	.w4(32'h3bb06a79),
	.w5(32'hbc97c0f6),
	.w6(32'hbcd0cd9b),
	.w7(32'h3c3f48f4),
	.w8(32'h3b4edd92),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb466cb),
	.w1(32'hba93c3bc),
	.w2(32'h3b4ad988),
	.w3(32'h3897cee3),
	.w4(32'hbc0ccf6f),
	.w5(32'hbb6d7362),
	.w6(32'hbc65655d),
	.w7(32'hbc470fca),
	.w8(32'hbb44b661),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba251511),
	.w1(32'h3ae9a8b6),
	.w2(32'h3d0ce605),
	.w3(32'h3a96f2bc),
	.w4(32'hbc9e5545),
	.w5(32'hbbebee78),
	.w6(32'h3bc18cc2),
	.w7(32'hbb588126),
	.w8(32'hbcae19b6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2924d7),
	.w1(32'hbcdc8a44),
	.w2(32'hbc0ca6d0),
	.w3(32'h3c1dfa76),
	.w4(32'h39fb1cd6),
	.w5(32'hbc00b20d),
	.w6(32'hba9226a5),
	.w7(32'h3b386be7),
	.w8(32'h3aa28f19),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dae2c),
	.w1(32'hba64a6fb),
	.w2(32'h398d2d78),
	.w3(32'hbb82d43b),
	.w4(32'hbb1d264c),
	.w5(32'hbc082019),
	.w6(32'hbb9bda9d),
	.w7(32'hb9902eee),
	.w8(32'hba6dd1ab),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ffc11),
	.w1(32'h3bf71136),
	.w2(32'h3d154023),
	.w3(32'hbb5c15c7),
	.w4(32'hbb8eeaa8),
	.w5(32'h3b63c270),
	.w6(32'hbc835940),
	.w7(32'h3c5aaaf9),
	.w8(32'hbd4646c1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78aa34),
	.w1(32'hbcccf416),
	.w2(32'h3c3f69cf),
	.w3(32'h3c304c6d),
	.w4(32'h3b178268),
	.w5(32'h3b4f6c2e),
	.w6(32'h3c7595c0),
	.w7(32'h3ba2d40c),
	.w8(32'h3bad9f6b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c756),
	.w1(32'h38682e57),
	.w2(32'hbd182ff5),
	.w3(32'hbc16b72d),
	.w4(32'h3c278b47),
	.w5(32'hbb5107c1),
	.w6(32'hb92c5a41),
	.w7(32'h3c2e9599),
	.w8(32'hbca50061),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d363635),
	.w1(32'hba4b7727),
	.w2(32'h3bf1b9c8),
	.w3(32'h3b6bef51),
	.w4(32'hbbfb3b3d),
	.w5(32'hba04f63f),
	.w6(32'hbb142fee),
	.w7(32'hbb467b6e),
	.w8(32'h3c5c6685),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc677bc1),
	.w1(32'hba8f1309),
	.w2(32'hb8bb1d8b),
	.w3(32'h38fa57e8),
	.w4(32'hbbdefb3a),
	.w5(32'h3c87eaf5),
	.w6(32'hbc929c34),
	.w7(32'hbb9b99f9),
	.w8(32'h3ad775c7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb3242),
	.w1(32'hbc325485),
	.w2(32'h3c9a0e73),
	.w3(32'h3c03358f),
	.w4(32'h3bdc6675),
	.w5(32'h3c880fdd),
	.w6(32'hbba4693c),
	.w7(32'hbc262662),
	.w8(32'h39b7adf5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8847),
	.w1(32'hbc7238ff),
	.w2(32'h3ca5eb4b),
	.w3(32'hbbc496dc),
	.w4(32'hbb9b1cb0),
	.w5(32'hbbd7fb99),
	.w6(32'h3c9506ca),
	.w7(32'hbcab3a8b),
	.w8(32'h3d58e1e9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2345e),
	.w1(32'h3be3ebf2),
	.w2(32'hbc4eb3a5),
	.w3(32'hbc82c4e1),
	.w4(32'h3c6c84c6),
	.w5(32'h3cc9bb71),
	.w6(32'hbcf7d85f),
	.w7(32'hbd1780d1),
	.w8(32'h3b056886),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd659428),
	.w1(32'h3b929c3c),
	.w2(32'hbbf6a97d),
	.w3(32'hba9c0ac1),
	.w4(32'hbbe5b3ae),
	.w5(32'h3b795663),
	.w6(32'h3cfa08de),
	.w7(32'h3cf1ebe3),
	.w8(32'hbbc1a98d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceb0c44),
	.w1(32'h3c99aed8),
	.w2(32'h3a186806),
	.w3(32'h3c8030f7),
	.w4(32'h3c12f80e),
	.w5(32'h3d18b387),
	.w6(32'hbc9e203a),
	.w7(32'hbcbe8f2f),
	.w8(32'h3c9d717f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc904362),
	.w1(32'hbbf0f196),
	.w2(32'h3d1fc86a),
	.w3(32'hbb653842),
	.w4(32'hbb367df5),
	.w5(32'h3c598512),
	.w6(32'h3ce4cbfb),
	.w7(32'hbc39ffef),
	.w8(32'hbc2e614e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6023e7),
	.w1(32'hb99ef2ab),
	.w2(32'h3c96e0cc),
	.w3(32'h3b3f2f36),
	.w4(32'hbc09c2cd),
	.w5(32'hb78861b9),
	.w6(32'h3cc54da6),
	.w7(32'hbc32eecc),
	.w8(32'hbca53159),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bfd8c),
	.w1(32'h3b064784),
	.w2(32'h3c6b39ed),
	.w3(32'h3b587c51),
	.w4(32'hbbfe478c),
	.w5(32'h3b9695a7),
	.w6(32'h3c2780ae),
	.w7(32'h3b5a9e9d),
	.w8(32'hbc36cdf2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc71159),
	.w1(32'hbc091242),
	.w2(32'h3c0c9335),
	.w3(32'hbb9c7565),
	.w4(32'h39476798),
	.w5(32'h3b9c0ab0),
	.w6(32'hbc77998c),
	.w7(32'h3c8f1257),
	.w8(32'h3ceeb890),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c7270),
	.w1(32'h3c39b89c),
	.w2(32'hbcc3b753),
	.w3(32'hbd12fc0d),
	.w4(32'hbafca0d1),
	.w5(32'hbc7653c1),
	.w6(32'h3cf1f437),
	.w7(32'h3d3bd3fc),
	.w8(32'hbd151950),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7a6481),
	.w1(32'h3c269e28),
	.w2(32'hbb43bc58),
	.w3(32'h3b21598d),
	.w4(32'h3c543cf2),
	.w5(32'h3b7d4681),
	.w6(32'hbc896ea4),
	.w7(32'h3b2ff935),
	.w8(32'h3a50d14c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4ca9b),
	.w1(32'h3bd72546),
	.w2(32'hb7c28e43),
	.w3(32'h3a3f9530),
	.w4(32'hbb095245),
	.w5(32'hbad342da),
	.w6(32'h3bfc147d),
	.w7(32'hba812751),
	.w8(32'hbaf21988),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97225b5),
	.w1(32'h3b22e5a1),
	.w2(32'h3ab169be),
	.w3(32'h3b0d26cd),
	.w4(32'h3c082ea1),
	.w5(32'h3b17c7cf),
	.w6(32'hbad2f35e),
	.w7(32'h3b77dca5),
	.w8(32'hb9dd7b90),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43c63a),
	.w1(32'hb9c66e06),
	.w2(32'hbb6f550d),
	.w3(32'h394771e4),
	.w4(32'hb8b93e8d),
	.w5(32'hbb51fed4),
	.w6(32'hbb882bf3),
	.w7(32'hbb5caaab),
	.w8(32'hbb8e39af),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ebfe1),
	.w1(32'hba2a9dce),
	.w2(32'h3b2926f0),
	.w3(32'hba3f16ad),
	.w4(32'h3b23ccb2),
	.w5(32'h3aea6da5),
	.w6(32'hba7af7c5),
	.w7(32'h39afd7ca),
	.w8(32'hba9b8f47),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba296e18),
	.w1(32'h3b3f63dd),
	.w2(32'hbb34839e),
	.w3(32'hba62f1a7),
	.w4(32'hbb67f39e),
	.w5(32'hbb8bb8e9),
	.w6(32'h3b6a9cf7),
	.w7(32'hbaab99c7),
	.w8(32'hbb094f76),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4174),
	.w1(32'h3b0a71f7),
	.w2(32'h3ad58813),
	.w3(32'hbafc6d8f),
	.w4(32'hbb3e72c1),
	.w5(32'h39fdf523),
	.w6(32'h3af4b1f6),
	.w7(32'hbb12b869),
	.w8(32'h3c28c5e7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83431),
	.w1(32'hbbcbb80a),
	.w2(32'h3a4af232),
	.w3(32'h3b84af36),
	.w4(32'h3c236df0),
	.w5(32'h3bfdc22e),
	.w6(32'hbad8b105),
	.w7(32'h3ba52277),
	.w8(32'h3af031a4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3871d2),
	.w1(32'hbba0aca7),
	.w2(32'hbc7209ad),
	.w3(32'hbbb12b3d),
	.w4(32'h3b18026a),
	.w5(32'h3b30fcf4),
	.w6(32'hb92865da),
	.w7(32'h3aee4511),
	.w8(32'hbbd070dd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae504d),
	.w1(32'h3b7cef09),
	.w2(32'h3c4d603d),
	.w3(32'h3beab694),
	.w4(32'h3c8d8654),
	.w5(32'h3c6f1dc7),
	.w6(32'hbbe69c85),
	.w7(32'h3c402043),
	.w8(32'h3c0fc54b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08b5be),
	.w1(32'h3c8ea067),
	.w2(32'hbac65840),
	.w3(32'h3c79657b),
	.w4(32'h3b8de382),
	.w5(32'h3b38cc06),
	.w6(32'h3c7aeb59),
	.w7(32'h3a99f2ef),
	.w8(32'hbbad5ff3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd9200),
	.w1(32'hbb042f7f),
	.w2(32'hbbd93657),
	.w3(32'hbb6ede29),
	.w4(32'h39830a31),
	.w5(32'h3aa1502c),
	.w6(32'hbb41207e),
	.w7(32'hba5b997c),
	.w8(32'hbb886ec6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa8982),
	.w1(32'hbb75e649),
	.w2(32'hbb226ce2),
	.w3(32'hbb21ff9c),
	.w4(32'hbb5820be),
	.w5(32'hbb911f61),
	.w6(32'hbbf6616b),
	.w7(32'hbba55327),
	.w8(32'hbb882ba1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81a368),
	.w1(32'hbae8e330),
	.w2(32'h3c81ab2f),
	.w3(32'hba5a8f4c),
	.w4(32'h3c834b65),
	.w5(32'h3c94a73e),
	.w6(32'hba619ce1),
	.w7(32'h3c8bea86),
	.w8(32'h3cbe3a4a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92edc7),
	.w1(32'h3b9214f7),
	.w2(32'h3b74cf98),
	.w3(32'h3bee8c4a),
	.w4(32'h3c7fda38),
	.w5(32'h3c1724c3),
	.w6(32'h3c16cb51),
	.w7(32'h3c136b86),
	.w8(32'h3b082cf3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d48fd),
	.w1(32'h3c606528),
	.w2(32'hbb6102e4),
	.w3(32'h3b4690bb),
	.w4(32'h3a8f14ce),
	.w5(32'hbb29833e),
	.w6(32'h3ba822d2),
	.w7(32'hbad8f6df),
	.w8(32'hbafb484f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24d968),
	.w1(32'hbb214672),
	.w2(32'h3b15a037),
	.w3(32'hb9c6f717),
	.w4(32'hbb835f69),
	.w5(32'hbb0bdeee),
	.w6(32'hba5bd7b0),
	.w7(32'hbb3ce387),
	.w8(32'hba1f01b7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac33894),
	.w1(32'h3af77645),
	.w2(32'h390cbecf),
	.w3(32'hbab8209b),
	.w4(32'h3aa8cab9),
	.w5(32'hb94fe5a9),
	.w6(32'hba079064),
	.w7(32'hba1e7634),
	.w8(32'hbb8ab83c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9397e1),
	.w1(32'hbb829b97),
	.w2(32'hbacba1ee),
	.w3(32'hbb619b7b),
	.w4(32'h3be14d9d),
	.w5(32'h3bc13359),
	.w6(32'hbbad12c2),
	.w7(32'h3ae3b995),
	.w8(32'hb9d4fc2f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d8a4),
	.w1(32'hbb4c320c),
	.w2(32'hbb2bccbf),
	.w3(32'hbb61c873),
	.w4(32'hbb414ff9),
	.w5(32'hbb0f07d7),
	.w6(32'hbbc6c31f),
	.w7(32'hbb298f28),
	.w8(32'hbacf04b6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b7eb5),
	.w1(32'hba2cc092),
	.w2(32'hbb368c95),
	.w3(32'hbb2c93bf),
	.w4(32'h3a7335a8),
	.w5(32'h3aa129ae),
	.w6(32'hbb92a2eb),
	.w7(32'hb99d980e),
	.w8(32'h3b0e90cb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a2c9d),
	.w1(32'h3afc6594),
	.w2(32'h38857a34),
	.w3(32'h3b9fdaa1),
	.w4(32'h3b885c65),
	.w5(32'h3be77991),
	.w6(32'hbb275d99),
	.w7(32'hbab2ae7b),
	.w8(32'h3b8df35f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d24ee),
	.w1(32'hbab7f91c),
	.w2(32'hbba1a6a4),
	.w3(32'h3b89d050),
	.w4(32'hbb9cd015),
	.w5(32'hbc1f84b3),
	.w6(32'h3b1a22f1),
	.w7(32'hbbe948d4),
	.w8(32'hbac95476),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06225f),
	.w1(32'hbaa40269),
	.w2(32'h3b4e741d),
	.w3(32'h3800ba94),
	.w4(32'h3b2cacb5),
	.w5(32'hbab5457a),
	.w6(32'h3b3f63a4),
	.w7(32'h3b637dba),
	.w8(32'hbaeaa698),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5f0aa),
	.w1(32'h3b2969b5),
	.w2(32'hbb59b6fc),
	.w3(32'h39eb94ff),
	.w4(32'h3a2a9075),
	.w5(32'h3b8e3e2e),
	.w6(32'h3a550601),
	.w7(32'hbb4a3d2b),
	.w8(32'h3aa3482d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d8ed),
	.w1(32'h3b9b0af8),
	.w2(32'hb993c290),
	.w3(32'h3ba4bfe7),
	.w4(32'h3af1e44d),
	.w5(32'hb9d9f58e),
	.w6(32'h3b7f6907),
	.w7(32'h3b9f0570),
	.w8(32'h3b43532b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0da2bd),
	.w1(32'hbbe5ed6d),
	.w2(32'h3aa17e94),
	.w3(32'hbbc0f7b8),
	.w4(32'h3b10436d),
	.w5(32'h3c158bac),
	.w6(32'h3aab3ab3),
	.w7(32'hbabd3384),
	.w8(32'h3c2005e2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c925cce),
	.w1(32'h3b2dae7f),
	.w2(32'hba6c5bf9),
	.w3(32'h3b8f2f89),
	.w4(32'h3a7b97a8),
	.w5(32'h3b66dffc),
	.w6(32'h3b2c2246),
	.w7(32'h3ac304dd),
	.w8(32'h39fc40ba),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68484d),
	.w1(32'hbb604431),
	.w2(32'hbad26448),
	.w3(32'hbb72b477),
	.w4(32'hbb3a2357),
	.w5(32'hbb1acd10),
	.w6(32'hbb41cdfe),
	.w7(32'hbb783610),
	.w8(32'hbb548b16),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e951f),
	.w1(32'hbb14c7c5),
	.w2(32'h3ad14ccb),
	.w3(32'hbae21493),
	.w4(32'hba844eae),
	.w5(32'h39a9e13e),
	.w6(32'hbb2f6b30),
	.w7(32'h3b4887f5),
	.w8(32'hbb4187c7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a125cbb),
	.w1(32'h3a527f4d),
	.w2(32'h3bf2dd84),
	.w3(32'h3ba610c7),
	.w4(32'h3b1c4f85),
	.w5(32'hba38fa4c),
	.w6(32'hbac8f0b8),
	.w7(32'hbaad2793),
	.w8(32'hba98cfc5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f99bb),
	.w1(32'h3bca0805),
	.w2(32'h3b2f0bdb),
	.w3(32'h3b5c49b7),
	.w4(32'hbaa94432),
	.w5(32'hbaaff638),
	.w6(32'h3b1297bc),
	.w7(32'hbb57a27f),
	.w8(32'h38b01882),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0ed45),
	.w1(32'hbc1c4566),
	.w2(32'hbab81adf),
	.w3(32'hbc15cab2),
	.w4(32'hbac97a2a),
	.w5(32'hbad8f54c),
	.w6(32'hbbe0ce4f),
	.w7(32'hbab97ae5),
	.w8(32'hbb7c8df2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fcbcd),
	.w1(32'hbb3f0301),
	.w2(32'h3aed3c25),
	.w3(32'hbae75cf0),
	.w4(32'hbb6394f3),
	.w5(32'hbb88824e),
	.w6(32'hbb48fb5b),
	.w7(32'h3a84276b),
	.w8(32'hbaa67610),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bc837),
	.w1(32'hbb4ea931),
	.w2(32'hbc1b0afb),
	.w3(32'hbbb2876d),
	.w4(32'hbc083b6e),
	.w5(32'hbaf782e0),
	.w6(32'hbba0364f),
	.w7(32'hbbf25493),
	.w8(32'h3b591051),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb9774),
	.w1(32'hbbeb057a),
	.w2(32'hbbc06824),
	.w3(32'hbb618ade),
	.w4(32'hbbdc0a24),
	.w5(32'hbbc8fa2c),
	.w6(32'hbae4e4b4),
	.w7(32'hbbf92978),
	.w8(32'hbc17932f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc667f9),
	.w1(32'hbb851c97),
	.w2(32'h396d0cf1),
	.w3(32'hbb73eecb),
	.w4(32'h3b1a97b0),
	.w5(32'hbb840bdb),
	.w6(32'hbb8b30ef),
	.w7(32'hba8c5d21),
	.w8(32'hbbdec783),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fc6b7),
	.w1(32'hbb59ba39),
	.w2(32'h3bf7bded),
	.w3(32'hbbbf86bf),
	.w4(32'hbb493f78),
	.w5(32'h3a84211b),
	.w6(32'hbb9c6742),
	.w7(32'h3ae5423e),
	.w8(32'h3bd6bf2c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65c5e0),
	.w1(32'h3b5771c0),
	.w2(32'h3b9bc44a),
	.w3(32'h3b8360d0),
	.w4(32'h3b804b60),
	.w5(32'h3bbaa927),
	.w6(32'h3b965c4f),
	.w7(32'h3bac58c1),
	.w8(32'h3bd50fae),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88248a),
	.w1(32'hba97f218),
	.w2(32'h3bec61d4),
	.w3(32'h3927d031),
	.w4(32'hba91328b),
	.w5(32'h3b143b27),
	.w6(32'hba2c28e0),
	.w7(32'h3b9b6d7f),
	.w8(32'hba9c491f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c070be1),
	.w1(32'h3b84b871),
	.w2(32'h3b326773),
	.w3(32'h3c03f076),
	.w4(32'hbc0eb2e5),
	.w5(32'hbb1b9c41),
	.w6(32'h3c0fed21),
	.w7(32'hbad4508c),
	.w8(32'h3b4332d5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba309535),
	.w1(32'h3a88ff41),
	.w2(32'h3b497fbf),
	.w3(32'hbae16d5e),
	.w4(32'h3c0aef9f),
	.w5(32'h3b378948),
	.w6(32'hbae65c34),
	.w7(32'h3b28dd12),
	.w8(32'h3b1c112a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8df05b),
	.w1(32'hbade4677),
	.w2(32'hba55ed6c),
	.w3(32'h3bc69edf),
	.w4(32'h3b1c83c3),
	.w5(32'h397ea3e0),
	.w6(32'hba77f94d),
	.w7(32'h3a9e6e33),
	.w8(32'hbadb3a6e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafde882),
	.w1(32'hba7818c0),
	.w2(32'hb9ebbd46),
	.w3(32'hb9830a63),
	.w4(32'hbb0cb25d),
	.w5(32'hba57b521),
	.w6(32'hbaf09698),
	.w7(32'h3a8ee513),
	.w8(32'hba8bf265),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec22e),
	.w1(32'h3b19bf62),
	.w2(32'hbadac8ee),
	.w3(32'h39c3f993),
	.w4(32'hb9f76e7e),
	.w5(32'hbac7a1fd),
	.w6(32'h3b775b73),
	.w7(32'hba3d5a98),
	.w8(32'hbb8a4f27),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb372bf),
	.w1(32'hbb892bef),
	.w2(32'hbb8dba35),
	.w3(32'hbb803eac),
	.w4(32'h3aa807a0),
	.w5(32'hbb374e98),
	.w6(32'hbbf15a04),
	.w7(32'hbbd48f1e),
	.w8(32'hbb9a8282),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cfa9c),
	.w1(32'h3c0e8a79),
	.w2(32'hb9fec641),
	.w3(32'hbb63bdf5),
	.w4(32'hbb780b20),
	.w5(32'hbaf5936f),
	.w6(32'hbb17c852),
	.w7(32'hbb293270),
	.w8(32'hbb0ab930),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b778d6),
	.w1(32'h3b054e8a),
	.w2(32'hba2ec101),
	.w3(32'hb9ed4ffb),
	.w4(32'hba018a55),
	.w5(32'hba8346b3),
	.w6(32'h3b61ffcb),
	.w7(32'hba4dcbdf),
	.w8(32'hbb07bd27),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36bbdd),
	.w1(32'hbb40d23f),
	.w2(32'hbbad23f0),
	.w3(32'hbb016271),
	.w4(32'hba1a45de),
	.w5(32'h3b8fd3f9),
	.w6(32'hbb67c50c),
	.w7(32'hba3c0d31),
	.w8(32'hba961e48),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe251bd),
	.w1(32'h3b719916),
	.w2(32'hbb7d67ee),
	.w3(32'hb7892e7f),
	.w4(32'hbbb5dd32),
	.w5(32'hbb56051c),
	.w6(32'hba52db48),
	.w7(32'hbba69249),
	.w8(32'hbbb4583e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf07b4b),
	.w1(32'hbbabb8d0),
	.w2(32'hbb047fcd),
	.w3(32'hbaa09ebe),
	.w4(32'hba93df6b),
	.w5(32'hbabb62b5),
	.w6(32'hbb8da00a),
	.w7(32'hba499788),
	.w8(32'hbb0f6596),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7b9b4),
	.w1(32'hbbdf3f58),
	.w2(32'h3b89d7d3),
	.w3(32'hbb82cc2f),
	.w4(32'h3b4b0a25),
	.w5(32'hbacf031d),
	.w6(32'hbb685edb),
	.w7(32'h3b1ef208),
	.w8(32'hbbc55876),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b577d34),
	.w1(32'h3ba51327),
	.w2(32'hbb1fa221),
	.w3(32'hba4ef209),
	.w4(32'hbb1e3419),
	.w5(32'hbb863e0d),
	.w6(32'hb920ffd4),
	.w7(32'hbb1daced),
	.w8(32'hbaeafb22),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule