module layer_10_featuremap_20(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fe83b),
	.w1(32'hbc1ef4a4),
	.w2(32'hbbd3fe6f),
	.w3(32'hbceac8e4),
	.w4(32'hbcf21d76),
	.w5(32'hbb448cfe),
	.w6(32'hba381828),
	.w7(32'hbca2196d),
	.w8(32'h3bdaf00e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc130cd3),
	.w1(32'hbc4b5951),
	.w2(32'hbcacc0ce),
	.w3(32'hbc4c19bd),
	.w4(32'hbcb7d1fd),
	.w5(32'hbd100252),
	.w6(32'hbb3659ff),
	.w7(32'hbc293c36),
	.w8(32'hbcb6825d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc976a71),
	.w1(32'hbbed1ab0),
	.w2(32'hbadfecad),
	.w3(32'hbce22817),
	.w4(32'hbc20a6fe),
	.w5(32'hbaef0057),
	.w6(32'hbccbadf4),
	.w7(32'hbc203116),
	.w8(32'h3b656a02),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03c8c2),
	.w1(32'hbb86bd31),
	.w2(32'h3c454c41),
	.w3(32'hbb90cd57),
	.w4(32'hbbca32f9),
	.w5(32'h3b15171d),
	.w6(32'hbbaf2c6e),
	.w7(32'hbb3e671f),
	.w8(32'hbb271a93),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39774a02),
	.w1(32'hbc0698e9),
	.w2(32'hbc2de23b),
	.w3(32'hbc3ebfb7),
	.w4(32'hbcd31d65),
	.w5(32'hbc82a9ee),
	.w6(32'hbc8f2426),
	.w7(32'hbc42f36c),
	.w8(32'hbcddd854),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0fe909),
	.w1(32'hbcbf6915),
	.w2(32'h3b3bf42d),
	.w3(32'hbd426439),
	.w4(32'hbcb82308),
	.w5(32'hbab7aff1),
	.w6(32'hbd138f5e),
	.w7(32'hbc7463d0),
	.w8(32'hbb08113a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37d862),
	.w1(32'h3a17d2ca),
	.w2(32'hbbe61b1d),
	.w3(32'h3bbe651d),
	.w4(32'hbaa8dcfa),
	.w5(32'h3ac912ec),
	.w6(32'h3b49ac28),
	.w7(32'hb96810b1),
	.w8(32'h38e6dce8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ef6e3),
	.w1(32'hbc2e09d3),
	.w2(32'h3a4d7c06),
	.w3(32'h3c40baa9),
	.w4(32'h3baef040),
	.w5(32'h3a9c9dde),
	.w6(32'hbb27ec7f),
	.w7(32'hbc301ae2),
	.w8(32'hbc3a6253),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a06bf),
	.w1(32'hbab0da2d),
	.w2(32'hba5737f0),
	.w3(32'hbbc2896c),
	.w4(32'hbc5aefe4),
	.w5(32'hbb700c5c),
	.w6(32'hbadf47db),
	.w7(32'h3b2cc8b0),
	.w8(32'hbbf07c64),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea1e6b),
	.w1(32'h3ca34351),
	.w2(32'hbb2c8309),
	.w3(32'h3c93653e),
	.w4(32'h3d03ca0b),
	.w5(32'hba386a49),
	.w6(32'h3c53bc3a),
	.w7(32'h3cd70466),
	.w8(32'h3983698c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3de35),
	.w1(32'h3bbeea0a),
	.w2(32'hbc1ae75a),
	.w3(32'h3ba57117),
	.w4(32'h3be1e3e8),
	.w5(32'hbb45f36d),
	.w6(32'h3b3c013c),
	.w7(32'h3b4e4c67),
	.w8(32'hbb6da374),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4899c),
	.w1(32'hbbb10e28),
	.w2(32'hbbffb815),
	.w3(32'h3b779ea4),
	.w4(32'hbb7b5407),
	.w5(32'hbbe016e1),
	.w6(32'h3c0d8a11),
	.w7(32'h3af3980f),
	.w8(32'hbb808fbd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadec527),
	.w1(32'hbb9fdb5a),
	.w2(32'hbc17e70b),
	.w3(32'h3b434258),
	.w4(32'h3a000a3e),
	.w5(32'hbbdf6af1),
	.w6(32'h3bb1a754),
	.w7(32'hb93737b3),
	.w8(32'h3b11897e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba897c5a),
	.w1(32'h3bba5407),
	.w2(32'h3b1dd587),
	.w3(32'h3b130dde),
	.w4(32'h3aa99d76),
	.w5(32'h3b887296),
	.w6(32'h3ad152f8),
	.w7(32'h3bbf8218),
	.w8(32'h3b187bd1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae255d2),
	.w1(32'hbb845e6c),
	.w2(32'h3b48a590),
	.w3(32'hbbf12b10),
	.w4(32'hbb7e5ce1),
	.w5(32'h3b053753),
	.w6(32'h3baeab33),
	.w7(32'h3c68d94e),
	.w8(32'hbbf7fbad),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf6f0c),
	.w1(32'h3b4c9600),
	.w2(32'hbbc9cb46),
	.w3(32'hbb0d3d47),
	.w4(32'h3ba76dbd),
	.w5(32'hbb8559ac),
	.w6(32'hbc286624),
	.w7(32'hbaf4c22b),
	.w8(32'hbbb6b0f2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56340c),
	.w1(32'h3babe34a),
	.w2(32'h3a558101),
	.w3(32'hb93de4b7),
	.w4(32'h3b86cc5c),
	.w5(32'h3b1ec538),
	.w6(32'h387a3b40),
	.w7(32'h3b372638),
	.w8(32'h3b846846),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6b159),
	.w1(32'hb9a4653d),
	.w2(32'hbc59a2d6),
	.w3(32'h3b73afe9),
	.w4(32'h395e3390),
	.w5(32'hbc3a50d6),
	.w6(32'hbb53504f),
	.w7(32'hbacedc77),
	.w8(32'hbc1e89b4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41185d),
	.w1(32'hb9f82616),
	.w2(32'hbbb810c9),
	.w3(32'h3b9370a9),
	.w4(32'hba3471e9),
	.w5(32'hbb483136),
	.w6(32'h3b240f42),
	.w7(32'hbc03abe8),
	.w8(32'h3ba34011),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b6131),
	.w1(32'hbc3cb1b6),
	.w2(32'hbbd25e83),
	.w3(32'hbbf6b6a4),
	.w4(32'hbc323273),
	.w5(32'h3a8ef7f2),
	.w6(32'h3c5c1b1f),
	.w7(32'h3b596459),
	.w8(32'hbb197ff1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0310fe),
	.w1(32'hbc0a3f95),
	.w2(32'h3ab49515),
	.w3(32'hbba3a634),
	.w4(32'hbc0f88be),
	.w5(32'h3c5ac379),
	.w6(32'hbb90fdc4),
	.w7(32'hbbbefbe8),
	.w8(32'h3b4b709f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dd2f9),
	.w1(32'h3c43a9a0),
	.w2(32'hbb0a7aea),
	.w3(32'h3c48c059),
	.w4(32'h3c317fb7),
	.w5(32'h3a1e81da),
	.w6(32'h3b4c5483),
	.w7(32'h3bebf935),
	.w8(32'h39fcf21a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc527440),
	.w1(32'hbc907c3f),
	.w2(32'hbc143343),
	.w3(32'hbc678276),
	.w4(32'hbc98dd70),
	.w5(32'hbadc1b6c),
	.w6(32'hba96e184),
	.w7(32'hbbc43bd9),
	.w8(32'hbba97b20),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ea6d7),
	.w1(32'h3a501a5c),
	.w2(32'h3ba69b49),
	.w3(32'h3b6d9c9c),
	.w4(32'h3b9b4b9c),
	.w5(32'h3bdff4b0),
	.w6(32'h3b929c6e),
	.w7(32'h3b886b85),
	.w8(32'h3bd5c375),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae902c0),
	.w1(32'h3c6b947d),
	.w2(32'h3b511e42),
	.w3(32'hbb4acb83),
	.w4(32'h3c379cd1),
	.w5(32'h3c5f3c0f),
	.w6(32'hba203f9e),
	.w7(32'h3bc67421),
	.w8(32'h3ca06b30),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd386c6),
	.w1(32'hbc1eb8a3),
	.w2(32'hbaae0f98),
	.w3(32'hbb59f400),
	.w4(32'hba804d8b),
	.w5(32'h3bf5191f),
	.w6(32'h3bbb1543),
	.w7(32'hba67fc42),
	.w8(32'h3bd3c217),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedd355),
	.w1(32'h3aa2be6f),
	.w2(32'h39b7d6e3),
	.w3(32'h3b8f2c04),
	.w4(32'hbba29944),
	.w5(32'hb98ae8b3),
	.w6(32'h3c0113ee),
	.w7(32'hbbc1e549),
	.w8(32'h3965e5f8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000a1b),
	.w1(32'h3accb5cf),
	.w2(32'hbbabfe78),
	.w3(32'hbb24bd6f),
	.w4(32'h3a98630f),
	.w5(32'hbc3b0a3d),
	.w6(32'hbaa33d7b),
	.w7(32'h3b176158),
	.w8(32'hbc490943),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb604cc),
	.w1(32'h3b2cb28b),
	.w2(32'hbbbd01a6),
	.w3(32'hbbb0ca9e),
	.w4(32'hbb5e7184),
	.w5(32'hbbbcd417),
	.w6(32'hbbbd20e3),
	.w7(32'hbaf5ed4a),
	.w8(32'hbb114822),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c3f51),
	.w1(32'h3bd4471c),
	.w2(32'h3bf6ae59),
	.w3(32'hbbf9c52e),
	.w4(32'h3bac2889),
	.w5(32'h3b512e3e),
	.w6(32'hbb272307),
	.w7(32'h3bacb3a1),
	.w8(32'h3bbc0f80),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60c14a),
	.w1(32'h3b6b3c5c),
	.w2(32'hbb84cf7b),
	.w3(32'hb9dce7dc),
	.w4(32'h3b44cfa0),
	.w5(32'h3a77faea),
	.w6(32'h3af7e4d5),
	.w7(32'h3b7a347a),
	.w8(32'hba49263a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe15ba4),
	.w1(32'hbaa2f28b),
	.w2(32'hbc2ec234),
	.w3(32'hbba2078b),
	.w4(32'h3bac96a4),
	.w5(32'hbc287122),
	.w6(32'hbbc6ce59),
	.w7(32'hbae66dc8),
	.w8(32'hb92be4e2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc486481),
	.w1(32'hbbcb279a),
	.w2(32'hbc17c99c),
	.w3(32'hbbc0a88f),
	.w4(32'h3b1d255d),
	.w5(32'hbc724717),
	.w6(32'hbadd0355),
	.w7(32'h3ba36b57),
	.w8(32'hbbd03e15),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a316a),
	.w1(32'h3b0110c3),
	.w2(32'h3b31028c),
	.w3(32'hbb92b353),
	.w4(32'h3ba59562),
	.w5(32'h3b4daec4),
	.w6(32'h3af82893),
	.w7(32'h3b805478),
	.w8(32'hbb4858d2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8cd36),
	.w1(32'hbc544740),
	.w2(32'hbaa63f83),
	.w3(32'hbc2f9789),
	.w4(32'hbc6f35d2),
	.w5(32'hbb4f3a25),
	.w6(32'hbc80ba8b),
	.w7(32'hbc4191ac),
	.w8(32'h3ade8f8c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc27e0a),
	.w1(32'h3b3f5bf8),
	.w2(32'hbc46e876),
	.w3(32'h3b96ca85),
	.w4(32'h3b4f728f),
	.w5(32'hbc06eac6),
	.w6(32'h3b23ab6c),
	.w7(32'h3ae704dd),
	.w8(32'hb9915215),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb794b0),
	.w1(32'h3c497387),
	.w2(32'hbccb875c),
	.w3(32'h3c7abc82),
	.w4(32'h3cd0e267),
	.w5(32'hbce1d16f),
	.w6(32'h3c04d8db),
	.w7(32'h3c708778),
	.w8(32'hbc8fe2bf),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2919e0),
	.w1(32'h3c40249d),
	.w2(32'h3b32a049),
	.w3(32'hbc1f595d),
	.w4(32'h3c41d5aa),
	.w5(32'h3b6ecf6c),
	.w6(32'hb9acccf2),
	.w7(32'h3c7f93de),
	.w8(32'h3bdfa0e6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40a953),
	.w1(32'h3c0013c8),
	.w2(32'h3b8f01c1),
	.w3(32'hbc6900c0),
	.w4(32'h3c01513d),
	.w5(32'h3ba5acc8),
	.w6(32'hb9164382),
	.w7(32'h3c497f6a),
	.w8(32'h3c4ea83e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb068c24),
	.w1(32'hbb445e7d),
	.w2(32'h3b243e8d),
	.w3(32'hbbfff714),
	.w4(32'hbbf9145b),
	.w5(32'h3bb04aae),
	.w6(32'hbaaad3f0),
	.w7(32'hbc008e9c),
	.w8(32'h3b489995),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025d34),
	.w1(32'hb9166aef),
	.w2(32'hbc2eb084),
	.w3(32'hbb44b789),
	.w4(32'h3a5fe37c),
	.w5(32'hbbf78752),
	.w6(32'hbab1a382),
	.w7(32'hba67c9f8),
	.w8(32'hbb96ae7d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6f7df),
	.w1(32'hba0677bf),
	.w2(32'hba3614d6),
	.w3(32'hbc287ec3),
	.w4(32'hbab9a222),
	.w5(32'h3aa3db39),
	.w6(32'hbb028714),
	.w7(32'hbb6f5152),
	.w8(32'h3b78970f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f02ad),
	.w1(32'h3b5741dc),
	.w2(32'hbac6577c),
	.w3(32'hbbd15c97),
	.w4(32'hba84f664),
	.w5(32'hbb144890),
	.w6(32'hbb9b8729),
	.w7(32'hbaae355a),
	.w8(32'hba54efdf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f26e1),
	.w1(32'hbbd8121f),
	.w2(32'h39bff858),
	.w3(32'h3b3a9d90),
	.w4(32'hbb1cfe24),
	.w5(32'h3a82aa83),
	.w6(32'h3ac6d9a8),
	.w7(32'hba7dee60),
	.w8(32'h3b8e15ac),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb633f27),
	.w1(32'hbb064756),
	.w2(32'hbbedc60e),
	.w3(32'hbbae68eb),
	.w4(32'hbb1dafc2),
	.w5(32'hbb515eea),
	.w6(32'hbbb8814c),
	.w7(32'h3b316eed),
	.w8(32'hbae13620),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc174ed6),
	.w1(32'hb8e914d7),
	.w2(32'hbbb88aea),
	.w3(32'hbbc2cad0),
	.w4(32'hbc063fb7),
	.w5(32'hbbc59e8a),
	.w6(32'hbbbba491),
	.w7(32'h37796117),
	.w8(32'h38e11f8c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25771e),
	.w1(32'hbc137ad6),
	.w2(32'h3aa036c0),
	.w3(32'hbc7ab46d),
	.w4(32'hbc2801d5),
	.w5(32'h3bac49de),
	.w6(32'hbc22b5ec),
	.w7(32'hbbba40b6),
	.w8(32'h3c14e84c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ca494),
	.w1(32'hbbeee7ed),
	.w2(32'hbc6f5a2f),
	.w3(32'h3b461580),
	.w4(32'hbb993ca0),
	.w5(32'hbc0b0793),
	.w6(32'hbaf76607),
	.w7(32'hbc2aede1),
	.w8(32'hbc196ad3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a300a0e),
	.w1(32'hbb002da2),
	.w2(32'hbbc59548),
	.w3(32'hb9090fd5),
	.w4(32'hbb680c2e),
	.w5(32'h3a6986fa),
	.w6(32'hbb24acba),
	.w7(32'hbb90820b),
	.w8(32'hbc15ec29),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16eeec),
	.w1(32'h3a7ffa7f),
	.w2(32'hbc1760ae),
	.w3(32'hbbadd867),
	.w4(32'hbb92eb16),
	.w5(32'hba410017),
	.w6(32'h3a9c238d),
	.w7(32'hbb954a02),
	.w8(32'hbb3d6126),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb134ce),
	.w1(32'hbbb96a77),
	.w2(32'h3c02ab8e),
	.w3(32'h3baa3e88),
	.w4(32'hbad24b7c),
	.w5(32'h3cccc9ac),
	.w6(32'hbb8628bb),
	.w7(32'hbbea27d2),
	.w8(32'h3c412320),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aafe4),
	.w1(32'hbb083ef5),
	.w2(32'hbc6aea9f),
	.w3(32'h3b18639b),
	.w4(32'hbc44fd91),
	.w5(32'h3a07c71a),
	.w6(32'hbbf71031),
	.w7(32'hbc519949),
	.w8(32'hbc395489),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacef24c),
	.w1(32'hbba4a663),
	.w2(32'hbbbadc7a),
	.w3(32'h3a36ceab),
	.w4(32'hbb8f4bd1),
	.w5(32'h3b19edf1),
	.w6(32'hbbc5ec3c),
	.w7(32'hbc0b3657),
	.w8(32'h3b033185),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f2b8e),
	.w1(32'hbbc0519f),
	.w2(32'hbca4fcd9),
	.w3(32'h3bdd044a),
	.w4(32'hbbb43b44),
	.w5(32'hbc854783),
	.w6(32'hba030189),
	.w7(32'hbc1aa982),
	.w8(32'hbbedb548),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b4567),
	.w1(32'h3afa85c7),
	.w2(32'hbba3e145),
	.w3(32'h3bf44a1a),
	.w4(32'hbaf76292),
	.w5(32'hbbcab59d),
	.w6(32'h3bbe8fbc),
	.w7(32'h3bd91bf9),
	.w8(32'hbaed8f32),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a5075),
	.w1(32'hbadb460b),
	.w2(32'h3b6e2c9a),
	.w3(32'hbb304ade),
	.w4(32'hbaa8997a),
	.w5(32'h3b90fd30),
	.w6(32'hbb8d4810),
	.w7(32'h3b9ecab4),
	.w8(32'h3c11567d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f7e2),
	.w1(32'h3943104e),
	.w2(32'hbc659a41),
	.w3(32'h3b76bc5f),
	.w4(32'h3a9169be),
	.w5(32'hbcc786d7),
	.w6(32'h3b1b26c7),
	.w7(32'hba7e8b3d),
	.w8(32'hbcd0b97a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b4ffa),
	.w1(32'hbacc99e8),
	.w2(32'hbae46a00),
	.w3(32'hbc95d1ab),
	.w4(32'hbb07e33d),
	.w5(32'hbb22c316),
	.w6(32'hbc4f9939),
	.w7(32'h3a418ff0),
	.w8(32'h3b8d8403),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385e7c2e),
	.w1(32'hbbc33a0c),
	.w2(32'hbc11a2ed),
	.w3(32'h3b2cae03),
	.w4(32'hbbb9dc15),
	.w5(32'hbc64f097),
	.w6(32'h3c1513f4),
	.w7(32'hb9a6c598),
	.w8(32'hbc5b14e3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc269dc2),
	.w1(32'hbba653f8),
	.w2(32'h3a584455),
	.w3(32'hbc49e2c4),
	.w4(32'hbbb70adc),
	.w5(32'hbbbeecf5),
	.w6(32'hbba8a733),
	.w7(32'hbb427150),
	.w8(32'hbc8041d1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde1514),
	.w1(32'hbb966aa4),
	.w2(32'hbc0fa812),
	.w3(32'hbc1d1193),
	.w4(32'hba95c12b),
	.w5(32'hbc40eb0c),
	.w6(32'hbc07c0bd),
	.w7(32'h3b05acd0),
	.w8(32'hbc18b79d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0313d5),
	.w1(32'hbba80188),
	.w2(32'hbc4ab212),
	.w3(32'hbb92c074),
	.w4(32'hbc015899),
	.w5(32'hbc6be6b5),
	.w6(32'hbb572001),
	.w7(32'hbb246b04),
	.w8(32'hbc92ef72),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2de2d3),
	.w1(32'hbb587584),
	.w2(32'hbb1092f2),
	.w3(32'hbaf6ddf7),
	.w4(32'h3b4dc4ea),
	.w5(32'hbb9c0922),
	.w6(32'hbbc70952),
	.w7(32'hb87efb04),
	.w8(32'h3b37676b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57f5e2),
	.w1(32'h3b88c70a),
	.w2(32'h3b3a2085),
	.w3(32'h3c1ddb5d),
	.w4(32'h3c3c974d),
	.w5(32'hbb9d2917),
	.w6(32'h3b709546),
	.w7(32'h3ac1ba9c),
	.w8(32'hbb9c98d9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac197d5),
	.w1(32'hbb9819ce),
	.w2(32'hbb5e04ba),
	.w3(32'hba792601),
	.w4(32'h38c9c5c7),
	.w5(32'hbba76db6),
	.w6(32'hb9689d5c),
	.w7(32'hbb901756),
	.w8(32'hbb38b2f5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b4864),
	.w1(32'hba84613d),
	.w2(32'hb89111a7),
	.w3(32'hbb86ee59),
	.w4(32'hba760e8a),
	.w5(32'hbb57e2eb),
	.w6(32'hbb20dd7f),
	.w7(32'hba70dc61),
	.w8(32'hba5dbe89),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb71df),
	.w1(32'hbc61664a),
	.w2(32'hbcea0be9),
	.w3(32'h3c1f9ab9),
	.w4(32'h39703f72),
	.w5(32'hbc6e202f),
	.w6(32'h3b1c6f0c),
	.w7(32'hba33c882),
	.w8(32'hbb9e4058),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca97f81),
	.w1(32'h3b882512),
	.w2(32'hbc0344bf),
	.w3(32'h3a924563),
	.w4(32'h3b5ba8f7),
	.w5(32'hbbf24b50),
	.w6(32'h3be2e86b),
	.w7(32'hbb6c8dd1),
	.w8(32'hbba56cb2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd47cf),
	.w1(32'hbaa6fcd9),
	.w2(32'hbb3648da),
	.w3(32'h3a979dce),
	.w4(32'hbaad5eee),
	.w5(32'hbaf003ea),
	.w6(32'h3aa32510),
	.w7(32'hbb3886b0),
	.w8(32'hbb270c7f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9eab9),
	.w1(32'h3c7e68e9),
	.w2(32'h3cba0763),
	.w3(32'hbbf6d959),
	.w4(32'h3c3b3510),
	.w5(32'h3d002d00),
	.w6(32'hbb29ac77),
	.w7(32'h3c43f43e),
	.w8(32'h3ce9949a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4de509),
	.w1(32'hbab7d9e7),
	.w2(32'hba4d5af7),
	.w3(32'h3c5aef5c),
	.w4(32'hbb84952a),
	.w5(32'hbc0b93be),
	.w6(32'h3baec53b),
	.w7(32'hbbf41939),
	.w8(32'hbbd6b967),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da100),
	.w1(32'h3a156435),
	.w2(32'hbb7837d8),
	.w3(32'hbbb1af70),
	.w4(32'hbac10ecd),
	.w5(32'hbc1c9535),
	.w6(32'hbbbc511b),
	.w7(32'h3aa71d84),
	.w8(32'hb7bfe0b5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc80a83),
	.w1(32'hba4e4b2f),
	.w2(32'h3afb3b64),
	.w3(32'hbc0da081),
	.w4(32'h3ac78a39),
	.w5(32'hbb8277f2),
	.w6(32'h3b5f1362),
	.w7(32'h3ba7670a),
	.w8(32'hba695688),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf12109),
	.w1(32'h39569633),
	.w2(32'hbb47d628),
	.w3(32'h3bb0aa99),
	.w4(32'h3b8df7ea),
	.w5(32'hbb616de7),
	.w6(32'h3b8007dd),
	.w7(32'h3ab8eedf),
	.w8(32'hbb27e31f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16aac8),
	.w1(32'hbb3b8aeb),
	.w2(32'hbc29076e),
	.w3(32'hbb981a9f),
	.w4(32'hbc05814a),
	.w5(32'hbc47b402),
	.w6(32'hbb8f80d3),
	.w7(32'hbc0a7ef7),
	.w8(32'hbc274270),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc217906),
	.w1(32'hbaebbb4e),
	.w2(32'hbbf9d1e8),
	.w3(32'hbbae4b08),
	.w4(32'h3bcf4dfe),
	.w5(32'h3b2e7a4b),
	.w6(32'hbaac05ee),
	.w7(32'h3bde8b11),
	.w8(32'h3a726e07),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce087e),
	.w1(32'hba4b46a8),
	.w2(32'hbc16935d),
	.w3(32'h3b314934),
	.w4(32'hba934866),
	.w5(32'hbbe5ef42),
	.w6(32'hbb14ff94),
	.w7(32'h3b57c803),
	.w8(32'hbc4ab33d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1baf14),
	.w1(32'h3aea4ad7),
	.w2(32'h3935dd15),
	.w3(32'hbae4c612),
	.w4(32'h3ae37278),
	.w5(32'hbba20530),
	.w6(32'hbac7f2b9),
	.w7(32'h3b8ea31a),
	.w8(32'h3af29c91),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4808a),
	.w1(32'hbb59cf34),
	.w2(32'hbb7c784b),
	.w3(32'hbba9e80e),
	.w4(32'hbb1578c1),
	.w5(32'hbb2e258c),
	.w6(32'hbbb7f5f0),
	.w7(32'hbc134f92),
	.w8(32'hbb12adbc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b181b4b),
	.w1(32'hbaae5e0d),
	.w2(32'h3a0cddd8),
	.w3(32'h3bb0cc97),
	.w4(32'hb932abec),
	.w5(32'h3c1ab5fc),
	.w6(32'h3b052f4b),
	.w7(32'h3aee6265),
	.w8(32'h3c0b48e6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac589a),
	.w1(32'hb9983226),
	.w2(32'hbc078bcd),
	.w3(32'h3c22467d),
	.w4(32'hbb4a82ab),
	.w5(32'hbc3ebd95),
	.w6(32'h3b957863),
	.w7(32'hbc00cf47),
	.w8(32'hbbcf6321),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab87cf),
	.w1(32'hbb5d084c),
	.w2(32'hbb7f41c6),
	.w3(32'hbba46a52),
	.w4(32'h3ab7c722),
	.w5(32'h3b49e01e),
	.w6(32'h3a47d242),
	.w7(32'h3b787b29),
	.w8(32'h3c029a5f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfff579),
	.w1(32'h3b1de155),
	.w2(32'hb956c4b0),
	.w3(32'h3af166e6),
	.w4(32'hbc366e99),
	.w5(32'hbae51fb5),
	.w6(32'h3bf1734c),
	.w7(32'hbb85d9ee),
	.w8(32'hbb2aebfd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc191a5f),
	.w1(32'hbc1f74c6),
	.w2(32'hbb9c17fb),
	.w3(32'hbc8e7f51),
	.w4(32'hbc22e89b),
	.w5(32'hbc20bbbc),
	.w6(32'hbc4c7845),
	.w7(32'hbbf53d14),
	.w8(32'hbc136f38),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99dff5),
	.w1(32'h3b533560),
	.w2(32'hbac6153f),
	.w3(32'hbb90bb91),
	.w4(32'h3b1ea03e),
	.w5(32'h38bb915b),
	.w6(32'h3c00021b),
	.w7(32'h3c1f72c9),
	.w8(32'hbc02e774),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e123a),
	.w1(32'h3b9c1ce3),
	.w2(32'hbc12280a),
	.w3(32'hbbf52077),
	.w4(32'hbbc26034),
	.w5(32'hbc7ee1c4),
	.w6(32'hbb2a9206),
	.w7(32'hbba4cd3e),
	.w8(32'hbc67ad2c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27d6b8),
	.w1(32'hbab793a4),
	.w2(32'hbb5d9db6),
	.w3(32'hbc35c957),
	.w4(32'hbab8b8e7),
	.w5(32'hb9646739),
	.w6(32'hbbf4b337),
	.w7(32'hb9661bb0),
	.w8(32'h3529f2dc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82bc9a),
	.w1(32'h3b15083e),
	.w2(32'hbc05b38b),
	.w3(32'hbb0ec3a1),
	.w4(32'hbaa886a2),
	.w5(32'hbad1c848),
	.w6(32'hbaf4de86),
	.w7(32'hbac7694a),
	.w8(32'h3b8bca34),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b7041),
	.w1(32'h3b75220f),
	.w2(32'hbadc956e),
	.w3(32'hbb39b607),
	.w4(32'hbc05adb3),
	.w5(32'h3a918ef6),
	.w6(32'h3ad4bd0a),
	.w7(32'hbc11fe22),
	.w8(32'hbb3449e0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac55ee),
	.w1(32'h3a7f1231),
	.w2(32'hbc1005be),
	.w3(32'h3b685f79),
	.w4(32'h399630a7),
	.w5(32'hbc08c9ee),
	.w6(32'h3bd80d92),
	.w7(32'h3a9acbdd),
	.w8(32'hbb6a18ba),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe90d4f),
	.w1(32'hb97efd26),
	.w2(32'h3c1e950b),
	.w3(32'hbb95ad75),
	.w4(32'h3b2f97ab),
	.w5(32'h3b3c8b98),
	.w6(32'h3b8c9a29),
	.w7(32'h3c03d9c6),
	.w8(32'h3b852835),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a835913),
	.w1(32'hbc1f4954),
	.w2(32'hbc56a546),
	.w3(32'h3b68aa6b),
	.w4(32'hbb8045b3),
	.w5(32'hbc0c574d),
	.w6(32'h3b122161),
	.w7(32'hba2313be),
	.w8(32'hbbbcc4b5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39958284),
	.w1(32'h3c2c4ba7),
	.w2(32'h3b8ed691),
	.w3(32'hbb08ea39),
	.w4(32'h3c1782c4),
	.w5(32'h3b3161b2),
	.w6(32'h3acb7e15),
	.w7(32'h3c1cc6ba),
	.w8(32'h3a66a94f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f39b9),
	.w1(32'hbbba091e),
	.w2(32'hbc64b893),
	.w3(32'h3a929c11),
	.w4(32'hbbacb41f),
	.w5(32'hbbbf5325),
	.w6(32'hbb4f657c),
	.w7(32'hbb75bb36),
	.w8(32'hbc0dbea9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94fd13),
	.w1(32'hbb765058),
	.w2(32'hbc084aa9),
	.w3(32'hba1cc03a),
	.w4(32'hbbbc9573),
	.w5(32'hbae073cc),
	.w6(32'h39efbb59),
	.w7(32'hb8a602fe),
	.w8(32'hbc1a62c0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03fbab),
	.w1(32'h3bfd0045),
	.w2(32'hb91ae786),
	.w3(32'hbc4081ad),
	.w4(32'h3bf9c4c2),
	.w5(32'h3beceab9),
	.w6(32'hbbf3dd3a),
	.w7(32'h3c29fe10),
	.w8(32'h3c2391dd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fbeb0),
	.w1(32'h3c0c05ea),
	.w2(32'hbbd7bf44),
	.w3(32'h3bc171c7),
	.w4(32'h3baf4b95),
	.w5(32'hbbcea176),
	.w6(32'h3bce279e),
	.w7(32'h3bb4ed7e),
	.w8(32'h3b3213d6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b7a9d),
	.w1(32'h3b7532fc),
	.w2(32'hbbeb8bf1),
	.w3(32'h3a7345af),
	.w4(32'hbb8ba6bb),
	.w5(32'hbc06586f),
	.w6(32'h3b4e4f0c),
	.w7(32'h3b3f6d8c),
	.w8(32'h3a9ceedf),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae162a),
	.w1(32'hbc067139),
	.w2(32'hbc54fc43),
	.w3(32'hba037286),
	.w4(32'hbb708022),
	.w5(32'hbb835135),
	.w6(32'h3ba90cd4),
	.w7(32'hbc07ec7e),
	.w8(32'hbb57f814),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60af88),
	.w1(32'h3c0b8cb6),
	.w2(32'hbc15f09d),
	.w3(32'h3b105063),
	.w4(32'h3c2d44fb),
	.w5(32'hbc8198da),
	.w6(32'hbb513c38),
	.w7(32'h3b8ab8ab),
	.w8(32'hbc7f8a23),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb802961),
	.w1(32'h3c79d735),
	.w2(32'h3c0e51a0),
	.w3(32'hbc2a8371),
	.w4(32'h3c3f50aa),
	.w5(32'h3c3e7ff4),
	.w6(32'h393e33e5),
	.w7(32'h3c756474),
	.w8(32'h3c50bfef),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb915d4d),
	.w1(32'h3b5a4bda),
	.w2(32'hbb2e6347),
	.w3(32'hbc7d5f91),
	.w4(32'h3ba857c7),
	.w5(32'h3ad80e3a),
	.w6(32'hbc03426e),
	.w7(32'h3ab43bb9),
	.w8(32'h3b93cfa1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b6131),
	.w1(32'h3be64609),
	.w2(32'hbb09e49c),
	.w3(32'h3c28a6a8),
	.w4(32'h3c6813ad),
	.w5(32'h3bd1c0e3),
	.w6(32'h3ba0b482),
	.w7(32'h3c17c034),
	.w8(32'h3c3e1cc3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c159b5d),
	.w1(32'h3a9fbccf),
	.w2(32'h3b8599a3),
	.w3(32'h3c1949c9),
	.w4(32'h3ac16050),
	.w5(32'h3c470cd0),
	.w6(32'h3bda7ed9),
	.w7(32'hbb9d2414),
	.w8(32'h3be55ca5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207f28),
	.w1(32'h3b08ce90),
	.w2(32'hbbf6e1f7),
	.w3(32'h3b864410),
	.w4(32'h3c1d4e2b),
	.w5(32'hbbae9b11),
	.w6(32'hbbd82164),
	.w7(32'hbb95c636),
	.w8(32'hbb3d3e52),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb618707),
	.w1(32'h3b95b989),
	.w2(32'hbb81eecb),
	.w3(32'h3bac52eb),
	.w4(32'h3c0f1abb),
	.w5(32'hbb9a613c),
	.w6(32'h3b7bd7be),
	.w7(32'h3bf1b4f6),
	.w8(32'hbb9253aa),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e7534),
	.w1(32'hbb189df0),
	.w2(32'hbb52a093),
	.w3(32'h3a4a58c8),
	.w4(32'hbbad2f75),
	.w5(32'hbb034627),
	.w6(32'hbb32b888),
	.w7(32'hbc07c6d2),
	.w8(32'h3aa923d9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76cb28),
	.w1(32'hbb4511b1),
	.w2(32'hbb62f116),
	.w3(32'h3744dd48),
	.w4(32'hbbaf7e5a),
	.w5(32'hbc306ade),
	.w6(32'hbb088179),
	.w7(32'hbbc2b89c),
	.w8(32'hbc167bfd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba431977),
	.w1(32'h3b84472a),
	.w2(32'hbb96f22c),
	.w3(32'h3a767406),
	.w4(32'hbaabefa6),
	.w5(32'hbc2083d2),
	.w6(32'h3c60e126),
	.w7(32'h3bcb26e4),
	.w8(32'hbb84fe9e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06d143),
	.w1(32'h3c075c40),
	.w2(32'hba27de31),
	.w3(32'hbc0ed8a6),
	.w4(32'h3b72c1a1),
	.w5(32'hbb2d23e1),
	.w6(32'hbba3498a),
	.w7(32'h3b41f7d0),
	.w8(32'h3a409cf5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fba66),
	.w1(32'hbb24d709),
	.w2(32'h3c4dbcd9),
	.w3(32'hbb780a6a),
	.w4(32'hba5b7161),
	.w5(32'h3c881025),
	.w6(32'hb9e3bb84),
	.w7(32'h3c484d2f),
	.w8(32'h3c8253be),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c8151),
	.w1(32'hbb29d37d),
	.w2(32'hbb957cd9),
	.w3(32'hba603697),
	.w4(32'hbc5f1398),
	.w5(32'h3bb09caf),
	.w6(32'hbbbddd91),
	.w7(32'hbc488597),
	.w8(32'h3c3c4c34),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca73332),
	.w1(32'h3c803e41),
	.w2(32'hba577446),
	.w3(32'h3c4158f5),
	.w4(32'h3baf7abd),
	.w5(32'hbc165cf0),
	.w6(32'h3c1fa6f0),
	.w7(32'h3bc6547a),
	.w8(32'hbbd0be26),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3990e4),
	.w1(32'hbbe258aa),
	.w2(32'hbc2e6987),
	.w3(32'hbc57a931),
	.w4(32'hbc49a598),
	.w5(32'hbc04beb1),
	.w6(32'hbbcb6f3e),
	.w7(32'hbbf4e17c),
	.w8(32'hbbc2cd7e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49b47e),
	.w1(32'h39074961),
	.w2(32'h3b68cb24),
	.w3(32'hbc4ab6bb),
	.w4(32'hbb297104),
	.w5(32'h3b84ed29),
	.w6(32'hbb3c217b),
	.w7(32'hbbc27c9e),
	.w8(32'h3b696853),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924de04),
	.w1(32'hbaf0037f),
	.w2(32'hba55bccb),
	.w3(32'hb91245c0),
	.w4(32'hbb98a481),
	.w5(32'h3a899929),
	.w6(32'hbb26b426),
	.w7(32'hbbc8e623),
	.w8(32'hbb84799d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb47578),
	.w1(32'hb97b8735),
	.w2(32'hbbfa559a),
	.w3(32'h3a730653),
	.w4(32'hbb8a11a6),
	.w5(32'hbc127eba),
	.w6(32'hbc0c8723),
	.w7(32'hbc471a9d),
	.w8(32'hbb60911e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc64dbb),
	.w1(32'hba866158),
	.w2(32'hbac955cb),
	.w3(32'hbb504bde),
	.w4(32'h3a8b65eb),
	.w5(32'hbb71c7b8),
	.w6(32'hbb437de6),
	.w7(32'hbab2a6a3),
	.w8(32'h3b307abf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66e0c2),
	.w1(32'hba2b8170),
	.w2(32'h3b390fcc),
	.w3(32'hbbd048c4),
	.w4(32'hba17d549),
	.w5(32'hbb65b225),
	.w6(32'h3a326ac8),
	.w7(32'h3ac8a4f5),
	.w8(32'hba8ce5bc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29162d),
	.w1(32'h3ab39371),
	.w2(32'hbb016554),
	.w3(32'hbc29e7f3),
	.w4(32'hb695a466),
	.w5(32'hba8ae139),
	.w6(32'hbb7b9b34),
	.w7(32'h3b130311),
	.w8(32'h3a83fb58),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04a9d1),
	.w1(32'hbb460c64),
	.w2(32'h3ad0fac7),
	.w3(32'hbaefc538),
	.w4(32'hbad9bb33),
	.w5(32'h3a3e12ce),
	.w6(32'hba8a1adb),
	.w7(32'h3a6b0393),
	.w8(32'h3a8ca7be),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c6fe5),
	.w1(32'h3ab16a82),
	.w2(32'hbb623dc8),
	.w3(32'h3b9d95dd),
	.w4(32'h3ae408e0),
	.w5(32'hbb29e9c9),
	.w6(32'h3b950a07),
	.w7(32'h3ad0abf6),
	.w8(32'hbb1a61a1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80dfca),
	.w1(32'h3bfac8de),
	.w2(32'h3b284beb),
	.w3(32'hbb6246b2),
	.w4(32'h3bf77879),
	.w5(32'hbb51c698),
	.w6(32'h392652e6),
	.w7(32'h3c1242df),
	.w8(32'h3a0d4be8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae10702),
	.w1(32'h3a87eb9e),
	.w2(32'hbbe06fe0),
	.w3(32'h3ab3e6d4),
	.w4(32'hbb4c85b8),
	.w5(32'hbc2049f8),
	.w6(32'h3ac21c87),
	.w7(32'h3a9c9097),
	.w8(32'hbc14254c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff0073),
	.w1(32'h3ab8d4ce),
	.w2(32'h3bf5d32d),
	.w3(32'hbc1717c9),
	.w4(32'hb9ad71e2),
	.w5(32'h3ca271a9),
	.w6(32'hbbeb760f),
	.w7(32'h3a6d0bd3),
	.w8(32'h3bf16279),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bc626),
	.w1(32'hbbb38e91),
	.w2(32'hbb6c2ddc),
	.w3(32'h3bdd5533),
	.w4(32'hbbb10aef),
	.w5(32'hba925dd9),
	.w6(32'h387cf826),
	.w7(32'hbb2f90f7),
	.w8(32'h3bc6cfa5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1116a),
	.w1(32'h3aafb317),
	.w2(32'h3b0dd0b5),
	.w3(32'h3c3361ca),
	.w4(32'h3a07513e),
	.w5(32'h3a766d38),
	.w6(32'h3c2c0fd4),
	.w7(32'hba8ac997),
	.w8(32'hbbf43194),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2bcbe),
	.w1(32'h3beef6a2),
	.w2(32'hbbff419b),
	.w3(32'h3c16897f),
	.w4(32'h3b2d7981),
	.w5(32'hbc992b43),
	.w6(32'hbb629f2f),
	.w7(32'hbba6d046),
	.w8(32'hbca6837a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0768),
	.w1(32'hbbd3f9b9),
	.w2(32'hbc8d4a94),
	.w3(32'hbb365e30),
	.w4(32'hbc06723a),
	.w5(32'hbc9e8b7c),
	.w6(32'h3b993e03),
	.w7(32'hba3031c1),
	.w8(32'hbc1193e8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcf94f),
	.w1(32'hbbee2fc9),
	.w2(32'hb9ee9f8d),
	.w3(32'hbc0e4644),
	.w4(32'hbc2bf72e),
	.w5(32'hbc2b0a66),
	.w6(32'h3a0ebec0),
	.w7(32'hbb8cb9e9),
	.w8(32'h3a424c9b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00c8bd),
	.w1(32'hb9ce557e),
	.w2(32'hba251ad6),
	.w3(32'hba86d0d3),
	.w4(32'h3aa3c4c3),
	.w5(32'hbb8142fb),
	.w6(32'hbb349944),
	.w7(32'hb946d4a3),
	.w8(32'hbb476d5a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc128e04),
	.w1(32'hbb804516),
	.w2(32'hbb62ff44),
	.w3(32'hbae87d62),
	.w4(32'hbb81c74a),
	.w5(32'hbb4d630a),
	.w6(32'hbc0f238f),
	.w7(32'hbc30ee11),
	.w8(32'h3babec14),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41b86a),
	.w1(32'hbb01e06a),
	.w2(32'hbbaccbd0),
	.w3(32'h3bd53ac3),
	.w4(32'hbb9b8744),
	.w5(32'hbb640d95),
	.w6(32'hbb55326e),
	.w7(32'hbbef2c82),
	.w8(32'hba785df2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ba710),
	.w1(32'hbc37c1d5),
	.w2(32'hbb972310),
	.w3(32'hbb118da2),
	.w4(32'hbc455cef),
	.w5(32'hbb53c787),
	.w6(32'h3b500dd2),
	.w7(32'hbbf8afce),
	.w8(32'h3ae5d289),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c36ec),
	.w1(32'hbbe0f983),
	.w2(32'hbcbebdb1),
	.w3(32'h3b94daa0),
	.w4(32'hbbcbe421),
	.w5(32'hbc31de2d),
	.w6(32'h3bb01438),
	.w7(32'hbb738947),
	.w8(32'hbc284332),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc484052),
	.w1(32'h3a0fc552),
	.w2(32'hbb6abd8d),
	.w3(32'hbbc29602),
	.w4(32'hbb10c771),
	.w5(32'hbc0ac2da),
	.w6(32'hbc372100),
	.w7(32'hbbd8406e),
	.w8(32'hba7ae50e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f05b0),
	.w1(32'hbb68a7aa),
	.w2(32'hbc0d5010),
	.w3(32'hbb5062e6),
	.w4(32'hbb9ff280),
	.w5(32'hbc0dbcca),
	.w6(32'h3b7f9432),
	.w7(32'h39bff0ff),
	.w8(32'hbc146aac),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d6ceb),
	.w1(32'hbb006ed0),
	.w2(32'hbbafcaae),
	.w3(32'hba6db0e4),
	.w4(32'hbae65c18),
	.w5(32'hbbcb68ea),
	.w6(32'h3b9e6434),
	.w7(32'h3ae7667f),
	.w8(32'hbb8ff6e6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69d789),
	.w1(32'h3b963f4f),
	.w2(32'hbb117f07),
	.w3(32'hbb1a9c53),
	.w4(32'h3b79f15f),
	.w5(32'hbb3bfc37),
	.w6(32'hba1de1c2),
	.w7(32'h3b3360c0),
	.w8(32'hbb2b3146),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2898b6),
	.w1(32'hbc567b12),
	.w2(32'hbbc5ea3e),
	.w3(32'hbb98c51f),
	.w4(32'hbbe3eb5c),
	.w5(32'hbbc51837),
	.w6(32'hbbee4ebd),
	.w7(32'hbc409978),
	.w8(32'hbbfbaab7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e66d4f),
	.w1(32'hba8e5e00),
	.w2(32'hbb909152),
	.w3(32'hbb21baea),
	.w4(32'hbb31c432),
	.w5(32'hbbc28cd0),
	.w6(32'hbaa5a77c),
	.w7(32'hba589d08),
	.w8(32'hbbebc5ca),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf45a),
	.w1(32'h3b85921d),
	.w2(32'h3c4c608b),
	.w3(32'hbca0b270),
	.w4(32'hbab206f1),
	.w5(32'h3c48df88),
	.w6(32'hbbd9415d),
	.w7(32'h3b5e31b5),
	.w8(32'h3c3be80c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb140675),
	.w1(32'h3b626f16),
	.w2(32'h39ca5116),
	.w3(32'hbbc06a8c),
	.w4(32'hba935ffb),
	.w5(32'hbad5efab),
	.w6(32'hba218d2a),
	.w7(32'h3ba78273),
	.w8(32'h3c1a63ff),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a958d76),
	.w1(32'hbad4eaf2),
	.w2(32'h39e0680a),
	.w3(32'h3b2372d5),
	.w4(32'h3a0a8ce0),
	.w5(32'hba4b4512),
	.w6(32'h3c035b10),
	.w7(32'h3b3d52e3),
	.w8(32'hbac04ed1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15bf36),
	.w1(32'h38f0a716),
	.w2(32'h3b32c2ba),
	.w3(32'hbafe46cc),
	.w4(32'h3a5f91a4),
	.w5(32'h3b8672cd),
	.w6(32'hba27a38e),
	.w7(32'h3b040d66),
	.w8(32'h3c1f8fa7),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf0235),
	.w1(32'hb9868239),
	.w2(32'hbba41943),
	.w3(32'h3bdd2d1b),
	.w4(32'hb992450b),
	.w5(32'hbb1220f6),
	.w6(32'h3c2bad94),
	.w7(32'h3b2b61ea),
	.w8(32'hbaacf07b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11ca4a),
	.w1(32'h3acf3bc8),
	.w2(32'hbab8a8be),
	.w3(32'hbbc91188),
	.w4(32'h3ac3214c),
	.w5(32'hbb5892f2),
	.w6(32'hbacd7702),
	.w7(32'h3bc9f940),
	.w8(32'h3bc21893),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb532504),
	.w1(32'h3a386f38),
	.w2(32'h3ad99f40),
	.w3(32'hbb6f25b9),
	.w4(32'h3bd3c3c3),
	.w5(32'h3be04a9c),
	.w6(32'hba8b6671),
	.w7(32'h3c1c4d87),
	.w8(32'h3b9f6ffe),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba699fd),
	.w1(32'hba33ab05),
	.w2(32'hbb45a78f),
	.w3(32'h3b67155b),
	.w4(32'hbae5fde6),
	.w5(32'hbbf68fe0),
	.w6(32'hbaf84c22),
	.w7(32'hbb85eba5),
	.w8(32'hbbaf7dc3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc043349),
	.w1(32'h3a375eaf),
	.w2(32'hbbf7bd88),
	.w3(32'hbb9f34f4),
	.w4(32'hbbc3f6b0),
	.w5(32'hbc09a6ef),
	.w6(32'h3b6c931f),
	.w7(32'h3b910da5),
	.w8(32'hbbe265fb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeafd92),
	.w1(32'h3be45abf),
	.w2(32'hbb6e7a46),
	.w3(32'h3a64f583),
	.w4(32'h3c07a3d8),
	.w5(32'hbbf7c8da),
	.w6(32'hba03ee9c),
	.w7(32'h3c0b7ecd),
	.w8(32'hbb1473bc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385d9e00),
	.w1(32'hb9c6e581),
	.w2(32'hbc58b864),
	.w3(32'h3b837dd0),
	.w4(32'h3b0f6132),
	.w5(32'hbc03f101),
	.w6(32'h3bc6a2b9),
	.w7(32'h3b07242b),
	.w8(32'hbbfc6ff9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76cc84),
	.w1(32'hbaaeae38),
	.w2(32'hbc36b5be),
	.w3(32'hbc29957c),
	.w4(32'h3925bddf),
	.w5(32'hbc24b9df),
	.w6(32'hbbad0d6a),
	.w7(32'h3a595a43),
	.w8(32'hbba298c7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f410a),
	.w1(32'h39f36391),
	.w2(32'hbb4b1835),
	.w3(32'hbc1c070e),
	.w4(32'hbb2951c7),
	.w5(32'h390cc145),
	.w6(32'h3b060659),
	.w7(32'h3b68b0c5),
	.w8(32'h3b004d7e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db069),
	.w1(32'hbb40a6c0),
	.w2(32'h3b0cb2c9),
	.w3(32'hba99f89a),
	.w4(32'h3afbc2c1),
	.w5(32'hba2fe4ae),
	.w6(32'hbb020a63),
	.w7(32'h3af3e8bb),
	.w8(32'h3b1c21e0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d25f6),
	.w1(32'h3ba7af69),
	.w2(32'hbc39206b),
	.w3(32'hba11f747),
	.w4(32'h3a80270c),
	.w5(32'hbb1c6790),
	.w6(32'h3aabd9ce),
	.w7(32'h3b95b15b),
	.w8(32'h3bd02668),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda8332),
	.w1(32'hbcd568b2),
	.w2(32'h3ba4ee10),
	.w3(32'h3a4c0269),
	.w4(32'h3b840755),
	.w5(32'hbc83b9c2),
	.w6(32'h3c06c20a),
	.w7(32'h3c416481),
	.w8(32'hbbbbe990),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fe61a),
	.w1(32'h3c022ac9),
	.w2(32'h3b06d78b),
	.w3(32'hbbff048c),
	.w4(32'h3b9e49a9),
	.w5(32'h3af38fc0),
	.w6(32'hbb9d6d75),
	.w7(32'hbb03abda),
	.w8(32'hba2bb04e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54665e),
	.w1(32'hb96a2460),
	.w2(32'h3c0964b2),
	.w3(32'hba117702),
	.w4(32'hba16cd4f),
	.w5(32'hbb722e5a),
	.w6(32'hbbaa01f4),
	.w7(32'hbb27bfa4),
	.w8(32'hbc70356e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4a7db),
	.w1(32'h3bf4c4b8),
	.w2(32'h3c8bba8b),
	.w3(32'hbb87332a),
	.w4(32'hbc3c734c),
	.w5(32'h3cb1e693),
	.w6(32'hbc902e92),
	.w7(32'hbc80c089),
	.w8(32'hbc1c70dd),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c968a72),
	.w1(32'h3bafb70a),
	.w2(32'hbc006116),
	.w3(32'h3cdbd921),
	.w4(32'h3c28eefe),
	.w5(32'hbbc74e39),
	.w6(32'hbc724f40),
	.w7(32'hbc94d164),
	.w8(32'hbc102f43),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe25ac7),
	.w1(32'hbb9c9115),
	.w2(32'h3b9edfb2),
	.w3(32'h3aabee1e),
	.w4(32'h3a5d5b85),
	.w5(32'hbc0b667a),
	.w6(32'hbb33a5c1),
	.w7(32'hbacad90f),
	.w8(32'hbc253652),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36ca20),
	.w1(32'hbc01d32a),
	.w2(32'hba6c9a95),
	.w3(32'hbc16b195),
	.w4(32'hbaf16540),
	.w5(32'h3a88d312),
	.w6(32'hbaeb1f42),
	.w7(32'hb82116c5),
	.w8(32'hbaffc9e9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb498056),
	.w1(32'hbb8d05a5),
	.w2(32'h3b588a06),
	.w3(32'h3b570d96),
	.w4(32'h3b1e4d34),
	.w5(32'h3b8be8db),
	.w6(32'h3ae902c4),
	.w7(32'hb999b834),
	.w8(32'h3b2b3a74),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d70a7),
	.w1(32'hba0dcdee),
	.w2(32'hbc837f3c),
	.w3(32'h3b5b770a),
	.w4(32'hbb990034),
	.w5(32'hbbba7abd),
	.w6(32'hb9df0b28),
	.w7(32'hbc2f00ed),
	.w8(32'hbc3f0ea9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc742210),
	.w1(32'hbc352e59),
	.w2(32'hbc8fdab4),
	.w3(32'h3bbe461a),
	.w4(32'h3b1f061d),
	.w5(32'h3c0d957f),
	.w6(32'hbb95b753),
	.w7(32'hbb7a4848),
	.w8(32'h3bff06c4),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbc912),
	.w1(32'hbc834416),
	.w2(32'hbc83583b),
	.w3(32'h3c73e918),
	.w4(32'h3c5684b7),
	.w5(32'hbc80d993),
	.w6(32'h3c7bcef2),
	.w7(32'h3bf1682d),
	.w8(32'h3aa26166),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9afa9),
	.w1(32'h3b2b8227),
	.w2(32'h3a05a10b),
	.w3(32'hbc809977),
	.w4(32'hbb7cc619),
	.w5(32'hbb30dbec),
	.w6(32'h3b8e0f37),
	.w7(32'h384a9489),
	.w8(32'hb9a1ad7d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8e4f2),
	.w1(32'h3ba0a51d),
	.w2(32'hbc4db236),
	.w3(32'h3898fdd4),
	.w4(32'h3bdfb949),
	.w5(32'hbb930c25),
	.w6(32'h3a6adc7b),
	.w7(32'h3b7988a6),
	.w8(32'hbba7b8cc),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48b535),
	.w1(32'hbba62d1e),
	.w2(32'hbbdecc6d),
	.w3(32'h3bff6bfd),
	.w4(32'hbb1bb61a),
	.w5(32'hbc8f5cbd),
	.w6(32'h3ae9fab9),
	.w7(32'hbc271c8c),
	.w8(32'hbbe56d27),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e81d6),
	.w1(32'h3b1035f6),
	.w2(32'hbc02d8d7),
	.w3(32'hbceda328),
	.w4(32'hbc479fdd),
	.w5(32'h38963bb6),
	.w6(32'hbc117930),
	.w7(32'hbc3b29c7),
	.w8(32'h3b697382),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc279c59),
	.w1(32'hbc011cb7),
	.w2(32'hbc6a456e),
	.w3(32'h3bbc4360),
	.w4(32'h3b284942),
	.w5(32'hbc13039c),
	.w6(32'h3c0e3993),
	.w7(32'h3b6de620),
	.w8(32'hbc019ea6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2221aa),
	.w1(32'hbbca7e11),
	.w2(32'hbb6148a0),
	.w3(32'h3af5194c),
	.w4(32'hbbd2963c),
	.w5(32'hbb14f232),
	.w6(32'h3b91b811),
	.w7(32'h3b8fcdfd),
	.w8(32'hbc38a51b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce2495),
	.w1(32'h3b8f1e2f),
	.w2(32'hbab3e71d),
	.w3(32'h3a8aefef),
	.w4(32'h3b4dd797),
	.w5(32'h3b182bf0),
	.w6(32'h3b3be307),
	.w7(32'h3a71fe7b),
	.w8(32'h3b8e4d41),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb148370),
	.w1(32'hbb5f9df3),
	.w2(32'hbc78dbc3),
	.w3(32'hbb85b8b2),
	.w4(32'hbbb6af8c),
	.w5(32'hbbaebba8),
	.w6(32'hbb8948c9),
	.w7(32'hbaf858b3),
	.w8(32'hbb38aec2),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc483bc4),
	.w1(32'hbbdcc5a8),
	.w2(32'hbb14c3a8),
	.w3(32'h3b74cbee),
	.w4(32'h3ba11b3e),
	.w5(32'h37c4c20a),
	.w6(32'h3c0ea577),
	.w7(32'h3a99b7e4),
	.w8(32'h3a6bda4e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb151a69),
	.w1(32'hbb64a768),
	.w2(32'hbb2c7d06),
	.w3(32'h3a8807db),
	.w4(32'hba37b422),
	.w5(32'hbcb39420),
	.w6(32'h3ae0d4ff),
	.w7(32'hba61c7dc),
	.w8(32'h3b1026cd),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc094f7d),
	.w1(32'hbbc3ecd5),
	.w2(32'hbac35e8a),
	.w3(32'hbcccbedb),
	.w4(32'hbc31a936),
	.w5(32'hbb8cf032),
	.w6(32'h39dbf639),
	.w7(32'hbb21ca22),
	.w8(32'hbc470f93),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb986de1),
	.w1(32'hbb955510),
	.w2(32'h3c8a32e6),
	.w3(32'h39f486a1),
	.w4(32'hbb6e3124),
	.w5(32'h3c4510aa),
	.w6(32'hbc2923fc),
	.w7(32'hbb2acd44),
	.w8(32'hbb6d1a65),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89ea6d),
	.w1(32'h3adcb3c7),
	.w2(32'hbac13c65),
	.w3(32'hbba53123),
	.w4(32'hbc89ac63),
	.w5(32'hbc0af2a0),
	.w6(32'hbc278e9d),
	.w7(32'hbc0515fb),
	.w8(32'hbbe28cbe),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2463e0),
	.w1(32'hbc3bb031),
	.w2(32'h3cabb1b9),
	.w3(32'hbb7ef8f5),
	.w4(32'hbc0fc2b8),
	.w5(32'hb885582a),
	.w6(32'hbc661b61),
	.w7(32'hbbb37238),
	.w8(32'hbc8fb9bc),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05acbd),
	.w1(32'h3ca1deaf),
	.w2(32'h3cc30064),
	.w3(32'hbb719e0c),
	.w4(32'hbc342408),
	.w5(32'hbc9e1a9f),
	.w6(32'hbc92bbd7),
	.w7(32'hbc62bc31),
	.w8(32'hbc867dde),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccceaa5),
	.w1(32'h3c3c5826),
	.w2(32'h3c9c6ede),
	.w3(32'hbcb7c6fd),
	.w4(32'hbc488699),
	.w5(32'h3bc834ac),
	.w6(32'hbc58d1d2),
	.w7(32'hbb385a00),
	.w8(32'hbbba7f54),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d070fe2),
	.w1(32'h3cf4c853),
	.w2(32'h3c7fa3b0),
	.w3(32'h3bf23fda),
	.w4(32'h3b99b2a1),
	.w5(32'hbb6801e9),
	.w6(32'hbb89f4f6),
	.w7(32'h3b99bce4),
	.w8(32'hbb5238fa),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becee68),
	.w1(32'h3b4429fe),
	.w2(32'hbc6d4f3b),
	.w3(32'h3b16164e),
	.w4(32'h3a1ba18b),
	.w5(32'hbc69377e),
	.w6(32'hbac68033),
	.w7(32'hbb3caf4c),
	.w8(32'hbbc313c0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59771e),
	.w1(32'hbc5020f5),
	.w2(32'hbb893710),
	.w3(32'hbb2762af),
	.w4(32'h3bcddbff),
	.w5(32'hbb6cd755),
	.w6(32'hba1f1330),
	.w7(32'h3c2b41d6),
	.w8(32'hbb1032f9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae1b99),
	.w1(32'h3b54f3b6),
	.w2(32'hbba4e337),
	.w3(32'h3a5cb463),
	.w4(32'h3b443deb),
	.w5(32'hbc36caa7),
	.w6(32'hb9f619b2),
	.w7(32'h3b2d1a55),
	.w8(32'h3c0cc62b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80f72d),
	.w1(32'hbc4f22f7),
	.w2(32'hbce4f6df),
	.w3(32'hbc1773f6),
	.w4(32'hbc3cce7f),
	.w5(32'hbcba817d),
	.w6(32'h3ca506f4),
	.w7(32'h3b9c00ea),
	.w8(32'hbc21e5e9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb94714),
	.w1(32'hbc350d40),
	.w2(32'hbbf3b6c4),
	.w3(32'hbc37d7e4),
	.w4(32'hbb3c9ca4),
	.w5(32'h3bca27e8),
	.w6(32'h3b8a8cfa),
	.w7(32'h3c3ca6da),
	.w8(32'h3b562cce),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b874cd2),
	.w1(32'hbad1d272),
	.w2(32'hbbb25ed8),
	.w3(32'h3bd02f11),
	.w4(32'h3ba5aea2),
	.w5(32'h3b5a7c3d),
	.w6(32'h3ae294d5),
	.w7(32'hbaf5b065),
	.w8(32'hbbb3e530),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45783b),
	.w1(32'hb9c2e404),
	.w2(32'hbb5ae8eb),
	.w3(32'h3a47852c),
	.w4(32'hbb987db3),
	.w5(32'hbbc54cd4),
	.w6(32'hbbc4cffb),
	.w7(32'hbbb81338),
	.w8(32'h3c1ad2f7),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d59f4),
	.w1(32'hba6c1f55),
	.w2(32'hbb1a4bc4),
	.w3(32'hbb95d199),
	.w4(32'h3a67ded2),
	.w5(32'h3bdbdb07),
	.w6(32'h3bfef94d),
	.w7(32'h3c6048d3),
	.w8(32'hbbf2a3be),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c3d65),
	.w1(32'hbaa52293),
	.w2(32'h3c0970ad),
	.w3(32'h3ae92bfc),
	.w4(32'hbb6d6c8a),
	.w5(32'h3bdde36b),
	.w6(32'hbaf8be92),
	.w7(32'h3b272552),
	.w8(32'hbbd243db),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c725e6b),
	.w1(32'h3ba08aee),
	.w2(32'hbc64bf62),
	.w3(32'h3c34b34d),
	.w4(32'h3b6d16db),
	.w5(32'hbbd329fa),
	.w6(32'hbb053710),
	.w7(32'hbb92e75e),
	.w8(32'hbbdf38b4),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c82d9),
	.w1(32'hbc508928),
	.w2(32'h3a8ea0df),
	.w3(32'h3ba9957b),
	.w4(32'hbb2ca257),
	.w5(32'hbb7ffeaa),
	.w6(32'h3b22ace4),
	.w7(32'hbb1bc6e3),
	.w8(32'h3ae508cb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe29c0a),
	.w1(32'h3a97009e),
	.w2(32'hbb1636bb),
	.w3(32'hbbf9632f),
	.w4(32'hbb3e661c),
	.w5(32'hbba49074),
	.w6(32'hbc3f03f9),
	.w7(32'hbb2babd9),
	.w8(32'hb97ab442),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6bf3a),
	.w1(32'hbc1d9ece),
	.w2(32'hbb9cc90e),
	.w3(32'hbbed4ec6),
	.w4(32'h3b7ab125),
	.w5(32'hbb7563a7),
	.w6(32'hbb392812),
	.w7(32'hbc142747),
	.w8(32'hba89a5d8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1730ce),
	.w1(32'hbc0ce997),
	.w2(32'hbc26a9e7),
	.w3(32'hb9dd19cf),
	.w4(32'hbbceb99e),
	.w5(32'hbbd60e66),
	.w6(32'h3aa94a3d),
	.w7(32'hbbaf4927),
	.w8(32'hbc2497c0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd65f32),
	.w1(32'h3b4ec248),
	.w2(32'h3bf31547),
	.w3(32'hbbacb222),
	.w4(32'hba5bb07a),
	.w5(32'h39b314f1),
	.w6(32'hbb4a2f2d),
	.w7(32'hbb49d5ba),
	.w8(32'hbc013f42),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30ab5e),
	.w1(32'h3b8cb2e6),
	.w2(32'hbb70d3a9),
	.w3(32'hbaae0d13),
	.w4(32'h3b1e533c),
	.w5(32'h3a3baa53),
	.w6(32'hbbb504ac),
	.w7(32'hbb11f8a9),
	.w8(32'hba485baa),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94ae28),
	.w1(32'hbb8b92a7),
	.w2(32'hbc1ff1e0),
	.w3(32'hbb8a4351),
	.w4(32'hbb19be86),
	.w5(32'hbb4b779e),
	.w6(32'hbbe45e85),
	.w7(32'hbb7bb60d),
	.w8(32'h3c001c04),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35a210),
	.w1(32'hbc1daed6),
	.w2(32'h3ad3a245),
	.w3(32'h3957a4b4),
	.w4(32'h3b9088d9),
	.w5(32'h38fe6f78),
	.w6(32'h3c78818e),
	.w7(32'h3c98a8cd),
	.w8(32'hbb07eeb9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3883d),
	.w1(32'hbafef607),
	.w2(32'hbc17acad),
	.w3(32'h38c003cb),
	.w4(32'h39705acc),
	.w5(32'hbc567851),
	.w6(32'hbb16b8d5),
	.w7(32'hbba6390d),
	.w8(32'hbc149df2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc722f70),
	.w1(32'hbc14b09b),
	.w2(32'h3a516edb),
	.w3(32'hbc6206ff),
	.w4(32'hbb6079bf),
	.w5(32'hbb4e45d8),
	.w6(32'hbc067938),
	.w7(32'h3b897f54),
	.w8(32'hbaef7643),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef83ec),
	.w1(32'h38871296),
	.w2(32'h3ab41614),
	.w3(32'hbb114696),
	.w4(32'hbb498cb9),
	.w5(32'hba9d021f),
	.w6(32'hbb9b414c),
	.w7(32'hba9b3fe2),
	.w8(32'hbc6dcefe),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7b841),
	.w1(32'hbb461990),
	.w2(32'h3a3625e9),
	.w3(32'hbc3902a1),
	.w4(32'hbcb3fcd2),
	.w5(32'hbbd47360),
	.w6(32'hbc1969e3),
	.w7(32'h3abbf99b),
	.w8(32'hba0713cd),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f9df3),
	.w1(32'h3c362ee9),
	.w2(32'h3acd7b00),
	.w3(32'hbc2f2cb0),
	.w4(32'h3b5f8e5a),
	.w5(32'h3bdc2c6e),
	.w6(32'hbad191ae),
	.w7(32'h3b35b5e9),
	.w8(32'h3be2db80),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c9e58),
	.w1(32'hb97f3a54),
	.w2(32'hbb229f77),
	.w3(32'h3c0cb4ee),
	.w4(32'h3b944a7e),
	.w5(32'h3b42ca0f),
	.w6(32'h3abbaa89),
	.w7(32'h3b0b24db),
	.w8(32'hbb450fe9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dfe52),
	.w1(32'h3b8c2134),
	.w2(32'hbb9f16d1),
	.w3(32'h3be2440a),
	.w4(32'h3b8ceb11),
	.w5(32'h39998944),
	.w6(32'h3b64888d),
	.w7(32'hb9b7f969),
	.w8(32'h3b05d74f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9532f9),
	.w1(32'hbb6cfd0d),
	.w2(32'hbbd9810c),
	.w3(32'h3bcfc626),
	.w4(32'h3b7b85a6),
	.w5(32'hba03ccee),
	.w6(32'h3bbb5320),
	.w7(32'h3b8cf773),
	.w8(32'hb9bf2a64),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f6f36),
	.w1(32'hbc906f46),
	.w2(32'hbc20916c),
	.w3(32'h3910b0d5),
	.w4(32'h3ba15730),
	.w5(32'hb9915fde),
	.w6(32'h3b7b2e04),
	.w7(32'hb9cd95d8),
	.w8(32'hb8b7e297),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba48873),
	.w1(32'hbc286032),
	.w2(32'hbc3f0c67),
	.w3(32'hbc20f01d),
	.w4(32'hbc098b92),
	.w5(32'hbc251dc9),
	.w6(32'h3b1a2f03),
	.w7(32'hbb1cbfdd),
	.w8(32'hbc3d2424),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe2e6d),
	.w1(32'hbac7be9d),
	.w2(32'hbc850e76),
	.w3(32'hbb5720d7),
	.w4(32'hbbc75a00),
	.w5(32'hbc12fca0),
	.w6(32'hbc346e0f),
	.w7(32'hbc371108),
	.w8(32'hbb383a59),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9455e1),
	.w1(32'hbc6f6abe),
	.w2(32'h3b2a33ac),
	.w3(32'h3b7f62e6),
	.w4(32'h3c643f73),
	.w5(32'h3af8d1d3),
	.w6(32'h3c2319b3),
	.w7(32'h3c572da8),
	.w8(32'hb8e9843c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24b986),
	.w1(32'hbc17bd8f),
	.w2(32'hbc08379e),
	.w3(32'h3bc6ba45),
	.w4(32'hb987685e),
	.w5(32'hbbf7ae2d),
	.w6(32'h3b8fcd8e),
	.w7(32'h3bc166f0),
	.w8(32'hbba97940),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9effc7),
	.w1(32'hb9db1e6d),
	.w2(32'h3c0eb716),
	.w3(32'hbb24b58c),
	.w4(32'hbaac4c24),
	.w5(32'hbb481c99),
	.w6(32'hbb5f5e19),
	.w7(32'hbad5b91f),
	.w8(32'hbc225983),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1909de),
	.w1(32'h39fc36ad),
	.w2(32'hbc3a4762),
	.w3(32'hbb81dc1c),
	.w4(32'hbbf6cc44),
	.w5(32'h3adaa84c),
	.w6(32'hbb90f05c),
	.w7(32'hbc420314),
	.w8(32'hbcaba562),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fad12),
	.w1(32'h3c108d0e),
	.w2(32'h3c573f7e),
	.w3(32'h3c4a362b),
	.w4(32'h3c19b4fd),
	.w5(32'h3b78d7af),
	.w6(32'hbc492d11),
	.w7(32'hbbb2eb6c),
	.w8(32'hbc55c4e9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfccbbd),
	.w1(32'h3c2f0506),
	.w2(32'hbc18b923),
	.w3(32'h3cc10690),
	.w4(32'h3bf3af47),
	.w5(32'hbc1fddee),
	.w6(32'hbba05f0b),
	.w7(32'hbbddddcb),
	.w8(32'hbc518e4f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd97381),
	.w1(32'hbc2c85e7),
	.w2(32'h3a7b5c03),
	.w3(32'hbbac7039),
	.w4(32'h3ae8a20c),
	.w5(32'h3ad6edab),
	.w6(32'hbb99145c),
	.w7(32'hba859464),
	.w8(32'h3a69f2d4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c340506),
	.w1(32'h3c990ed7),
	.w2(32'h3ad24031),
	.w3(32'h3bd4d800),
	.w4(32'h3c8d6967),
	.w5(32'h3b972e4b),
	.w6(32'h3baa5457),
	.w7(32'h3c5e73ce),
	.w8(32'h3c1a8349),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd20b31),
	.w1(32'h3a9bb786),
	.w2(32'hbaee923c),
	.w3(32'hbba4b166),
	.w4(32'h3b06316c),
	.w5(32'h396a76ff),
	.w6(32'h3b1fa2bc),
	.w7(32'h3bd612e2),
	.w8(32'h3ac9a350),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb846926),
	.w1(32'hbb04f06e),
	.w2(32'hbb0cde25),
	.w3(32'hba408df0),
	.w4(32'hba5c205b),
	.w5(32'hba5c6aab),
	.w6(32'hbba86b6f),
	.w7(32'hbbcab4ff),
	.w8(32'hb9806d1f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30483b),
	.w1(32'h3bffe202),
	.w2(32'h3c130403),
	.w3(32'h3bbbfee2),
	.w4(32'h3bc59c4b),
	.w5(32'hbc15cedf),
	.w6(32'hbbfa5129),
	.w7(32'hbbbe5a70),
	.w8(32'hbc1a4bb7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb68a43),
	.w1(32'h3ac37d9c),
	.w2(32'h3b2f8d77),
	.w3(32'hbc21f35a),
	.w4(32'hbc5f40ae),
	.w5(32'h3b1608a6),
	.w6(32'hbc0a91e6),
	.w7(32'hbc1bde9c),
	.w8(32'hbbd0ead8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be36b74),
	.w1(32'h3b22af0e),
	.w2(32'h3c789b96),
	.w3(32'hbb20c5c9),
	.w4(32'h374a2976),
	.w5(32'hbb8a394a),
	.w6(32'hbc0e82c1),
	.w7(32'hbc026574),
	.w8(32'hbc9d6fa4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96e75b),
	.w1(32'h3b438b0f),
	.w2(32'hbc121175),
	.w3(32'hbc59d0aa),
	.w4(32'hbc60d6f5),
	.w5(32'h3b934206),
	.w6(32'hbc380655),
	.w7(32'hbc5f5cfe),
	.w8(32'h3b531b53),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdda8df),
	.w1(32'h39268576),
	.w2(32'hbc60e442),
	.w3(32'h3aca3fda),
	.w4(32'h3980efac),
	.w5(32'hbc93f02a),
	.w6(32'h39ab7ad2),
	.w7(32'hbb781e12),
	.w8(32'hbb3f9dbe),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9338c1),
	.w1(32'hbc255764),
	.w2(32'h3adc42c2),
	.w3(32'hbc6fd97c),
	.w4(32'hbc0fd58f),
	.w5(32'hbc053ca1),
	.w6(32'hbb03e8c6),
	.w7(32'hba105e4e),
	.w8(32'hbbf714d0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace5ad0),
	.w1(32'hbb8d4817),
	.w2(32'hbcc41114),
	.w3(32'hbc593328),
	.w4(32'hbb8e72f7),
	.w5(32'hbc012e52),
	.w6(32'hbc54aca2),
	.w7(32'hb9989e9b),
	.w8(32'hba055919),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3cd50),
	.w1(32'hbc75c6d3),
	.w2(32'h39f3ea3b),
	.w3(32'h3b82ef21),
	.w4(32'h3c0b0b04),
	.w5(32'hbba3111d),
	.w6(32'h3c1883ab),
	.w7(32'h3bfd8b72),
	.w8(32'hbc78517b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ceeaf),
	.w1(32'h3c0edac0),
	.w2(32'hbb87dc10),
	.w3(32'h3b98a2d9),
	.w4(32'hbb9bf98f),
	.w5(32'hbab7e268),
	.w6(32'hbba19709),
	.w7(32'hbbede9d3),
	.w8(32'h3b0a8675),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb869e0),
	.w1(32'hbc32b424),
	.w2(32'hba746980),
	.w3(32'h3bd13a09),
	.w4(32'h3a2e044a),
	.w5(32'hbba17653),
	.w6(32'hb993050c),
	.w7(32'hb6932ee5),
	.w8(32'hbba211f3),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc115196),
	.w1(32'hbc3c4074),
	.w2(32'hbb0c7741),
	.w3(32'h3b5475ea),
	.w4(32'h39838694),
	.w5(32'h3ad22913),
	.w6(32'h3bd04711),
	.w7(32'hbb2d99ba),
	.w8(32'hbb7f3ad5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248a41),
	.w1(32'hbc04fc0d),
	.w2(32'hbc83e128),
	.w3(32'h39824fda),
	.w4(32'hbb821e32),
	.w5(32'hbc5a3f34),
	.w6(32'hba8226b2),
	.w7(32'hbb56668e),
	.w8(32'h3b1a3f0e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9bd97),
	.w1(32'hbc5a7ecd),
	.w2(32'h3ad93b16),
	.w3(32'hbca73743),
	.w4(32'hbc97e2e5),
	.w5(32'hbae64ad0),
	.w6(32'hbaa329dd),
	.w7(32'hbc00c7d5),
	.w8(32'hbc057068),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b020293),
	.w1(32'h3b431e57),
	.w2(32'h3c4f3bec),
	.w3(32'hbc18b95c),
	.w4(32'hbbc17963),
	.w5(32'hbc5cf73b),
	.w6(32'hbc63a476),
	.w7(32'hbb7df06b),
	.w8(32'hbbbf35f9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79a691),
	.w1(32'h3a25879e),
	.w2(32'hbc29a60f),
	.w3(32'hbc8d02c6),
	.w4(32'hbc8db836),
	.w5(32'h3b94af2e),
	.w6(32'hbbb6624a),
	.w7(32'hbadf0a60),
	.w8(32'h3c209740),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d2b72),
	.w1(32'hbb12a15c),
	.w2(32'h3bf64929),
	.w3(32'hbb321111),
	.w4(32'h3af9be4a),
	.w5(32'h3c0958eb),
	.w6(32'hbb9f1b8e),
	.w7(32'hbb882597),
	.w8(32'h3c5bc480),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d1482),
	.w1(32'hbc46474d),
	.w2(32'h3a1d7b2a),
	.w3(32'h3c85daad),
	.w4(32'h3ba3b3f0),
	.w5(32'h3c2ea041),
	.w6(32'h3c9dd044),
	.w7(32'h3bd73b9e),
	.w8(32'hbbbf3e72),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72fe1b),
	.w1(32'h3bfee4cc),
	.w2(32'hbb8064e3),
	.w3(32'h3c0a0c57),
	.w4(32'hbbd6e2c2),
	.w5(32'hbcb9ea40),
	.w6(32'hbc45c17e),
	.w7(32'hbc7744a1),
	.w8(32'hbc165d7b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1f66d),
	.w1(32'hba0c7001),
	.w2(32'hbb83386a),
	.w3(32'hbcace324),
	.w4(32'hbca11fe8),
	.w5(32'hbbc4505f),
	.w6(32'hbc3a71e3),
	.w7(32'hbc6db283),
	.w8(32'hbaf8f8fb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb548833),
	.w1(32'hbb5f0224),
	.w2(32'hbc79ba7d),
	.w3(32'hbc9a92aa),
	.w4(32'hbcad8089),
	.w5(32'h3a837b02),
	.w6(32'h3b16db92),
	.w7(32'h3ae4861f),
	.w8(32'h3c52554e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6a16a),
	.w1(32'hbc1e1660),
	.w2(32'h3c73e3bc),
	.w3(32'hbbd0339c),
	.w4(32'hb9f2d92b),
	.w5(32'h3bc0f453),
	.w6(32'h3c0973fa),
	.w7(32'h3c328618),
	.w8(32'hbc17f4a6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3d88c),
	.w1(32'h3c1d64a3),
	.w2(32'hbc9bff46),
	.w3(32'h3bece97f),
	.w4(32'h3b706f4e),
	.w5(32'h3b8f3533),
	.w6(32'hbc3161db),
	.w7(32'hbbd269cd),
	.w8(32'h3bbb91b9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ce497),
	.w1(32'hbc8b8a72),
	.w2(32'h3c40cfac),
	.w3(32'h3abf8383),
	.w4(32'hb9f68e4c),
	.w5(32'hbb1f6407),
	.w6(32'h3bbf6257),
	.w7(32'h3a51c8e6),
	.w8(32'hbc09b784),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdd281),
	.w1(32'h3bd39fa2),
	.w2(32'hbc08714d),
	.w3(32'hbc2d47fb),
	.w4(32'hbc04c180),
	.w5(32'hbc04d59d),
	.w6(32'hbc5e895d),
	.w7(32'hbc2bbf25),
	.w8(32'hbc179a49),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48c3a0),
	.w1(32'hbc222d02),
	.w2(32'hbb8a6a03),
	.w3(32'hbc19859c),
	.w4(32'hb9c07192),
	.w5(32'hbb726c7c),
	.w6(32'h3a5f7a2b),
	.w7(32'hbbc8e19b),
	.w8(32'h3ab1084a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e6e4),
	.w1(32'hbbbb751e),
	.w2(32'h3b920be6),
	.w3(32'h3a449572),
	.w4(32'h3ac05f19),
	.w5(32'h3b55fb64),
	.w6(32'hbaa5b579),
	.w7(32'h3b969ec7),
	.w8(32'h3a5f4e54),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d1e0b),
	.w1(32'h3b2cf34a),
	.w2(32'h3b2e0517),
	.w3(32'h3adbbfba),
	.w4(32'h3b4315c9),
	.w5(32'hb8e6cd9d),
	.w6(32'hb9d8bd24),
	.w7(32'h39ffa1bb),
	.w8(32'hba9d7866),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c1a47),
	.w1(32'h3ba2a7a7),
	.w2(32'hbbda74bf),
	.w3(32'hba516b07),
	.w4(32'h3aa0227c),
	.w5(32'h3b697761),
	.w6(32'hbac708d4),
	.w7(32'h3a7290e5),
	.w8(32'hbae31b74),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bfd72),
	.w1(32'hbb8393c2),
	.w2(32'hbc33fadc),
	.w3(32'h3be1b377),
	.w4(32'h3c078cb5),
	.w5(32'hbb82c3ee),
	.w6(32'h3b38b971),
	.w7(32'h3b8a5a22),
	.w8(32'h3a119a1a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc510470),
	.w1(32'hbc3dc419),
	.w2(32'h3c8bfae2),
	.w3(32'hba7be15c),
	.w4(32'h3a3e3e66),
	.w5(32'h3c0d747b),
	.w6(32'h3b85bcf7),
	.w7(32'h3bc8674d),
	.w8(32'hbb89ed40),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30a532),
	.w1(32'hbc04a0c3),
	.w2(32'hbc5ac912),
	.w3(32'hbc29cd2b),
	.w4(32'hbc59550e),
	.w5(32'hbaac50fe),
	.w6(32'hbc7fea44),
	.w7(32'hbbf26a4b),
	.w8(32'h3b9196a1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb118e2d),
	.w1(32'hbb20f88a),
	.w2(32'hbaeb7b87),
	.w3(32'hbb3922a4),
	.w4(32'hb9dc0c43),
	.w5(32'hbbc398ca),
	.w6(32'hb9123988),
	.w7(32'hbb60ee9c),
	.w8(32'hbb5cb2e7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b3443),
	.w1(32'hba42ca10),
	.w2(32'h3bb4c524),
	.w3(32'hbbf61f26),
	.w4(32'h3b84ac71),
	.w5(32'hbaccb3be),
	.w6(32'hbc03fdf4),
	.w7(32'hbb95be44),
	.w8(32'hbc1c596e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule