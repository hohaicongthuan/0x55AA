module layer_8_featuremap_58(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8d1c),
	.w1(32'hb89c2fd4),
	.w2(32'hb994502f),
	.w3(32'h3a926498),
	.w4(32'h396318ac),
	.w5(32'hb8cc382a),
	.w6(32'h3a184369),
	.w7(32'h39c6e4b2),
	.w8(32'hba5378ab),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabab900),
	.w1(32'hb99d61ff),
	.w2(32'hb981c820),
	.w3(32'hba841ab1),
	.w4(32'h39cca982),
	.w5(32'h39913132),
	.w6(32'hba9ee9b0),
	.w7(32'hb93d6012),
	.w8(32'hb98c8c54),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8661c),
	.w1(32'hb8a88c01),
	.w2(32'hb9956d07),
	.w3(32'hbaa6b530),
	.w4(32'h39e18444),
	.w5(32'h3999e422),
	.w6(32'hbaa79347),
	.w7(32'h3911bae5),
	.w8(32'hba7c2801),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba022a3c),
	.w1(32'h3a772e72),
	.w2(32'hb965a991),
	.w3(32'h39ff0f3a),
	.w4(32'h3af00992),
	.w5(32'h3a998617),
	.w6(32'hb97de4de),
	.w7(32'hba8c0deb),
	.w8(32'h37f00bc9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d6a77),
	.w1(32'hba67e4e2),
	.w2(32'hba448cab),
	.w3(32'h370c7dcc),
	.w4(32'h39b1357e),
	.w5(32'hb89ac54c),
	.w6(32'hba30c100),
	.w7(32'hb93fff02),
	.w8(32'h3a11a0fd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa72810),
	.w1(32'hb9aebdbd),
	.w2(32'hb91ea339),
	.w3(32'hb9f2adf7),
	.w4(32'h3a14a06c),
	.w5(32'h39d49c68),
	.w6(32'hba107fff),
	.w7(32'h3a71b801),
	.w8(32'hbad2f3d2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed7f25),
	.w1(32'h3996121d),
	.w2(32'h39ca5f3c),
	.w3(32'h3947475b),
	.w4(32'h390a957e),
	.w5(32'h395fe7ce),
	.w6(32'hb8cb188f),
	.w7(32'h38ac3807),
	.w8(32'h39dc4850),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacb51f),
	.w1(32'hba858036),
	.w2(32'hba24a73a),
	.w3(32'hba432475),
	.w4(32'h3a490c97),
	.w5(32'h3a097082),
	.w6(32'hbad48609),
	.w7(32'hba374afb),
	.w8(32'hba86551f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c7895),
	.w1(32'hba85b943),
	.w2(32'hba6819f8),
	.w3(32'h39294f12),
	.w4(32'h39b111d8),
	.w5(32'hb8e27f94),
	.w6(32'hb9b0b04c),
	.w7(32'hb996f2e5),
	.w8(32'hbab7cca1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195f9a),
	.w1(32'h3a20ed1e),
	.w2(32'hba971ee1),
	.w3(32'h3aed04c7),
	.w4(32'h3b168595),
	.w5(32'h3b0acd13),
	.w6(32'hbabec3c5),
	.w7(32'hb979461c),
	.w8(32'hb9003d6c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c38be4),
	.w1(32'hba0dd974),
	.w2(32'hbad3c7bd),
	.w3(32'h3a37d7e1),
	.w4(32'hba061f19),
	.w5(32'hba9e8284),
	.w6(32'h39bc9201),
	.w7(32'hb9aa83cf),
	.w8(32'hba6273cc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399de236),
	.w1(32'h399816d7),
	.w2(32'hb6cb9ca6),
	.w3(32'h3a3f93a5),
	.w4(32'h3a3e198c),
	.w5(32'h39ab89ad),
	.w6(32'h37913dc6),
	.w7(32'h398e3c85),
	.w8(32'h38255d08),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a0a72),
	.w1(32'h389fd029),
	.w2(32'h3995892e),
	.w3(32'hba20e721),
	.w4(32'h3a44ea2b),
	.w5(32'h3a4ca0f6),
	.w6(32'hbac9870d),
	.w7(32'hb91ddd5c),
	.w8(32'h3ac66742),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5feade),
	.w1(32'h3a1c7c4f),
	.w2(32'h3ac109db),
	.w3(32'h3aaa79fe),
	.w4(32'h3a8180b2),
	.w5(32'h3ab7f924),
	.w6(32'h3adeabe3),
	.w7(32'h3b1c6a1d),
	.w8(32'h3a048bf6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a196cda),
	.w1(32'h39c07378),
	.w2(32'h3a3b6f89),
	.w3(32'h3a749a72),
	.w4(32'h3a553ce0),
	.w5(32'h3a51719b),
	.w6(32'h3a0fdb12),
	.w7(32'h3a444923),
	.w8(32'hb83b883c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd6296),
	.w1(32'hb92c35e2),
	.w2(32'h3710a242),
	.w3(32'hba0602b4),
	.w4(32'hb9bbab9a),
	.w5(32'hb7cf6fb8),
	.w6(32'hb94d08d2),
	.w7(32'hb92fcb3f),
	.w8(32'h39dd52f1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5d9f3),
	.w1(32'h3a93b43b),
	.w2(32'hba30058b),
	.w3(32'h39b4cd98),
	.w4(32'h3ac26263),
	.w5(32'hb8d8cee9),
	.w6(32'h3a8f3d4f),
	.w7(32'h3a01c032),
	.w8(32'hba31d37a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d84ce6),
	.w1(32'h3a351ff2),
	.w2(32'h3a65a2e6),
	.w3(32'h39176bf4),
	.w4(32'h3aa31578),
	.w5(32'h3ab9770d),
	.w6(32'hba2d34fe),
	.w7(32'h3a2957fd),
	.w8(32'h38b67717),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba196e8a),
	.w1(32'hbb4b3f10),
	.w2(32'hbbb6d4b2),
	.w3(32'hba49ba14),
	.w4(32'hbb2eaa41),
	.w5(32'hbb8ccb1b),
	.w6(32'hbadf6b07),
	.w7(32'hb9d47990),
	.w8(32'hbb7d4748),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb166035),
	.w1(32'hbb9737db),
	.w2(32'hbbece251),
	.w3(32'hbb0669cc),
	.w4(32'hbb25b884),
	.w5(32'hbb798ba4),
	.w6(32'hba6590e4),
	.w7(32'hba804d6e),
	.w8(32'hbb583b27),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fb175),
	.w1(32'hbaabe4c9),
	.w2(32'hbab4a08b),
	.w3(32'hba4f4a9a),
	.w4(32'hba76d2f9),
	.w5(32'hbad1e262),
	.w6(32'hba7617f6),
	.w7(32'hb9f51735),
	.w8(32'hba8061cb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8c460),
	.w1(32'h3a8bb9f0),
	.w2(32'h3a95deb8),
	.w3(32'h3a89fb97),
	.w4(32'h3afdfd46),
	.w5(32'h3b019f13),
	.w6(32'h3960a025),
	.w7(32'h3a9c4e2e),
	.w8(32'h3ac6904f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71c2101),
	.w1(32'hbb1a96b5),
	.w2(32'hbb34b9fa),
	.w3(32'hb9faabbb),
	.w4(32'hbb0bd624),
	.w5(32'hbb06bf5e),
	.w6(32'h3aa6e1e3),
	.w7(32'h3a1cfebb),
	.w8(32'hbb192b6d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30e399),
	.w1(32'hb92924ee),
	.w2(32'h3980c269),
	.w3(32'h3a99753b),
	.w4(32'h3a2fca8a),
	.w5(32'h3a7a993f),
	.w6(32'h399aedc1),
	.w7(32'h3a38212a),
	.w8(32'hbaec7d03),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e1f11),
	.w1(32'hbae60d37),
	.w2(32'hbb3e69ad),
	.w3(32'hbad3f997),
	.w4(32'hbb078a7f),
	.w5(32'hbb2ca212),
	.w6(32'hbafbc0c2),
	.w7(32'hbb1b9d3c),
	.w8(32'hba916360),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf9482),
	.w1(32'hbae29a28),
	.w2(32'hbab7c1d4),
	.w3(32'hba08ef79),
	.w4(32'hbaacbf79),
	.w5(32'hba4cc554),
	.w6(32'h3b140c5e),
	.w7(32'h3afab00d),
	.w8(32'h3905b361),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddb501),
	.w1(32'hba286764),
	.w2(32'h39852405),
	.w3(32'hba517e7e),
	.w4(32'hba489928),
	.w5(32'h396e5378),
	.w6(32'h3a4065d1),
	.w7(32'h3ac560f9),
	.w8(32'hb9c8c7d4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b86f3),
	.w1(32'hb9393ae5),
	.w2(32'hbb613fc6),
	.w3(32'h3b921a6a),
	.w4(32'hbac0db63),
	.w5(32'hbb0630fa),
	.w6(32'hbad4e9a1),
	.w7(32'hbbfa7043),
	.w8(32'hbc13c13c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9adf6e),
	.w1(32'hbb26aae5),
	.w2(32'hb9ff333c),
	.w3(32'hbb17c60c),
	.w4(32'hba9acef8),
	.w5(32'hba5842fd),
	.w6(32'h3a4a23cc),
	.w7(32'h3a856993),
	.w8(32'hba3ea5a4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c08658),
	.w1(32'hb8f66175),
	.w2(32'hb981790c),
	.w3(32'hb95a1c53),
	.w4(32'h393f544e),
	.w5(32'hb91b5ac8),
	.w6(32'hba443817),
	.w7(32'hb98b9f04),
	.w8(32'h3a0429b5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2badd9),
	.w1(32'h392d1bc6),
	.w2(32'hbb46bbcd),
	.w3(32'hb9a4ad73),
	.w4(32'h3aa79e54),
	.w5(32'hba5a453d),
	.w6(32'h39d31e76),
	.w7(32'hb9887841),
	.w8(32'hba8d9e38),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa71d26),
	.w1(32'hb9a8a09d),
	.w2(32'h39f9e9b2),
	.w3(32'hbab9e452),
	.w4(32'hba515b53),
	.w5(32'hb9fe8eb8),
	.w6(32'hba5140c9),
	.w7(32'h3999a2a6),
	.w8(32'h3aad1e4e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf79c7),
	.w1(32'h3b0fc2a3),
	.w2(32'h3a493ed1),
	.w3(32'h3aecde3d),
	.w4(32'h3b3a86fb),
	.w5(32'h3af7549c),
	.w6(32'h3b1120c1),
	.w7(32'h3a65b61d),
	.w8(32'h39abc318),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba364e96),
	.w1(32'hba281102),
	.w2(32'hbacb6257),
	.w3(32'hbaaeab3e),
	.w4(32'hbad9d17e),
	.w5(32'hba45405c),
	.w6(32'hb977c1cc),
	.w7(32'hb9456838),
	.w8(32'h3ab76f85),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905efff),
	.w1(32'h3a9b179e),
	.w2(32'h3a7814da),
	.w3(32'h39bea50e),
	.w4(32'h3acc4b9f),
	.w5(32'h3a38734c),
	.w6(32'hb903d484),
	.w7(32'h3b040807),
	.w8(32'hbacaa65d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb892f122),
	.w1(32'hba955b82),
	.w2(32'hba68f9f3),
	.w3(32'hb95ec5c2),
	.w4(32'hba843956),
	.w5(32'hba3237f9),
	.w6(32'hba1f120a),
	.w7(32'hb902ee4d),
	.w8(32'hbaf93786),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3f0d6),
	.w1(32'hba96d26e),
	.w2(32'hbacac33f),
	.w3(32'hba986d08),
	.w4(32'hbab2b60a),
	.w5(32'hbaa5b9e5),
	.w6(32'hba77ca15),
	.w7(32'hbad08f45),
	.w8(32'hb9ed11a6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5e325),
	.w1(32'hb9f54f96),
	.w2(32'h398d286f),
	.w3(32'hb9e78239),
	.w4(32'h3956a084),
	.w5(32'h3a465986),
	.w6(32'hba571a5c),
	.w7(32'hb8d4e314),
	.w8(32'h3ac83090),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60c289),
	.w1(32'h398ab4ad),
	.w2(32'h3a7cef38),
	.w3(32'h3ace5b6a),
	.w4(32'h3ab65d41),
	.w5(32'h3aa025f9),
	.w6(32'h3a0d9cb3),
	.w7(32'h3a796c0e),
	.w8(32'hb9d136bf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926f7df),
	.w1(32'h395327cb),
	.w2(32'h38143e74),
	.w3(32'hb9ea3b96),
	.w4(32'hb98e422b),
	.w5(32'hb9b014ed),
	.w6(32'hb8d89724),
	.w7(32'hb98ad178),
	.w8(32'h39b0b83c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb174c6e),
	.w1(32'hbac27aed),
	.w2(32'hba760961),
	.w3(32'hbb1b5322),
	.w4(32'hbadf264e),
	.w5(32'hba74bf27),
	.w6(32'hbb30e808),
	.w7(32'hbaae31f1),
	.w8(32'hbb1a3ddc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972ef4c),
	.w1(32'hb809b5f3),
	.w2(32'hba0c8a81),
	.w3(32'hb928e994),
	.w4(32'hb83c468d),
	.w5(32'hba06a279),
	.w6(32'hb9252a2a),
	.w7(32'hb911a887),
	.w8(32'hba1bc809),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9697239),
	.w1(32'hb91787cc),
	.w2(32'hb90087a9),
	.w3(32'hb98697ca),
	.w4(32'hb912862e),
	.w5(32'hb8f05037),
	.w6(32'hb96ab6c5),
	.w7(32'hb8f009cc),
	.w8(32'hb8fdd754),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ca234),
	.w1(32'hba074956),
	.w2(32'hba91d263),
	.w3(32'h38e70f3b),
	.w4(32'hb9a47650),
	.w5(32'hba43a2da),
	.w6(32'h384aa70d),
	.w7(32'hb9478cf4),
	.w8(32'hba46f75f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e580b2),
	.w1(32'hba99cf0b),
	.w2(32'hbb27a084),
	.w3(32'h3a67c1a2),
	.w4(32'hb8fe6780),
	.w5(32'hbab42432),
	.w6(32'h3a6e178f),
	.w7(32'h3a040bfe),
	.w8(32'hba88d225),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c8c19),
	.w1(32'h39d0b7a3),
	.w2(32'h39cfa7ed),
	.w3(32'hb80d5ed6),
	.w4(32'h39408874),
	.w5(32'h392e0398),
	.w6(32'hb8dd4364),
	.w7(32'h3947e42e),
	.w8(32'h385c9950),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376fbc1d),
	.w1(32'h3715363c),
	.w2(32'h3811e7dd),
	.w3(32'h36d0066a),
	.w4(32'h36153d92),
	.w5(32'h37be0530),
	.w6(32'h3772fcdc),
	.w7(32'h37188999),
	.w8(32'h38054ac8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8774e7a),
	.w1(32'hbab8b311),
	.w2(32'hbb269ce1),
	.w3(32'h39d6b926),
	.w4(32'hb9e4d0e5),
	.w5(32'hbac10b4c),
	.w6(32'h3a4e009e),
	.w7(32'h3999062e),
	.w8(32'hba73d42e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba435c05),
	.w1(32'hb90e0461),
	.w2(32'hba6caf7c),
	.w3(32'hb9aeef13),
	.w4(32'h39d4dbf0),
	.w5(32'hb9a5dfa1),
	.w6(32'hba27df90),
	.w7(32'h37bc8038),
	.w8(32'hba36b662),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391144af),
	.w1(32'h39d818f9),
	.w2(32'h38a7e07c),
	.w3(32'hb7bf335e),
	.w4(32'h393900d1),
	.w5(32'h38d50b78),
	.w6(32'hb80eb3f8),
	.w7(32'h391c442a),
	.w8(32'h37f451e5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac01a47),
	.w1(32'hb89d3cfe),
	.w2(32'h3a99939d),
	.w3(32'h3853769e),
	.w4(32'h3a90ef88),
	.w5(32'h3b068edc),
	.w6(32'hb8158438),
	.w7(32'h3a27b856),
	.w8(32'h3adb9295),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a7d9),
	.w1(32'hbb90d610),
	.w2(32'hbc05f0f4),
	.w3(32'hbb35912d),
	.w4(32'hbb554d21),
	.w5(32'hbbc9bc0e),
	.w6(32'hbb2df554),
	.w7(32'hbb30326e),
	.w8(32'hbbcadd34),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad039b5),
	.w1(32'hbb259988),
	.w2(32'hbb5f28e2),
	.w3(32'hb9c1b9bb),
	.w4(32'hba8bda2e),
	.w5(32'hbb04dc43),
	.w6(32'hb99f8f0e),
	.w7(32'hba635936),
	.w8(32'hbafe533a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab8531),
	.w1(32'h39e27e21),
	.w2(32'h3884a77e),
	.w3(32'h3a057624),
	.w4(32'h3a38ab58),
	.w5(32'h399a4569),
	.w6(32'h3780dfcc),
	.w7(32'h3a160a22),
	.w8(32'hb98d2cda),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381cdf91),
	.w1(32'h3603ee73),
	.w2(32'h3833d421),
	.w3(32'h379fb5e7),
	.w4(32'hb7913218),
	.w5(32'h37e44fd3),
	.w6(32'h3826cd5b),
	.w7(32'h36cddb61),
	.w8(32'h3858f1d9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c85f0a),
	.w1(32'hba568973),
	.w2(32'hbaad9c09),
	.w3(32'h395da3e5),
	.w4(32'hba8846d4),
	.w5(32'hba903a21),
	.w6(32'hb9c9eafb),
	.w7(32'hba440ff0),
	.w8(32'hba958873),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fbbc6),
	.w1(32'hb9e340e8),
	.w2(32'hba9a9355),
	.w3(32'hb9c2af26),
	.w4(32'hb92fa62a),
	.w5(32'hba6f9c81),
	.w6(32'hba206d8a),
	.w7(32'hb9b7809b),
	.w8(32'hbaa7ea66),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac64dc9),
	.w1(32'hbabe92da),
	.w2(32'hbafd414e),
	.w3(32'hbb076886),
	.w4(32'hba89da09),
	.w5(32'hbadaea75),
	.w6(32'hbaff1c6b),
	.w7(32'hba8be96d),
	.w8(32'hbae90af4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9388672),
	.w1(32'hb9fb1a8d),
	.w2(32'hba7f3240),
	.w3(32'hb91dd01f),
	.w4(32'hba30992c),
	.w5(32'hba9ac727),
	.w6(32'hba2ac5c5),
	.w7(32'hba350022),
	.w8(32'hba8f72ae),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd0eb8),
	.w1(32'hb9fc30ec),
	.w2(32'hba030220),
	.w3(32'hba27b325),
	.w4(32'hba0c63f0),
	.w5(32'hb9fa1baf),
	.w6(32'hba5e9908),
	.w7(32'hba1a168a),
	.w8(32'hba1d97d4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1166ac),
	.w1(32'hba388e70),
	.w2(32'hba2a0269),
	.w3(32'hba242bd1),
	.w4(32'hba20dad1),
	.w5(32'hba189ce9),
	.w6(32'hba27a26e),
	.w7(32'hba2f6d58),
	.w8(32'hba08d818),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38683058),
	.w1(32'h37c751be),
	.w2(32'hb7fb9fc8),
	.w3(32'h385e778c),
	.w4(32'h3708aa29),
	.w5(32'hb78fa284),
	.w6(32'h37402585),
	.w7(32'h370cb0a1),
	.w8(32'hb715c986),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba462c94),
	.w1(32'hba3a61c0),
	.w2(32'hbaeb9853),
	.w3(32'h3a077ead),
	.w4(32'h3a3ce22a),
	.w5(32'hb9db748d),
	.w6(32'hb9815985),
	.w7(32'hb93816b7),
	.w8(32'hbabd8890),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a4aa1),
	.w1(32'hb8d58a22),
	.w2(32'hba4ecaa6),
	.w3(32'hba1469f4),
	.w4(32'h39f4f090),
	.w5(32'h37cbbe89),
	.w6(32'hb9d25744),
	.w7(32'h39dd6623),
	.w8(32'hb9978c41),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05a2d9),
	.w1(32'h39bbe9df),
	.w2(32'hb935ebb0),
	.w3(32'h3a7fd4d4),
	.w4(32'h3a728ce3),
	.w5(32'h39fa6fee),
	.w6(32'h3a61c56d),
	.w7(32'h3a2bc83e),
	.w8(32'h399521f3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba361019),
	.w1(32'hba552209),
	.w2(32'hba75110d),
	.w3(32'hba6833ff),
	.w4(32'hba87cea1),
	.w5(32'hba8991f6),
	.w6(32'hba670ff3),
	.w7(32'hba833202),
	.w8(32'hba99b3ac),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabf880),
	.w1(32'hb9c81065),
	.w2(32'hba7619b8),
	.w3(32'hba4a3655),
	.w4(32'h3a1e467c),
	.w5(32'h389bb3aa),
	.w6(32'hba38c973),
	.w7(32'h3929ccda),
	.w8(32'hb98f31e7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf709c),
	.w1(32'hba0bf4b8),
	.w2(32'hba897136),
	.w3(32'hba0545c3),
	.w4(32'hba376085),
	.w5(32'hba8e5a5a),
	.w6(32'hba87e6fd),
	.w7(32'hba64dec0),
	.w8(32'hbaa6c954),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5b01d),
	.w1(32'hb9d548dc),
	.w2(32'hb9d0f8bf),
	.w3(32'hb9770d25),
	.w4(32'hb9640468),
	.w5(32'hb9672bf8),
	.w6(32'hb962facc),
	.w7(32'hb917d5a0),
	.w8(32'hb90540be),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25267c),
	.w1(32'hbaf866d0),
	.w2(32'hbb7adcfe),
	.w3(32'h39f3f94c),
	.w4(32'hbad821ae),
	.w5(32'hbb53e8bd),
	.w6(32'h3a8d3a4b),
	.w7(32'hb8f75d20),
	.w8(32'hbb104cf9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387c687a),
	.w1(32'h389a925f),
	.w2(32'h38bd551f),
	.w3(32'h38b5b0e9),
	.w4(32'h38f326c4),
	.w5(32'h3907cb28),
	.w6(32'h38acb232),
	.w7(32'h38e5504a),
	.w8(32'h390e3e78),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35fa40),
	.w1(32'hba38ffa2),
	.w2(32'hbaeba7e8),
	.w3(32'h38b9d13a),
	.w4(32'h391083ee),
	.w5(32'hbaabf2e2),
	.w6(32'hb9c3b36d),
	.w7(32'hb97a301b),
	.w8(32'hbacd6ea6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37895eba),
	.w1(32'hb861a170),
	.w2(32'hb7870f97),
	.w3(32'hb84708d0),
	.w4(32'hb8913381),
	.w5(32'h37f35575),
	.w6(32'hb87f8043),
	.w7(32'hb85756f7),
	.w8(32'h3622d2d2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba928878),
	.w1(32'hb9a87292),
	.w2(32'hba18f8c7),
	.w3(32'hba5cd6fd),
	.w4(32'hb9410814),
	.w5(32'hb90e1daa),
	.w6(32'hbaaab60c),
	.w7(32'hba8a6e5c),
	.w8(32'hba78f349),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371ed029),
	.w1(32'h36fec7a6),
	.w2(32'h376d095e),
	.w3(32'h36f27e02),
	.w4(32'h369da6e7),
	.w5(32'h370cbc76),
	.w6(32'h37270380),
	.w7(32'h36ac362c),
	.w8(32'h37386815),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad67c9a),
	.w1(32'hbac5b922),
	.w2(32'hbb2d8fc5),
	.w3(32'hbad4bda3),
	.w4(32'hbaa4b9ba),
	.w5(32'hbb1e5c92),
	.w6(32'hbaff2998),
	.w7(32'hbac1e984),
	.w8(32'hbb2dda73),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb805988c),
	.w1(32'hb84957f4),
	.w2(32'hb8811a19),
	.w3(32'hb87d7b9a),
	.w4(32'hb86532f0),
	.w5(32'hb875af1c),
	.w6(32'hb813c797),
	.w7(32'hb82ac398),
	.w8(32'hb82e9fe6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9654ed2),
	.w1(32'hba964f7d),
	.w2(32'hbb10a1cd),
	.w3(32'h3a06b417),
	.w4(32'hb9e903cb),
	.w5(32'hbabb0ff0),
	.w6(32'h398fd53a),
	.w7(32'hb911638f),
	.w8(32'hbab7e8ac),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90131d0),
	.w1(32'hb9efc37f),
	.w2(32'hba291dc7),
	.w3(32'hb9c1466c),
	.w4(32'hb9eaaadf),
	.w5(32'hb9bb2608),
	.w6(32'hb98e7d40),
	.w7(32'hba4db8c2),
	.w8(32'hba37ae74),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d69cee),
	.w1(32'hb981fd2c),
	.w2(32'hb9ef8695),
	.w3(32'hb9145b35),
	.w4(32'hb97fe04c),
	.w5(32'hb9db5725),
	.w6(32'hb9582600),
	.w7(32'hb95f3872),
	.w8(32'hb9e7fbf8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc9d6f),
	.w1(32'h3765a4ea),
	.w2(32'h38396ee6),
	.w3(32'h3774d742),
	.w4(32'h371d9a85),
	.w5(32'h384dc219),
	.w6(32'h37aedb0d),
	.w7(32'h37f31c6a),
	.w8(32'h388063ab),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba806d37),
	.w1(32'hba13e828),
	.w2(32'hba72e662),
	.w3(32'hb9ffebea),
	.w4(32'hb991699c),
	.w5(32'hba1a9581),
	.w6(32'hb9f723ac),
	.w7(32'hb99d51ce),
	.w8(32'hba312844),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3859710f),
	.w1(32'hba4c1463),
	.w2(32'hbac5a036),
	.w3(32'h3a7664bc),
	.w4(32'h3882e9eb),
	.w5(32'hba37c034),
	.w6(32'h3a82efb0),
	.w7(32'h398a2f63),
	.w8(32'hba7f414e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6f327),
	.w1(32'hba9c559c),
	.w2(32'hbb4a5917),
	.w3(32'hbb0457c9),
	.w4(32'hb977d115),
	.w5(32'hbb13da51),
	.w6(32'hbb201099),
	.w7(32'hbaa449cb),
	.w8(32'hbb8244f5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a3bb9),
	.w1(32'hbb0414a1),
	.w2(32'hbb8431cf),
	.w3(32'h3a6b5d73),
	.w4(32'hb937b8f8),
	.w5(32'hbb193326),
	.w6(32'h3a998caf),
	.w7(32'h388bd8fc),
	.w8(32'hbb01ef7f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c84d4),
	.w1(32'hbb0e53f1),
	.w2(32'hbb40d1d9),
	.w3(32'hb9c0fc4f),
	.w4(32'hba859a83),
	.w5(32'hbafb73cc),
	.w6(32'h3923a5da),
	.w7(32'hbabe14c8),
	.w8(32'hbad818fc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39056b96),
	.w1(32'h38ba9f45),
	.w2(32'h398962a9),
	.w3(32'h388043f7),
	.w4(32'hb6ff48e9),
	.w5(32'h394c0942),
	.w6(32'h388124ce),
	.w7(32'h3875eceb),
	.w8(32'h3967d645),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ef5c7a),
	.w1(32'h3755d456),
	.w2(32'h384e4a1e),
	.w3(32'h3727f1ca),
	.w4(32'hb6e203e8),
	.w5(32'h37fd0516),
	.w6(32'h379f72a2),
	.w7(32'h36bd04e7),
	.w8(32'h383067b1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902cdec),
	.w1(32'h38c56e4a),
	.w2(32'h389bb679),
	.w3(32'h390914ff),
	.w4(32'h38a353e6),
	.w5(32'h37828926),
	.w6(32'h38946d61),
	.w7(32'h381ab80b),
	.w8(32'hb6d01e88),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d578ac),
	.w1(32'hba056805),
	.w2(32'hba4a720f),
	.w3(32'h3a23dfca),
	.w4(32'h3985bd98),
	.w5(32'hb96749aa),
	.w6(32'h39d2a29c),
	.w7(32'hb72d1017),
	.w8(32'hb9bffc9c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04ed4e),
	.w1(32'hb9199c2a),
	.w2(32'hb98ce06f),
	.w3(32'hb99f57a2),
	.w4(32'hb90f6d37),
	.w5(32'hb9bc4dfa),
	.w6(32'hba093b9e),
	.w7(32'hb9bce8e4),
	.w8(32'hba138963),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915ea8e),
	.w1(32'h39e558ff),
	.w2(32'hb9798d85),
	.w3(32'h39c51439),
	.w4(32'h3a14c0ae),
	.w5(32'hb867cf0f),
	.w6(32'h39a3c5cf),
	.w7(32'h39e8a149),
	.w8(32'hb92ac128),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38c680),
	.w1(32'h39ab46dc),
	.w2(32'hba3647c2),
	.w3(32'hb71e01d7),
	.w4(32'h3a90d90c),
	.w5(32'hb8c4b457),
	.w6(32'hba17758c),
	.w7(32'h39bde3ab),
	.w8(32'hba3741b3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98168bc),
	.w1(32'hb9138a2c),
	.w2(32'hba96dccb),
	.w3(32'h3a4eca2c),
	.w4(32'h3a8f3cd5),
	.w5(32'hb5ebb8d0),
	.w6(32'h395f2001),
	.w7(32'h39a4b201),
	.w8(32'hba47f2ef),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1e5a2),
	.w1(32'h3a0a5a5b),
	.w2(32'h39c43e7c),
	.w3(32'h3a0bb11d),
	.w4(32'h3a02d47e),
	.w5(32'h39c5c36d),
	.w6(32'h39957569),
	.w7(32'h39bee4b7),
	.w8(32'hb71deaa9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968df4c),
	.w1(32'h3839ec67),
	.w2(32'hba90e516),
	.w3(32'h3a6047ba),
	.w4(32'h3a1d10c9),
	.w5(32'hba0dfa1b),
	.w6(32'h3a0428db),
	.w7(32'h39f57665),
	.w8(32'hba87d9fc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03dc98),
	.w1(32'hbb2ff10f),
	.w2(32'hbb7db612),
	.w3(32'hb9573d85),
	.w4(32'hb9e16851),
	.w5(32'hbb053cee),
	.w6(32'hba2eee5c),
	.w7(32'hba699df4),
	.w8(32'hbb23e528),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37da253a),
	.w1(32'h3780b3d5),
	.w2(32'h387f77ae),
	.w3(32'h378afd04),
	.w4(32'h369c8b1f),
	.w5(32'h38501813),
	.w6(32'h37f4b651),
	.w7(32'h378a8238),
	.w8(32'h386d652a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907dc40),
	.w1(32'h38aea57e),
	.w2(32'h39789a0d),
	.w3(32'h38900243),
	.w4(32'h3751a59b),
	.w5(32'h39320695),
	.w6(32'h38ea5c98),
	.w7(32'h38845419),
	.w8(32'h3968fe49),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38798ba2),
	.w1(32'h3822f716),
	.w2(32'h390033a0),
	.w3(32'h37d62f41),
	.w4(32'hb4863280),
	.w5(32'h38b5fed2),
	.w6(32'h385ceeab),
	.w7(32'h37f45a1e),
	.w8(32'h38f5ab26),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379e7ff4),
	.w1(32'h37559e86),
	.w2(32'hb9001cfa),
	.w3(32'h38508d55),
	.w4(32'h381cf046),
	.w5(32'hb8a5dafa),
	.w6(32'hb74a9803),
	.w7(32'h360baac3),
	.w8(32'hb8df294e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9685bb6),
	.w1(32'h38fabc39),
	.w2(32'hb89242e8),
	.w3(32'h399c4318),
	.w4(32'h3998c527),
	.w5(32'h39af76d4),
	.w6(32'h39996e23),
	.w7(32'h3971cf12),
	.w8(32'hb9180f2f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e331b),
	.w1(32'hb9d7c8f0),
	.w2(32'hba469b2a),
	.w3(32'hb9dedb6f),
	.w4(32'hb7e090d6),
	.w5(32'hba0a4f7b),
	.w6(32'hba544016),
	.w7(32'hba03f775),
	.w8(32'hba57c427),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9deb0c),
	.w1(32'hb9654f9e),
	.w2(32'hba5e9518),
	.w3(32'hba7f6ae4),
	.w4(32'h3935b9af),
	.w5(32'hb9cb6bfb),
	.w6(32'hba93c735),
	.w7(32'hb9778274),
	.w8(32'hba3fe6ab),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c594c2),
	.w1(32'h39235ce8),
	.w2(32'hba060274),
	.w3(32'hb9b589f1),
	.w4(32'h399f0b77),
	.w5(32'hb9d0af46),
	.w6(32'hba102588),
	.w7(32'hb7cf651a),
	.w8(32'hbc0ed3d6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f2801),
	.w1(32'hbbdffd26),
	.w2(32'hbc21a3f5),
	.w3(32'h3b045390),
	.w4(32'h3aae034b),
	.w5(32'h39c77445),
	.w6(32'hbb0f9fc7),
	.w7(32'h3a423cc2),
	.w8(32'h3b244c63),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71db84),
	.w1(32'h3bd88d58),
	.w2(32'h3b883cf1),
	.w3(32'h3c006639),
	.w4(32'hbc1bd153),
	.w5(32'hbcc9e542),
	.w6(32'hba4a2ac3),
	.w7(32'h3c733f3f),
	.w8(32'hbc011a38),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d2157),
	.w1(32'hbb944efa),
	.w2(32'hbb9a54a1),
	.w3(32'hbaaeb379),
	.w4(32'hbbd48a61),
	.w5(32'hb8d170da),
	.w6(32'h3b013296),
	.w7(32'h3abb7542),
	.w8(32'hbae124f1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b316b19),
	.w1(32'hbb4a30a0),
	.w2(32'hbb5fd4b7),
	.w3(32'h3b1d5720),
	.w4(32'hbba5a9e8),
	.w5(32'hbb693cbd),
	.w6(32'h3b2a84b6),
	.w7(32'h3b6d4793),
	.w8(32'hbc437212),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb661082),
	.w1(32'hbbd6d944),
	.w2(32'hbc42a119),
	.w3(32'h3b84fc63),
	.w4(32'hbb875b13),
	.w5(32'hbb4c1c71),
	.w6(32'hbc3b4546),
	.w7(32'hbbe088fa),
	.w8(32'hbcc27f9a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd434d21),
	.w1(32'h3c0b0a37),
	.w2(32'hbd7ceca5),
	.w3(32'hbd005311),
	.w4(32'hbd177670),
	.w5(32'hbc80fb46),
	.w6(32'hbd13a216),
	.w7(32'hbd2f8353),
	.w8(32'h3c65cdf8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c274ce7),
	.w1(32'hbb6ece65),
	.w2(32'hbc46f4b4),
	.w3(32'hbbc432af),
	.w4(32'hbc2c3638),
	.w5(32'hbc113c69),
	.w6(32'h3c38f9bb),
	.w7(32'hbc195300),
	.w8(32'hbc0a7679),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc742ece),
	.w1(32'hbbe8948a),
	.w2(32'h3c0c3fec),
	.w3(32'h3c2c64ee),
	.w4(32'h3ca354d9),
	.w5(32'h3c3f70d6),
	.w6(32'hbc947c2d),
	.w7(32'h3ba1f916),
	.w8(32'hbb942de7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac94087),
	.w1(32'hbb6f064e),
	.w2(32'hbbd17236),
	.w3(32'h38e371f9),
	.w4(32'hbb93d78a),
	.w5(32'hbbcdd1fb),
	.w6(32'hba8b7e71),
	.w7(32'hba8619d2),
	.w8(32'h39a4d25c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd162a7),
	.w1(32'h3aee4b30),
	.w2(32'h3ac4309f),
	.w3(32'h3b46f2b8),
	.w4(32'hba9aff93),
	.w5(32'h3a9d2991),
	.w6(32'h3b8c3aca),
	.w7(32'h3b482255),
	.w8(32'hbb081ed2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c102c8f),
	.w1(32'hbb031876),
	.w2(32'hb96235a0),
	.w3(32'h3b69d4e8),
	.w4(32'hbb94cca4),
	.w5(32'h3bd928b9),
	.w6(32'h3bd60cc2),
	.w7(32'h3badfb1f),
	.w8(32'h3c924e85),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17744a),
	.w1(32'hbc50f6f7),
	.w2(32'h3c695de5),
	.w3(32'hbc3b7838),
	.w4(32'hbc831dd4),
	.w5(32'h3cccea46),
	.w6(32'hbcec395f),
	.w7(32'hbc7839d1),
	.w8(32'hbc4d5145),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd113c),
	.w1(32'hbbfad70a),
	.w2(32'hba19a5b4),
	.w3(32'h3c511759),
	.w4(32'h3c5cddfe),
	.w5(32'h3ae9afb8),
	.w6(32'hbc7be745),
	.w7(32'hbaa6b02f),
	.w8(32'hbc82bc7e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fe961),
	.w1(32'h3cb20736),
	.w2(32'hbbbd4c98),
	.w3(32'hbc5f1298),
	.w4(32'hbd0dda86),
	.w5(32'hbbb2c1c4),
	.w6(32'hbc9214c5),
	.w7(32'h3b3891f4),
	.w8(32'hbba1edb4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23d1cc),
	.w1(32'hbac04542),
	.w2(32'hba3385e8),
	.w3(32'hbc2d2f66),
	.w4(32'h3b62854c),
	.w5(32'h3bf22714),
	.w6(32'hbcb730d8),
	.w7(32'hbc0aec30),
	.w8(32'hbc175c19),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc592c32),
	.w1(32'h3b2c16a1),
	.w2(32'hbc14392d),
	.w3(32'hbc6def02),
	.w4(32'hbc726ef2),
	.w5(32'hbbddf406),
	.w6(32'hbc89d7bf),
	.w7(32'hbc551800),
	.w8(32'h3c84a5bb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6be27),
	.w1(32'h3bf7cdc8),
	.w2(32'hbc80a9e9),
	.w3(32'hbb8f6fd0),
	.w4(32'h3cc097d6),
	.w5(32'hbb988c6d),
	.w6(32'h3ce6bd7f),
	.w7(32'hbbaab9c4),
	.w8(32'h3b8f8914),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2458b),
	.w1(32'hbc5750c8),
	.w2(32'hbbf6ac2d),
	.w3(32'h3bbede74),
	.w4(32'hbb38230a),
	.w5(32'h3b960165),
	.w6(32'h3a747fea),
	.w7(32'h3b0c80cc),
	.w8(32'hbacfaeb0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ba341),
	.w1(32'h3c0b9806),
	.w2(32'hbbb7cfe9),
	.w3(32'hbc3074ea),
	.w4(32'hbbc06ddb),
	.w5(32'hbc421784),
	.w6(32'h3a0cbaa8),
	.w7(32'hbb672d04),
	.w8(32'h3bba045e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05f66b),
	.w1(32'h3b9f8804),
	.w2(32'hbcc584a1),
	.w3(32'hbd03bafd),
	.w4(32'hbca02899),
	.w5(32'hbd100fde),
	.w6(32'hbcff7bf5),
	.w7(32'hbce0f212),
	.w8(32'hbac991e8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3de64),
	.w1(32'hbbf6fab8),
	.w2(32'hbc66ab20),
	.w3(32'hb9176b85),
	.w4(32'hbb222bdd),
	.w5(32'h3b82150e),
	.w6(32'hbc1dac58),
	.w7(32'hbc0c204b),
	.w8(32'h3b1946f1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03d4a7),
	.w1(32'hbbeedb07),
	.w2(32'hbc1061da),
	.w3(32'h3bf5c3bc),
	.w4(32'hbb9c9943),
	.w5(32'hbc4c1b5d),
	.w6(32'h3b605b05),
	.w7(32'h3b39a40a),
	.w8(32'hbc2a57a2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69f0a9),
	.w1(32'hbc3148dd),
	.w2(32'hba8bde80),
	.w3(32'hbb5ddbec),
	.w4(32'h3c6c4302),
	.w5(32'h3c52853f),
	.w6(32'h3d171fa0),
	.w7(32'hba39ced4),
	.w8(32'hbc0f1892),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule