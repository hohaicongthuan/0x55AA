module layer_8_featuremap_4(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0540af),
	.w1(32'h3afad4d4),
	.w2(32'h3c5191fc),
	.w3(32'h39f2b9fa),
	.w4(32'h3bca728e),
	.w5(32'h3c8e2f8f),
	.w6(32'hbb92bb75),
	.w7(32'h3b0800ff),
	.w8(32'h3be8d33a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac234f),
	.w1(32'h3b87a162),
	.w2(32'h3bff6677),
	.w3(32'h3c3efe98),
	.w4(32'h3ba45151),
	.w5(32'h3c252c86),
	.w6(32'h3b8f4ed7),
	.w7(32'hbace6388),
	.w8(32'hbabd442b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf55772),
	.w1(32'h3bde777c),
	.w2(32'h3c444e61),
	.w3(32'h3bc53454),
	.w4(32'h3c11caa9),
	.w5(32'h3c5b3cd4),
	.w6(32'hbba88aa4),
	.w7(32'h3b9022b3),
	.w8(32'h3baf0856),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37f3aa),
	.w1(32'h3c2615fb),
	.w2(32'h3c954f1c),
	.w3(32'h3c448d00),
	.w4(32'h3c1a8e4c),
	.w5(32'h3c8fddc9),
	.w6(32'h3b7a731b),
	.w7(32'hba1ebcea),
	.w8(32'h3b6a5e9b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86e1df),
	.w1(32'hbad80fb8),
	.w2(32'h3be9807d),
	.w3(32'h3c741e09),
	.w4(32'h3c1c7656),
	.w5(32'h3c9af79d),
	.w6(32'h3ab6b1ae),
	.w7(32'hbad31174),
	.w8(32'h3af78f71),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b845482),
	.w1(32'hbb99022f),
	.w2(32'h3a66c0b6),
	.w3(32'h3c84c07f),
	.w4(32'hbb0396bf),
	.w5(32'hbb975fdb),
	.w6(32'h3b0cdfcd),
	.w7(32'h3c1eaef5),
	.w8(32'h3bce89c5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9f9cb),
	.w1(32'hbbb3c34c),
	.w2(32'hbb730b33),
	.w3(32'hbb320d49),
	.w4(32'hbc31a837),
	.w5(32'hbc0ca4a7),
	.w6(32'h3b5bedb1),
	.w7(32'hbc43ca7e),
	.w8(32'hbc3ac91e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf22efb),
	.w1(32'hbb108875),
	.w2(32'h3a1fe764),
	.w3(32'hbb9d0317),
	.w4(32'h3b9941e8),
	.w5(32'h3c130be8),
	.w6(32'hbc0085ec),
	.w7(32'h3bdcad56),
	.w8(32'h3c59eab2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be11cc3),
	.w1(32'hbbb8b1f3),
	.w2(32'hbbd3cc33),
	.w3(32'h3a400c50),
	.w4(32'hbb673eeb),
	.w5(32'hbb94876a),
	.w6(32'h3c063d04),
	.w7(32'hb98ab03c),
	.w8(32'hba4d7130),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96cc01),
	.w1(32'hbbc5813f),
	.w2(32'h3b89762a),
	.w3(32'hbb6aab82),
	.w4(32'hbc26727a),
	.w5(32'hb822bb43),
	.w6(32'h3a44200e),
	.w7(32'h3bcb500c),
	.w8(32'h3bdf9a25),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b036),
	.w1(32'hb883d94b),
	.w2(32'hbb2007f1),
	.w3(32'h3ba2ce2b),
	.w4(32'hbaf3c834),
	.w5(32'hbb323bcc),
	.w6(32'h3bc3efed),
	.w7(32'hbaab9a06),
	.w8(32'h39047b65),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16cca),
	.w1(32'h39c304b9),
	.w2(32'h3b329b7d),
	.w3(32'hbbe26238),
	.w4(32'h39eab1f7),
	.w5(32'hb99ceb5d),
	.w6(32'hbba2ddf8),
	.w7(32'h3a4aba0f),
	.w8(32'h3ba8c989),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45b35f),
	.w1(32'hbc1440b8),
	.w2(32'h3ae8c594),
	.w3(32'h3bbdaea1),
	.w4(32'hbbef69dd),
	.w5(32'h3b3b39f0),
	.w6(32'hbaf84b77),
	.w7(32'hbc29f6e4),
	.w8(32'hbad59098),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc17db5),
	.w1(32'h3acd17ad),
	.w2(32'h3b9f49f5),
	.w3(32'h3abdf97e),
	.w4(32'h3c156546),
	.w5(32'h3c6dd839),
	.w6(32'hbc732311),
	.w7(32'h3c10b3a5),
	.w8(32'h3c9f9d35),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb3a26),
	.w1(32'h3a9a1158),
	.w2(32'h39fd1667),
	.w3(32'h3c1e7cd7),
	.w4(32'h3abb471b),
	.w5(32'hba1ec05f),
	.w6(32'h3c7db9a5),
	.w7(32'h3b99f3e1),
	.w8(32'h3a9d5d5d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52197c),
	.w1(32'hbab6c6d2),
	.w2(32'hbb126a77),
	.w3(32'h39807632),
	.w4(32'hbaf51cdc),
	.w5(32'hbb6fdc9a),
	.w6(32'h3ac66334),
	.w7(32'h3c9e9bb1),
	.w8(32'h3c893637),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab5709),
	.w1(32'h3c486da6),
	.w2(32'h3bc71ba6),
	.w3(32'hbb02f803),
	.w4(32'h3c1651d9),
	.w5(32'hbb448685),
	.w6(32'h3c3c61c3),
	.w7(32'h3b0cde18),
	.w8(32'hbb52c26f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39c7ad),
	.w1(32'h3a1921e9),
	.w2(32'h3aab68b9),
	.w3(32'hbc2e9ce2),
	.w4(32'h3b3f62c8),
	.w5(32'h3bb00c3c),
	.w6(32'hbc586591),
	.w7(32'h3ba620e9),
	.w8(32'h3c0c355f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb062fc4),
	.w1(32'h3a4b82af),
	.w2(32'h3c258bd5),
	.w3(32'h3abe1d5d),
	.w4(32'hbae16d6a),
	.w5(32'h3c36a7e9),
	.w6(32'h3b81aac3),
	.w7(32'h3b2ae88e),
	.w8(32'h3c465810),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8085f9),
	.w1(32'hbba51bbe),
	.w2(32'hbaebd443),
	.w3(32'h3b81bd79),
	.w4(32'hbbf8777d),
	.w5(32'hbb9a5c9c),
	.w6(32'h3b98d7ed),
	.w7(32'hbbbaabd6),
	.w8(32'hbb9042d3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb55d9),
	.w1(32'hbb1f8beb),
	.w2(32'h3ba4f0db),
	.w3(32'hbb064e19),
	.w4(32'h3b037dcc),
	.w5(32'h3c2a6be2),
	.w6(32'hbb209553),
	.w7(32'h3b84a892),
	.w8(32'h3c72567f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9a54a),
	.w1(32'h3c557410),
	.w2(32'h3c7f3b72),
	.w3(32'h3bbf262a),
	.w4(32'h3ca89b7b),
	.w5(32'h3c8aa534),
	.w6(32'h3c10e1c7),
	.w7(32'h3c88ef19),
	.w8(32'h3ca2b9fa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b019c),
	.w1(32'hba5830ba),
	.w2(32'hb985d24f),
	.w3(32'h3c3070f2),
	.w4(32'hbc4978ea),
	.w5(32'hbbdb1062),
	.w6(32'h3c5ca5ba),
	.w7(32'h3b4f3d13),
	.w8(32'h3c6c4e77),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cedc8),
	.w1(32'hbb8ec35b),
	.w2(32'hba09c4d6),
	.w3(32'h3c0e53c1),
	.w4(32'hbc21ac45),
	.w5(32'hbbd402c1),
	.w6(32'h3c0e2405),
	.w7(32'hbc3748f5),
	.w8(32'hbc11cb2b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96522f),
	.w1(32'h3b1558f8),
	.w2(32'hbb4e4300),
	.w3(32'hbb93cc3d),
	.w4(32'hbab5be4f),
	.w5(32'hbb8394bb),
	.w6(32'hbc04b99a),
	.w7(32'hbc2c9672),
	.w8(32'hbc71f7ac),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4448dc),
	.w1(32'hbaf73ed6),
	.w2(32'hbb40017b),
	.w3(32'hbb178884),
	.w4(32'hba980f7e),
	.w5(32'hbb879156),
	.w6(32'hbc149f59),
	.w7(32'h3c812d80),
	.w8(32'h3bc0a47d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2546dc),
	.w1(32'h3b20b75f),
	.w2(32'h3b8ac9d3),
	.w3(32'hbb6c8a09),
	.w4(32'h3b4bdaca),
	.w5(32'h3bd866d9),
	.w6(32'h3beabf5c),
	.w7(32'h3b7aa959),
	.w8(32'h3bf90818),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72c66e),
	.w1(32'h3b8c71ed),
	.w2(32'h3b7bda01),
	.w3(32'h3b54c6d0),
	.w4(32'hbba40723),
	.w5(32'h399ec504),
	.w6(32'h3b799772),
	.w7(32'h37b6ceef),
	.w8(32'hba24bf61),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3c3c7),
	.w1(32'hb9c3c49e),
	.w2(32'hbb0853e5),
	.w3(32'h3b04ab0f),
	.w4(32'h3be8adac),
	.w5(32'h3ba1ce61),
	.w6(32'hbab43f5a),
	.w7(32'h3c2cdd6b),
	.w8(32'h3be459f9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2ca56),
	.w1(32'h390ba859),
	.w2(32'hbaa5dff2),
	.w3(32'h3b6ba57e),
	.w4(32'h3853e7ae),
	.w5(32'hba1b3a5d),
	.w6(32'h3c226126),
	.w7(32'hb8b6be78),
	.w8(32'hba957743),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fbad1),
	.w1(32'hbc1889a9),
	.w2(32'hbbfe968e),
	.w3(32'hbaaf58dc),
	.w4(32'hbc152d90),
	.w5(32'hbc4b6ed6),
	.w6(32'hbaef2f33),
	.w7(32'hbb9c21be),
	.w8(32'hbbaf72ad),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc450e),
	.w1(32'hb9516fb3),
	.w2(32'h3917f6e1),
	.w3(32'hbc715dac),
	.w4(32'hbaa6fcc7),
	.w5(32'hbafe7b7d),
	.w6(32'hbc0f09b7),
	.w7(32'hbaceecd2),
	.w8(32'hbb29f240),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0eab27),
	.w1(32'hba50fad0),
	.w2(32'hbb003162),
	.w3(32'hbb2d1f93),
	.w4(32'h38c80827),
	.w5(32'hb643241f),
	.w6(32'hbb497904),
	.w7(32'h3a14fd52),
	.w8(32'h3acbaef0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b0d74),
	.w1(32'h3a0d0c2f),
	.w2(32'h3911ba70),
	.w3(32'hba77c3ce),
	.w4(32'h3b0428f5),
	.w5(32'hb93792c5),
	.w6(32'h3944d261),
	.w7(32'h3c261a91),
	.w8(32'h3b266a15),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3309e),
	.w1(32'h3adb86c3),
	.w2(32'h3aee473c),
	.w3(32'hbb6c5349),
	.w4(32'h3ba31232),
	.w5(32'h3b9297a2),
	.w6(32'hbba4683f),
	.w7(32'h3bd81a0e),
	.w8(32'h3bfc5960),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2616bb),
	.w1(32'h394e91dc),
	.w2(32'h3b3a6b75),
	.w3(32'h3a54ac0a),
	.w4(32'h3bf3ea0a),
	.w5(32'h3c2feab6),
	.w6(32'h3b7cf936),
	.w7(32'h3c0903c7),
	.w8(32'h3c4b01fb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a869e68),
	.w1(32'hbc1a4292),
	.w2(32'h3bb99ee9),
	.w3(32'h3b899746),
	.w4(32'hbabfc9a3),
	.w5(32'h3b189978),
	.w6(32'h3bee9d05),
	.w7(32'h3c0ea87d),
	.w8(32'h3c11bba2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c573df5),
	.w1(32'hbc71adb9),
	.w2(32'hbc240c5e),
	.w3(32'h3c72cb5c),
	.w4(32'hbcbc0d16),
	.w5(32'hbc478b3b),
	.w6(32'h3c95123c),
	.w7(32'hbcaa6262),
	.w8(32'hbca12299),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c6f79),
	.w1(32'hbbbb038c),
	.w2(32'hbbc30952),
	.w3(32'hbbf2f2fe),
	.w4(32'hbbe0dd14),
	.w5(32'hbc6d6140),
	.w6(32'hbb14a01c),
	.w7(32'h3b04059f),
	.w8(32'hbb79afe5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4335c),
	.w1(32'hb6b73243),
	.w2(32'h39fecede),
	.w3(32'hbb91ae95),
	.w4(32'hbb1e4378),
	.w5(32'h399c85c2),
	.w6(32'h3bc173d8),
	.w7(32'hbb41812b),
	.w8(32'h3a852f80),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9597f8f),
	.w1(32'hba3bf9c0),
	.w2(32'hbb232ddf),
	.w3(32'hbb1d11e7),
	.w4(32'hba7f7c11),
	.w5(32'hbac168ce),
	.w6(32'hbb21ef06),
	.w7(32'hba4884f7),
	.w8(32'h3a8385a1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0b959),
	.w1(32'hb916bbd2),
	.w2(32'h3b093eeb),
	.w3(32'hba5a9655),
	.w4(32'h3abf1ddb),
	.w5(32'h3b9066d0),
	.w6(32'hbc07dc80),
	.w7(32'h3864ec22),
	.w8(32'h3bb4a440),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06628c),
	.w1(32'hbb834c4e),
	.w2(32'hbbf71199),
	.w3(32'h3a98155a),
	.w4(32'h3a3fedb8),
	.w5(32'hbb24d09e),
	.w6(32'h3b168740),
	.w7(32'h3af4edd8),
	.w8(32'hb986c6d0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf84480),
	.w1(32'hbafefeac),
	.w2(32'hbaee66fa),
	.w3(32'hbac8fe44),
	.w4(32'hbaaa0cd2),
	.w5(32'hba7c195e),
	.w6(32'h3b2a0f19),
	.w7(32'hbb4130bc),
	.w8(32'hbac20525),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae663e9),
	.w1(32'h3abbcb38),
	.w2(32'h3c2fd688),
	.w3(32'hba95b25f),
	.w4(32'hbb5a4144),
	.w5(32'h3b47f9c0),
	.w6(32'h3b98f0b5),
	.w7(32'hbbbb0127),
	.w8(32'h3a9a48d7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cd721),
	.w1(32'hb9931a96),
	.w2(32'h39f20826),
	.w3(32'h3cb6db63),
	.w4(32'hbb77e12f),
	.w5(32'hbae53814),
	.w6(32'h3c693a7f),
	.w7(32'hba9aafbc),
	.w8(32'hba09a439),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaf451),
	.w1(32'hb6d1015d),
	.w2(32'h3b312e46),
	.w3(32'hbb483f4e),
	.w4(32'h3a9fde58),
	.w5(32'hbbc5801e),
	.w6(32'h3a4703f4),
	.w7(32'h39dc9471),
	.w8(32'hbaf7fe18),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8ac3c),
	.w1(32'hb9f928d6),
	.w2(32'h3bde5fda),
	.w3(32'hbca7c0f8),
	.w4(32'hbafd9106),
	.w5(32'hbb74454d),
	.w6(32'hbca7a343),
	.w7(32'hbb733aa4),
	.w8(32'h3b121639),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e9adc),
	.w1(32'h3ae18d39),
	.w2(32'h3a82a302),
	.w3(32'h3a1b3683),
	.w4(32'h3a612ad5),
	.w5(32'h39aff242),
	.w6(32'h3a3b965c),
	.w7(32'h3abebb91),
	.w8(32'h38d856df),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1332ac),
	.w1(32'hbb88ee1e),
	.w2(32'hbbe02dd7),
	.w3(32'h3a264805),
	.w4(32'h3b57fcd9),
	.w5(32'hbb48e363),
	.w6(32'h3a8eee75),
	.w7(32'h3b0a552e),
	.w8(32'h3b6f8fb9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc073019),
	.w1(32'h3a20e656),
	.w2(32'h3b6b4929),
	.w3(32'hbc5646fc),
	.w4(32'hbb0ad4c5),
	.w5(32'h3a028e3a),
	.w6(32'h3b2e5d26),
	.w7(32'hba96558c),
	.w8(32'hba6ea700),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81f747),
	.w1(32'hbb03764b),
	.w2(32'hbbb13b9a),
	.w3(32'h3ae79c35),
	.w4(32'h3aabc6f4),
	.w5(32'hbb04afd8),
	.w6(32'hb9e639e8),
	.w7(32'h3ae570f7),
	.w8(32'hba676f89),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0937b5),
	.w1(32'h3b1dfcd2),
	.w2(32'h3b0a1a3e),
	.w3(32'hbb722e93),
	.w4(32'h3bb7bbfc),
	.w5(32'h3ab4222b),
	.w6(32'hba4c22f9),
	.w7(32'h3b0b7888),
	.w8(32'hb9ee9a65),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12176b),
	.w1(32'hbac8ec27),
	.w2(32'h3be1917c),
	.w3(32'h3c42500f),
	.w4(32'hbc29885b),
	.w5(32'h3a50a3fc),
	.w6(32'h3ac15f18),
	.w7(32'hbb437b5c),
	.w8(32'h3b70abaa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc060f9),
	.w1(32'h3b62d31f),
	.w2(32'h3bb66130),
	.w3(32'h3b4e2ed8),
	.w4(32'hbc4931e3),
	.w5(32'hbbceaedf),
	.w6(32'h3ab47324),
	.w7(32'hbcb6d52c),
	.w8(32'hbbe786c8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39dcbf),
	.w1(32'h3b1b55ca),
	.w2(32'h3af70f36),
	.w3(32'hbb09f73e),
	.w4(32'h3bc2cf4d),
	.w5(32'h3bf7d660),
	.w6(32'hbaec8c4b),
	.w7(32'h3bf41646),
	.w8(32'h3c334f5d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a64aa),
	.w1(32'hb9005cc3),
	.w2(32'h39256f92),
	.w3(32'h3ad378e0),
	.w4(32'h3a1f8d37),
	.w5(32'hbae1fbac),
	.w6(32'h3b97fd73),
	.w7(32'h3b1c9634),
	.w8(32'h3a876725),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0f965),
	.w1(32'hb736ae46),
	.w2(32'h3b6243d2),
	.w3(32'h3ab53215),
	.w4(32'hbbfb1761),
	.w5(32'hbb12211a),
	.w6(32'h3b574a5d),
	.w7(32'hbb0e1d50),
	.w8(32'h3b0cef38),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188fce),
	.w1(32'hbba14f0a),
	.w2(32'hbbaaaa41),
	.w3(32'hbbbf4f90),
	.w4(32'hbb5bcfbc),
	.w5(32'hbb8fbd14),
	.w6(32'hbb6b1bc9),
	.w7(32'hbaac387a),
	.w8(32'hbb1d9db0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba148c5),
	.w1(32'hbbdfbf78),
	.w2(32'hbafca3a4),
	.w3(32'hbb7986c0),
	.w4(32'hbc81e0e9),
	.w5(32'hbc33e4fd),
	.w6(32'hbb129053),
	.w7(32'hbc849e26),
	.w8(32'hbc3a0558),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba9d95),
	.w1(32'h391d1c0b),
	.w2(32'h3c173b34),
	.w3(32'hbbd6d378),
	.w4(32'h3b09eb39),
	.w5(32'h3c81b50b),
	.w6(32'hba8cd3fe),
	.w7(32'h3cdd9bfd),
	.w8(32'h3d368911),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc822ffc),
	.w1(32'hbb1db1d5),
	.w2(32'hba459b89),
	.w3(32'hbc66efbd),
	.w4(32'hbaf1d5cf),
	.w5(32'hbc72ea8a),
	.w6(32'h3c1c013a),
	.w7(32'hbb8e3700),
	.w8(32'hbca41971),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61e117),
	.w1(32'hbb26b6a1),
	.w2(32'hbb1fc267),
	.w3(32'hbb9a6d96),
	.w4(32'hb8bf3fc5),
	.w5(32'hba9d7fc1),
	.w6(32'hbbf9d92a),
	.w7(32'h3aa136ec),
	.w8(32'h39396925),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02cd20),
	.w1(32'hbc8a585d),
	.w2(32'hbb7e0f0b),
	.w3(32'h39083fc0),
	.w4(32'hbaa50908),
	.w5(32'h3a8ed596),
	.w6(32'h3acbc39e),
	.w7(32'h3c622846),
	.w8(32'h3c731b74),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba308cc),
	.w1(32'hbb8613c1),
	.w2(32'h3b9c7c09),
	.w3(32'hbbe078cf),
	.w4(32'h3b3c5406),
	.w5(32'h3c976614),
	.w6(32'h3a26d869),
	.w7(32'h3beeabc5),
	.w8(32'h3ce85e3f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf596c9),
	.w1(32'hbb5a809c),
	.w2(32'hbb8f134f),
	.w3(32'hbb0182ac),
	.w4(32'h3b8fed3a),
	.w5(32'h3b416852),
	.w6(32'h3bb45d09),
	.w7(32'h3ba06060),
	.w8(32'h3bc30818),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00df3),
	.w1(32'hba15d379),
	.w2(32'hba136170),
	.w3(32'h3a2d8f33),
	.w4(32'h3c0889bf),
	.w5(32'h3c04d8e5),
	.w6(32'h3b81e4c8),
	.w7(32'h3c4152c3),
	.w8(32'h3c7620c8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892bfa),
	.w1(32'hbbe542f0),
	.w2(32'hbb1e9e44),
	.w3(32'h3b959d40),
	.w4(32'h3be88696),
	.w5(32'h3c235ed9),
	.w6(32'h3c431cda),
	.w7(32'h3c3df2d6),
	.w8(32'h3c8b43e8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc88fc8),
	.w1(32'hbc2136cb),
	.w2(32'hbbb78b50),
	.w3(32'h3b911436),
	.w4(32'hbb864034),
	.w5(32'h3b85b8e2),
	.w6(32'h3c8032d5),
	.w7(32'h3b8e5fa2),
	.w8(32'h3c8f1de2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d6a2a),
	.w1(32'hbcbd0dbd),
	.w2(32'hbcc77cf3),
	.w3(32'hbbed1d6d),
	.w4(32'hbc9593cf),
	.w5(32'hbcb7691a),
	.w6(32'h3b824848),
	.w7(32'hbc49ec81),
	.w8(32'hbc512b70),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc448a3a),
	.w1(32'h3b2a5ce1),
	.w2(32'h3c011122),
	.w3(32'hbc900df8),
	.w4(32'h3bed7baa),
	.w5(32'h3c60d0b2),
	.w6(32'hbc392484),
	.w7(32'h3b901ae5),
	.w8(32'h3bf658f0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7821d8),
	.w1(32'hbb62f84d),
	.w2(32'hbc1c52f0),
	.w3(32'h3c0218c6),
	.w4(32'hbc41914c),
	.w5(32'hbcbd3c7e),
	.w6(32'h3b1f3796),
	.w7(32'hbc022326),
	.w8(32'hbbb95eee),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba952a79),
	.w1(32'hba63ec7f),
	.w2(32'hbb06a832),
	.w3(32'hbc0fd729),
	.w4(32'hbb3dfb2f),
	.w5(32'hbb8bc797),
	.w6(32'hbc15ab9d),
	.w7(32'hba078391),
	.w8(32'hbb28d9cb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ee1a2),
	.w1(32'hbb489ca4),
	.w2(32'hbbceaad2),
	.w3(32'hbb8f646c),
	.w4(32'hbb7c6c4e),
	.w5(32'hbc724a4a),
	.w6(32'hbac91ece),
	.w7(32'hbc328f53),
	.w8(32'hbc983c77),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35fc30),
	.w1(32'h3a067d72),
	.w2(32'h3c03896e),
	.w3(32'hbc5a032f),
	.w4(32'h3bc1fdc7),
	.w5(32'h3c2c764f),
	.w6(32'hbc52cc3f),
	.w7(32'h3bc6031c),
	.w8(32'h3c428118),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b764770),
	.w1(32'hbba283f6),
	.w2(32'h3b94e727),
	.w3(32'h3c161d2e),
	.w4(32'hba9938f7),
	.w5(32'h3c95f290),
	.w6(32'h3c23eed9),
	.w7(32'hbbf93cda),
	.w8(32'h3c2c8be4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb87c73),
	.w1(32'hbbdbb973),
	.w2(32'hbbc2c9cc),
	.w3(32'hb9b898f8),
	.w4(32'h3b14cab6),
	.w5(32'hbc643bb6),
	.w6(32'hbb16a830),
	.w7(32'h3c24fdaf),
	.w8(32'h3b13af51),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77ba23),
	.w1(32'h3b351c49),
	.w2(32'h3b7fb4ce),
	.w3(32'hbc3c9498),
	.w4(32'h3b1b5d54),
	.w5(32'h3b816cec),
	.w6(32'hbba7ed91),
	.w7(32'h39ee2255),
	.w8(32'h3b8657e9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b114920),
	.w1(32'h3aea3b4b),
	.w2(32'h398d6208),
	.w3(32'h3b607f81),
	.w4(32'h3b2f0c96),
	.w5(32'h3b1dd90e),
	.w6(32'h3b943714),
	.w7(32'h3b9b9854),
	.w8(32'h3bcdbd8c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aedd0),
	.w1(32'hbc02394e),
	.w2(32'hbc18f9fb),
	.w3(32'hbb05b0e5),
	.w4(32'hbbb5a0e9),
	.w5(32'hbc0a72c1),
	.w6(32'hba946db1),
	.w7(32'hbb96b588),
	.w8(32'hbb9fcc4b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ff497),
	.w1(32'hbc63f05f),
	.w2(32'hbb7188cd),
	.w3(32'hbb5296c9),
	.w4(32'hbc800ef7),
	.w5(32'hbb62f243),
	.w6(32'hba4a3ca5),
	.w7(32'hbbc5c65b),
	.w8(32'h3bb375c7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc03e64),
	.w1(32'hbbac4af6),
	.w2(32'hbb985fde),
	.w3(32'hbc41d83c),
	.w4(32'hbba72d9e),
	.w5(32'hbb45777e),
	.w6(32'hbc25390d),
	.w7(32'hbba03161),
	.w8(32'hbb8113e2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba3073),
	.w1(32'hbb305be7),
	.w2(32'hbc8a9181),
	.w3(32'hbb7b319c),
	.w4(32'hbc6c62aa),
	.w5(32'hbc80db21),
	.w6(32'hbb41263b),
	.w7(32'hbc0000df),
	.w8(32'hbc8ba619),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8910af),
	.w1(32'hbb0cb55c),
	.w2(32'hba5cd3e2),
	.w3(32'hbce721fc),
	.w4(32'h3962c651),
	.w5(32'h3a9b65bd),
	.w6(32'hbc87f8a9),
	.w7(32'hba572403),
	.w8(32'hbb1e841e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b5483),
	.w1(32'hbc20dc0c),
	.w2(32'hbbec0fc9),
	.w3(32'hba59e54c),
	.w4(32'hbc1ddef5),
	.w5(32'hbbe26167),
	.w6(32'hbb6a8dfd),
	.w7(32'hbc133acb),
	.w8(32'hbb0de96f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841ed4),
	.w1(32'h3b47f24a),
	.w2(32'h3b83d8fd),
	.w3(32'hba19a887),
	.w4(32'h39a2dcf6),
	.w5(32'h3c10137a),
	.w6(32'h3b448a9b),
	.w7(32'h3be16ab7),
	.w8(32'hb78191dc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b0e99),
	.w1(32'h3b2558fd),
	.w2(32'hbca4ae58),
	.w3(32'h3c48eccd),
	.w4(32'hbbefaa74),
	.w5(32'hbce15283),
	.w6(32'h3c166515),
	.w7(32'hbc6a9d80),
	.w8(32'hbcc5b94e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb67212),
	.w1(32'hbb9aec02),
	.w2(32'h3b26f3fd),
	.w3(32'hbcb3a2f7),
	.w4(32'hba726ba8),
	.w5(32'h3bc83479),
	.w6(32'hbccadba8),
	.w7(32'hbb7eb8b6),
	.w8(32'h3b3920aa),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a72b4),
	.w1(32'hbb8d0dca),
	.w2(32'h3b8e6216),
	.w3(32'h3bbbc992),
	.w4(32'h3bde43dd),
	.w5(32'h3cc94298),
	.w6(32'h3b734dfe),
	.w7(32'h3bf40d51),
	.w8(32'h3c88c819),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1067a1),
	.w1(32'h3b9a2b36),
	.w2(32'h3b47c08d),
	.w3(32'h3c9a3dbc),
	.w4(32'h3c3d50ca),
	.w5(32'h3c3b7572),
	.w6(32'h3b81a2f3),
	.w7(32'h3c2132ee),
	.w8(32'h3bf049d8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b310a3c),
	.w1(32'hbb58f4b8),
	.w2(32'h3bc98ce4),
	.w3(32'h3be4a16f),
	.w4(32'hb9d71369),
	.w5(32'h3c39ba62),
	.w6(32'hb97d4fc5),
	.w7(32'hbb62c521),
	.w8(32'h3c173590),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962c9ac),
	.w1(32'h3d4bf7a3),
	.w2(32'h3d74e355),
	.w3(32'h3b9b68ff),
	.w4(32'h3d851e06),
	.w5(32'h3d9a9c56),
	.w6(32'h3b28f2d5),
	.w7(32'h3d1d5377),
	.w8(32'h3d533ced),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d20f79d),
	.w1(32'hbaa98e8d),
	.w2(32'hbbc5cce1),
	.w3(32'h3d699a2f),
	.w4(32'hbbd061f4),
	.w5(32'hbc030fa0),
	.w6(32'h3d28cc03),
	.w7(32'hbb8cf445),
	.w8(32'hbbccc224),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91df22),
	.w1(32'hbab17ae2),
	.w2(32'hb901acb9),
	.w3(32'hbbe739f5),
	.w4(32'hb8e7505c),
	.w5(32'h3ac47fbd),
	.w6(32'hbb805d93),
	.w7(32'h3a9382be),
	.w8(32'h3ac40253),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26cd62),
	.w1(32'h3d224beb),
	.w2(32'h3d945bed),
	.w3(32'hba2075e8),
	.w4(32'h3d5e036c),
	.w5(32'h3db0265e),
	.w6(32'h3ae2080e),
	.w7(32'h3d34dd80),
	.w8(32'h3d8a2d48),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d502bde),
	.w1(32'h3a220d3f),
	.w2(32'h3b87a9f4),
	.w3(32'h3d8b29a7),
	.w4(32'h3b0a851b),
	.w5(32'h3baf1ef7),
	.w6(32'h3d31eee1),
	.w7(32'h39580f88),
	.w8(32'h3b8436c9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b141545),
	.w1(32'hbb6829e4),
	.w2(32'hba7d7c97),
	.w3(32'h3b8a1961),
	.w4(32'hbb2848c2),
	.w5(32'hb8ee9606),
	.w6(32'h3bb1a092),
	.w7(32'hbba9363c),
	.w8(32'hbb71f87e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15f47c),
	.w1(32'hbc17767d),
	.w2(32'hbc220cf4),
	.w3(32'hba9d7f3b),
	.w4(32'hbb526f98),
	.w5(32'hbb1e6eff),
	.w6(32'hbb865cf6),
	.w7(32'hbaa4ceec),
	.w8(32'h3b8b9677),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc612bea),
	.w1(32'hbb4d8e14),
	.w2(32'hbb85e86b),
	.w3(32'hbc9bb9db),
	.w4(32'hbbaacde7),
	.w5(32'hbbfaae0a),
	.w6(32'hbc36f74a),
	.w7(32'hbb7e8b7b),
	.w8(32'hbbc056b0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60fb4f),
	.w1(32'h3b068cb7),
	.w2(32'h3b9912ec),
	.w3(32'hbbca9a0a),
	.w4(32'h39f77791),
	.w5(32'h3c05e1f0),
	.w6(32'hbba1043f),
	.w7(32'h3b8d186b),
	.w8(32'h3b9b87c9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a31bf1),
	.w1(32'hbae53a17),
	.w2(32'h3b59e00e),
	.w3(32'h3ac91eb2),
	.w4(32'hbbd86d35),
	.w5(32'hbbf90088),
	.w6(32'h3bcaa096),
	.w7(32'hbc5b61d3),
	.w8(32'hbc499130),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aa2d1),
	.w1(32'hbc82e94a),
	.w2(32'hbc5ba71b),
	.w3(32'hbba56e65),
	.w4(32'hbae52667),
	.w5(32'hbc2104d5),
	.w6(32'hbc1ed702),
	.w7(32'hbafd3a98),
	.w8(32'hbb7ff5c2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36f88d),
	.w1(32'hbb97f864),
	.w2(32'h3aa89403),
	.w3(32'hbb868a9a),
	.w4(32'h3b977ed3),
	.w5(32'hbb4c919d),
	.w6(32'h3ad0413d),
	.w7(32'h3b553895),
	.w8(32'hbc267da5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe21cd),
	.w1(32'hbb33f2a1),
	.w2(32'hba70c85f),
	.w3(32'h3c009f73),
	.w4(32'hbbe626a5),
	.w5(32'hbc008673),
	.w6(32'h3b0eca5b),
	.w7(32'hbc0ad14c),
	.w8(32'hbc2c7fdb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94e39c),
	.w1(32'h3b83e667),
	.w2(32'h3bb46909),
	.w3(32'hbc8995d2),
	.w4(32'h3b19a453),
	.w5(32'h3a2c576a),
	.w6(32'hbca63d63),
	.w7(32'h3a07426c),
	.w8(32'h3b6e45c9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b28de),
	.w1(32'hbb121f0b),
	.w2(32'hbafcf8c1),
	.w3(32'h3b5e4132),
	.w4(32'hbb1f477e),
	.w5(32'hbb4357d6),
	.w6(32'h39ad75fd),
	.w7(32'hbb5ab5fa),
	.w8(32'hbb2c1222),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a00ad),
	.w1(32'h3bbb155e),
	.w2(32'h3b8e0e5a),
	.w3(32'hbab497ad),
	.w4(32'h3bb0a3c5),
	.w5(32'h3b7f8b7e),
	.w6(32'hbab34028),
	.w7(32'h3baed5b9),
	.w8(32'h3b8764c8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59fed1),
	.w1(32'hbbd014d0),
	.w2(32'hba98bbd3),
	.w3(32'h3b3dd01f),
	.w4(32'hb90a6a2f),
	.w5(32'h3bd041c4),
	.w6(32'h3b22a536),
	.w7(32'hbc0d8112),
	.w8(32'hbc0394ec),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae80e81),
	.w1(32'hbbeb8885),
	.w2(32'hbb3e0afa),
	.w3(32'hb72f60b0),
	.w4(32'hbb85a826),
	.w5(32'hbbf08bc5),
	.w6(32'h3bfd08f8),
	.w7(32'hbb181fdb),
	.w8(32'hbbc3ad1f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc643fd8),
	.w1(32'hbc5c47cb),
	.w2(32'h3ad82b1f),
	.w3(32'h3b2c63b0),
	.w4(32'h3b1ebc03),
	.w5(32'h3bb79c68),
	.w6(32'hbc001e42),
	.w7(32'h3ac8b37f),
	.w8(32'h3b2ebb31),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d06f0),
	.w1(32'hbc6cf197),
	.w2(32'hbca9f552),
	.w3(32'h3b795350),
	.w4(32'hbcf432d1),
	.w5(32'hbcce57c5),
	.w6(32'hb997419b),
	.w7(32'hbcd7196a),
	.w8(32'hbcbc1301),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc872e92),
	.w1(32'hbc912f8a),
	.w2(32'hbc1d3ef7),
	.w3(32'hbcd35a70),
	.w4(32'hbc86ef43),
	.w5(32'h3baddb5a),
	.w6(32'hbc88be31),
	.w7(32'hbc9b2253),
	.w8(32'hba84051b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf24c),
	.w1(32'h3a2b7edd),
	.w2(32'h3b50bbc1),
	.w3(32'hbb594d20),
	.w4(32'h3b79ba04),
	.w5(32'h3bc8a014),
	.w6(32'hbbdfba23),
	.w7(32'h3b8ce7d2),
	.w8(32'h3bcad612),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad645eb),
	.w1(32'hbabcb98c),
	.w2(32'h3b997b6c),
	.w3(32'h3b625a71),
	.w4(32'hbb87e232),
	.w5(32'hb9eee96f),
	.w6(32'h3acde2dd),
	.w7(32'h3b3afae9),
	.w8(32'h3c309522),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae30ec6),
	.w1(32'hbbea9316),
	.w2(32'hbbe451a7),
	.w3(32'hbac1dfff),
	.w4(32'hbbcd93c4),
	.w5(32'hbb953d93),
	.w6(32'h3b8c9fed),
	.w7(32'hbb292412),
	.w8(32'hbb0d0a13),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb914f7a),
	.w1(32'h3ab4e5e3),
	.w2(32'h3ac60fa0),
	.w3(32'hbac4e412),
	.w4(32'h3ab7a55c),
	.w5(32'h3a44857b),
	.w6(32'hbb3583b5),
	.w7(32'h3b2cbc3b),
	.w8(32'h3b1e2336),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1338f7),
	.w1(32'h3ca6e344),
	.w2(32'h3d21b4df),
	.w3(32'hba0d067e),
	.w4(32'h3d395ad9),
	.w5(32'h3d9cee83),
	.w6(32'h3a8eb6a2),
	.w7(32'h3d1cf8a3),
	.w8(32'h3d6d4aed),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d39f5de),
	.w1(32'h3b89a5df),
	.w2(32'h3bbe63ea),
	.w3(32'h3d863297),
	.w4(32'hbc144273),
	.w5(32'hbcbae0ee),
	.w6(32'h3d2bcd3d),
	.w7(32'hbc2f94ee),
	.w8(32'hbcd4147b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a55af),
	.w1(32'h3a79344e),
	.w2(32'hbb9449fe),
	.w3(32'hbc1642ac),
	.w4(32'hbafc3b4f),
	.w5(32'hbb86ade0),
	.w6(32'hbc269ab2),
	.w7(32'h3c0c1747),
	.w8(32'hbaedc97f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51edf5),
	.w1(32'hbb6aca04),
	.w2(32'hbaf8a586),
	.w3(32'hbcb9f07b),
	.w4(32'hbb737dcb),
	.w5(32'hbab0e0d5),
	.w6(32'hbc6089a5),
	.w7(32'hbb851be9),
	.w8(32'hba844dc3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9582d0),
	.w1(32'h3bcc0f9f),
	.w2(32'h3babd427),
	.w3(32'hbb71faf4),
	.w4(32'h3c0c2460),
	.w5(32'h3be43f13),
	.w6(32'hbb46cc17),
	.w7(32'h3bc88a94),
	.w8(32'h3bac6490),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dee9e),
	.w1(32'h3b845fb3),
	.w2(32'hbb2339b7),
	.w3(32'h3b2e3751),
	.w4(32'h3b6b2712),
	.w5(32'hbad8660c),
	.w6(32'h3b1f5b05),
	.w7(32'h3b323702),
	.w8(32'hbc0c1199),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf216c9),
	.w1(32'hbb324d55),
	.w2(32'hbb800787),
	.w3(32'hbbd1d0d0),
	.w4(32'hbabfba87),
	.w5(32'hbaf00428),
	.w6(32'hbc2a0a96),
	.w7(32'hbb1afa2a),
	.w8(32'hbb3f6714),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e74fb),
	.w1(32'hbbb2a5d8),
	.w2(32'hbc298f9c),
	.w3(32'hbb544fd3),
	.w4(32'hbbd9d43a),
	.w5(32'h3c40c423),
	.w6(32'hbb833b8a),
	.w7(32'hbab46ae0),
	.w8(32'h3bdb4c92),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f07fe),
	.w1(32'h3b046108),
	.w2(32'h3c0f25d2),
	.w3(32'h3b12fe21),
	.w4(32'h3b85e018),
	.w5(32'h3bfec2f5),
	.w6(32'hbb305b6b),
	.w7(32'h3c01d974),
	.w8(32'h3c862ead),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4132a),
	.w1(32'hbc5250b9),
	.w2(32'h39aaa21e),
	.w3(32'h3c3539aa),
	.w4(32'hbc0a4447),
	.w5(32'h3ba07a48),
	.w6(32'h3ca1a92d),
	.w7(32'hbbba08b8),
	.w8(32'h3b9f935d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ce88),
	.w1(32'h3c093d88),
	.w2(32'h3bbef7f9),
	.w3(32'hbc26781e),
	.w4(32'h3c259a45),
	.w5(32'h3bd74e95),
	.w6(32'hbb97076f),
	.w7(32'h3c37aac1),
	.w8(32'h3c02b14f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a7274),
	.w1(32'hbbc24696),
	.w2(32'hbc9a00ca),
	.w3(32'h3b71780f),
	.w4(32'hbc7427fa),
	.w5(32'hbc82e078),
	.w6(32'h3ba70422),
	.w7(32'h3b3e2423),
	.w8(32'hbb916d0c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule