module layer_8_featuremap_19(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7e09a),
	.w1(32'hbb97a53b),
	.w2(32'h3beefa48),
	.w3(32'h3b956b0c),
	.w4(32'h3d31e5bd),
	.w5(32'h3bf0781c),
	.w6(32'h3a0414c7),
	.w7(32'h3b8998b0),
	.w8(32'h3c7b9740),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1adfa),
	.w1(32'hbb3db22a),
	.w2(32'hbb74a921),
	.w3(32'h3cb010a6),
	.w4(32'h3b6fe139),
	.w5(32'hba818beb),
	.w6(32'h3c2739ff),
	.w7(32'h3bec25cb),
	.w8(32'h3cf047af),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978cd6),
	.w1(32'h3c810f39),
	.w2(32'h3c753452),
	.w3(32'h3b9d2962),
	.w4(32'hb9a7bf89),
	.w5(32'h3a22eced),
	.w6(32'hbab48a38),
	.w7(32'hbc3461ed),
	.w8(32'h3ae77419),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2a652),
	.w1(32'hbc4cce0e),
	.w2(32'h3bcb4a69),
	.w3(32'h3baf2334),
	.w4(32'hb8c76f69),
	.w5(32'h3c405acd),
	.w6(32'h3bb53eae),
	.w7(32'h3ceb623a),
	.w8(32'hbb4a2a0e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e9389),
	.w1(32'hbc06ffd2),
	.w2(32'hbbd5c901),
	.w3(32'h3c0b739c),
	.w4(32'hbc35378b),
	.w5(32'hba3e2e63),
	.w6(32'hbcd87064),
	.w7(32'h3beb7b81),
	.w8(32'h3bc3d13e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c845b43),
	.w1(32'hbc676450),
	.w2(32'h3b8e0770),
	.w3(32'h3ce5bedf),
	.w4(32'h3cc96fc4),
	.w5(32'hbc1db148),
	.w6(32'h3c219133),
	.w7(32'h3c9ea7e0),
	.w8(32'hbc2d8b79),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba85a58),
	.w1(32'h3b93631b),
	.w2(32'h39e09273),
	.w3(32'h3c2b7702),
	.w4(32'h3c403518),
	.w5(32'hbc7b9172),
	.w6(32'hb91547e9),
	.w7(32'hbb04b5b5),
	.w8(32'h3c191a2f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be24b),
	.w1(32'h3ba8611c),
	.w2(32'hbb960827),
	.w3(32'h3c2eff67),
	.w4(32'h3c267ab2),
	.w5(32'h3b44c1c6),
	.w6(32'hbb8b2824),
	.w7(32'h3c6253b8),
	.w8(32'hbc578c47),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3450c3),
	.w1(32'h3b405579),
	.w2(32'h3b45b2cc),
	.w3(32'h3c2b681f),
	.w4(32'h3ae47b9b),
	.w5(32'h3c5717ab),
	.w6(32'hba8d0906),
	.w7(32'h3bd1d0fe),
	.w8(32'h3aeeeced),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba854c71),
	.w1(32'hb8564fab),
	.w2(32'hbbb3563c),
	.w3(32'hb8f1034f),
	.w4(32'h3a966927),
	.w5(32'h3c2e934f),
	.w6(32'hbbdd4312),
	.w7(32'hbb92185e),
	.w8(32'hbbcf4093),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc890aa9),
	.w1(32'h3c14c982),
	.w2(32'h3c536be7),
	.w3(32'hbaf368f2),
	.w4(32'hbac3a2ee),
	.w5(32'h3ce37149),
	.w6(32'h3c24f401),
	.w7(32'hbbd362f5),
	.w8(32'h3bb145a1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87aff7),
	.w1(32'h3a1f4892),
	.w2(32'hb8ca495f),
	.w3(32'h3c2adbb3),
	.w4(32'h3b94c53b),
	.w5(32'h3bb052fd),
	.w6(32'h3b57f3aa),
	.w7(32'hbb690adc),
	.w8(32'h3ba502cd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb970de),
	.w1(32'h3c36493d),
	.w2(32'h3b6b2a2c),
	.w3(32'h3ae01543),
	.w4(32'h3bc79a66),
	.w5(32'hbb889c2f),
	.w6(32'hbb8aa7b4),
	.w7(32'hbd34f164),
	.w8(32'hbb78179b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c168ec2),
	.w1(32'hbc0b79ae),
	.w2(32'hb8c4d8c4),
	.w3(32'hbc30725e),
	.w4(32'hbb39acfa),
	.w5(32'h3c8012e9),
	.w6(32'hba312bf8),
	.w7(32'hbd6f5013),
	.w8(32'hbadf383b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e9793),
	.w1(32'h3c1b3f8b),
	.w2(32'hba215ff8),
	.w3(32'hbc646ab3),
	.w4(32'h3bab4945),
	.w5(32'hbca3cf2b),
	.w6(32'hbd49a359),
	.w7(32'hbb85adaf),
	.w8(32'h3bfa1da9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e383e),
	.w1(32'h3c0512a7),
	.w2(32'h3bd85ce8),
	.w3(32'hba4e2cb4),
	.w4(32'hbb02ccde),
	.w5(32'h3d7d3435),
	.w6(32'h3b4ed8e9),
	.w7(32'h3bee999b),
	.w8(32'hbb96c794),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce85b24),
	.w1(32'h3bfe80da),
	.w2(32'hbb1f02ab),
	.w3(32'h3cfcad01),
	.w4(32'hbc17e9eb),
	.w5(32'hbd0c2dea),
	.w6(32'h3c307739),
	.w7(32'hbaad4dea),
	.w8(32'hbb8c87b5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc5d31),
	.w1(32'h3c308c82),
	.w2(32'h3ae883fa),
	.w3(32'h3c25b1b8),
	.w4(32'hbbe152af),
	.w5(32'hbc0cb371),
	.w6(32'h3d45fd4a),
	.w7(32'h3bc59ba6),
	.w8(32'hbb86237b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc903b5),
	.w1(32'hbbfddf61),
	.w2(32'h3c06bff2),
	.w3(32'h3abfdacb),
	.w4(32'hbc452134),
	.w5(32'hbb6e407e),
	.w6(32'h3c5c9ecb),
	.w7(32'h3b5a4067),
	.w8(32'hbb34f475),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac949d9),
	.w1(32'h3bfe7f88),
	.w2(32'h3bf7f3e1),
	.w3(32'h3be166d0),
	.w4(32'hbd31fe08),
	.w5(32'h3c7e28f8),
	.w6(32'hbb89ac57),
	.w7(32'h3d65f80a),
	.w8(32'h3bbd41a4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e9b6f),
	.w1(32'h3b1b1ff2),
	.w2(32'hbb828691),
	.w3(32'h3b3ae457),
	.w4(32'hbd5923c3),
	.w5(32'hbc180287),
	.w6(32'hbb6edb9c),
	.w7(32'hbb81b2aa),
	.w8(32'hbbad0e4e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9485b6),
	.w1(32'hbc1711de),
	.w2(32'hbbd34a99),
	.w3(32'hbbacacef),
	.w4(32'hbb1a1913),
	.w5(32'h3b46e7d8),
	.w6(32'hbbd5d85f),
	.w7(32'h3a499661),
	.w8(32'h3c0b4e11),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9f2d),
	.w1(32'h3d671702),
	.w2(32'hbc1c15e3),
	.w3(32'hb99e51b5),
	.w4(32'hbb6a5020),
	.w5(32'h3baabf94),
	.w6(32'hbb5668ac),
	.w7(32'hbc01089d),
	.w8(32'h3c8de285),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40df15),
	.w1(32'hbb15615b),
	.w2(32'hbb5d93bb),
	.w3(32'hbb03e55c),
	.w4(32'hbb8faae7),
	.w5(32'hbbb60434),
	.w6(32'hbb3eb154),
	.w7(32'hbb618d8c),
	.w8(32'h3c49d5a0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb2f9),
	.w1(32'h3b907b77),
	.w2(32'h3c504fb0),
	.w3(32'h3b0354a3),
	.w4(32'hbc3eeee6),
	.w5(32'h3c68e713),
	.w6(32'h3bc17005),
	.w7(32'hbc1c1f9f),
	.w8(32'hbbfd995f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bed41),
	.w1(32'h3baecb0f),
	.w2(32'h3c20b785),
	.w3(32'h3c9a7ef4),
	.w4(32'h3b6edd3a),
	.w5(32'h3b55762c),
	.w6(32'hbb08130c),
	.w7(32'h3c0a3fe8),
	.w8(32'hbb0ef115),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ddd83),
	.w1(32'h3c6e435f),
	.w2(32'h3baa5064),
	.w3(32'hbc1293d7),
	.w4(32'h3b0770e2),
	.w5(32'hbd1ace6b),
	.w6(32'h3c19552c),
	.w7(32'hbbda1541),
	.w8(32'h3b462339),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd16aa0),
	.w1(32'hbc5d3d90),
	.w2(32'hbbc2c5ca),
	.w3(32'hbaf0da99),
	.w4(32'hba54ae2c),
	.w5(32'hbd5186b7),
	.w6(32'h3c07a6aa),
	.w7(32'hbbf29232),
	.w8(32'h3a0edff3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c2c64),
	.w1(32'hbc4517ba),
	.w2(32'h3b8b3981),
	.w3(32'hbab55bde),
	.w4(32'hbd2c9fb3),
	.w5(32'hbb6b3e87),
	.w6(32'hbb3f9eeb),
	.w7(32'h3c03634c),
	.w8(32'hba104beb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c6431),
	.w1(32'hba36724d),
	.w2(32'hbade09b4),
	.w3(32'h3bd55420),
	.w4(32'h3b303573),
	.w5(32'h3bcc3f94),
	.w6(32'hbb72d406),
	.w7(32'h3be3bf48),
	.w8(32'h3bb9ee05),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d581cc8),
	.w1(32'h3cd6e31b),
	.w2(32'hbc0394f3),
	.w3(32'hbb81c228),
	.w4(32'h3c15c95a),
	.w5(32'hba989c84),
	.w6(32'h3cc6c71e),
	.w7(32'h3bd9c3b7),
	.w8(32'hbb05ac19),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf04306),
	.w1(32'h3c0c3fe9),
	.w2(32'hbbbf0c83),
	.w3(32'hbb7624c7),
	.w4(32'h3d294dc7),
	.w5(32'h3bac47c7),
	.w6(32'h3bb76194),
	.w7(32'h3c18abf5),
	.w8(32'h3adb3f20),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefdca9),
	.w1(32'h3a50b6ea),
	.w2(32'hbc1ffd12),
	.w3(32'hbb654f09),
	.w4(32'h3c3f00bb),
	.w5(32'h3b420784),
	.w6(32'hbb969db0),
	.w7(32'hbba5b523),
	.w8(32'h3c0f57a5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf183),
	.w1(32'h3bc5279f),
	.w2(32'hbd1859d0),
	.w3(32'hbb2c84bf),
	.w4(32'hbb6c2dbe),
	.w5(32'h3d445983),
	.w6(32'hbab42c39),
	.w7(32'h3bd94e17),
	.w8(32'h3bd0960e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5752cd),
	.w1(32'h3b209835),
	.w2(32'hbd38cc36),
	.w3(32'h3b9c8140),
	.w4(32'hbb45d2f8),
	.w5(32'hbb50dc52),
	.w6(32'h3c2773ad),
	.w7(32'h3b154068),
	.w8(32'hbb4d15bc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e24f),
	.w1(32'hbba10d89),
	.w2(32'hbb2ab9a9),
	.w3(32'hbb8d85fe),
	.w4(32'hbbb6fa8b),
	.w5(32'h39eef713),
	.w6(32'h3c7fd0b2),
	.w7(32'hbbff7cb7),
	.w8(32'hbbb1b349),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24dfe6),
	.w1(32'hba33b60d),
	.w2(32'hbb3fe712),
	.w3(32'h3bec09f4),
	.w4(32'hbb30e0b6),
	.w5(32'hbbd36910),
	.w6(32'hbad10458),
	.w7(32'h3d4a541f),
	.w8(32'hbbd9c643),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba26705),
	.w1(32'hbad59609),
	.w2(32'hbb741dd5),
	.w3(32'h3c73e114),
	.w4(32'hbb2363af),
	.w5(32'hbb42d41e),
	.w6(32'h3c25c670),
	.w7(32'hbb009ca7),
	.w8(32'hbb44b9ae),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d28aa),
	.w1(32'h3ae17b70),
	.w2(32'hbc232d0b),
	.w3(32'h3c2bb9e3),
	.w4(32'h3ba54e23),
	.w5(32'hbc056418),
	.w6(32'hbb569231),
	.w7(32'h3b773111),
	.w8(32'h3c31dba0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46ea05),
	.w1(32'h3c830557),
	.w2(32'h3b4ec523),
	.w3(32'hbbd7e6a5),
	.w4(32'hbae88bcf),
	.w5(32'h3bed8705),
	.w6(32'h3bf6d366),
	.w7(32'h3ba05e37),
	.w8(32'h3c0eef54),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55f2ab),
	.w1(32'hbc01614e),
	.w2(32'h3ab8a7b9),
	.w3(32'hbad3d383),
	.w4(32'h3c05c262),
	.w5(32'hbbaf195a),
	.w6(32'hbb7ff148),
	.w7(32'h3c4985fc),
	.w8(32'h3ada75b8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc925cbf),
	.w1(32'hbc0b456f),
	.w2(32'hbb446c9d),
	.w3(32'hbb91f3f5),
	.w4(32'h3b7f4ad3),
	.w5(32'hbc0bdf7f),
	.w6(32'h3b9c4eeb),
	.w7(32'hba5b88c9),
	.w8(32'hbb059291),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca21d27),
	.w1(32'h3c4b5b94),
	.w2(32'hbc604cbf),
	.w3(32'hb8b7941f),
	.w4(32'hbbb9e75b),
	.w5(32'h3a836ac7),
	.w6(32'h3c241584),
	.w7(32'hbc1d5087),
	.w8(32'h3b0c14bc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb733d9b),
	.w1(32'hbbb73107),
	.w2(32'h3ad777e9),
	.w3(32'hbbb8c436),
	.w4(32'h3b96603e),
	.w5(32'h3c609a4a),
	.w6(32'hbbf7c0a0),
	.w7(32'hbc3a85b8),
	.w8(32'hbb722197),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae00578),
	.w1(32'hb9ca6752),
	.w2(32'h3b51cee6),
	.w3(32'h3a5fe469),
	.w4(32'h3c7039f4),
	.w5(32'hba001a9f),
	.w6(32'h3cd0b28a),
	.w7(32'h3c1019b5),
	.w8(32'hb9769f07),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf2c8),
	.w1(32'hba9a340e),
	.w2(32'h3c8ca1a5),
	.w3(32'hb9e2cdd1),
	.w4(32'h3b01343c),
	.w5(32'h3c0ab4cb),
	.w6(32'hbcfbe3b3),
	.w7(32'h3c5bb273),
	.w8(32'hbae6ba70),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6bfd3),
	.w1(32'h3b1920c6),
	.w2(32'h3cc600bd),
	.w3(32'hbc910460),
	.w4(32'hbac643ad),
	.w5(32'h3ae2fcac),
	.w6(32'h3c2281df),
	.w7(32'hbbaab642),
	.w8(32'hbad288a4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9269a28),
	.w1(32'hbbbfa224),
	.w2(32'h3b691c7e),
	.w3(32'hbbbfeb49),
	.w4(32'hba0edda6),
	.w5(32'hbbc7e70e),
	.w6(32'h3ba6e0d0),
	.w7(32'h3c9a7176),
	.w8(32'hbc7f3142),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d2f3f),
	.w1(32'h3b18cd2a),
	.w2(32'hbb021cf7),
	.w3(32'h3cb08aff),
	.w4(32'h3987a8c5),
	.w5(32'h3c16e014),
	.w6(32'h3b8f7f96),
	.w7(32'hbb2738c9),
	.w8(32'hbc7c7d39),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b602849),
	.w1(32'hbabc96a8),
	.w2(32'h3b8f4435),
	.w3(32'hba004106),
	.w4(32'h3becbb05),
	.w5(32'h3bb4b4ff),
	.w6(32'hbb82e079),
	.w7(32'hbac5ecc0),
	.w8(32'hbb8588a2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3754c4),
	.w1(32'hbb514b25),
	.w2(32'hba1f5aa0),
	.w3(32'hbb14fcb4),
	.w4(32'hbba1b6f2),
	.w5(32'h3cba196a),
	.w6(32'h3aaf1604),
	.w7(32'hbb548d72),
	.w8(32'hba656687),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd258c7),
	.w1(32'h3c2fe237),
	.w2(32'hbb04c85b),
	.w3(32'hbc0e3733),
	.w4(32'h3c07cecf),
	.w5(32'hbc2c3923),
	.w6(32'hbacd5913),
	.w7(32'hba602130),
	.w8(32'h390c560e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c406533),
	.w1(32'h3ba9e9aa),
	.w2(32'h3a98b1f7),
	.w3(32'hbbce3330),
	.w4(32'h3a5e0552),
	.w5(32'hbbc0896b),
	.w6(32'hbbaa34f3),
	.w7(32'hb7125172),
	.w8(32'h3bc10db2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95b7a0),
	.w1(32'h3aff942d),
	.w2(32'hbb8c536a),
	.w3(32'h3bc92866),
	.w4(32'h3c6d7c51),
	.w5(32'h3c28e2e7),
	.w6(32'hbb1f5da5),
	.w7(32'h3c403948),
	.w8(32'h3a0e7c5c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc8eca),
	.w1(32'hba0d02a6),
	.w2(32'h3cb4c8c7),
	.w3(32'h3c63f06b),
	.w4(32'hbb0a7e15),
	.w5(32'h3c86e95f),
	.w6(32'hbbd6bc08),
	.w7(32'hb74a466d),
	.w8(32'hbb1de6c0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13009b),
	.w1(32'h3bc75ffe),
	.w2(32'hbc827228),
	.w3(32'h3c9b81d9),
	.w4(32'hbb2cb3b1),
	.w5(32'hbcac93d2),
	.w6(32'hbd23be72),
	.w7(32'hbcd7edb0),
	.w8(32'hbba65ec2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd15f2f),
	.w1(32'h3b58c14c),
	.w2(32'hbc3e912a),
	.w3(32'hbba8b0c1),
	.w4(32'hbbe62bea),
	.w5(32'h37171bf7),
	.w6(32'hba0babc4),
	.w7(32'hbc1cb4fa),
	.w8(32'h3c126b33),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d093b80),
	.w1(32'h3ce94ae5),
	.w2(32'hbcc59b0f),
	.w3(32'h37d7c324),
	.w4(32'hbc3b9d64),
	.w5(32'h3c91d4fe),
	.w6(32'h3c6af323),
	.w7(32'hbd307cea),
	.w8(32'hbc396785),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd94e),
	.w1(32'hbd060014),
	.w2(32'hbba73878),
	.w3(32'hbd0516a6),
	.w4(32'hbce6f084),
	.w5(32'hbbd9a6de),
	.w6(32'hbaa067ac),
	.w7(32'h3c8f57f4),
	.w8(32'h3ceb66a0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44a6cb),
	.w1(32'hba919d8f),
	.w2(32'hbc2a44b0),
	.w3(32'hbb909092),
	.w4(32'h3c5194be),
	.w5(32'hbb5c8ed7),
	.w6(32'hbc3c3d7f),
	.w7(32'h3c365374),
	.w8(32'h3d2cce13),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0b4b),
	.w1(32'hbb2fe5f1),
	.w2(32'hbc3e9118),
	.w3(32'h3bff9512),
	.w4(32'hbc1706fa),
	.w5(32'hbc0774d3),
	.w6(32'hbd238886),
	.w7(32'hba82b8ba),
	.w8(32'hbc4b9d84),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1efad),
	.w1(32'h3d94b928),
	.w2(32'h3b5b73bf),
	.w3(32'hbc22c9c5),
	.w4(32'h3bf3e400),
	.w5(32'hbc554379),
	.w6(32'hbc2f038f),
	.w7(32'hbc7e3a11),
	.w8(32'hbca46fad),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01d94a),
	.w1(32'h3ac044c8),
	.w2(32'hbcac8e29),
	.w3(32'hbc3e7e68),
	.w4(32'hba2003c8),
	.w5(32'hbd1f96bb),
	.w6(32'hbc26ec52),
	.w7(32'hbb75778e),
	.w8(32'hbb3bf579),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc466235),
	.w1(32'hbc891b24),
	.w2(32'h3c81391c),
	.w3(32'h3d17f256),
	.w4(32'h3d672e5d),
	.w5(32'hbb4f96d6),
	.w6(32'hbc11e5ff),
	.w7(32'h3a9230f7),
	.w8(32'h3b2ca876),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c522f64),
	.w1(32'h3a871019),
	.w2(32'hbc905b6a),
	.w3(32'h3bb5b722),
	.w4(32'h39ad8cd2),
	.w5(32'hbb85d4cf),
	.w6(32'hbd177257),
	.w7(32'h3d622705),
	.w8(32'h379171ff),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a550519),
	.w1(32'hbbe9d7e4),
	.w2(32'h3a438f22),
	.w3(32'hb9d9ad8b),
	.w4(32'h3c147d36),
	.w5(32'h3c4348c0),
	.w6(32'hbc7168da),
	.w7(32'hbbde9448),
	.w8(32'hbaa7a606),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000ff1),
	.w1(32'hbcab189f),
	.w2(32'hbbd8f069),
	.w3(32'h3d37c052),
	.w4(32'hbc37e165),
	.w5(32'h3b571e25),
	.w6(32'h3c04cc58),
	.w7(32'hb9d09ef2),
	.w8(32'h3d1fe2cb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09453f),
	.w1(32'h3c6ae43a),
	.w2(32'hbb3de1aa),
	.w3(32'h3c267c93),
	.w4(32'hbba204fc),
	.w5(32'h3c7366a5),
	.w6(32'h3c663160),
	.w7(32'hbb2e9ee8),
	.w8(32'h3b32094b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b206384),
	.w1(32'h3c22ec0b),
	.w2(32'hbb37ff54),
	.w3(32'hbc3cacd7),
	.w4(32'hbc64d319),
	.w5(32'h3d1e2869),
	.w6(32'hbc943eb2),
	.w7(32'h3a1aa480),
	.w8(32'h383adfce),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e1cf3),
	.w1(32'hbaa0aff9),
	.w2(32'h3a83cb3b),
	.w3(32'hbacee435),
	.w4(32'h3b94d27a),
	.w5(32'hba4a36b3),
	.w6(32'hba167f6a),
	.w7(32'h3955f250),
	.w8(32'hbadbd740),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b19f2),
	.w1(32'h391794a6),
	.w2(32'hba9e6e3b),
	.w3(32'h39ecd114),
	.w4(32'h3c359f74),
	.w5(32'hb7946276),
	.w6(32'h3a4f762f),
	.w7(32'h3a5fd393),
	.w8(32'h3b8e74b2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f3b33),
	.w1(32'hba8a972f),
	.w2(32'h3b0b4570),
	.w3(32'h3b6811d2),
	.w4(32'hb8a03f2f),
	.w5(32'h3a69205c),
	.w6(32'h38b78ba4),
	.w7(32'h3b0a5a6b),
	.w8(32'hbac1b68e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a060638),
	.w1(32'hb7b5156a),
	.w2(32'hbbd4c755),
	.w3(32'h38c7cfd3),
	.w4(32'hba90b1b7),
	.w5(32'h3a0bb343),
	.w6(32'hba8c4aca),
	.w7(32'hbaaf1aca),
	.w8(32'hbb598bc1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb799f84),
	.w1(32'h3b4bcccd),
	.w2(32'h3a5b980f),
	.w3(32'hbab8d41e),
	.w4(32'h3a9a52b9),
	.w5(32'hba9afbd9),
	.w6(32'hba87de75),
	.w7(32'h39ff1802),
	.w8(32'hbab4c234),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a50c0),
	.w1(32'hbabeb8a1),
	.w2(32'h3b60aedd),
	.w3(32'hbb8cfc3c),
	.w4(32'h3b8a126f),
	.w5(32'h3a417892),
	.w6(32'hbb0fe6b8),
	.w7(32'h3ab3e885),
	.w8(32'h3a721351),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8320d1b),
	.w1(32'h3a1da39c),
	.w2(32'hba3f5887),
	.w3(32'hbb0523c2),
	.w4(32'hba4cbfaa),
	.w5(32'hb93752a8),
	.w6(32'h3a5cc6f7),
	.w7(32'hbb097323),
	.w8(32'h3a445a0a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa522f),
	.w1(32'h3bc22ee5),
	.w2(32'hbb2525ac),
	.w3(32'hba5f00f9),
	.w4(32'hbba7a220),
	.w5(32'hb9dccd26),
	.w6(32'hb9b5dcf2),
	.w7(32'hbac369b8),
	.w8(32'h3b43a2de),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b069677),
	.w1(32'h3bca3448),
	.w2(32'hba13233a),
	.w3(32'h3a7c3fbc),
	.w4(32'h3b197972),
	.w5(32'h3aa8822c),
	.w6(32'hba32e6bd),
	.w7(32'h3981cf28),
	.w8(32'hbbe4b765),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f91eb5),
	.w1(32'h3a62785f),
	.w2(32'h3a376452),
	.w3(32'h3b06768a),
	.w4(32'hbadf5ca7),
	.w5(32'hb88667f9),
	.w6(32'h3b38e4fb),
	.w7(32'hb7da746b),
	.w8(32'h3add14a5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba66ed),
	.w1(32'h39cb49ca),
	.w2(32'hb9d7c317),
	.w3(32'h39d391e9),
	.w4(32'hba04fb7b),
	.w5(32'hbb06e848),
	.w6(32'hbbcef951),
	.w7(32'hb9efe044),
	.w8(32'hba8cf0d5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f74c1e),
	.w1(32'hbae85038),
	.w2(32'h39f47568),
	.w3(32'h39b961f8),
	.w4(32'hbad7f1c0),
	.w5(32'hbaabd4f0),
	.w6(32'h38181c45),
	.w7(32'hbadafc0f),
	.w8(32'hba3218cf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8064f83),
	.w1(32'h3b1f91dc),
	.w2(32'hb9e77d4f),
	.w3(32'h3ab8d520),
	.w4(32'h3a0590f7),
	.w5(32'hba592391),
	.w6(32'hb9e6fb12),
	.w7(32'hba7fc268),
	.w8(32'hba9bf303),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1495be),
	.w1(32'h39b18ca8),
	.w2(32'h3a39b834),
	.w3(32'h3ae5d6b1),
	.w4(32'h3a84d8cd),
	.w5(32'h39eb8f45),
	.w6(32'hbad90594),
	.w7(32'hbbb5ab76),
	.w8(32'hb9a4c006),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c6d51),
	.w1(32'h3b00223c),
	.w2(32'hbd1709f4),
	.w3(32'hbaa29463),
	.w4(32'hba12fc56),
	.w5(32'h3b1b2148),
	.w6(32'hbbe29017),
	.w7(32'h3c8d2165),
	.w8(32'h3ba27fad),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c92bf),
	.w1(32'hbc2a449d),
	.w2(32'hbc0a7a9a),
	.w3(32'h3d5d4b88),
	.w4(32'hbc16bf4c),
	.w5(32'hbc66538a),
	.w6(32'hbc805c8a),
	.w7(32'hbb86376d),
	.w8(32'hbd08288f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2ed36),
	.w1(32'h3b943fdc),
	.w2(32'hbbc9808c),
	.w3(32'hbc71f60d),
	.w4(32'hbca21176),
	.w5(32'hbcc26f14),
	.w6(32'hbc90cab7),
	.w7(32'hbbb6bbe0),
	.w8(32'hbbd4a9c8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbb70d),
	.w1(32'hbb866825),
	.w2(32'h3cce9c5b),
	.w3(32'hbb87cb2a),
	.w4(32'h3cb4f19f),
	.w5(32'hbc2bac0f),
	.w6(32'h3c8ec0b0),
	.w7(32'hbc336958),
	.w8(32'hbc475557),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc25cbc),
	.w1(32'hbcce008f),
	.w2(32'h3bdb84b2),
	.w3(32'hbc4c6b56),
	.w4(32'h3b299481),
	.w5(32'h3a96c989),
	.w6(32'h3c3eeaa2),
	.w7(32'h3dc3c8bf),
	.w8(32'hbaa4c1dc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc042aac),
	.w1(32'hbc40214d),
	.w2(32'hbc88b125),
	.w3(32'h3bed8e5c),
	.w4(32'h3ba3172c),
	.w5(32'hbb23c5b6),
	.w6(32'hbb3609aa),
	.w7(32'h3ad5493f),
	.w8(32'h3b862210),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16f57c),
	.w1(32'hbba13c86),
	.w2(32'hbc034624),
	.w3(32'h3c9a89c9),
	.w4(32'hbba86a4e),
	.w5(32'hbb12c8d0),
	.w6(32'hbd2f967f),
	.w7(32'hbb3832c4),
	.w8(32'hbbb0ff3f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0de92e),
	.w1(32'hbb8ac372),
	.w2(32'hbc09cb0d),
	.w3(32'h3a3a7ebe),
	.w4(32'h3ca6d54a),
	.w5(32'hbbd76ce9),
	.w6(32'hbb8f6147),
	.w7(32'h3d27af7b),
	.w8(32'hbbb1d554),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a863e65),
	.w1(32'hbbeee103),
	.w2(32'h3cbf1d56),
	.w3(32'h3d115a2b),
	.w4(32'h3b30cca4),
	.w5(32'h3ce5334c),
	.w6(32'h3cc16dd1),
	.w7(32'hbc32bff4),
	.w8(32'hbc2602fc),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b502def),
	.w1(32'hba3b92b2),
	.w2(32'h3d26565f),
	.w3(32'hbb9779d4),
	.w4(32'h3c1ef04d),
	.w5(32'hbccd2b29),
	.w6(32'hba2678c4),
	.w7(32'hbc0accff),
	.w8(32'hbc301b6a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb388700),
	.w1(32'hbb3fc668),
	.w2(32'hbb8e9a80),
	.w3(32'hbc725fb5),
	.w4(32'h3d399cd0),
	.w5(32'h3d20076e),
	.w6(32'hbc89cd8f),
	.w7(32'hbb796b8d),
	.w8(32'hbc1d4304),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d198),
	.w1(32'hbae3e122),
	.w2(32'hbc2e705e),
	.w3(32'h3c310667),
	.w4(32'hbc4bd9b1),
	.w5(32'hbc037feb),
	.w6(32'hbce3da84),
	.w7(32'h3c39098c),
	.w8(32'hbc900eae),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca74cd6),
	.w1(32'h3a820bb7),
	.w2(32'h3c8c23da),
	.w3(32'hbc0cef10),
	.w4(32'hbc26b955),
	.w5(32'h3bc7716d),
	.w6(32'hbd02bc2d),
	.w7(32'h3b8e2e22),
	.w8(32'hbc46b083),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda6c7a),
	.w1(32'h3d60ad4d),
	.w2(32'hbc5db577),
	.w3(32'h3bf4d0f2),
	.w4(32'hbbd46c9f),
	.w5(32'h393b09f0),
	.w6(32'h3c35cf10),
	.w7(32'hbc4ff5c0),
	.w8(32'h3d22b490),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3556a),
	.w1(32'h3b64e129),
	.w2(32'h3c158cbe),
	.w3(32'hbc192203),
	.w4(32'h3c4a2bb4),
	.w5(32'hbc2dfeb0),
	.w6(32'hbc1d2871),
	.w7(32'hbc28532c),
	.w8(32'h3a1adbad),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6aac2),
	.w1(32'hbbb1faba),
	.w2(32'hbb4621aa),
	.w3(32'h3bdc6d02),
	.w4(32'hbcc4c29d),
	.w5(32'hbb830187),
	.w6(32'hbabce66c),
	.w7(32'hbc871b55),
	.w8(32'hbcd72faa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dac9f),
	.w1(32'h3c4040c2),
	.w2(32'h3aa3d7b4),
	.w3(32'h3c7f0c10),
	.w4(32'hbc5b3f98),
	.w5(32'h3bbc01a3),
	.w6(32'h3c8fb3da),
	.w7(32'hbc4e9b45),
	.w8(32'hbc3915e4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886f6f8),
	.w1(32'hbc031cf7),
	.w2(32'h3d06702c),
	.w3(32'hbc1e01f9),
	.w4(32'hbaeee8ff),
	.w5(32'h3c369bfd),
	.w6(32'h3c2283e7),
	.w7(32'h3b3a632c),
	.w8(32'hbbb6360b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcb1d8),
	.w1(32'h3cd1efe1),
	.w2(32'h396b3633),
	.w3(32'h3d193ce6),
	.w4(32'h3d120a47),
	.w5(32'hba8ecc1b),
	.w6(32'hbb272c4f),
	.w7(32'h3bc58615),
	.w8(32'h3b9460ba),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba668ff3),
	.w1(32'h3bd7f86b),
	.w2(32'h3c9fbc8d),
	.w3(32'h3bd00b11),
	.w4(32'h3d17bb98),
	.w5(32'hbb24c110),
	.w6(32'hbc0426bb),
	.w7(32'h3ccc2b71),
	.w8(32'h3c1c1916),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba266267),
	.w1(32'hbb4891ef),
	.w2(32'h3b8af9c3),
	.w3(32'h3c953209),
	.w4(32'hbbb71281),
	.w5(32'hbd435c8d),
	.w6(32'hbb6cbd20),
	.w7(32'h3c582ab6),
	.w8(32'hbbb3e21e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931bb7e),
	.w1(32'hba892e61),
	.w2(32'h3b83a6be),
	.w3(32'hbbc08e03),
	.w4(32'h3c8b0a05),
	.w5(32'hbb598dab),
	.w6(32'hbc3b6543),
	.w7(32'hbb8c7500),
	.w8(32'hbc112f60),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d89c0b2),
	.w1(32'hbc533393),
	.w2(32'h3a54ce12),
	.w3(32'h3d2352d6),
	.w4(32'hbb646ad8),
	.w5(32'hbb3f298f),
	.w6(32'h3accbe2c),
	.w7(32'hbb7d9f9c),
	.w8(32'hbb6e4fe9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04aa52),
	.w1(32'hbc0c4fa1),
	.w2(32'h3c6fd95f),
	.w3(32'hbb6bd940),
	.w4(32'h3cad5729),
	.w5(32'hbbc35f61),
	.w6(32'hbaa119ce),
	.w7(32'h3c45050d),
	.w8(32'hbbd51148),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee670b),
	.w1(32'h3c1ba876),
	.w2(32'h3d10fc31),
	.w3(32'h3be46426),
	.w4(32'hbc5f15df),
	.w5(32'hbade034f),
	.w6(32'h3c157ca2),
	.w7(32'hbaa93127),
	.w8(32'hbbe077ed),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2a7d8),
	.w1(32'h3c867b4a),
	.w2(32'hbacf5abb),
	.w3(32'h3c34a6cb),
	.w4(32'h3c458fd6),
	.w5(32'hbc2d5f20),
	.w6(32'h3c914db4),
	.w7(32'hbaadb025),
	.w8(32'hbc0b8483),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95e8a2),
	.w1(32'h36c38fc0),
	.w2(32'hbc0ec943),
	.w3(32'h386686a4),
	.w4(32'hbba28678),
	.w5(32'h3c6de998),
	.w6(32'hbba43daa),
	.w7(32'h3b072035),
	.w8(32'h3c3f7618),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2054ad),
	.w1(32'h3d3bbfa5),
	.w2(32'h3c9b758d),
	.w3(32'hbb980466),
	.w4(32'hbc263075),
	.w5(32'h3b924ab8),
	.w6(32'hbb521ec9),
	.w7(32'h3ba0f22d),
	.w8(32'hbb492e51),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392de270),
	.w1(32'h3b7c7392),
	.w2(32'hbb7dd942),
	.w3(32'hbc299d8e),
	.w4(32'h3c118d4f),
	.w5(32'h3ae3bef8),
	.w6(32'hba8288e3),
	.w7(32'h3d21b340),
	.w8(32'hba9e7477),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fdcd9),
	.w1(32'hbc035842),
	.w2(32'hbc3de8f3),
	.w3(32'h3aa488ab),
	.w4(32'h3c3b5afb),
	.w5(32'hbb374729),
	.w6(32'h3bf97e31),
	.w7(32'h3d750d30),
	.w8(32'h3adb5a34),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0999fc),
	.w1(32'hbab84253),
	.w2(32'hbb725cb8),
	.w3(32'hbc1a7d25),
	.w4(32'hbb0c6e04),
	.w5(32'h3ba246f4),
	.w6(32'h3d1cf7f3),
	.w7(32'hba9c90e5),
	.w8(32'hbbabb42c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cacb982),
	.w1(32'hbc8ed027),
	.w2(32'hbcda79dc),
	.w3(32'hbc509575),
	.w4(32'hbd00ae28),
	.w5(32'h3b73ff6e),
	.w6(32'hbd2fc103),
	.w7(32'hbb83f9c8),
	.w8(32'h3b52929e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87a48c),
	.w1(32'h3b95a7e0),
	.w2(32'hbca213ab),
	.w3(32'h3be939f5),
	.w4(32'hbbc921f2),
	.w5(32'h3bdf2d1e),
	.w6(32'hbbd45f11),
	.w7(32'h3c07a1c5),
	.w8(32'h39f77658),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d225d8a),
	.w1(32'h3cb2c572),
	.w2(32'h3a3f6b30),
	.w3(32'h3c7a61e0),
	.w4(32'hbc28683a),
	.w5(32'h3b18a2e8),
	.w6(32'h3a1301cb),
	.w7(32'h3ba02e12),
	.w8(32'hbb1c1a81),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122cee),
	.w1(32'hbc0f4fdc),
	.w2(32'hbc75285d),
	.w3(32'h3c6d3ace),
	.w4(32'hbc35d510),
	.w5(32'hbb98ff84),
	.w6(32'hbba50145),
	.w7(32'hbc906f1d),
	.w8(32'hbb284bca),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb866c0c),
	.w1(32'hbc51cdf7),
	.w2(32'h3b65e354),
	.w3(32'hbb8a80eb),
	.w4(32'hb9a6da37),
	.w5(32'hbbb0ead9),
	.w6(32'hbc004f51),
	.w7(32'h341f2b26),
	.w8(32'h3d138bc4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e0256),
	.w1(32'hbb63f0fe),
	.w2(32'hbc90b075),
	.w3(32'h3c29334d),
	.w4(32'hbba2a488),
	.w5(32'h3b11edbb),
	.w6(32'hbb136630),
	.w7(32'h3c955ffc),
	.w8(32'h3ce47d42),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0a03f),
	.w1(32'hbc723a6c),
	.w2(32'hb7dcad67),
	.w3(32'hbc2744c6),
	.w4(32'h3ae6f09c),
	.w5(32'hbbcb88f4),
	.w6(32'hbc95413a),
	.w7(32'hbad04f7a),
	.w8(32'h3c8e01fc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cb9aa),
	.w1(32'h3b863b13),
	.w2(32'h3bf2202b),
	.w3(32'h3bfbf68b),
	.w4(32'hbc328467),
	.w5(32'hba1b2cc2),
	.w6(32'hbc879fb9),
	.w7(32'h3bb74daf),
	.w8(32'h3c9fb4f6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba616e19),
	.w1(32'hbc52d28d),
	.w2(32'hbca2d47c),
	.w3(32'hbc83fcbc),
	.w4(32'h3b75c48a),
	.w5(32'hb9ca0658),
	.w6(32'h3b279d07),
	.w7(32'h398e61b2),
	.w8(32'hbcbf0642),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8ad66),
	.w1(32'hbb35bf71),
	.w2(32'h3bf1b0cb),
	.w3(32'hbc36e629),
	.w4(32'h3d854793),
	.w5(32'hbb8f1207),
	.w6(32'hbcd7124a),
	.w7(32'hbca6b05f),
	.w8(32'hbb3ab7fd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb61105),
	.w1(32'h3aa07d6a),
	.w2(32'h3caefdb5),
	.w3(32'h3cce5a7a),
	.w4(32'hbbe99ab9),
	.w5(32'hbbca9b38),
	.w6(32'h3ccc6325),
	.w7(32'hbc177de7),
	.w8(32'hbb2ac23d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45613b),
	.w1(32'h3ca13e59),
	.w2(32'hbbe11ac6),
	.w3(32'h3c64dfa1),
	.w4(32'h3836e7a4),
	.w5(32'hbc2d4a36),
	.w6(32'h3c0f690e),
	.w7(32'hbb9d9841),
	.w8(32'h3c95434d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c915d84),
	.w1(32'hbb28f520),
	.w2(32'h3c9923bd),
	.w3(32'hbcb5a96a),
	.w4(32'hbc7f4911),
	.w5(32'hbc3929e8),
	.w6(32'hbbcb38ed),
	.w7(32'h3807cb12),
	.w8(32'h3b13fc46),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0526c7),
	.w1(32'h3aac03f4),
	.w2(32'h3b6c656a),
	.w3(32'hbc188cb4),
	.w4(32'hbc8293ee),
	.w5(32'h3cc0643f),
	.w6(32'hbc80a504),
	.w7(32'hbc05f1ed),
	.w8(32'h3b4a8be3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule