module layer_10_featuremap_277(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43bd58),
	.w1(32'h3c25b2f5),
	.w2(32'h3be1f05f),
	.w3(32'h3bb60fb2),
	.w4(32'h3c107982),
	.w5(32'hbc2dc8ed),
	.w6(32'h3bbe3ed8),
	.w7(32'h3c0b2a42),
	.w8(32'hbbbccc85),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39baf2e7),
	.w1(32'hbb5bdc78),
	.w2(32'hbc3d66e0),
	.w3(32'hbaf59cbe),
	.w4(32'hbbefac5c),
	.w5(32'hbb30b0cb),
	.w6(32'hbbb42d27),
	.w7(32'hbc449449),
	.w8(32'hbbd64cce),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b341ed2),
	.w1(32'h3b74fc46),
	.w2(32'hbba38bcd),
	.w3(32'hbb40412f),
	.w4(32'h3b28b73a),
	.w5(32'hbbd25479),
	.w6(32'h3c0b67ab),
	.w7(32'hbbc46bb0),
	.w8(32'hbc1d3466),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6e413),
	.w1(32'hbb96693f),
	.w2(32'hbbe385f6),
	.w3(32'hbc09800f),
	.w4(32'hbbf5830d),
	.w5(32'h3b0987c2),
	.w6(32'hbbc0b94a),
	.w7(32'hbc17f3f0),
	.w8(32'hbaec34de),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed8277),
	.w1(32'hbb205ad1),
	.w2(32'h3b58bc53),
	.w3(32'hbaa45708),
	.w4(32'h3b27aa0a),
	.w5(32'h3b9e9be0),
	.w6(32'hbbbf9049),
	.w7(32'hbc06a439),
	.w8(32'hba3dbd72),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b951e6),
	.w1(32'hba81a7d8),
	.w2(32'h3a8d37d7),
	.w3(32'h3a779df0),
	.w4(32'hba8f21a9),
	.w5(32'hba2e99d4),
	.w6(32'hbb8883c1),
	.w7(32'hbb60c37b),
	.w8(32'hbbc8761f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb62a44),
	.w1(32'hbbc96846),
	.w2(32'hbb64b472),
	.w3(32'hba124506),
	.w4(32'hbbd556b4),
	.w5(32'h3c20f7b1),
	.w6(32'hbb6ff738),
	.w7(32'hbb7bdd79),
	.w8(32'h3c83d941),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb96c9a),
	.w1(32'h3cd3ba34),
	.w2(32'h3bcd33e0),
	.w3(32'h3c88e407),
	.w4(32'h3cab117e),
	.w5(32'h3ba36142),
	.w6(32'h3d2f51f3),
	.w7(32'h3c87117f),
	.w8(32'hbb14a690),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a146347),
	.w1(32'hbb3743aa),
	.w2(32'h3abdcf96),
	.w3(32'hbb2c9744),
	.w4(32'hbab36444),
	.w5(32'h3acf89f3),
	.w6(32'hbbad4877),
	.w7(32'hba52cda8),
	.w8(32'hba8a450b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb290e30),
	.w1(32'hbabc7ae6),
	.w2(32'hbae5c545),
	.w3(32'hbb41d3aa),
	.w4(32'hbad0db1f),
	.w5(32'hbb10e792),
	.w6(32'hbbc04870),
	.w7(32'hbbc4ef58),
	.w8(32'hbc3dbd76),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6ddaa),
	.w1(32'h3983e48f),
	.w2(32'hbb2e464f),
	.w3(32'hbbb648aa),
	.w4(32'hbb2c2801),
	.w5(32'hb8f457b4),
	.w6(32'hba919db7),
	.w7(32'hbb0b8af8),
	.w8(32'h3acae5bb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1ddb3),
	.w1(32'h3c551549),
	.w2(32'h3b5d5b49),
	.w3(32'h3be466de),
	.w4(32'h3bdf04b5),
	.w5(32'hb9df0615),
	.w6(32'h3c1e15d3),
	.w7(32'h3bdace92),
	.w8(32'h3c09cafb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6d74e),
	.w1(32'h3c244ec8),
	.w2(32'h3c217e51),
	.w3(32'h3bb5b685),
	.w4(32'h3c1ebfb6),
	.w5(32'hbb8421d5),
	.w6(32'h3c07310c),
	.w7(32'h3b54fa0f),
	.w8(32'hbb002945),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96935a),
	.w1(32'hbb406a05),
	.w2(32'h3b1a2477),
	.w3(32'h3a465ebd),
	.w4(32'h3b12f79d),
	.w5(32'hbc0881ee),
	.w6(32'hbb8b519e),
	.w7(32'h3b055fee),
	.w8(32'hbc60ee73),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ac757),
	.w1(32'hbc2fa7cc),
	.w2(32'hbbb761a8),
	.w3(32'hbc3387a3),
	.w4(32'hbc1b6846),
	.w5(32'hbabc9999),
	.w6(32'hbc83281a),
	.w7(32'hbc31f949),
	.w8(32'hbb1bf08f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23dd9d),
	.w1(32'hbb2e3344),
	.w2(32'h3af49043),
	.w3(32'hbb769371),
	.w4(32'hbc0e3afa),
	.w5(32'h3b9c1b0a),
	.w6(32'hbc1ebf00),
	.w7(32'hbb6b14b3),
	.w8(32'hbb07d225),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d47c2d),
	.w1(32'hbacb433e),
	.w2(32'h3bb4ae52),
	.w3(32'h3bfe541d),
	.w4(32'h3a2b5b94),
	.w5(32'h3b833172),
	.w6(32'h3a29d46f),
	.w7(32'hba8ffa55),
	.w8(32'h3b386c2b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2084),
	.w1(32'h3a044f92),
	.w2(32'h3a8605f1),
	.w3(32'hbbc81902),
	.w4(32'hbb7428b3),
	.w5(32'hbb314a7a),
	.w6(32'hbb91684c),
	.w7(32'hbb704cf6),
	.w8(32'hbbaaaaec),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc176498),
	.w1(32'hbc038c8c),
	.w2(32'hbbadbf00),
	.w3(32'hbb9e6dfe),
	.w4(32'hb7d9cf50),
	.w5(32'hba5b7bba),
	.w6(32'hba1eee55),
	.w7(32'hbb3a2fa6),
	.w8(32'hbbd8ba5a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0fbd4),
	.w1(32'hbb1835a1),
	.w2(32'h3bd0420d),
	.w3(32'h3ac2ca44),
	.w4(32'h3b9bb70e),
	.w5(32'hbbc2f300),
	.w6(32'hbc927946),
	.w7(32'hbab80dcd),
	.w8(32'hbb202088),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9d003),
	.w1(32'hbbe7ff3d),
	.w2(32'hbb1d2704),
	.w3(32'hbbe82fb6),
	.w4(32'hbb97b267),
	.w5(32'h39dbfe8b),
	.w6(32'hbc6b52e8),
	.w7(32'hbb775952),
	.w8(32'hbb0e426c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb093ac5),
	.w1(32'h3aae693a),
	.w2(32'h39b9a862),
	.w3(32'h3a3ed985),
	.w4(32'hbadb6c4e),
	.w5(32'h3adb09e4),
	.w6(32'h3abed15f),
	.w7(32'hbad5f682),
	.w8(32'hbab79d5d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb92d49),
	.w1(32'h3b0e6fca),
	.w2(32'hba3e8ea9),
	.w3(32'hbb78c29e),
	.w4(32'hbb9ce03f),
	.w5(32'hbbbb0883),
	.w6(32'hbbdf433a),
	.w7(32'hbac61768),
	.w8(32'hbb982ca4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac55003),
	.w1(32'hbad424fe),
	.w2(32'hbbd34d60),
	.w3(32'hbae3bdcf),
	.w4(32'hbaee2419),
	.w5(32'hbb971ae5),
	.w6(32'h3bd94139),
	.w7(32'hbaccc014),
	.w8(32'hba445b9f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46ee68),
	.w1(32'hbaf12269),
	.w2(32'hbb27befc),
	.w3(32'hba5ed201),
	.w4(32'h3b1893ce),
	.w5(32'hbb165af1),
	.w6(32'h3b76c524),
	.w7(32'hbb05356a),
	.w8(32'hbc2fd65e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc519415),
	.w1(32'hbc143702),
	.w2(32'h3ac945f9),
	.w3(32'hbb97226b),
	.w4(32'hbc1cbde5),
	.w5(32'h3b293d1b),
	.w6(32'hbc0ade12),
	.w7(32'hbb348475),
	.w8(32'h3adb21ec),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb869d),
	.w1(32'h3b3d4d62),
	.w2(32'h3b4e653b),
	.w3(32'hb9bcae30),
	.w4(32'h3a73da32),
	.w5(32'h3c0b4fc9),
	.w6(32'h3b5194bb),
	.w7(32'h3b429fbb),
	.w8(32'h3b8e2eca),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdda029),
	.w1(32'hbaf9b9d3),
	.w2(32'h3b99f154),
	.w3(32'hbad99028),
	.w4(32'h3b3e36d1),
	.w5(32'h39bb8114),
	.w6(32'hbc5feb00),
	.w7(32'hbb920f25),
	.w8(32'hb9fe65b4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eb390),
	.w1(32'h3b0894b6),
	.w2(32'h3b5b5045),
	.w3(32'hbb4a95dd),
	.w4(32'h3ab7e45c),
	.w5(32'h37fef1d9),
	.w6(32'hbbe23cf6),
	.w7(32'h3a8c7bdb),
	.w8(32'h3b31381c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b2ea),
	.w1(32'hbb61621a),
	.w2(32'hbbabc112),
	.w3(32'h3b1fb92c),
	.w4(32'h3aba52f1),
	.w5(32'hbb82cee0),
	.w6(32'hba6d2aff),
	.w7(32'hbad6eea4),
	.w8(32'h3b9c1c77),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad79f09),
	.w1(32'hbb811b4a),
	.w2(32'h3b80e3fe),
	.w3(32'h3c072afe),
	.w4(32'hb92e23ac),
	.w5(32'h3a555ebf),
	.w6(32'h3be4a3c7),
	.w7(32'hbc085c94),
	.w8(32'hbc1c1a08),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a610567),
	.w1(32'hb9d61cdd),
	.w2(32'h3b70d983),
	.w3(32'hbaceed4b),
	.w4(32'hbb3ac91a),
	.w5(32'hbb9e5702),
	.w6(32'hbc49e584),
	.w7(32'hbbc9fa81),
	.w8(32'hbb4ccc4a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ff176),
	.w1(32'hbbb47351),
	.w2(32'h3bc731a0),
	.w3(32'hba293a70),
	.w4(32'h3b3287bd),
	.w5(32'h3bce0bee),
	.w6(32'h3c46c0bd),
	.w7(32'h3aa17284),
	.w8(32'h3bbb6ba3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca6f3),
	.w1(32'hbb2ef0ad),
	.w2(32'hbae35d00),
	.w3(32'h3a0ad8c6),
	.w4(32'h3a60b71d),
	.w5(32'h3b7370f7),
	.w6(32'hbb771116),
	.w7(32'h3b327722),
	.w8(32'h3b0f3fb1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd8083),
	.w1(32'hbb32af07),
	.w2(32'h3bb4a59c),
	.w3(32'hbb814c2e),
	.w4(32'h3ac37972),
	.w5(32'hbbc6aa92),
	.w6(32'hbc5d0686),
	.w7(32'h3af19c7f),
	.w8(32'hbb62c86c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf7061),
	.w1(32'hbbaf0ce3),
	.w2(32'hba39b2d9),
	.w3(32'hbbbdceef),
	.w4(32'hbab8ccd8),
	.w5(32'hbbbd4116),
	.w6(32'h39fa4326),
	.w7(32'h3b0d7535),
	.w8(32'h38802796),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b019c),
	.w1(32'hbb819678),
	.w2(32'h3a341acd),
	.w3(32'hbb1dd041),
	.w4(32'h3b4993ca),
	.w5(32'h3bc4d211),
	.w6(32'hbbcd015a),
	.w7(32'hbc16c22f),
	.w8(32'hbb4184ef),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfd530),
	.w1(32'hba93c2bf),
	.w2(32'h3b589de3),
	.w3(32'h39bf9d7a),
	.w4(32'hbbb6ad88),
	.w5(32'h3b67ee1f),
	.w6(32'hbadde4fd),
	.w7(32'h3aa4bb2a),
	.w8(32'h3b4fe8c8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0eb11),
	.w1(32'h3c04a3ad),
	.w2(32'hbb6d3090),
	.w3(32'h3ab65c6f),
	.w4(32'h3bc5e207),
	.w5(32'hbb2183e5),
	.w6(32'h3a87173a),
	.w7(32'hb95782bc),
	.w8(32'hbafe917f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e4eda),
	.w1(32'h3b653c98),
	.w2(32'hbbd21629),
	.w3(32'h3b71b2cf),
	.w4(32'hbc707bbb),
	.w5(32'hba759625),
	.w6(32'h3a5d2991),
	.w7(32'hbb7e3f15),
	.w8(32'hbaae3074),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9431341),
	.w1(32'h3b7f543f),
	.w2(32'h3af0d5db),
	.w3(32'hbbc8ea13),
	.w4(32'hbbcefb0f),
	.w5(32'h3b166c3a),
	.w6(32'hbb7a2cbd),
	.w7(32'h3c043770),
	.w8(32'hbb62a3ba),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb416518),
	.w1(32'hbb14d33f),
	.w2(32'h3a2b9cc7),
	.w3(32'hb8ea68fe),
	.w4(32'hb92b0006),
	.w5(32'hba765c4a),
	.w6(32'hba6f2c8b),
	.w7(32'hbacae736),
	.w8(32'hb9722730),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaadb10),
	.w1(32'hba82fdef),
	.w2(32'hbbc1e4bd),
	.w3(32'hbc0be878),
	.w4(32'hbc23e9fe),
	.w5(32'h3b18e837),
	.w6(32'hbbc287fd),
	.w7(32'hbaa0a6b2),
	.w8(32'hbb1b698a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23c255),
	.w1(32'hbb9064bb),
	.w2(32'hbbea1506),
	.w3(32'hbc220776),
	.w4(32'hbbb29476),
	.w5(32'hbc425df7),
	.w6(32'hbbd7440f),
	.w7(32'hbbbda836),
	.w8(32'hbc404799),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeecc30),
	.w1(32'hbba376b7),
	.w2(32'hbc030685),
	.w3(32'hbbff0c96),
	.w4(32'hbbd5cbbb),
	.w5(32'hba6cedbe),
	.w6(32'hbc1f14be),
	.w7(32'hbbf1d730),
	.w8(32'hbb83cce3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb431209),
	.w1(32'hbb291ada),
	.w2(32'hbb8f6a47),
	.w3(32'h3b425c94),
	.w4(32'h3b8936ba),
	.w5(32'hbbfad3c9),
	.w6(32'hb99c83bf),
	.w7(32'hbbc7226b),
	.w8(32'hbbc4870c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbced2c5),
	.w1(32'hbb46740f),
	.w2(32'hbbb3fae0),
	.w3(32'hbbc917f8),
	.w4(32'hba2cac22),
	.w5(32'h3b746f90),
	.w6(32'hbaf01001),
	.w7(32'hbbb6f7e3),
	.w8(32'hba7d97c1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390953fb),
	.w1(32'h3ad66edb),
	.w2(32'h3b156c0e),
	.w3(32'hb982c3a3),
	.w4(32'hbbc31b81),
	.w5(32'h3a28b0d9),
	.w6(32'hbab96a08),
	.w7(32'hbbb70dc0),
	.w8(32'h3bc29db9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c423f4c),
	.w1(32'h3c1a4cc8),
	.w2(32'h3ae11f41),
	.w3(32'h3bb95116),
	.w4(32'h3c34d474),
	.w5(32'hb9ecd6f8),
	.w6(32'h3c2b6920),
	.w7(32'h3b3b6841),
	.w8(32'hbbb72a5f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901826),
	.w1(32'hbb415843),
	.w2(32'hba8a0134),
	.w3(32'hbabccefa),
	.w4(32'hbb563676),
	.w5(32'hba697163),
	.w6(32'hbc05fa88),
	.w7(32'hbb968ef5),
	.w8(32'h3a5fad1f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f457),
	.w1(32'hbc568233),
	.w2(32'hba626630),
	.w3(32'hbb88361d),
	.w4(32'h3828ef27),
	.w5(32'hbaf71693),
	.w6(32'hbb45ca40),
	.w7(32'hbb1b5737),
	.w8(32'h394aac7f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80cd74),
	.w1(32'h3b7c15db),
	.w2(32'hbb13549e),
	.w3(32'hbbad400c),
	.w4(32'hbaa57292),
	.w5(32'hbba22519),
	.w6(32'hbbc2f2a1),
	.w7(32'hbba1010b),
	.w8(32'hbbd3f9f4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81d68f),
	.w1(32'h3ace4da3),
	.w2(32'hbb82ba71),
	.w3(32'hbba9eb69),
	.w4(32'h3aed0526),
	.w5(32'h3c100c92),
	.w6(32'h3b537608),
	.w7(32'h3b63a16d),
	.w8(32'h3bdbd413),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0de9bf),
	.w1(32'hbb93e656),
	.w2(32'hbbd32d3b),
	.w3(32'hbaa1edf8),
	.w4(32'h3b648093),
	.w5(32'h3b711dfb),
	.w6(32'hbb4a73e7),
	.w7(32'h3b2f8f66),
	.w8(32'hbbb4e999),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86dc32),
	.w1(32'h3b771a32),
	.w2(32'h3b8df11a),
	.w3(32'h3a896e0a),
	.w4(32'hba7529a4),
	.w5(32'h3a5e52c7),
	.w6(32'hbc38664b),
	.w7(32'hbaa465d5),
	.w8(32'hbae4ad87),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24832f),
	.w1(32'hbb213095),
	.w2(32'h3b53161c),
	.w3(32'hbb59e5be),
	.w4(32'h3ad583ad),
	.w5(32'hb78e8214),
	.w6(32'hbc909ccf),
	.w7(32'hbb586f17),
	.w8(32'hbaf00ad7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18bace),
	.w1(32'hbb2dd934),
	.w2(32'h3be7b19b),
	.w3(32'hbb888671),
	.w4(32'h397e47a5),
	.w5(32'hbb78a4e5),
	.w6(32'hbc100f8c),
	.w7(32'h3bbd45cb),
	.w8(32'hba8a5657),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64925f),
	.w1(32'hba043752),
	.w2(32'hbb9c85ea),
	.w3(32'hbad8f2d8),
	.w4(32'hb92bfb0b),
	.w5(32'h3bb0884e),
	.w6(32'h3b875f54),
	.w7(32'h3aa604ad),
	.w8(32'hbb8958d8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77cd82),
	.w1(32'hbb630916),
	.w2(32'h3af6a100),
	.w3(32'h39522e89),
	.w4(32'hbacd4794),
	.w5(32'h3bb3787e),
	.w6(32'hbc24db9f),
	.w7(32'hba517f2b),
	.w8(32'h3b4c8ea1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff1e5a),
	.w1(32'h3bdd9989),
	.w2(32'h3b7bb6a8),
	.w3(32'h3c100992),
	.w4(32'h3adb7ad5),
	.w5(32'h3a565d77),
	.w6(32'h3be47ef5),
	.w7(32'h3beaada4),
	.w8(32'hbbb16a72),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0af0cf),
	.w1(32'h3aed3d0c),
	.w2(32'hb9f37877),
	.w3(32'hbbcd7506),
	.w4(32'hbaffa244),
	.w5(32'hbc0eade9),
	.w6(32'hbc4eaefd),
	.w7(32'hbb9b9c6b),
	.w8(32'hbc2b3d86),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc168c15),
	.w1(32'hbc428319),
	.w2(32'hbbf04d44),
	.w3(32'hbbedb24a),
	.w4(32'hbbc52b83),
	.w5(32'h3ad394e4),
	.w6(32'hbc30e5de),
	.w7(32'hbc0205a6),
	.w8(32'hbb9b8235),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f03dc),
	.w1(32'h3b36f32d),
	.w2(32'hb778e319),
	.w3(32'hba24773b),
	.w4(32'hba3afede),
	.w5(32'h3abab2fa),
	.w6(32'hbbea1455),
	.w7(32'hbb61c9fa),
	.w8(32'h3b9020bd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa695c6),
	.w1(32'hbb752810),
	.w2(32'h3b67d791),
	.w3(32'hbba03513),
	.w4(32'h3988d61c),
	.w5(32'h3b2e860c),
	.w6(32'hbc2a9f4e),
	.w7(32'h3bcaf018),
	.w8(32'hbb6a7231),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b821436),
	.w1(32'hbb473ea8),
	.w2(32'h3b084177),
	.w3(32'hbb7d21d2),
	.w4(32'hbb78bab9),
	.w5(32'h3b546ab1),
	.w6(32'hbc660d56),
	.w7(32'hbb372f75),
	.w8(32'hbbe025f7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c088a),
	.w1(32'h3c4d9f97),
	.w2(32'h3b422415),
	.w3(32'h39dda108),
	.w4(32'h3a26963b),
	.w5(32'h3a644725),
	.w6(32'hbbb2b854),
	.w7(32'h3ab7f3af),
	.w8(32'hbbd208da),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b7612),
	.w1(32'h3c0057ef),
	.w2(32'h3a175c95),
	.w3(32'hbb478151),
	.w4(32'h3b6e5cec),
	.w5(32'h3bd67a96),
	.w6(32'h3b7be87f),
	.w7(32'h3a48ce83),
	.w8(32'h3bf824b0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d3569e),
	.w1(32'hbabb4167),
	.w2(32'h39d20a84),
	.w3(32'h3a9935f5),
	.w4(32'h3b6f1a19),
	.w5(32'hbb21336f),
	.w6(32'h3bad00c1),
	.w7(32'h3b7f063c),
	.w8(32'hbb6592d3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc7bbd),
	.w1(32'hbbf2410b),
	.w2(32'hba8f72a9),
	.w3(32'h3a39bd22),
	.w4(32'h3bbd6eb8),
	.w5(32'hbbae865d),
	.w6(32'hbbb09f8e),
	.w7(32'h3ba0c5fd),
	.w8(32'hbbe99834),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a0c1c),
	.w1(32'hbc39729a),
	.w2(32'hbc294eab),
	.w3(32'hbc094ec3),
	.w4(32'hbb746b26),
	.w5(32'hba6fea82),
	.w6(32'h3912907e),
	.w7(32'hbb40c2ce),
	.w8(32'hbb6f21db),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997131c),
	.w1(32'hba300999),
	.w2(32'h3ac4aa68),
	.w3(32'hbb5575d1),
	.w4(32'hba7d17a2),
	.w5(32'h3a89611d),
	.w6(32'h3a1d04cc),
	.w7(32'hba32d068),
	.w8(32'hbb12395c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d3fd1),
	.w1(32'h3c1c7322),
	.w2(32'h3b811b3c),
	.w3(32'h3c1d7069),
	.w4(32'h3b94f66a),
	.w5(32'h3b3d1a26),
	.w6(32'h3c873cfe),
	.w7(32'h3c0bcdaa),
	.w8(32'h3c28af0c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac774a2),
	.w1(32'h3abb223e),
	.w2(32'hbb815094),
	.w3(32'hbace241f),
	.w4(32'hb930df2c),
	.w5(32'hbb92cada),
	.w6(32'h3b86d3c1),
	.w7(32'hbb149146),
	.w8(32'hba7e254c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf6fa6),
	.w1(32'hbb20812f),
	.w2(32'hbbdab564),
	.w3(32'hbaec1676),
	.w4(32'h3a499285),
	.w5(32'h3b91c025),
	.w6(32'hbc12df18),
	.w7(32'hba89727d),
	.w8(32'hbbd8b3d3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba3d8c),
	.w1(32'h3be23673),
	.w2(32'h3ba58f82),
	.w3(32'hbb98b9cf),
	.w4(32'hbb76ea72),
	.w5(32'h3aca02c7),
	.w6(32'hbb849b67),
	.w7(32'h3b5b8ca2),
	.w8(32'h3bd011b2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bc351),
	.w1(32'h3ac58dfb),
	.w2(32'hba7ff278),
	.w3(32'h3b4b38a6),
	.w4(32'h3ba2692c),
	.w5(32'h3b3f1d94),
	.w6(32'h3a9b3f47),
	.w7(32'h3b9cdcb5),
	.w8(32'h3a06019e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb708343),
	.w1(32'h3b85c076),
	.w2(32'hba151bac),
	.w3(32'hbbd80be6),
	.w4(32'hbb530978),
	.w5(32'hbc333ad3),
	.w6(32'h3ad5f2ba),
	.w7(32'h3bd0212f),
	.w8(32'hbbdf5438),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47ddea),
	.w1(32'hbbc51258),
	.w2(32'hbbf6af37),
	.w3(32'hbc3a7fd1),
	.w4(32'hbc23a37a),
	.w5(32'h3b22417c),
	.w6(32'hbbeccb43),
	.w7(32'hbc2c7469),
	.w8(32'hbb188442),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aa2aa),
	.w1(32'h3af6c948),
	.w2(32'hb9268941),
	.w3(32'h3c1851ae),
	.w4(32'h3c5d3629),
	.w5(32'h3b5b9d09),
	.w6(32'h3bfb91b3),
	.w7(32'hb941f3b8),
	.w8(32'hbb0abaf3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202d41),
	.w1(32'hbaac931d),
	.w2(32'h3b6a46dc),
	.w3(32'hba106e02),
	.w4(32'h3a497e7d),
	.w5(32'h3bcbb34b),
	.w6(32'hbb53e949),
	.w7(32'hbbf02225),
	.w8(32'h3b835d01),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e105f),
	.w1(32'h3bbf486a),
	.w2(32'h3b4d42d1),
	.w3(32'h3c19b0ba),
	.w4(32'h3c4cbac8),
	.w5(32'h3a441363),
	.w6(32'h3a184146),
	.w7(32'h3c177335),
	.w8(32'h3b9151ae),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a488d10),
	.w1(32'hba3e18fe),
	.w2(32'h3af81274),
	.w3(32'hba9d117a),
	.w4(32'h3b539150),
	.w5(32'hbad55937),
	.w6(32'h3a856969),
	.w7(32'h3b3f34d3),
	.w8(32'hbaf9a952),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2add58),
	.w1(32'hbbb858d4),
	.w2(32'hbb9139e3),
	.w3(32'h3b183843),
	.w4(32'h3a2f4089),
	.w5(32'h37da0a20),
	.w6(32'h3bac5c52),
	.w7(32'hbb44478b),
	.w8(32'h3c243c90),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d8d5),
	.w1(32'h3c445e1a),
	.w2(32'h3c74ebe4),
	.w3(32'h3c4be8cf),
	.w4(32'h3bff339b),
	.w5(32'h3adceb8c),
	.w6(32'h3c9d79c0),
	.w7(32'h3c8f6565),
	.w8(32'h3b13564f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb192b0b),
	.w1(32'h3b930dc7),
	.w2(32'h3b82716e),
	.w3(32'h3abf8cd6),
	.w4(32'hbb5fea4a),
	.w5(32'hba138001),
	.w6(32'h39f8edba),
	.w7(32'hbb4c729f),
	.w8(32'hbbdd56fc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0054ac),
	.w1(32'hbb949150),
	.w2(32'hbae5e7af),
	.w3(32'hbb63c91e),
	.w4(32'h3a1890da),
	.w5(32'h38f60755),
	.w6(32'hbbab3161),
	.w7(32'hbb64d61b),
	.w8(32'hbb2cb4b6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcbd04),
	.w1(32'hbc0cf41c),
	.w2(32'hbc3b77ca),
	.w3(32'hbbdafaf3),
	.w4(32'hbb6fe8d8),
	.w5(32'h3bc4ad5b),
	.w6(32'hbaff8531),
	.w7(32'hbc33745e),
	.w8(32'hba8d3afe),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66d261),
	.w1(32'h3b9b1339),
	.w2(32'h3b3695ea),
	.w3(32'h3b07fe83),
	.w4(32'h3b386824),
	.w5(32'h3a9e20b5),
	.w6(32'hbc2f8eb2),
	.w7(32'hbb9be7de),
	.w8(32'hbbd2ccf2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe71c12),
	.w1(32'hbc09bc7b),
	.w2(32'hb88830dd),
	.w3(32'hbb6150d5),
	.w4(32'hbbd25d6f),
	.w5(32'h3b6b93da),
	.w6(32'hbc1b3b16),
	.w7(32'hbbdf8a4a),
	.w8(32'h3a906a5f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa07bf3),
	.w1(32'hba56da7f),
	.w2(32'h3b6c7663),
	.w3(32'h3ae69369),
	.w4(32'hbc129c47),
	.w5(32'h3aeab67f),
	.w6(32'h3ba9596c),
	.w7(32'hba428de3),
	.w8(32'hba668284),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb788b6),
	.w1(32'hbb38f4a1),
	.w2(32'hbab3acc5),
	.w3(32'h3bc368bc),
	.w4(32'h3b79a20d),
	.w5(32'hbb2b7f53),
	.w6(32'h3b84658f),
	.w7(32'h3bc87bc5),
	.w8(32'hba277360),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d06b1),
	.w1(32'hbc15b096),
	.w2(32'hba826486),
	.w3(32'hbba61120),
	.w4(32'hbb5ba210),
	.w5(32'hbba8a88d),
	.w6(32'hbb904371),
	.w7(32'hbaae73bd),
	.w8(32'hbc3dc01d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb6388),
	.w1(32'hbc349d29),
	.w2(32'hba3f44b1),
	.w3(32'hbc2b74e2),
	.w4(32'hbb8388a6),
	.w5(32'hbaaf87be),
	.w6(32'hbc7fafdc),
	.w7(32'hbb2833f3),
	.w8(32'hb94ece16),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399343d7),
	.w1(32'hbb34aee5),
	.w2(32'hbb15685f),
	.w3(32'hbab33857),
	.w4(32'h3b756e8d),
	.w5(32'h3b079c0f),
	.w6(32'h3a9e287a),
	.w7(32'h3b5d3593),
	.w8(32'h392ea6f5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88dbe1),
	.w1(32'h39e75fd0),
	.w2(32'h3ac5b518),
	.w3(32'h3aa54ba8),
	.w4(32'hbb9f3125),
	.w5(32'h3b0b0154),
	.w6(32'h3b8824d5),
	.w7(32'h3b86d31b),
	.w8(32'hba6f0cd6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4722b8),
	.w1(32'h3ba918cf),
	.w2(32'h3b807537),
	.w3(32'hbbe67c42),
	.w4(32'hbc4d15f3),
	.w5(32'hbb3449cb),
	.w6(32'hbbb35f26),
	.w7(32'hbb12cd68),
	.w8(32'h3afc7244),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf049c),
	.w1(32'hbac7c6ca),
	.w2(32'hbc1e0f52),
	.w3(32'h3beeb1b5),
	.w4(32'h3a460743),
	.w5(32'hbb4f3557),
	.w6(32'hbb975e4f),
	.w7(32'hbb49bb1b),
	.w8(32'h3ab368e3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3327d7),
	.w1(32'hbbd8924b),
	.w2(32'h3a8c58a6),
	.w3(32'hba787168),
	.w4(32'hbb0f6a8b),
	.w5(32'hbbd543d2),
	.w6(32'hbbc28c60),
	.w7(32'h3bbdbacf),
	.w8(32'hb97a99e8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb556a1f),
	.w1(32'h3bd7decc),
	.w2(32'hbbce4088),
	.w3(32'h3be0b6b6),
	.w4(32'hbb3a9f45),
	.w5(32'h3c24d5f8),
	.w6(32'h3b760d62),
	.w7(32'hbc53dbe1),
	.w8(32'h3cc449a0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b127b),
	.w1(32'hba6226af),
	.w2(32'hbba30055),
	.w3(32'hbb063077),
	.w4(32'h3a27329a),
	.w5(32'h3c4d5630),
	.w6(32'hb9ec835d),
	.w7(32'hbb6fb88f),
	.w8(32'h3cc8173d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b73a3),
	.w1(32'h3c1891c6),
	.w2(32'hbc0dc8c0),
	.w3(32'h3b864e73),
	.w4(32'hbb068035),
	.w5(32'h3c29df4d),
	.w6(32'hbbdc9d7c),
	.w7(32'hbcc2760f),
	.w8(32'h3b825bd4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb95f5),
	.w1(32'hbb85745c),
	.w2(32'hbbff1c90),
	.w3(32'h3ae294fd),
	.w4(32'hbb6a0d3d),
	.w5(32'hbba325de),
	.w6(32'hbb7a3fcc),
	.w7(32'h3b501a39),
	.w8(32'hbbb3729e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5d955),
	.w1(32'hbb064abc),
	.w2(32'hbb7eb0ab),
	.w3(32'hbbb21b0c),
	.w4(32'hbb0d2385),
	.w5(32'h3c914790),
	.w6(32'h3a9e1c90),
	.w7(32'hbb56608b),
	.w8(32'h3d0c239a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d029fc4),
	.w1(32'h3af512d1),
	.w2(32'hbc75a581),
	.w3(32'hbc0b7a50),
	.w4(32'hbc2d4dbf),
	.w5(32'h3b473d47),
	.w6(32'hbb9568a5),
	.w7(32'hbd0e7cd6),
	.w8(32'h3bfb2e35),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1efd95),
	.w1(32'hba869da6),
	.w2(32'hbbe4a0ab),
	.w3(32'h3bd54d5c),
	.w4(32'hbb7a9f4b),
	.w5(32'hbbcbb9f3),
	.w6(32'hbb75bf68),
	.w7(32'hbbf9d2a4),
	.w8(32'hbbddbb6f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05be24),
	.w1(32'hbb7c4f90),
	.w2(32'hbb9cc70e),
	.w3(32'h3b1e1f52),
	.w4(32'hbb306e6a),
	.w5(32'hbc3e841a),
	.w6(32'h3b41f7a5),
	.w7(32'hbb86cd17),
	.w8(32'hbbc3d956),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaa742),
	.w1(32'hbba68916),
	.w2(32'h3ac01620),
	.w3(32'hbbe25bd4),
	.w4(32'hba4118c2),
	.w5(32'h3ace7d38),
	.w6(32'h3a8b0ed6),
	.w7(32'h3aa5ff37),
	.w8(32'h3b9b72f2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52d1a9),
	.w1(32'hbba0d3e1),
	.w2(32'hbc3b0687),
	.w3(32'hb9f97b8c),
	.w4(32'hbbce457a),
	.w5(32'h3b9397d5),
	.w6(32'h3864b542),
	.w7(32'hbbfd045f),
	.w8(32'h3c7be070),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3b375),
	.w1(32'h3c1c3727),
	.w2(32'hbc1fffb2),
	.w3(32'h3c195f0c),
	.w4(32'hbc096abe),
	.w5(32'hbc7d1a0e),
	.w6(32'h3b979e75),
	.w7(32'hbc8d4832),
	.w8(32'hbc9d52a1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d9536),
	.w1(32'hbbc4b441),
	.w2(32'hbb7e4e8d),
	.w3(32'hbb786152),
	.w4(32'hbb0e3d29),
	.w5(32'h3a81ffa6),
	.w6(32'hbbc79c93),
	.w7(32'hbb301d93),
	.w8(32'h3bebb5f0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f9794),
	.w1(32'h3b2026cc),
	.w2(32'hbc1eefb7),
	.w3(32'hbb4698c7),
	.w4(32'hbb52cf2a),
	.w5(32'hbb0408d8),
	.w6(32'hbb523613),
	.w7(32'hbbef4ad3),
	.w8(32'hbbec278a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a31ba),
	.w1(32'hbb274485),
	.w2(32'hbb893968),
	.w3(32'hbabae3d5),
	.w4(32'hb9dd15b3),
	.w5(32'hbc80d14e),
	.w6(32'h3ba117d7),
	.w7(32'hbc0f3c67),
	.w8(32'hbcae1616),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81d9d9),
	.w1(32'hbac7b0ba),
	.w2(32'h3c1cfe15),
	.w3(32'h3c06a77e),
	.w4(32'h3c16d657),
	.w5(32'hbb1c260a),
	.w6(32'h3bc12e1d),
	.w7(32'h3c6aa191),
	.w8(32'h3a742927),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb337223),
	.w1(32'hbb127f61),
	.w2(32'h3bb1e845),
	.w3(32'h39b61c61),
	.w4(32'h398dd4a3),
	.w5(32'h3b8a77a5),
	.w6(32'hbc40873e),
	.w7(32'hbb0983a4),
	.w8(32'h3bfb4979),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7aca2),
	.w1(32'h3c9ba381),
	.w2(32'hbaff3231),
	.w3(32'h3ae47a8d),
	.w4(32'hbc3b92ef),
	.w5(32'hbb5092d6),
	.w6(32'h3c8a188d),
	.w7(32'hbc640dee),
	.w8(32'hbbfa2091),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af34c56),
	.w1(32'hbb1a26ec),
	.w2(32'hbc0b503a),
	.w3(32'h39c0f74f),
	.w4(32'hbb0ab186),
	.w5(32'h3ada0c67),
	.w6(32'h3b410ecc),
	.w7(32'hbc16e2b8),
	.w8(32'hba620e31),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8fca0),
	.w1(32'hbaac3597),
	.w2(32'hba8828cf),
	.w3(32'h3a32687d),
	.w4(32'hba8cb7f5),
	.w5(32'h3ad9a6d9),
	.w6(32'h3aa4d928),
	.w7(32'h39cd2005),
	.w8(32'h3ba8bba8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c003e5f),
	.w1(32'hbc2a5723),
	.w2(32'hbc770976),
	.w3(32'hbb63fb68),
	.w4(32'h3b3e50cb),
	.w5(32'h3ac3c26f),
	.w6(32'hbc50e0a8),
	.w7(32'hbb32e64c),
	.w8(32'h3c1206f6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387743e2),
	.w1(32'hbb89c447),
	.w2(32'hbb75382a),
	.w3(32'hb9297802),
	.w4(32'hbbdf81d4),
	.w5(32'h3c2a7653),
	.w6(32'hbb586da1),
	.w7(32'hbc2b1c12),
	.w8(32'h3ca0e9a0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d14d8),
	.w1(32'h3bbb1778),
	.w2(32'hbc8d7380),
	.w3(32'h3af6927b),
	.w4(32'hbc26881a),
	.w5(32'h39b585a8),
	.w6(32'hbbde358a),
	.w7(32'hbd255183),
	.w8(32'hbc5dc4ca),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2573c),
	.w1(32'hbae4fc64),
	.w2(32'hbbdee19f),
	.w3(32'hbc076737),
	.w4(32'h3b4566e0),
	.w5(32'h3b15db06),
	.w6(32'hbb80db83),
	.w7(32'hb9e5d0ec),
	.w8(32'hbb85d625),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb386c06),
	.w1(32'hbbfa79dc),
	.w2(32'h3c0978a9),
	.w3(32'hbc09343d),
	.w4(32'h3c22f42c),
	.w5(32'hbbb5aa47),
	.w6(32'hbc165c22),
	.w7(32'h3c22a05c),
	.w8(32'hbc713d6c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51bb8a),
	.w1(32'hbc2f04ca),
	.w2(32'h3bf6a54a),
	.w3(32'h3ba0a99d),
	.w4(32'h3c639eae),
	.w5(32'hbc1f9e4a),
	.w6(32'hba2068b3),
	.w7(32'h3cd6be5b),
	.w8(32'hbc80c450),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03db5),
	.w1(32'h3a7cdf93),
	.w2(32'h3c56d0ad),
	.w3(32'h3ada90ae),
	.w4(32'h3b588e67),
	.w5(32'h37e9f9af),
	.w6(32'h3915c46a),
	.w7(32'h3c77e99d),
	.w8(32'hbc1b03e1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0db773),
	.w1(32'hbb826259),
	.w2(32'h3bec9027),
	.w3(32'hbc05b746),
	.w4(32'h3a12dc4c),
	.w5(32'hbb4fff2e),
	.w6(32'h3bc43e43),
	.w7(32'h3c971a8b),
	.w8(32'hbbf10ff0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeecb6),
	.w1(32'hbc1515c6),
	.w2(32'hbbbf7530),
	.w3(32'hba01b6d1),
	.w4(32'hbb057f35),
	.w5(32'h3c46ec0c),
	.w6(32'hb7cee4ae),
	.w7(32'h3a591a4d),
	.w8(32'h3c4aba89),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b634b94),
	.w1(32'h3b2cd8af),
	.w2(32'hbb860956),
	.w3(32'h3ad3cf16),
	.w4(32'hbc746764),
	.w5(32'hba31d887),
	.w6(32'h3bcbae27),
	.w7(32'hbb86a8ff),
	.w8(32'hbb424e4b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f48f0),
	.w1(32'h3ae4081d),
	.w2(32'h3b8e7bd2),
	.w3(32'hba4758a8),
	.w4(32'h3b549e8b),
	.w5(32'hbc0bd17f),
	.w6(32'h3c802e6c),
	.w7(32'hba1e5309),
	.w8(32'hbc16de21),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38304c),
	.w1(32'hbba79b7f),
	.w2(32'h3ac7f38f),
	.w3(32'h3a72a6fb),
	.w4(32'h3c108a57),
	.w5(32'h3a92bfb3),
	.w6(32'hba768ad0),
	.w7(32'h3c105995),
	.w8(32'hbb6549ae),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4131b),
	.w1(32'h39e40e26),
	.w2(32'h3c2df4cf),
	.w3(32'h3bbf9dce),
	.w4(32'h3bb71750),
	.w5(32'h3a2fb446),
	.w6(32'h3c212784),
	.w7(32'h3c5c2f2e),
	.w8(32'h3bef0391),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d35d6),
	.w1(32'h3a27e288),
	.w2(32'h39396554),
	.w3(32'hba8402e3),
	.w4(32'hba788d97),
	.w5(32'h3c28a3b5),
	.w6(32'h3ac5bd7d),
	.w7(32'hbb41738a),
	.w8(32'h3c68c731),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15eb66),
	.w1(32'h39164ddd),
	.w2(32'hbc725988),
	.w3(32'hba765506),
	.w4(32'hbc68e203),
	.w5(32'h3c138544),
	.w6(32'h3ac4f225),
	.w7(32'hbc8a723b),
	.w8(32'h3c04ca1c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29563f),
	.w1(32'hbc5b3504),
	.w2(32'h3bd9cf2f),
	.w3(32'hbc92016b),
	.w4(32'h3a09ffa0),
	.w5(32'hbb963837),
	.w6(32'hbc6b6336),
	.w7(32'h3abdd24f),
	.w8(32'hbbfcbde1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194065),
	.w1(32'hbc05d522),
	.w2(32'hbc5a700b),
	.w3(32'hbb30086f),
	.w4(32'hbc24ce0f),
	.w5(32'h3b0b6b94),
	.w6(32'hbb92d6c9),
	.w7(32'hbc56ab36),
	.w8(32'h3af0d8a2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a5515),
	.w1(32'hbb45425d),
	.w2(32'hbb884a40),
	.w3(32'hbb97a6db),
	.w4(32'hbc272cf9),
	.w5(32'hbaf030c5),
	.w6(32'hbb01668d),
	.w7(32'hbb86d9b5),
	.w8(32'hbb69be87),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8556fc),
	.w1(32'hbb8f8dd1),
	.w2(32'hbc45426b),
	.w3(32'h3c0da4fb),
	.w4(32'h3c33f22e),
	.w5(32'hbb8ecbf9),
	.w6(32'h3b946c19),
	.w7(32'h3b1e3fc8),
	.w8(32'hbc5bf5c9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc475eb9),
	.w1(32'hbba7c78f),
	.w2(32'h3beb4afc),
	.w3(32'hb9943888),
	.w4(32'h3bece4c4),
	.w5(32'hbad3be85),
	.w6(32'hbb74d598),
	.w7(32'h3c068a4e),
	.w8(32'hbb2c195f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc00c10),
	.w1(32'hbbbef9ad),
	.w2(32'hbc4b73fd),
	.w3(32'hbb5d0a69),
	.w4(32'hbc2f8258),
	.w5(32'h3b38d1a6),
	.w6(32'hbb6e222d),
	.w7(32'hbc4809e5),
	.w8(32'h3b437b06),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf25be),
	.w1(32'hbc436de5),
	.w2(32'hbc96c55b),
	.w3(32'hbb9a6000),
	.w4(32'hbc1af7e2),
	.w5(32'h3b3291bd),
	.w6(32'hbc01ff51),
	.w7(32'hbc7ecff0),
	.w8(32'h3bed7179),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99f7a6),
	.w1(32'hbbe25c1c),
	.w2(32'h39f7571d),
	.w3(32'hbb33bf1b),
	.w4(32'hba797f8b),
	.w5(32'hbc916147),
	.w6(32'hbc2a9b3d),
	.w7(32'hbbc4a160),
	.w8(32'hbcf6f7f3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1ea2a),
	.w1(32'hbc08d55b),
	.w2(32'h3caf1e0b),
	.w3(32'hbba113ee),
	.w4(32'h3cc53e79),
	.w5(32'hbbf601af),
	.w6(32'hbc15f3ff),
	.w7(32'h3d08d3bb),
	.w8(32'hbb22913f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb640a41),
	.w1(32'hbbc60fcc),
	.w2(32'h3ac4a93a),
	.w3(32'hbc07bc11),
	.w4(32'hbb124557),
	.w5(32'hb8d22b32),
	.w6(32'h3c008d46),
	.w7(32'hbb38b2ea),
	.w8(32'h3a660528),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe5be2),
	.w1(32'hb968ea4f),
	.w2(32'hbc01d45b),
	.w3(32'hbb9cada8),
	.w4(32'hbb949849),
	.w5(32'hbb821e16),
	.w6(32'hbb179178),
	.w7(32'hbb7a374d),
	.w8(32'hb936ab73),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a836fe0),
	.w1(32'hbc08dc7f),
	.w2(32'hba676cd2),
	.w3(32'hbb95340a),
	.w4(32'hbb500518),
	.w5(32'hba3c2657),
	.w6(32'hbbb1341e),
	.w7(32'h3bc96f9f),
	.w8(32'hbbaf4a46),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29c57b),
	.w1(32'hbc2614b9),
	.w2(32'hbbde5cc4),
	.w3(32'h3beeae9c),
	.w4(32'h3b257f8e),
	.w5(32'hbaa75886),
	.w6(32'h39a70acc),
	.w7(32'hba8e9475),
	.w8(32'hba3d9824),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae278b5),
	.w1(32'hbb3e7d67),
	.w2(32'h3a9e51ca),
	.w3(32'hbbca90c2),
	.w4(32'h38a93a85),
	.w5(32'h3c3cae5f),
	.w6(32'hbb4471cf),
	.w7(32'hbb2665ce),
	.w8(32'h3cc545b4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c691c03),
	.w1(32'hbb44b7c4),
	.w2(32'hbc91c6c7),
	.w3(32'h3a9f0f83),
	.w4(32'hbc3c254a),
	.w5(32'h3b29dd74),
	.w6(32'hbbb1fa1e),
	.w7(32'hbcb7ab0a),
	.w8(32'h3a33fec0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39563e60),
	.w1(32'hbb465ebb),
	.w2(32'hba875877),
	.w3(32'hbb26ca21),
	.w4(32'hbb953153),
	.w5(32'hb994a048),
	.w6(32'h3b0b52f8),
	.w7(32'hbb8a83db),
	.w8(32'hba88778d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b085f50),
	.w1(32'h3b25c0be),
	.w2(32'h3c5e2590),
	.w3(32'hb8ae8367),
	.w4(32'h3adbacc1),
	.w5(32'h3c1392fe),
	.w6(32'h3ae60d0c),
	.w7(32'h3c88e493),
	.w8(32'h3c3f7206),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be94757),
	.w1(32'h3aeeee10),
	.w2(32'hbc3e5eb7),
	.w3(32'h3a83ea6e),
	.w4(32'hbc3dfe3a),
	.w5(32'hbb84979e),
	.w6(32'hb995d5e5),
	.w7(32'hbc728e34),
	.w8(32'hbb8cbf8f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e676b),
	.w1(32'h3b598303),
	.w2(32'h3b59ee60),
	.w3(32'h38ef1e43),
	.w4(32'hba9751dc),
	.w5(32'hbb4f0967),
	.w6(32'h3ae6ff19),
	.w7(32'hb8f1e12f),
	.w8(32'hbc2f4ac5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb041c1c),
	.w1(32'hba79dd43),
	.w2(32'h3bbaaf76),
	.w3(32'h3a6f744e),
	.w4(32'h3c538e2b),
	.w5(32'hbacd021a),
	.w6(32'h3c0a6cd6),
	.w7(32'h3c1b82a6),
	.w8(32'hbb48bc08),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39917),
	.w1(32'h3b6434ee),
	.w2(32'hbb870713),
	.w3(32'hbb18e4ee),
	.w4(32'hbb4968bc),
	.w5(32'h3b530fae),
	.w6(32'hbc0cc19e),
	.w7(32'hbb22edb1),
	.w8(32'h3c0d6d1d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b652e47),
	.w1(32'h38ce677b),
	.w2(32'hbc1236ed),
	.w3(32'hba689100),
	.w4(32'hbc003455),
	.w5(32'hbadab1b1),
	.w6(32'hbb405434),
	.w7(32'hbbf902c9),
	.w8(32'h3b13fe66),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9d624),
	.w1(32'h3a12bcfc),
	.w2(32'hbbb91513),
	.w3(32'h3b0520dd),
	.w4(32'h39aa10d2),
	.w5(32'hbc3f4e2e),
	.w6(32'hbb148c15),
	.w7(32'hbb80b150),
	.w8(32'hbc943371),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca78d8e),
	.w1(32'hbba64c21),
	.w2(32'h3c176fc4),
	.w3(32'hbb717acf),
	.w4(32'h3c115cdc),
	.w5(32'h39a24885),
	.w6(32'hbbdd575a),
	.w7(32'h3c3f5e8d),
	.w8(32'h3b51994d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d75b),
	.w1(32'hbbb18977),
	.w2(32'hbb18e20e),
	.w3(32'hbaee9d62),
	.w4(32'hbbd8e53d),
	.w5(32'h3b19a696),
	.w6(32'h3bc17a37),
	.w7(32'hb9aec34f),
	.w8(32'h3a4058b3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c9461),
	.w1(32'h3b5487e8),
	.w2(32'h3b7e70fe),
	.w3(32'h3ba29a5d),
	.w4(32'h3b954a2c),
	.w5(32'h3b337c06),
	.w6(32'h3c19146b),
	.w7(32'h3b71ef12),
	.w8(32'h3b447a4d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2dade),
	.w1(32'h3bc622f2),
	.w2(32'h3bf31e01),
	.w3(32'hbb414412),
	.w4(32'h3c0842eb),
	.w5(32'hba714c78),
	.w6(32'hbb84d889),
	.w7(32'h3c3ebc76),
	.w8(32'h3a26acb9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98fa22),
	.w1(32'h3c01194a),
	.w2(32'h3c2d9038),
	.w3(32'h3ba39bf6),
	.w4(32'h3add4cd9),
	.w5(32'h3c03c184),
	.w6(32'h3ae9a70c),
	.w7(32'h3c12cd69),
	.w8(32'h3c1e07fb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c222e53),
	.w1(32'h3bd5a9af),
	.w2(32'h3bdc3716),
	.w3(32'h3b879d7b),
	.w4(32'h3b220f46),
	.w5(32'hbac8fa2b),
	.w6(32'h3c4d62b3),
	.w7(32'hbbb023c5),
	.w8(32'hba1f3e45),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1e4a4),
	.w1(32'hbbb97987),
	.w2(32'h3a0f9215),
	.w3(32'hbb977833),
	.w4(32'h3a0c839d),
	.w5(32'hbbc38455),
	.w6(32'h3abad129),
	.w7(32'hbb001163),
	.w8(32'hbba81a4b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45e063),
	.w1(32'hbaa4c5bd),
	.w2(32'hba3b45bf),
	.w3(32'hbb7c4cb5),
	.w4(32'hbbdc3e58),
	.w5(32'hbbbd9545),
	.w6(32'hbb6f54ed),
	.w7(32'hbb5c1486),
	.w8(32'hba29c425),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a8e59),
	.w1(32'h3bf11599),
	.w2(32'h3b261f68),
	.w3(32'h38face23),
	.w4(32'h3be2c930),
	.w5(32'h3b4b735a),
	.w6(32'h3bc9f190),
	.w7(32'h3c309e07),
	.w8(32'h3bb15d33),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f7379),
	.w1(32'hbbd03f70),
	.w2(32'hbbe8d64f),
	.w3(32'h3a4290bf),
	.w4(32'h3c129b46),
	.w5(32'hbba7536a),
	.w6(32'hbc468df4),
	.w7(32'hbbb36d97),
	.w8(32'hbb63086b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb785b3a),
	.w1(32'hba279c0f),
	.w2(32'hbc0a5808),
	.w3(32'hba49bb1b),
	.w4(32'hbc19deef),
	.w5(32'hbc42d252),
	.w6(32'h39d371d4),
	.w7(32'hbba2b860),
	.w8(32'hbc2f9ce1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9a54),
	.w1(32'h3b89bd5f),
	.w2(32'h3ba8315e),
	.w3(32'hbb752cab),
	.w4(32'h3b6a8af0),
	.w5(32'h3c5206d6),
	.w6(32'hba89c353),
	.w7(32'h3ca3db64),
	.w8(32'h3cede080),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c7882),
	.w1(32'h3b2f3e16),
	.w2(32'hbc875640),
	.w3(32'hbbda3025),
	.w4(32'hbc4b6c4d),
	.w5(32'hbbc8f013),
	.w6(32'hbb9da875),
	.w7(32'hbcf7652d),
	.w8(32'hbb07f975),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb513414),
	.w1(32'h3c171520),
	.w2(32'h3bb5727f),
	.w3(32'h3ac48ae9),
	.w4(32'h3c20715c),
	.w5(32'h3bd5a1e0),
	.w6(32'h3c239a46),
	.w7(32'h3c4a4ae7),
	.w8(32'h3c01f6b9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb5302),
	.w1(32'h3a96e0cc),
	.w2(32'hbc72f523),
	.w3(32'h3b684f4b),
	.w4(32'hbc56ae23),
	.w5(32'h3b90e147),
	.w6(32'h3b8289b1),
	.w7(32'hbc600ebd),
	.w8(32'h3bc75f83),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aafb9),
	.w1(32'h3b79ae37),
	.w2(32'hbad63556),
	.w3(32'hbb781bd2),
	.w4(32'hbc04fc64),
	.w5(32'h39c46b34),
	.w6(32'hbb86f06a),
	.w7(32'hbc34b060),
	.w8(32'h3bfd7a8f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eb669),
	.w1(32'hbbb36697),
	.w2(32'hbafa1df6),
	.w3(32'h3b580454),
	.w4(32'hb9d562fc),
	.w5(32'h3c90cceb),
	.w6(32'hba93fa01),
	.w7(32'hbb30425e),
	.w8(32'h3d028471),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8105c),
	.w1(32'h3c2bda6d),
	.w2(32'hbc9e41df),
	.w3(32'h3b721fdb),
	.w4(32'hbc1d849d),
	.w5(32'h3c40c6f5),
	.w6(32'h3a469cf1),
	.w7(32'hbd12fe2c),
	.w8(32'h3c760b38),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd5055),
	.w1(32'hbb3526f6),
	.w2(32'hbc3b6148),
	.w3(32'h3b16bed2),
	.w4(32'hbb6e72ce),
	.w5(32'h3c328755),
	.w6(32'h3b41f025),
	.w7(32'hbc021eec),
	.w8(32'h3cc305ae),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6afbca),
	.w1(32'hbb9d1d1a),
	.w2(32'hbc788487),
	.w3(32'hbc387d23),
	.w4(32'hbc288b8e),
	.w5(32'hbc0bc633),
	.w6(32'hbc45fa2f),
	.w7(32'hbcc40e6f),
	.w8(32'hbcb16001),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fa994),
	.w1(32'hbb179d1f),
	.w2(32'h3c7b01fa),
	.w3(32'h389accca),
	.w4(32'h3c77f586),
	.w5(32'hbc766d7c),
	.w6(32'hb97477c5),
	.w7(32'h3cc5710c),
	.w8(32'hbccddcfc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97bb5b),
	.w1(32'h3bfc7134),
	.w2(32'h3cc2bc48),
	.w3(32'hbb4a4163),
	.w4(32'h3c89cca2),
	.w5(32'h3bfbad2c),
	.w6(32'h3afa3a5c),
	.w7(32'h3ced7410),
	.w8(32'h3c114033),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfce5c7),
	.w1(32'h3aac22d7),
	.w2(32'hbc037507),
	.w3(32'h3b13e911),
	.w4(32'hbc1eed28),
	.w5(32'h3bd613f8),
	.w6(32'h3b942888),
	.w7(32'hbc3a132d),
	.w8(32'hbbc9256a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32b6fe),
	.w1(32'hbbf2a590),
	.w2(32'h3b8acaa9),
	.w3(32'hbc0b2d69),
	.w4(32'h3c6f5a5a),
	.w5(32'h3b8393f0),
	.w6(32'hbb96ed5c),
	.w7(32'h3bbce241),
	.w8(32'h3be8de1a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05eab3),
	.w1(32'h3997ac61),
	.w2(32'hbc36bc08),
	.w3(32'hbb692cbd),
	.w4(32'hbc4d646d),
	.w5(32'hbac0f66d),
	.w6(32'hbbe6e143),
	.w7(32'hbc7cd800),
	.w8(32'h3b060319),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982e58e),
	.w1(32'h3933304e),
	.w2(32'hbc378972),
	.w3(32'hbc38d656),
	.w4(32'hbb82da9d),
	.w5(32'hbb941347),
	.w6(32'hbbe54e3c),
	.w7(32'hbc27cde2),
	.w8(32'hbb3d3ffe),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac14ba4),
	.w1(32'h3ab6e0fd),
	.w2(32'h3c0dccc3),
	.w3(32'h397095ba),
	.w4(32'h3bd95817),
	.w5(32'h3c03d114),
	.w6(32'hba05b4d0),
	.w7(32'h3b3d9256),
	.w8(32'h3ac45f8a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad45554),
	.w1(32'hbb7b8081),
	.w2(32'hbb476c2d),
	.w3(32'h3aef391f),
	.w4(32'hbbf78021),
	.w5(32'h3ad1b4dd),
	.w6(32'h3b4616d1),
	.w7(32'hbb81d68f),
	.w8(32'hbb6b504c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ef9ca),
	.w1(32'hbbe9727c),
	.w2(32'hba91f39a),
	.w3(32'h3b5e0d89),
	.w4(32'h3a090293),
	.w5(32'hbbe8e506),
	.w6(32'h3beeec2b),
	.w7(32'h3b86db46),
	.w8(32'hbbe555f9),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22d2db),
	.w1(32'hbb57a7f7),
	.w2(32'h390f791f),
	.w3(32'h395c50a2),
	.w4(32'h3abf5e35),
	.w5(32'hbb535510),
	.w6(32'h3badbd0d),
	.w7(32'h3b943697),
	.w8(32'hbae55235),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba151229),
	.w1(32'hbc228703),
	.w2(32'hbb50f66e),
	.w3(32'hbbeeb55f),
	.w4(32'hb9d5c6c8),
	.w5(32'h3bedb0f0),
	.w6(32'hbb2005e7),
	.w7(32'hbb054416),
	.w8(32'h3ba84ce4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09b385),
	.w1(32'h3b18be88),
	.w2(32'hbaa56c75),
	.w3(32'h3b896881),
	.w4(32'hbb6d9606),
	.w5(32'h3c66e101),
	.w6(32'h3b87e3f7),
	.w7(32'hbb076fd4),
	.w8(32'h3c8eee77),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d5600),
	.w1(32'hbbf7c88d),
	.w2(32'hbb91f73b),
	.w3(32'h3b0241f0),
	.w4(32'h3b0133a2),
	.w5(32'hbba4b1eb),
	.w6(32'hbc9cf45f),
	.w7(32'hbbe7d519),
	.w8(32'hba8d8b69),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5af9b6),
	.w1(32'h3b808974),
	.w2(32'hb9f2c93c),
	.w3(32'hbaf71cb1),
	.w4(32'h3ad435ef),
	.w5(32'h3b798042),
	.w6(32'hba7eee50),
	.w7(32'h3b9a1262),
	.w8(32'h3c06c0b6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1df0fa),
	.w1(32'hbb96f84b),
	.w2(32'hbbc469f9),
	.w3(32'hba83174e),
	.w4(32'hbc09caaf),
	.w5(32'hbb48256b),
	.w6(32'h3b2b264a),
	.w7(32'hbad64734),
	.w8(32'hbc335fc3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3d850),
	.w1(32'hbb975526),
	.w2(32'hba1acd3e),
	.w3(32'hbb663a21),
	.w4(32'h3b5f037d),
	.w5(32'hbad5c0d8),
	.w6(32'hbc04bbe6),
	.w7(32'h39735f06),
	.w8(32'hbaa66cc3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6759ab),
	.w1(32'h39dea15b),
	.w2(32'h3a7aa23f),
	.w3(32'h3b1aef61),
	.w4(32'h3b9aa1ea),
	.w5(32'h3bc99a70),
	.w6(32'h3c2cda1f),
	.w7(32'h3b7a75d0),
	.w8(32'hba9d9b08),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ce329),
	.w1(32'hb945f3a5),
	.w2(32'h3b5b1268),
	.w3(32'h3aedc521),
	.w4(32'hbbf01e5a),
	.w5(32'h3bd08c7b),
	.w6(32'h3c14d2c4),
	.w7(32'h3a4cd18b),
	.w8(32'h3b683688),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccacc5),
	.w1(32'hbaa02edd),
	.w2(32'hbc0c3d8f),
	.w3(32'hba049d89),
	.w4(32'hbb236ae4),
	.w5(32'h36ea0ad3),
	.w6(32'hbc0c964e),
	.w7(32'hbae70b39),
	.w8(32'h3a408223),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb46ef5),
	.w1(32'hbb21bdd6),
	.w2(32'hbc571ce9),
	.w3(32'h3a23ef8c),
	.w4(32'hbb365206),
	.w5(32'hbb5072d0),
	.w6(32'h3ad5068a),
	.w7(32'hba9b284d),
	.w8(32'hbc6b7a33),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60d4dd),
	.w1(32'hbc13c1ad),
	.w2(32'h3c1e5291),
	.w3(32'hbb147368),
	.w4(32'h3bcd8036),
	.w5(32'hb96e3ea5),
	.w6(32'hbc26187f),
	.w7(32'h3c443bcc),
	.w8(32'hbbd6f9bc),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b770732),
	.w1(32'hbc25cd7b),
	.w2(32'hbaee1ede),
	.w3(32'hbc462180),
	.w4(32'hbb530612),
	.w5(32'hbc187572),
	.w6(32'h39fcbaeb),
	.w7(32'hba71e393),
	.w8(32'h3bcfafc4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f228b),
	.w1(32'hbb632361),
	.w2(32'hbb7fa167),
	.w3(32'h3b905db7),
	.w4(32'hbbadd64a),
	.w5(32'h3b372bd3),
	.w6(32'h3c06d0ba),
	.w7(32'hbc5cca9e),
	.w8(32'h3c1f5569),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdba88f),
	.w1(32'hbb02ff98),
	.w2(32'hbc3264d9),
	.w3(32'hbae618ba),
	.w4(32'hbbef1738),
	.w5(32'hbba81f17),
	.w6(32'hbc0a30a1),
	.w7(32'hbc942fa6),
	.w8(32'h3a785319),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d4c80),
	.w1(32'h3b9c9179),
	.w2(32'h3983e6f6),
	.w3(32'h3b7fc6ab),
	.w4(32'h3c1d3462),
	.w5(32'hbc272c2b),
	.w6(32'hba68d543),
	.w7(32'h3c65a8ff),
	.w8(32'hbc1dc5a9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9cad6),
	.w1(32'hba436232),
	.w2(32'h3b9307d5),
	.w3(32'hba690c40),
	.w4(32'h3b16aa90),
	.w5(32'hbbfc3708),
	.w6(32'hbc1a1534),
	.w7(32'h3bc594db),
	.w8(32'hbc168b40),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc205c93),
	.w1(32'hbb3a7219),
	.w2(32'h3bec798e),
	.w3(32'hba16164c),
	.w4(32'h3c01469b),
	.w5(32'hbb83fffa),
	.w6(32'h3aacac78),
	.w7(32'h3c4b814b),
	.w8(32'hbb9ade30),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd2412),
	.w1(32'hbc202c0c),
	.w2(32'hbc4fcefe),
	.w3(32'hba78f1d5),
	.w4(32'hbb532dfb),
	.w5(32'hbc85657b),
	.w6(32'hbb4fecdf),
	.w7(32'hbbd4bfdc),
	.w8(32'hbcaaa90b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc786cc6),
	.w1(32'hbb218c6d),
	.w2(32'h3cbe28ce),
	.w3(32'hbbb0f629),
	.w4(32'h3ca9ddfb),
	.w5(32'hbb1ff92e),
	.w6(32'hbba9e538),
	.w7(32'h3cf276fa),
	.w8(32'h3b05af69),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d4650),
	.w1(32'h39b963fa),
	.w2(32'hbb6964bc),
	.w3(32'hbaa984ff),
	.w4(32'h3b117894),
	.w5(32'h3c3482c9),
	.w6(32'hbb358417),
	.w7(32'h3ab31f1a),
	.w8(32'h3cdc8219),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5db687),
	.w1(32'hbbc8dc5f),
	.w2(32'hbc623eba),
	.w3(32'hbbb0b6b8),
	.w4(32'hbc3fbb3c),
	.w5(32'h3bfd2cb9),
	.w6(32'h3ad80f0a),
	.w7(32'hbcc37577),
	.w8(32'h3c2fb97d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb97d71),
	.w1(32'h3b12f636),
	.w2(32'hbb0b8835),
	.w3(32'hba3eec73),
	.w4(32'h3b1153dd),
	.w5(32'hbc1f8d8f),
	.w6(32'hbc0df028),
	.w7(32'hbbbc8708),
	.w8(32'hbc81efab),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9003cd),
	.w1(32'hbbcd2878),
	.w2(32'hbb82aed4),
	.w3(32'hbb5100ed),
	.w4(32'h3990f0fe),
	.w5(32'hbc3a1569),
	.w6(32'hbb2e85e3),
	.w7(32'h3b68ca59),
	.w8(32'hbc011097),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbb9fd),
	.w1(32'h3bc7b9c6),
	.w2(32'h3be90b11),
	.w3(32'hbb6a86d9),
	.w4(32'h3b998ba2),
	.w5(32'hbc1e26ce),
	.w6(32'hbb17e050),
	.w7(32'hbb4fa71f),
	.w8(32'hbc2db000),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee4e7f),
	.w1(32'h3b635463),
	.w2(32'h3bb22f52),
	.w3(32'hbb0307e7),
	.w4(32'hbb10b5b9),
	.w5(32'h3b25a660),
	.w6(32'h3b199345),
	.w7(32'h3b575857),
	.w8(32'h3b9435cf),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c68c4),
	.w1(32'hb96c835d),
	.w2(32'hbc116272),
	.w3(32'hbb79dd48),
	.w4(32'hbb3c5306),
	.w5(32'h3ba0db25),
	.w6(32'h3bf41737),
	.w7(32'hba45216b),
	.w8(32'hba433d43),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba469b82),
	.w1(32'hbb660629),
	.w2(32'hbb97e38f),
	.w3(32'hbabdd185),
	.w4(32'hbb8a80fe),
	.w5(32'hbb50b705),
	.w6(32'hbb51b569),
	.w7(32'h3a05f85f),
	.w8(32'hbb8b706d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf407d0),
	.w1(32'hba90ed4f),
	.w2(32'h3ac1ff57),
	.w3(32'hbb99529c),
	.w4(32'h3a1f6c33),
	.w5(32'h3bc2615b),
	.w6(32'hb9fdf1a2),
	.w7(32'h3b8c1097),
	.w8(32'h3c194252),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89b0c6),
	.w1(32'hba341abd),
	.w2(32'hbbede4b4),
	.w3(32'h3aafd91f),
	.w4(32'hb9af088b),
	.w5(32'hbaa5393c),
	.w6(32'h3b8875d4),
	.w7(32'h3c0bbd53),
	.w8(32'h3b319f72),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c164721),
	.w1(32'hbb9090d1),
	.w2(32'hbc2b5749),
	.w3(32'hbb8f4683),
	.w4(32'hbb620c4b),
	.w5(32'hba30c38e),
	.w6(32'hba5fd596),
	.w7(32'hbc4ee83d),
	.w8(32'hbb3ef09d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53bb38),
	.w1(32'hbb886390),
	.w2(32'hba5edbd2),
	.w3(32'hba84aad4),
	.w4(32'h3b1d855c),
	.w5(32'hbb6dfbf7),
	.w6(32'hbb878577),
	.w7(32'h3b92dd30),
	.w8(32'hbbc686f6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9ed78),
	.w1(32'hbba727a3),
	.w2(32'hbb960cf9),
	.w3(32'hbb8029bb),
	.w4(32'hbbb80798),
	.w5(32'h3abf61aa),
	.w6(32'hbb51206a),
	.w7(32'hbb84cc83),
	.w8(32'hbb38bb2b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4f990),
	.w1(32'hbb105be7),
	.w2(32'h3b1628b1),
	.w3(32'h3b6b837e),
	.w4(32'h3c1a4ed8),
	.w5(32'hbb765349),
	.w6(32'h3aaeff61),
	.w7(32'hba4af4ae),
	.w8(32'hbc2a14a8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf4f4c),
	.w1(32'h3c008d1f),
	.w2(32'h3ca02032),
	.w3(32'hb8a1104c),
	.w4(32'h3c4ff7fc),
	.w5(32'h3be22054),
	.w6(32'h3c8286a3),
	.w7(32'h3c310efd),
	.w8(32'h3c75450f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b875e25),
	.w1(32'hbbf6c126),
	.w2(32'hbb29c235),
	.w3(32'hbc154688),
	.w4(32'hbc091427),
	.w5(32'h3ba726d3),
	.w6(32'hbc0faa86),
	.w7(32'hbbf70c80),
	.w8(32'h3956e590),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1054d4),
	.w1(32'hbbef7067),
	.w2(32'h3b88f1a7),
	.w3(32'hbc2427c1),
	.w4(32'h3bf19aab),
	.w5(32'h38fc586b),
	.w6(32'hbb4c2b9d),
	.w7(32'h3b679504),
	.w8(32'hba6ac2d9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b5be7),
	.w1(32'hbbe87c3d),
	.w2(32'hbbaea27c),
	.w3(32'hbc1a938b),
	.w4(32'hbbfbd6e4),
	.w5(32'hb93b10ea),
	.w6(32'hbc291621),
	.w7(32'hbba6cb29),
	.w8(32'h3b71d46f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc8311),
	.w1(32'h3b0ddd15),
	.w2(32'hbac20804),
	.w3(32'hb98d4549),
	.w4(32'hbb02c2d3),
	.w5(32'h3c21ddbc),
	.w6(32'h3bac3d3a),
	.w7(32'h39923d6f),
	.w8(32'h3c8198d4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be93b9b),
	.w1(32'h3b1d646f),
	.w2(32'hbb93a18d),
	.w3(32'hbb7843d6),
	.w4(32'hbc80ed90),
	.w5(32'h3c21fcf8),
	.w6(32'hbb7eff95),
	.w7(32'hbc80f4ea),
	.w8(32'h3c66ad62),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87b578),
	.w1(32'h3b49d553),
	.w2(32'hbb7fd7eb),
	.w3(32'h3c009594),
	.w4(32'h3bcb3d46),
	.w5(32'hbb102a46),
	.w6(32'hbb6ca584),
	.w7(32'hbc650675),
	.w8(32'h3af9e838),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc39ebf),
	.w1(32'h3a2b27c7),
	.w2(32'h3b5c9590),
	.w3(32'hbc1bf139),
	.w4(32'h3be188eb),
	.w5(32'hbb063453),
	.w6(32'h3c09f764),
	.w7(32'h3c0e7ed9),
	.w8(32'h3ae72b75),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd1744),
	.w1(32'h3904a770),
	.w2(32'h3b130dca),
	.w3(32'h3a08606d),
	.w4(32'h3b44cbd8),
	.w5(32'h39c02566),
	.w6(32'h3bf1799e),
	.w7(32'h3c0c211f),
	.w8(32'h3a3b5411),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8eeb7),
	.w1(32'h3a81f038),
	.w2(32'hbaba15fa),
	.w3(32'hb9aeaf34),
	.w4(32'hbb061260),
	.w5(32'h3916175a),
	.w6(32'hbb1f1924),
	.w7(32'hbb84f4d1),
	.w8(32'hbb874717),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab98b5d),
	.w1(32'hbb0c6f9d),
	.w2(32'hba613ce8),
	.w3(32'hbb3994fe),
	.w4(32'h3ad22a47),
	.w5(32'hbb9960d5),
	.w6(32'hbbd073df),
	.w7(32'hbb2d9ce3),
	.w8(32'hbacf5476),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89e5c6),
	.w1(32'h3c01c548),
	.w2(32'h3c124a12),
	.w3(32'hbb96db96),
	.w4(32'hbbc490d1),
	.w5(32'h3a3ca98c),
	.w6(32'hba76b9c7),
	.w7(32'h3bb1c0a9),
	.w8(32'hbac21ef1),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb368418),
	.w1(32'hba2d2392),
	.w2(32'hba990a43),
	.w3(32'hbb20399e),
	.w4(32'hbb75810f),
	.w5(32'hbb9fdb2b),
	.w6(32'hbb8b9e1f),
	.w7(32'hbb748e51),
	.w8(32'hbb5c4cf0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a724aee),
	.w1(32'h3b9ddeca),
	.w2(32'h3b3b54a3),
	.w3(32'hba28d3fd),
	.w4(32'hba297f01),
	.w5(32'hbac5c687),
	.w6(32'h3b840135),
	.w7(32'h3b2758dc),
	.w8(32'h3adb11c5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a64c),
	.w1(32'hbbae11aa),
	.w2(32'h3b97c48e),
	.w3(32'h3c134281),
	.w4(32'h3c1985c0),
	.w5(32'h3acd0b65),
	.w6(32'h3c6e8384),
	.w7(32'h3c84ac68),
	.w8(32'h3ba0785b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b3723),
	.w1(32'h3b4fb7d9),
	.w2(32'hba1119da),
	.w3(32'h3b5aa56f),
	.w4(32'h3b8b6daf),
	.w5(32'hbae3a6fe),
	.w6(32'h3a36f1d6),
	.w7(32'h39a5eb3b),
	.w8(32'hb982ac58),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f80ac),
	.w1(32'hbbaa39e0),
	.w2(32'hbb9fca89),
	.w3(32'h3a670fda),
	.w4(32'hb7e9a1e9),
	.w5(32'hbb27cc60),
	.w6(32'hbb8baa61),
	.w7(32'hbaf6b22d),
	.w8(32'hbc177ee8),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b258566),
	.w1(32'h3b9d9a2d),
	.w2(32'h3acbc2a4),
	.w3(32'hbb0b1759),
	.w4(32'hb9f53cdd),
	.w5(32'hbbe71020),
	.w6(32'hbbe29244),
	.w7(32'hbc2393eb),
	.w8(32'h3b19f3a9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82aeb9),
	.w1(32'hbb9a22d1),
	.w2(32'hbb25f027),
	.w3(32'hbba43858),
	.w4(32'hbb1f4568),
	.w5(32'hba8625ed),
	.w6(32'h3bcf8b98),
	.w7(32'h3bf0f82b),
	.w8(32'h3a4321e4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2afb4),
	.w1(32'h3c35dea7),
	.w2(32'h3c2c1d05),
	.w3(32'hb9b9ac06),
	.w4(32'h3b90bdde),
	.w5(32'h3bf6d071),
	.w6(32'h3c1d1351),
	.w7(32'h3b9d66c6),
	.w8(32'h390c5fce),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b741f08),
	.w1(32'h3bb5f584),
	.w2(32'h3be59dcc),
	.w3(32'h3b044d37),
	.w4(32'hbaf57292),
	.w5(32'h3abeef02),
	.w6(32'hb976229e),
	.w7(32'h3bad6e07),
	.w8(32'hbb215c53),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca100e),
	.w1(32'h3b13114f),
	.w2(32'h3b9085a2),
	.w3(32'h39b27601),
	.w4(32'h3ac78228),
	.w5(32'hbb44bb10),
	.w6(32'h3a0fd179),
	.w7(32'h3aa50151),
	.w8(32'h3ae00411),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb744868),
	.w1(32'h3ad94ffe),
	.w2(32'hbb6b2d3d),
	.w3(32'h3928e362),
	.w4(32'hbb6c18bb),
	.w5(32'h3b724d56),
	.w6(32'h3bc3c1a4),
	.w7(32'h3b06e8c2),
	.w8(32'h3b9b526a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc128dd1),
	.w1(32'hbbdc666f),
	.w2(32'hbbb04649),
	.w3(32'hb9379889),
	.w4(32'hba809c13),
	.w5(32'hb92f0b6e),
	.w6(32'h3b951210),
	.w7(32'h3b3ef568),
	.w8(32'hbb1e1d93),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b29fe),
	.w1(32'h3a67e3af),
	.w2(32'h3ac3acfb),
	.w3(32'h3b912d28),
	.w4(32'h3b063463),
	.w5(32'h3b316ee5),
	.w6(32'hb98c366f),
	.w7(32'h3b14d233),
	.w8(32'h3b711dd9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cc6b3),
	.w1(32'h3bb0dce6),
	.w2(32'h3ae196e6),
	.w3(32'hb8be58ec),
	.w4(32'hba8a7ae4),
	.w5(32'h3c257a29),
	.w6(32'h3b949b87),
	.w7(32'h3bcbabb0),
	.w8(32'h3c23fab8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d2864),
	.w1(32'h3bffb7df),
	.w2(32'h3bb36366),
	.w3(32'h3c6dcecd),
	.w4(32'h3c5355fa),
	.w5(32'hbb91830e),
	.w6(32'h3c3dab1c),
	.w7(32'h3bc1e482),
	.w8(32'hbb424143),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4834),
	.w1(32'hbb3fe819),
	.w2(32'h3b1be5d0),
	.w3(32'hbb876b78),
	.w4(32'hbb118eaa),
	.w5(32'hbaa2be22),
	.w6(32'h3ab06c1e),
	.w7(32'h3a182bbf),
	.w8(32'h3bb376c3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd68875),
	.w1(32'hbab825d0),
	.w2(32'hbbebfee9),
	.w3(32'h3b025e24),
	.w4(32'hbb0b4fd8),
	.w5(32'hbc61bef1),
	.w6(32'h3c171e4c),
	.w7(32'h3b2d606f),
	.w8(32'hbc07e4f9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31fa9c),
	.w1(32'hbbe71891),
	.w2(32'hbbb6df7d),
	.w3(32'hbc489b02),
	.w4(32'hbc10a2f8),
	.w5(32'h3a6b6b7a),
	.w6(32'hbbae3341),
	.w7(32'hbb02792b),
	.w8(32'hbba3a095),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae61b29),
	.w1(32'hbb416a88),
	.w2(32'hba3ed358),
	.w3(32'hba9eb737),
	.w4(32'hbb779fab),
	.w5(32'h3b790dfa),
	.w6(32'hbbb28d2d),
	.w7(32'hbb88a34f),
	.w8(32'h3ba58cd5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37ba8e),
	.w1(32'h3a7d5f31),
	.w2(32'h3bea8b1f),
	.w3(32'h3b07ed08),
	.w4(32'h3b99202a),
	.w5(32'hbc15fb78),
	.w6(32'hbb025b80),
	.w7(32'h3bde1d33),
	.w8(32'hbad2983e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1073ee),
	.w1(32'h3b0a9dbb),
	.w2(32'hb9e805f5),
	.w3(32'hbcae5b29),
	.w4(32'hbc45a2c0),
	.w5(32'h397b0bec),
	.w6(32'hbc8a5f93),
	.w7(32'hbb0d16db),
	.w8(32'hba8116bb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7da407),
	.w1(32'hbb33fc2f),
	.w2(32'h3ae92e66),
	.w3(32'hba28e1d4),
	.w4(32'h3b8e72ae),
	.w5(32'hbc2ee358),
	.w6(32'hbbf6eb97),
	.w7(32'h3a579fa8),
	.w8(32'hbc1f263f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8981c3),
	.w1(32'hbb00ab6f),
	.w2(32'hba8227f0),
	.w3(32'hbc7f4e0b),
	.w4(32'hbc226061),
	.w5(32'h3860c4c3),
	.w6(32'hbcb38730),
	.w7(32'hbc26729d),
	.w8(32'h3ae9da90),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4b7f5),
	.w1(32'h3b8884e6),
	.w2(32'h3b8e4c4e),
	.w3(32'hbaf9551b),
	.w4(32'hba354542),
	.w5(32'h3aca4640),
	.w6(32'hbb2c1258),
	.w7(32'h391bc98d),
	.w8(32'hbb9c07f6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c361280),
	.w1(32'h3c28e58d),
	.w2(32'h3c6b83a3),
	.w3(32'h3856df04),
	.w4(32'h3b6bf4ca),
	.w5(32'hbaa415ca),
	.w6(32'hbc219399),
	.w7(32'hbbfc6e29),
	.w8(32'hbaabb7a2),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeadce2),
	.w1(32'h3a696da8),
	.w2(32'hbb5f6b40),
	.w3(32'h3b857475),
	.w4(32'h3b396167),
	.w5(32'hba8e8bec),
	.w6(32'h3b404baa),
	.w7(32'h3b0f878d),
	.w8(32'hbb8908a9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule