module layer_10_featuremap_339(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f1ae3),
	.w1(32'h3c479488),
	.w2(32'h3c03cb98),
	.w3(32'hba0d7fbf),
	.w4(32'h3b985f98),
	.w5(32'h3c38d53d),
	.w6(32'h3c2e2af6),
	.w7(32'h3c1e3347),
	.w8(32'h3a6fb3e3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988b5ba),
	.w1(32'hbb981233),
	.w2(32'hbc41a27f),
	.w3(32'h3bbe542f),
	.w4(32'h3b9477ef),
	.w5(32'hba8d3ad2),
	.w6(32'hbb376a2c),
	.w7(32'hbc1a48b3),
	.w8(32'hbc078915),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25b0bf),
	.w1(32'h3a9db116),
	.w2(32'hba607f44),
	.w3(32'hbba07367),
	.w4(32'hbb909cc5),
	.w5(32'hba93bb2b),
	.w6(32'hb907722e),
	.w7(32'h3b1bfd53),
	.w8(32'hbb96cd6e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddd880),
	.w1(32'hbb130209),
	.w2(32'h39060278),
	.w3(32'hbabe0a2e),
	.w4(32'hbabdbd73),
	.w5(32'h3a1f2ee0),
	.w6(32'hbb9942f0),
	.w7(32'hbb507346),
	.w8(32'hbb87132a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31d601),
	.w1(32'hbc1fb6fb),
	.w2(32'hbc2110fe),
	.w3(32'hbc0a32c7),
	.w4(32'hbbf72eeb),
	.w5(32'hbb856d2c),
	.w6(32'hbbd05531),
	.w7(32'hbc2b857b),
	.w8(32'hbb4eb3f7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b37b0),
	.w1(32'hba595604),
	.w2(32'h3990ff3b),
	.w3(32'hbae2b61a),
	.w4(32'hbb0cc5cf),
	.w5(32'h3a763952),
	.w6(32'h3a24bd38),
	.w7(32'hba4021d5),
	.w8(32'hbb9aa00d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8079ef),
	.w1(32'h3af2a0a8),
	.w2(32'h3a41c66a),
	.w3(32'h3ba5e814),
	.w4(32'h3b0d8797),
	.w5(32'hbb50545f),
	.w6(32'h3b5a6976),
	.w7(32'h3afa6ab2),
	.w8(32'hbac18f32),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e6552),
	.w1(32'h3b2ef0d6),
	.w2(32'h3c8d3e09),
	.w3(32'hbb97ffa6),
	.w4(32'h390a7a16),
	.w5(32'h3b8d7e4d),
	.w6(32'hbb315eac),
	.w7(32'h3c17a12f),
	.w8(32'h3bc545e9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad61a4),
	.w1(32'h3b467bfa),
	.w2(32'h3b7bbad9),
	.w3(32'h3b41bd66),
	.w4(32'h3b1c8a72),
	.w5(32'hbba9ae97),
	.w6(32'h3ade081c),
	.w7(32'h3b0f998a),
	.w8(32'hbb11fa99),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7f681),
	.w1(32'h3ae05329),
	.w2(32'hb86349d8),
	.w3(32'hbad9eceb),
	.w4(32'hba71311a),
	.w5(32'hbb3a74de),
	.w6(32'h3b4cfaf1),
	.w7(32'h3b1b2c9a),
	.w8(32'hbbcbe91d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9ac78),
	.w1(32'hbb8d7486),
	.w2(32'hbb76293c),
	.w3(32'hbbcc9f54),
	.w4(32'hbbb63e00),
	.w5(32'h38d61815),
	.w6(32'hbb40f0f8),
	.w7(32'hbb376ec8),
	.w8(32'h3a2f5b34),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba547b18),
	.w1(32'hba663a03),
	.w2(32'h3baeebf7),
	.w3(32'h3acf98fc),
	.w4(32'h39b850b3),
	.w5(32'hbbcd0e71),
	.w6(32'h3a0d202a),
	.w7(32'h3b55abe3),
	.w8(32'hb884f32c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd40637),
	.w1(32'hb928ab32),
	.w2(32'hbb40af4d),
	.w3(32'hbbfe30c8),
	.w4(32'h3b817c77),
	.w5(32'h3b9d7793),
	.w6(32'hbabd02ce),
	.w7(32'h3ab5b06d),
	.w8(32'h3b9dbe83),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53d538),
	.w1(32'hbb13e402),
	.w2(32'hbb6f1df6),
	.w3(32'h3ba1c46c),
	.w4(32'h3ae3ec39),
	.w5(32'hb9c6505f),
	.w6(32'h3aaa6f57),
	.w7(32'hbb8f043a),
	.w8(32'hba7a93ba),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca0052),
	.w1(32'hbb9e6fc1),
	.w2(32'hbac852d3),
	.w3(32'h3aeb5dd4),
	.w4(32'hbb53fa2b),
	.w5(32'h3c1db80d),
	.w6(32'hbb2d7a8a),
	.w7(32'hbba89207),
	.w8(32'h3aaf3781),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad512a8),
	.w1(32'h3b15b757),
	.w2(32'h3b841903),
	.w3(32'h3b044af0),
	.w4(32'h3b7cf9b8),
	.w5(32'h3b4bbcb9),
	.w6(32'hbb50dde1),
	.w7(32'hbafefd98),
	.w8(32'h3b0c66f7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77080f),
	.w1(32'hbb96aa10),
	.w2(32'h3aa8b3dc),
	.w3(32'h3b2987db),
	.w4(32'h3bbdc826),
	.w5(32'h3bab3ace),
	.w6(32'hbb2e49ea),
	.w7(32'hba90c5a4),
	.w8(32'h3b2b3f9b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6f791),
	.w1(32'hbab7eefc),
	.w2(32'h3b94c2eb),
	.w3(32'h3ad4379b),
	.w4(32'h3bc98718),
	.w5(32'h3c2e588f),
	.w6(32'hba1c0611),
	.w7(32'h3c10bfa7),
	.w8(32'h3c8c1158),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb11a2),
	.w1(32'h39ce2d02),
	.w2(32'h3ba1dc9c),
	.w3(32'h3abd7093),
	.w4(32'h3b2c47f2),
	.w5(32'h3bb4e8c0),
	.w6(32'hba05ffc7),
	.w7(32'h3bfac253),
	.w8(32'h3bf197d6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b237d60),
	.w1(32'hbaa8566d),
	.w2(32'hbb4a0422),
	.w3(32'h3b872851),
	.w4(32'h3b63f0a4),
	.w5(32'h3c30f813),
	.w6(32'hbb1b2ec4),
	.w7(32'hbb7bf528),
	.w8(32'h3b8bf1ac),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac018b7),
	.w1(32'hbb8c275a),
	.w2(32'hbae7c96e),
	.w3(32'h3b5268b8),
	.w4(32'h3bdf7de1),
	.w5(32'h39a46729),
	.w6(32'hbb9506ae),
	.w7(32'hbad88c3b),
	.w8(32'hba79d7ca),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14a076),
	.w1(32'hbac171a6),
	.w2(32'h3907878d),
	.w3(32'h3b4eba1a),
	.w4(32'h3b28ef74),
	.w5(32'hb90ee162),
	.w6(32'hb9f0cb80),
	.w7(32'h3ad0019f),
	.w8(32'hbb2b8efa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bcf8c),
	.w1(32'hbc578df9),
	.w2(32'h3b03a22f),
	.w3(32'hbba471ad),
	.w4(32'hbb3d8310),
	.w5(32'h3c61d4a2),
	.w6(32'hbb957fff),
	.w7(32'h3b8dfed3),
	.w8(32'h3c2a9f53),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bee25),
	.w1(32'h3b96d05a),
	.w2(32'h3b15cac5),
	.w3(32'hba0799ee),
	.w4(32'h3bb1c834),
	.w5(32'hbb40a8cd),
	.w6(32'h3b5f0240),
	.w7(32'h39bb7b7c),
	.w8(32'hbb11960d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2c171),
	.w1(32'h3b769ac7),
	.w2(32'hbb907d81),
	.w3(32'hbb4ce603),
	.w4(32'hbb884ea4),
	.w5(32'hbbc62da0),
	.w6(32'hbb03f972),
	.w7(32'hbbe58172),
	.w8(32'hbc068c95),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7a60),
	.w1(32'hbbd76cb3),
	.w2(32'h3b4e1e6b),
	.w3(32'h3a78135a),
	.w4(32'hbb28bc78),
	.w5(32'hba3d719c),
	.w6(32'hbb51309c),
	.w7(32'hbb3d1e39),
	.w8(32'hbb41d18e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb518de4),
	.w1(32'hbb2a5da3),
	.w2(32'hbb16e373),
	.w3(32'hba98ad44),
	.w4(32'hbb3335fd),
	.w5(32'hb993887d),
	.w6(32'hbafd5d68),
	.w7(32'hbb4d569c),
	.w8(32'h3b4d4154),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb674c8),
	.w1(32'h3c373025),
	.w2(32'h3b73cd85),
	.w3(32'h3b60e09a),
	.w4(32'h3bb1f223),
	.w5(32'hbb5966b8),
	.w6(32'h3bcb40e3),
	.w7(32'h3a819608),
	.w8(32'hbc185ee3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9832fe0),
	.w1(32'hba8a44a8),
	.w2(32'hb945a469),
	.w3(32'h3aebb52b),
	.w4(32'hba84cc8b),
	.w5(32'hb9f9796a),
	.w6(32'hbb4443f5),
	.w7(32'hbb08f808),
	.w8(32'hbadc04a0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e3a61),
	.w1(32'h3ae5a631),
	.w2(32'hbb93f03a),
	.w3(32'hb911670c),
	.w4(32'hbaabb99e),
	.w5(32'hbbb39b6c),
	.w6(32'hba95160d),
	.w7(32'hbc2f5e41),
	.w8(32'hbc0abe46),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e2d1a),
	.w1(32'h3a0bf1b4),
	.w2(32'h37c3ed5b),
	.w3(32'h3b3560a7),
	.w4(32'hbb988ceb),
	.w5(32'hb9b77e60),
	.w6(32'h3bbaf082),
	.w7(32'h395ef272),
	.w8(32'h3ad7fc81),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58521a),
	.w1(32'hbb11eacd),
	.w2(32'hbabfaf3c),
	.w3(32'h3b906326),
	.w4(32'h3babf6a5),
	.w5(32'hbaefa704),
	.w6(32'h3b029037),
	.w7(32'h3ba42537),
	.w8(32'hbb2cc8aa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc189f50),
	.w1(32'hbbc276d2),
	.w2(32'hb9eb53b4),
	.w3(32'h39ab5dd4),
	.w4(32'hbb8af563),
	.w5(32'h3c0f93d1),
	.w6(32'hbbb79464),
	.w7(32'hbafd4fb2),
	.w8(32'h3ab3f123),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb315321),
	.w1(32'hbaacc4a2),
	.w2(32'hbb5e5a77),
	.w3(32'h3bdcc063),
	.w4(32'h3b2fd931),
	.w5(32'hb9fa3ebf),
	.w6(32'h3ad7d808),
	.w7(32'hbbba5960),
	.w8(32'hbb681504),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fe48c),
	.w1(32'hb9d0c818),
	.w2(32'h3aee608d),
	.w3(32'hbabf1c34),
	.w4(32'hb99aa890),
	.w5(32'h3aee1b7a),
	.w6(32'hbb910ff0),
	.w7(32'hbadd7a65),
	.w8(32'hbb0fa4d9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67033c),
	.w1(32'hba33016f),
	.w2(32'h3a73b18b),
	.w3(32'h3ae21a1a),
	.w4(32'hb98c4453),
	.w5(32'h3c0533d5),
	.w6(32'hbb1ef908),
	.w7(32'hb9951ca8),
	.w8(32'h3b77a3f3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cae9d),
	.w1(32'hbbeb3876),
	.w2(32'h3b1567e1),
	.w3(32'h3c0a22d3),
	.w4(32'hbbf57038),
	.w5(32'h3b8d4999),
	.w6(32'h3b1753d0),
	.w7(32'hbb6e82f7),
	.w8(32'h3b80852d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399232e6),
	.w1(32'hbaafc1e1),
	.w2(32'hbc14ccd3),
	.w3(32'h3bbd1adf),
	.w4(32'hbb065fd0),
	.w5(32'h3a69efc0),
	.w6(32'h3b5d3263),
	.w7(32'hbbfc59c1),
	.w8(32'hbbc5c681),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ab1bd),
	.w1(32'h3c38b73c),
	.w2(32'hbbae7e85),
	.w3(32'h3c6ac498),
	.w4(32'h3bc441f6),
	.w5(32'hbc5e97bc),
	.w6(32'h3c4bd40e),
	.w7(32'h3af0e13f),
	.w8(32'hbcaff895),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06f6d3),
	.w1(32'hbbf83049),
	.w2(32'hbc490ea4),
	.w3(32'hb9e309f4),
	.w4(32'hbb3f4215),
	.w5(32'h3acf3e07),
	.w6(32'hbb9e631e),
	.w7(32'hbc08fb15),
	.w8(32'h3ae29bbf),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4f985),
	.w1(32'h39fd6bee),
	.w2(32'h3b533c75),
	.w3(32'h3b66fb0c),
	.w4(32'h3b61cf82),
	.w5(32'hbbb0d641),
	.w6(32'h3b395332),
	.w7(32'h3b7292a7),
	.w8(32'hbbd4ba0c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ae73),
	.w1(32'hbbd6e83c),
	.w2(32'h3a381f0c),
	.w3(32'hbb9ea663),
	.w4(32'hbbb01f98),
	.w5(32'h3b0d1c38),
	.w6(32'hbb72fbd9),
	.w7(32'hbb2e4993),
	.w8(32'h3bb88cef),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be18d3f),
	.w1(32'h3b326405),
	.w2(32'h3944e879),
	.w3(32'hbab2ca1e),
	.w4(32'hbbc58de4),
	.w5(32'hb9ae3940),
	.w6(32'hb9b2d253),
	.w7(32'hbad6d323),
	.w8(32'hbb541a12),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe27777),
	.w1(32'hbbde6096),
	.w2(32'hbb954585),
	.w3(32'hbc4aa508),
	.w4(32'hbbb92405),
	.w5(32'h3b71c7a2),
	.w6(32'hbbe6978a),
	.w7(32'hbb94acff),
	.w8(32'h3c056da9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c56cb),
	.w1(32'hb8fc17aa),
	.w2(32'hbb4757a9),
	.w3(32'h3ad590f8),
	.w4(32'hba94d7d1),
	.w5(32'hbb5c9067),
	.w6(32'h3b4bfd10),
	.w7(32'h38e19a58),
	.w8(32'hbb2b400a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80058ea),
	.w1(32'h3b8a6c16),
	.w2(32'h3c046b07),
	.w3(32'hbb387a2e),
	.w4(32'h3b282de6),
	.w5(32'hbb0fc4fc),
	.w6(32'h3bd3bdf5),
	.w7(32'h3bf4ea1b),
	.w8(32'hbacb083f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6438a),
	.w1(32'hba9faf10),
	.w2(32'hba846287),
	.w3(32'hb9dd8b71),
	.w4(32'hb780d1a2),
	.w5(32'h3b0a9e64),
	.w6(32'hb9c419e9),
	.w7(32'hb7bdb54b),
	.w8(32'h3b70bcff),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3603f6),
	.w1(32'h3b08d1a7),
	.w2(32'h3c362350),
	.w3(32'h3b991a30),
	.w4(32'h3c50e137),
	.w5(32'h3b2a3031),
	.w6(32'h3b2ce29b),
	.w7(32'h3c853aea),
	.w8(32'h3c861a3f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09c171),
	.w1(32'h3a67b044),
	.w2(32'hbb87f4f6),
	.w3(32'hbc153be4),
	.w4(32'hbb9e8123),
	.w5(32'h3bb7ab1f),
	.w6(32'h3b106fd8),
	.w7(32'hbb5b4d75),
	.w8(32'h3a8c11e9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3645b3),
	.w1(32'h3a6cf4a6),
	.w2(32'h3b8abfaa),
	.w3(32'h3bc40687),
	.w4(32'h3bb6e19c),
	.w5(32'hbc56d85f),
	.w6(32'h3b406a3c),
	.w7(32'h3bbac955),
	.w8(32'hbbf27db2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab6c05),
	.w1(32'h3aca265a),
	.w2(32'h3ad32973),
	.w3(32'hbb8917b3),
	.w4(32'h37914220),
	.w5(32'h39b4c1be),
	.w6(32'h3b5b7d28),
	.w7(32'h3af37bbb),
	.w8(32'hb9911490),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ee7a4),
	.w1(32'hbb65bb1c),
	.w2(32'hbb8df6ed),
	.w3(32'hbb3b6044),
	.w4(32'hbb8a9ede),
	.w5(32'h3af7a672),
	.w6(32'hbba8b75f),
	.w7(32'hbbabc3cf),
	.w8(32'hbb4c34cc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a4634),
	.w1(32'h3b27bc4e),
	.w2(32'h3a16d283),
	.w3(32'hbae95003),
	.w4(32'h3b4928ff),
	.w5(32'h3b229628),
	.w6(32'h3b7c8336),
	.w7(32'h3bb7a62c),
	.w8(32'hbb2fe900),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc461bfb),
	.w1(32'hbc04d235),
	.w2(32'hb968f025),
	.w3(32'hbba0cd16),
	.w4(32'hb9dcb49d),
	.w5(32'h3c4cf779),
	.w6(32'hbb68f019),
	.w7(32'h3b84959d),
	.w8(32'h3c55c23a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc4817),
	.w1(32'hbb725529),
	.w2(32'hbb78db78),
	.w3(32'hba6947db),
	.w4(32'h3a772698),
	.w5(32'h3b6d9757),
	.w6(32'hbb56264b),
	.w7(32'hbb55eb9d),
	.w8(32'h3b4c4aed),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1988e5),
	.w1(32'hbab52f88),
	.w2(32'hba3784b7),
	.w3(32'h3afa5449),
	.w4(32'hbb23dccf),
	.w5(32'h3b879ba1),
	.w6(32'hbadc28fe),
	.w7(32'hbba4cf65),
	.w8(32'h3bd61f13),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90db9f),
	.w1(32'h3b4f2f8a),
	.w2(32'h3bbe2169),
	.w3(32'h3bcffd74),
	.w4(32'h3ba2dc66),
	.w5(32'h3b3cfe47),
	.w6(32'h3b43986b),
	.w7(32'h3b9e15d4),
	.w8(32'hb9c7672a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ad72e),
	.w1(32'h390f60b1),
	.w2(32'hbbb89a38),
	.w3(32'hb9bca7fe),
	.w4(32'h381a9913),
	.w5(32'h3bb012ea),
	.w6(32'h37dc4efa),
	.w7(32'hbb54cb00),
	.w8(32'h39e92b76),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0332),
	.w1(32'h3a298e41),
	.w2(32'h3b86059b),
	.w3(32'h3be90128),
	.w4(32'h3b6b71bf),
	.w5(32'h3ac4e3c9),
	.w6(32'h3b6719f1),
	.w7(32'h3badfd87),
	.w8(32'h3c3fa57a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be093ec),
	.w1(32'h3bd38cdb),
	.w2(32'h3ba96bd9),
	.w3(32'h3ad3993c),
	.w4(32'h3a92236a),
	.w5(32'h3bc9db40),
	.w6(32'h3c2a15d2),
	.w7(32'h3c190de1),
	.w8(32'h3bbbc5c8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70ea47),
	.w1(32'h3b8dd349),
	.w2(32'h3bf93c3b),
	.w3(32'h3ab3d08b),
	.w4(32'h3b42d17b),
	.w5(32'h3b91cabd),
	.w6(32'h3b60d1d3),
	.w7(32'h3b87fb8e),
	.w8(32'h3b6360cb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdd1f7),
	.w1(32'hbb38e418),
	.w2(32'h3bf015c9),
	.w3(32'hbb8dc25a),
	.w4(32'h3b8f690c),
	.w5(32'h3b93cc24),
	.w6(32'h3ad12a5b),
	.w7(32'h3bacfaa3),
	.w8(32'h3b8fc6da),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4592b5),
	.w1(32'hbb614c67),
	.w2(32'hbb0449d2),
	.w3(32'hb9729458),
	.w4(32'h3a7ac3f7),
	.w5(32'hba0eaf0f),
	.w6(32'h3a3446a2),
	.w7(32'hb9a71040),
	.w8(32'hbb497662),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ab957),
	.w1(32'hbb367fa2),
	.w2(32'hbb3bc7b1),
	.w3(32'hbaebb391),
	.w4(32'hbac7c0f3),
	.w5(32'h3b40060e),
	.w6(32'hbb4ea2a6),
	.w7(32'hbb531226),
	.w8(32'hbac6784c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2407),
	.w1(32'hbb6f47a4),
	.w2(32'hbae16816),
	.w3(32'h3ad7e70b),
	.w4(32'h3b7fb0e6),
	.w5(32'h3bad0e02),
	.w6(32'hbb8df059),
	.w7(32'hbb16861c),
	.w8(32'h3a8b28f9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cc579),
	.w1(32'h3a6c0056),
	.w2(32'hba966212),
	.w3(32'h3b66705f),
	.w4(32'h3b7f618b),
	.w5(32'hbad8281b),
	.w6(32'h3aa5285e),
	.w7(32'hbac15761),
	.w8(32'hbbc1f135),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5eae),
	.w1(32'h3c0ab03f),
	.w2(32'h3c616a28),
	.w3(32'hbbfb5b21),
	.w4(32'hbb23bf36),
	.w5(32'hba7c21f7),
	.w6(32'hbaf75196),
	.w7(32'h3a4ade9e),
	.w8(32'h3a7ab68a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31cec6),
	.w1(32'hbb541e71),
	.w2(32'hbb99da8c),
	.w3(32'hbc2626e9),
	.w4(32'hbc1baf2c),
	.w5(32'hbb630d51),
	.w6(32'hbb260ff1),
	.w7(32'hba0f0c4f),
	.w8(32'h3a950c91),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc83be5),
	.w1(32'hbb04c37d),
	.w2(32'hba56f107),
	.w3(32'hbab2f00d),
	.w4(32'h3a108915),
	.w5(32'h3ba97458),
	.w6(32'hbb3643c6),
	.w7(32'h3a4af27e),
	.w8(32'h3c0e0fe5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adda030),
	.w1(32'h3b2770f5),
	.w2(32'hbbbbe3f5),
	.w3(32'h3b49644f),
	.w4(32'h3b3adb26),
	.w5(32'hbb255f9d),
	.w6(32'h3b689768),
	.w7(32'hbb97e79b),
	.w8(32'hbc0f1a99),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe97b0),
	.w1(32'hbb0eaa08),
	.w2(32'hbb0091c8),
	.w3(32'h394a8551),
	.w4(32'hbae0937c),
	.w5(32'h3b0c2b2c),
	.w6(32'hbaf4cef2),
	.w7(32'hbb25125d),
	.w8(32'h3a5f7d9b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2fdac),
	.w1(32'h3b06abbb),
	.w2(32'h3bd82ad6),
	.w3(32'h3ba732d8),
	.w4(32'h3ba1bcae),
	.w5(32'h3b58a331),
	.w6(32'hbae08306),
	.w7(32'h386b1b89),
	.w8(32'h3be0d616),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba112344),
	.w1(32'h3a6f01fc),
	.w2(32'hba145e8a),
	.w3(32'h3b81683c),
	.w4(32'h3afa0c80),
	.w5(32'h3bb210fa),
	.w6(32'h3b1e4452),
	.w7(32'h3b9fadae),
	.w8(32'h3ac74188),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0595ca),
	.w1(32'hbb98acca),
	.w2(32'hbbb54f5a),
	.w3(32'h3b160152),
	.w4(32'hba39d8ec),
	.w5(32'h3bb75931),
	.w6(32'hba1c9502),
	.w7(32'hbbd782ae),
	.w8(32'h3b1970a1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d9397),
	.w1(32'h3ace0a75),
	.w2(32'hbad2f7ea),
	.w3(32'hbb11dbef),
	.w4(32'hbaf4d0e9),
	.w5(32'hbb9b0688),
	.w6(32'hbade5fe1),
	.w7(32'hbb6c30f7),
	.w8(32'h3a832d87),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacff812),
	.w1(32'hbb6107ca),
	.w2(32'hbafc53f0),
	.w3(32'hbb90e8eb),
	.w4(32'hbbd6a8d1),
	.w5(32'h3c005292),
	.w6(32'h37a462bb),
	.w7(32'hbaad508e),
	.w8(32'h3bbb7f65),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a964953),
	.w1(32'hbadf31be),
	.w2(32'h3b32a137),
	.w3(32'hbb27b0f2),
	.w4(32'hbb0aca2d),
	.w5(32'h3c04b04d),
	.w6(32'h3af90935),
	.w7(32'h3bcb95b0),
	.w8(32'h3c03c1a1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24dfb7),
	.w1(32'h3b3c7308),
	.w2(32'hb8f5798f),
	.w3(32'h3bd4474d),
	.w4(32'h3b6dfb8b),
	.w5(32'hbadc4d2a),
	.w6(32'h3b771503),
	.w7(32'h3a78d483),
	.w8(32'hbb811f50),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea5b54),
	.w1(32'h3b832ec3),
	.w2(32'h3b1ad02c),
	.w3(32'h3ad751d2),
	.w4(32'h3b952d2a),
	.w5(32'h3aec9e9b),
	.w6(32'h3b1b2abc),
	.w7(32'h3b8f32fc),
	.w8(32'h3a721d71),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf56aa3),
	.w1(32'h383c0bd4),
	.w2(32'h3bd8ee31),
	.w3(32'hbb07c397),
	.w4(32'h3ad2ba12),
	.w5(32'hbad0d1ff),
	.w6(32'h3a54a437),
	.w7(32'hbb2ed654),
	.w8(32'hbb04b59d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c027cb7),
	.w1(32'h3b8f69c9),
	.w2(32'h3ba9806c),
	.w3(32'hba1ca909),
	.w4(32'h3ade5f26),
	.w5(32'h3b3e35a1),
	.w6(32'h3a47e421),
	.w7(32'h3b19436b),
	.w8(32'h3bb58e4b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927f2d3),
	.w1(32'h3add1d97),
	.w2(32'h3b2d256d),
	.w3(32'h39bec62a),
	.w4(32'h3a8405d4),
	.w5(32'h3b108f48),
	.w6(32'h3b9fb09c),
	.w7(32'h3b978991),
	.w8(32'h3b8f7593),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae766fb),
	.w1(32'h3b07e7dd),
	.w2(32'hba1da7ad),
	.w3(32'hbade31a0),
	.w4(32'h3b2895b2),
	.w5(32'hbb37225d),
	.w6(32'h3b9b08bb),
	.w7(32'h3b5a7ac1),
	.w8(32'hbb851a29),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbe615),
	.w1(32'hbc0362d4),
	.w2(32'hbc3160a7),
	.w3(32'hba26adc5),
	.w4(32'hbbfd2aff),
	.w5(32'h3a41347d),
	.w6(32'hbbdfd5c7),
	.w7(32'hbc296e32),
	.w8(32'h3a75b779),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fc525),
	.w1(32'h3b6dbc31),
	.w2(32'h3ac9cc28),
	.w3(32'h3901aed8),
	.w4(32'h3a9fc50d),
	.w5(32'h3a6efe71),
	.w6(32'h3b7645e3),
	.w7(32'h3b09c2ff),
	.w8(32'h3a1d3a07),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc96924),
	.w1(32'h3b4b1c51),
	.w2(32'h3bb828dc),
	.w3(32'h3b057939),
	.w4(32'h3bc5ecb0),
	.w5(32'h3a34dd87),
	.w6(32'h3c3746ac),
	.w7(32'h3c26c7da),
	.w8(32'hba775439),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bf633),
	.w1(32'hb9dc2e8f),
	.w2(32'hbb433869),
	.w3(32'hbb060b43),
	.w4(32'hbb83cccf),
	.w5(32'hbaacba1d),
	.w6(32'hb8c52274),
	.w7(32'hbb4657b6),
	.w8(32'hbaa27450),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b9dc5),
	.w1(32'hb9a18341),
	.w2(32'hbaf063e5),
	.w3(32'hbaab505b),
	.w4(32'hbaf9a693),
	.w5(32'h382cb5ec),
	.w6(32'hba829d68),
	.w7(32'hbb47e584),
	.w8(32'hbb84b504),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb646de1),
	.w1(32'hbb931968),
	.w2(32'hbae71c65),
	.w3(32'hba7ca2e6),
	.w4(32'hbae63621),
	.w5(32'hbbd8e10a),
	.w6(32'hbb97e0f0),
	.w7(32'hbb67149c),
	.w8(32'hbc018b16),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacc048),
	.w1(32'hb9fcc392),
	.w2(32'h3b866041),
	.w3(32'hbb0252b5),
	.w4(32'h3ba375c2),
	.w5(32'h3b941397),
	.w6(32'h3b077e21),
	.w7(32'h3b6c1436),
	.w8(32'h3afd9afc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47f4d3),
	.w1(32'hba2090f0),
	.w2(32'hbc0c9fa7),
	.w3(32'h3bbc3cf3),
	.w4(32'h3adb3b4c),
	.w5(32'hbbbd60bc),
	.w6(32'hb9693ef3),
	.w7(32'hbc1c84aa),
	.w8(32'hbc40457c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d491),
	.w1(32'hba579cc6),
	.w2(32'h3bad6a4e),
	.w3(32'hba413570),
	.w4(32'hba650d94),
	.w5(32'h3ab784d1),
	.w6(32'hbb661b8b),
	.w7(32'hbb47f3a4),
	.w8(32'hbbe901fb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47663b),
	.w1(32'hbc3b35a1),
	.w2(32'hbc83d36d),
	.w3(32'hbb12b2fc),
	.w4(32'hbc18b267),
	.w5(32'hbbff0e9e),
	.w6(32'hbbdc6bf8),
	.w7(32'hbc61e554),
	.w8(32'hbc1d0f10),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68583e),
	.w1(32'h37acfd78),
	.w2(32'h3aee512c),
	.w3(32'hb9527db6),
	.w4(32'hba0fac48),
	.w5(32'h3b4094c6),
	.w6(32'hba8ece0a),
	.w7(32'hba97292e),
	.w8(32'h3bfa832c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b3f9c),
	.w1(32'h3c01f6da),
	.w2(32'h3c08b31b),
	.w3(32'h3b21a319),
	.w4(32'h3b1a00de),
	.w5(32'h38e94258),
	.w6(32'h3b996132),
	.w7(32'h3b3c9e3c),
	.w8(32'hba3c3028),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12f599),
	.w1(32'h3bd6a3c8),
	.w2(32'hba7b19eb),
	.w3(32'h3b5ced6c),
	.w4(32'hbb8a59d5),
	.w5(32'hbb938570),
	.w6(32'hbb60397b),
	.w7(32'hbb0a6dab),
	.w8(32'hbbef2cfa),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba946ec3),
	.w1(32'hbae0692d),
	.w2(32'hbbb679f0),
	.w3(32'h3b4a32c3),
	.w4(32'h3b47b4fe),
	.w5(32'h3ab4f1b3),
	.w6(32'h3b1977a7),
	.w7(32'h3aff1e64),
	.w8(32'h3b9d0f2f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76a374),
	.w1(32'hbb9fa179),
	.w2(32'h3bb7b9b0),
	.w3(32'h3c502cf5),
	.w4(32'h3bd0d61f),
	.w5(32'h3c228950),
	.w6(32'h3b87d4b9),
	.w7(32'h3c041403),
	.w8(32'h3c46abe3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a058f47),
	.w1(32'h3bc64252),
	.w2(32'h3c05eb46),
	.w3(32'h3bd2f50d),
	.w4(32'h3bd2a141),
	.w5(32'h3b5d4862),
	.w6(32'h3be81e48),
	.w7(32'h3b6db0c6),
	.w8(32'hbb5bba82),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaca6e),
	.w1(32'hbbe45874),
	.w2(32'hbb6c2610),
	.w3(32'hbbc8ce44),
	.w4(32'hbc7d5405),
	.w5(32'h3ba072f7),
	.w6(32'hbc0faf53),
	.w7(32'hbbed27f3),
	.w8(32'h3c8053b8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bc6e0),
	.w1(32'h3a3283cb),
	.w2(32'hbc992859),
	.w3(32'hbb008383),
	.w4(32'hbc2b2e9f),
	.w5(32'hbc115d7a),
	.w6(32'h3bd85123),
	.w7(32'hbc9b3586),
	.w8(32'hbc0bcc2f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb739d3),
	.w1(32'h3a696f73),
	.w2(32'h3c6786c7),
	.w3(32'h3ab234eb),
	.w4(32'hbb8617ae),
	.w5(32'hbb37c803),
	.w6(32'h3bd685a9),
	.w7(32'h3a7c8c3e),
	.w8(32'hbc3dafc3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc84f72),
	.w1(32'h3c39a26d),
	.w2(32'h3c1ad17e),
	.w3(32'h3b6ca681),
	.w4(32'h3b7ce8fa),
	.w5(32'h3baf36fb),
	.w6(32'h3ca6580b),
	.w7(32'h3c73f94d),
	.w8(32'hb8d03016),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5324b8),
	.w1(32'hba291a8f),
	.w2(32'hbb2c4c84),
	.w3(32'hbb7ba848),
	.w4(32'hbba4b8ef),
	.w5(32'h3b5bb3c9),
	.w6(32'hbc35d3f5),
	.w7(32'h3b6288b2),
	.w8(32'h3bd75956),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad03ec1),
	.w1(32'hbc0fcb6b),
	.w2(32'hbc0692d3),
	.w3(32'h3c26f895),
	.w4(32'hbc6d0d81),
	.w5(32'h3be90a24),
	.w6(32'h3c66f0b5),
	.w7(32'hbb0b13ed),
	.w8(32'h3b1d5d32),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0999a8),
	.w1(32'h3af1a59f),
	.w2(32'h3aa9bb56),
	.w3(32'hbbbb424c),
	.w4(32'hba91d028),
	.w5(32'h3a87deac),
	.w6(32'hbc05ea7b),
	.w7(32'hba8ee594),
	.w8(32'h3c10908d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb37f66),
	.w1(32'hbc6b69d6),
	.w2(32'hbc2e94bb),
	.w3(32'hbc23b2df),
	.w4(32'hbbff2d92),
	.w5(32'h3b87713f),
	.w6(32'hbc1fa6a1),
	.w7(32'hbc25d005),
	.w8(32'h3b169ffc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8941b),
	.w1(32'h3b78a5c4),
	.w2(32'hbb3c846a),
	.w3(32'h39bc6834),
	.w4(32'hbb2cfca1),
	.w5(32'h3c3be25a),
	.w6(32'h3c00423b),
	.w7(32'hbb581208),
	.w8(32'h3c4df5f7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c050861),
	.w1(32'h3c013f8a),
	.w2(32'h3c2ee73a),
	.w3(32'h3c3ca742),
	.w4(32'h3c415797),
	.w5(32'h3ba863e0),
	.w6(32'h3ba475c3),
	.w7(32'h3c0212be),
	.w8(32'h3b40d88c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8df0e5),
	.w1(32'hbb73dd54),
	.w2(32'hbad8c1c6),
	.w3(32'hbb6e43c8),
	.w4(32'h3aaf3e07),
	.w5(32'hbb0a3496),
	.w6(32'hbc129f02),
	.w7(32'hbbe8919d),
	.w8(32'hbbe7c4c9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04d9d6),
	.w1(32'h3b824652),
	.w2(32'hbbdf6762),
	.w3(32'h3ba9dcff),
	.w4(32'hbba2e8a7),
	.w5(32'hbbf30806),
	.w6(32'h3bcf08ee),
	.w7(32'hbb6c12fd),
	.w8(32'hbc4f54e7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbabcc7),
	.w1(32'h390bd064),
	.w2(32'h3cb6985b),
	.w3(32'hbc2ff756),
	.w4(32'h3c643b95),
	.w5(32'h3a0923e9),
	.w6(32'hbb484bdf),
	.w7(32'h3cceaf17),
	.w8(32'hbb664ee7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbae812),
	.w1(32'h3b18c1eb),
	.w2(32'h3c012a49),
	.w3(32'h3c14e62c),
	.w4(32'h3bdedda9),
	.w5(32'h3b690cba),
	.w6(32'h3b64c942),
	.w7(32'h3b8d4009),
	.w8(32'hb9a40461),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ce7ee),
	.w1(32'h3c570c83),
	.w2(32'h3c2e2848),
	.w3(32'h3a15e497),
	.w4(32'h3cbf4d9e),
	.w5(32'h3c0313ac),
	.w6(32'hbbb83ca7),
	.w7(32'h3cb284d9),
	.w8(32'h3b3ec446),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba097c5b),
	.w1(32'hbb6403ef),
	.w2(32'hbb31d8b9),
	.w3(32'hbb7572f9),
	.w4(32'hbaee87e8),
	.w5(32'h3afc7c76),
	.w6(32'hbad5a466),
	.w7(32'hbb663d1b),
	.w8(32'h3a5bdfa3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2585e1),
	.w1(32'hbb2d38e6),
	.w2(32'h3c9d1189),
	.w3(32'hbbe0a920),
	.w4(32'h3aa8259f),
	.w5(32'h39cbfaf4),
	.w6(32'hbc00f852),
	.w7(32'h3bb605c9),
	.w8(32'h3a57bf04),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b981ebb),
	.w1(32'h39ac966a),
	.w2(32'hbae76f89),
	.w3(32'hbb77c9e8),
	.w4(32'hbba32cef),
	.w5(32'hb9157e72),
	.w6(32'hbb8168db),
	.w7(32'hbb90331f),
	.w8(32'h3bf89141),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8786d),
	.w1(32'hbbe6506f),
	.w2(32'hbc5bc513),
	.w3(32'hbb5bf12a),
	.w4(32'hbbe1c0db),
	.w5(32'hb988fb3e),
	.w6(32'h37cee684),
	.w7(32'hbc35e302),
	.w8(32'hbba68831),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8723b),
	.w1(32'hbc148365),
	.w2(32'hbc4fd971),
	.w3(32'hbba02d84),
	.w4(32'hbbbfecd7),
	.w5(32'h3b9c5e61),
	.w6(32'hbb85a800),
	.w7(32'hbc179c9b),
	.w8(32'hbaf62067),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aa8d5),
	.w1(32'h3bf3136d),
	.w2(32'h3bef4d0d),
	.w3(32'h3c1c98f8),
	.w4(32'h3c13611b),
	.w5(32'h3a93186f),
	.w6(32'h3c07be16),
	.w7(32'h3c4322f3),
	.w8(32'hbb0a5cc4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d1bee),
	.w1(32'h3b83b73c),
	.w2(32'h3c9ca4f1),
	.w3(32'hbc51b9be),
	.w4(32'h3c64e434),
	.w5(32'hbb341936),
	.w6(32'hbc81b9b0),
	.w7(32'h3cebaddc),
	.w8(32'hbc06c65c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cd110),
	.w1(32'hbbf7e9a2),
	.w2(32'h3c25d35c),
	.w3(32'hbb6e2ee4),
	.w4(32'h3ba56ebc),
	.w5(32'h38f812fb),
	.w6(32'hbbde3d1e),
	.w7(32'h3c57bdf1),
	.w8(32'h3bbb9f86),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45b7a5),
	.w1(32'hbb6802ad),
	.w2(32'hbb936444),
	.w3(32'h3b0d8c04),
	.w4(32'h38e4e507),
	.w5(32'hbbb03897),
	.w6(32'h3a6e0f81),
	.w7(32'hbbe5c49c),
	.w8(32'hbc6431ac),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d6b9c),
	.w1(32'hbb8acd33),
	.w2(32'h3b12cac3),
	.w3(32'hbb6899cf),
	.w4(32'hba5d3819),
	.w5(32'hba87e2e0),
	.w6(32'hba5569be),
	.w7(32'h3b222957),
	.w8(32'h3b899f1b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab66e7f),
	.w1(32'h3a5b3921),
	.w2(32'hba112dd2),
	.w3(32'hbafa3d5a),
	.w4(32'h3a3620d8),
	.w5(32'hbb20d10d),
	.w6(32'h3aa50101),
	.w7(32'h3b0cf82c),
	.w8(32'hba9cc7b5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31b08d),
	.w1(32'hbb9a8040),
	.w2(32'h3b9ebceb),
	.w3(32'h3b8387cd),
	.w4(32'h3c845a47),
	.w5(32'hbab09417),
	.w6(32'hbb014aa8),
	.w7(32'h3c936bac),
	.w8(32'hb88f6649),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9cb5c),
	.w1(32'h3b61adb7),
	.w2(32'h37ab92d4),
	.w3(32'hbaa41cca),
	.w4(32'hbb926cd7),
	.w5(32'hbad68188),
	.w6(32'h3b77e0a1),
	.w7(32'h391f1dff),
	.w8(32'hbb343347),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac91452),
	.w1(32'hbc22c219),
	.w2(32'h3c3730a4),
	.w3(32'hbbdaa1ac),
	.w4(32'h3c1c9885),
	.w5(32'h3b7fe533),
	.w6(32'hbc005892),
	.w7(32'h3c323e48),
	.w8(32'h3b96691d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4902e3),
	.w1(32'hba92785f),
	.w2(32'h3c001f8e),
	.w3(32'hba42ac30),
	.w4(32'h3c29402f),
	.w5(32'h3acd5231),
	.w6(32'hbbc7b691),
	.w7(32'h3be134a1),
	.w8(32'h3aa2dd3c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af82e5b),
	.w1(32'h3afd54c7),
	.w2(32'h3b0bfbd2),
	.w3(32'hbaab8fc6),
	.w4(32'hbb234b5e),
	.w5(32'h3b20ba24),
	.w6(32'h3b8a01bc),
	.w7(32'h3aa1d527),
	.w8(32'h3c6738bf),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4ba49),
	.w1(32'hbc28b2e2),
	.w2(32'hba8c5113),
	.w3(32'hbbf4288c),
	.w4(32'hbc6b9aa4),
	.w5(32'h3b9f0080),
	.w6(32'hbb741d3b),
	.w7(32'hbc3ad515),
	.w8(32'h3c0dcc89),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b950859),
	.w1(32'h3b09b180),
	.w2(32'hbb51b8fa),
	.w3(32'hba63791d),
	.w4(32'hbb3642fd),
	.w5(32'hbc5de03c),
	.w6(32'h3b7fef4c),
	.w7(32'hbbbe950c),
	.w8(32'hbc5ab05b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15c1df),
	.w1(32'hbad3b1ec),
	.w2(32'hba87faa4),
	.w3(32'h3abfc915),
	.w4(32'h3b2bef92),
	.w5(32'h3b4b7f39),
	.w6(32'h3c0e09bf),
	.w7(32'h3bcd1b72),
	.w8(32'h3ba47cc7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0829fe),
	.w1(32'h3a7a9b69),
	.w2(32'hbb0bf521),
	.w3(32'h3a3ecc5f),
	.w4(32'hb9cc7f73),
	.w5(32'hbb102893),
	.w6(32'h39932955),
	.w7(32'hbb91d3fa),
	.w8(32'hbb556c4a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95622a),
	.w1(32'hbae9f8c1),
	.w2(32'hba7868d6),
	.w3(32'hbc120e2b),
	.w4(32'hbbc16a80),
	.w5(32'h3c2622ca),
	.w6(32'hb9a660b2),
	.w7(32'h3a9384e1),
	.w8(32'h3c279ddf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5500d),
	.w1(32'h3a1bef5b),
	.w2(32'hbb5dd71a),
	.w3(32'h3bb4e9ce),
	.w4(32'hb8c48ea6),
	.w5(32'hb9dc2323),
	.w6(32'h394d8f8f),
	.w7(32'hbb8d77ab),
	.w8(32'hbb560902),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadd3d5),
	.w1(32'hbadd528e),
	.w2(32'h3a585a6d),
	.w3(32'hbaa535e4),
	.w4(32'hbb050725),
	.w5(32'h3b392131),
	.w6(32'hbb9b139f),
	.w7(32'hbb9967a6),
	.w8(32'h3b773f5d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b3e18),
	.w1(32'h3b3afdd9),
	.w2(32'h3bb1e3fc),
	.w3(32'hbb0bf356),
	.w4(32'h3b85de83),
	.w5(32'h3b9d81f0),
	.w6(32'h3b406515),
	.w7(32'h3b66e696),
	.w8(32'h3c305c28),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998767c),
	.w1(32'hbb99a73c),
	.w2(32'hbc1f6c6b),
	.w3(32'hbb88813f),
	.w4(32'hbb770c9c),
	.w5(32'hbb04bb34),
	.w6(32'h3aa0bc3b),
	.w7(32'hbb9e9255),
	.w8(32'hbb4c2fe4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b674b89),
	.w1(32'h3bc7fa34),
	.w2(32'hb9ec5a93),
	.w3(32'h3b0fdaa0),
	.w4(32'h3bd09f9f),
	.w5(32'hbb823612),
	.w6(32'hba401491),
	.w7(32'h3c4b0cc3),
	.w8(32'hbbbf015a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c9648),
	.w1(32'hb97712bb),
	.w2(32'h3afdaa79),
	.w3(32'hbbbcef05),
	.w4(32'hba5e1322),
	.w5(32'hbbd9d963),
	.w6(32'hbc1e914c),
	.w7(32'hba94cb61),
	.w8(32'hbbdda87f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9010133),
	.w1(32'h3cac2841),
	.w2(32'h3b9afb84),
	.w3(32'h3c711918),
	.w4(32'h3bfdaa27),
	.w5(32'hbc0e5d49),
	.w6(32'h3d1a213b),
	.w7(32'h3c9fc858),
	.w8(32'hbc4fb432),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6abaea),
	.w1(32'h3b9feeda),
	.w2(32'hbb02f5a6),
	.w3(32'h3aec6ce7),
	.w4(32'hbb8981d0),
	.w5(32'hba018045),
	.w6(32'h3b8c9307),
	.w7(32'hbb34c84c),
	.w8(32'hb934125f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71e357),
	.w1(32'h3bb630dd),
	.w2(32'h3b808787),
	.w3(32'h3b3cf297),
	.w4(32'h3be1fa5d),
	.w5(32'h3b0d22a1),
	.w6(32'h3c416108),
	.w7(32'h3bffe9e3),
	.w8(32'h3ae3def9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f6d09),
	.w1(32'h3acd8606),
	.w2(32'hba84cd7d),
	.w3(32'h3adf0307),
	.w4(32'hbb95a37f),
	.w5(32'hbb094185),
	.w6(32'h3af44de3),
	.w7(32'hbbbf535c),
	.w8(32'h39eb6e59),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0a8d8),
	.w1(32'hbab3049f),
	.w2(32'hbb20fca4),
	.w3(32'hbab49947),
	.w4(32'hbba53181),
	.w5(32'h3a5d1a05),
	.w6(32'hbb40745a),
	.w7(32'hba8bf2ce),
	.w8(32'hbb71b501),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2020d7),
	.w1(32'h3bec476d),
	.w2(32'hbab29ab2),
	.w3(32'h3b992f96),
	.w4(32'hbb518234),
	.w5(32'hbad40cc2),
	.w6(32'h3ab3cd08),
	.w7(32'h3b31de4a),
	.w8(32'hbb40db00),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39c6ef),
	.w1(32'hbc14d6ec),
	.w2(32'h3bcaae06),
	.w3(32'h39fd66bb),
	.w4(32'h3cad4057),
	.w5(32'hba9b6817),
	.w6(32'hbc0fbab5),
	.w7(32'h3c8e1b0a),
	.w8(32'hbb1a1965),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac334fb),
	.w1(32'hbb3c0e36),
	.w2(32'hb935cbd4),
	.w3(32'hbbf69212),
	.w4(32'hbb24ad73),
	.w5(32'h3b6a7c0a),
	.w6(32'hbbd497e4),
	.w7(32'h3b7c2a96),
	.w8(32'h3b61b3a5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b026d65),
	.w1(32'h3bb26691),
	.w2(32'hba796260),
	.w3(32'hba4c4a72),
	.w4(32'hbac13b53),
	.w5(32'hbb0973f9),
	.w6(32'hbaf0626f),
	.w7(32'hbb3930fb),
	.w8(32'hbc321e8c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57e862),
	.w1(32'h3c403db9),
	.w2(32'h3bbb5010),
	.w3(32'h3b2654e8),
	.w4(32'h3c6d6b4c),
	.w5(32'hbb1eb458),
	.w6(32'h3bdbce41),
	.w7(32'h3ca95866),
	.w8(32'hb8f57e6b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbce2d0),
	.w1(32'hbb22dcf6),
	.w2(32'h3c0ce9b3),
	.w3(32'h3be59aea),
	.w4(32'h3bdd9126),
	.w5(32'h3c7a67cc),
	.w6(32'h3bae6d28),
	.w7(32'h3c5ba755),
	.w8(32'h3c351686),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f8a2a),
	.w1(32'hbb3c54ea),
	.w2(32'h3cb21026),
	.w3(32'h3c5bfe6b),
	.w4(32'hbc5c9523),
	.w5(32'hbb99e2ed),
	.w6(32'h3c07cfc1),
	.w7(32'h3a723bda),
	.w8(32'hbb42d9c0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae53598),
	.w1(32'h3c1b9360),
	.w2(32'hbb03a9e2),
	.w3(32'h3b4cd338),
	.w4(32'hbb44433f),
	.w5(32'h3ae1ede6),
	.w6(32'h3c303713),
	.w7(32'hbb6c9bc1),
	.w8(32'h3bfdcabf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eb332),
	.w1(32'h3a9ed37d),
	.w2(32'h3bb1f933),
	.w3(32'h3af25251),
	.w4(32'h3b2c16a7),
	.w5(32'h3b5fa43f),
	.w6(32'h3c01c4dd),
	.w7(32'h3a6d8865),
	.w8(32'hbb5516e2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60ed7d),
	.w1(32'hbbfc8dd8),
	.w2(32'hbb091312),
	.w3(32'hbbc99128),
	.w4(32'hb9ffa0c6),
	.w5(32'h3ba5a040),
	.w6(32'hbc559e00),
	.w7(32'hbbe37428),
	.w8(32'hbbc61ff6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc599d00),
	.w1(32'hbb5284bd),
	.w2(32'h3c1e6f73),
	.w3(32'h3ca0830c),
	.w4(32'h3c16641e),
	.w5(32'hbb188997),
	.w6(32'h3cd9c9ec),
	.w7(32'h3cc0e1f8),
	.w8(32'hbb9c0a85),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadada4f),
	.w1(32'hbc082b0e),
	.w2(32'hbb35f663),
	.w3(32'hbbed90da),
	.w4(32'hbae97489),
	.w5(32'hba7ce342),
	.w6(32'hbb811fb4),
	.w7(32'h3b1c113e),
	.w8(32'h3b400897),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb125c8),
	.w1(32'h3baf6a37),
	.w2(32'hbc37a225),
	.w3(32'h3bf507b5),
	.w4(32'h3b6ddb32),
	.w5(32'h3bcc82aa),
	.w6(32'h3b14c4af),
	.w7(32'hbc29645a),
	.w8(32'h3c6e03a7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb837675d),
	.w1(32'hbbd53388),
	.w2(32'hbb886a4f),
	.w3(32'h3bc52bc6),
	.w4(32'hbb69d914),
	.w5(32'h3b8f5c1e),
	.w6(32'h3b0ea472),
	.w7(32'hbba6aa79),
	.w8(32'h3c0850ed),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c95c9),
	.w1(32'hbc6cc075),
	.w2(32'h3c1554f8),
	.w3(32'hbc1adb03),
	.w4(32'hbb7d8881),
	.w5(32'h3aceee51),
	.w6(32'hbc3baa3b),
	.w7(32'h3ac66d68),
	.w8(32'h3bc041a2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f9075),
	.w1(32'hba5c1dab),
	.w2(32'h3b89673d),
	.w3(32'hb90b0187),
	.w4(32'h3b3f5560),
	.w5(32'hbb323de6),
	.w6(32'h3a5655bd),
	.w7(32'h3c0e3c93),
	.w8(32'hbc365d53),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bdf4d),
	.w1(32'hbb83fa82),
	.w2(32'h3c8e2757),
	.w3(32'h3bb9fbf7),
	.w4(32'hbb8e94c4),
	.w5(32'h3b9397cd),
	.w6(32'h3c9ab553),
	.w7(32'h3c6fa5c4),
	.w8(32'hbb8abbaf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ba2ab),
	.w1(32'hbc2ad606),
	.w2(32'h3abbb23a),
	.w3(32'hba8831d6),
	.w4(32'hbb4064f8),
	.w5(32'h3bc36a0e),
	.w6(32'hbc7c8a5b),
	.w7(32'hbbd84c86),
	.w8(32'h3bdc5f56),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1afc95),
	.w1(32'h3a3a3df7),
	.w2(32'hbbe1150c),
	.w3(32'h3b95ce9b),
	.w4(32'hbba7a180),
	.w5(32'hbbbd0dbb),
	.w6(32'h3bb1c986),
	.w7(32'hbaf4b40f),
	.w8(32'hba8e5926),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49b1f5),
	.w1(32'h3a82888a),
	.w2(32'hba239437),
	.w3(32'h3acd93cc),
	.w4(32'h3aeee553),
	.w5(32'hbaaf9651),
	.w6(32'h3bd12c63),
	.w7(32'h3acd1476),
	.w8(32'hbb3d680e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70e356),
	.w1(32'hba18dc26),
	.w2(32'hbaaf5f95),
	.w3(32'h3a0f8f3d),
	.w4(32'h3b57acd0),
	.w5(32'h3a3c3035),
	.w6(32'h3b8488f8),
	.w7(32'h3b41d7df),
	.w8(32'h3a254d83),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadedfa0),
	.w1(32'hba050c44),
	.w2(32'hbc068996),
	.w3(32'hbac5a1c4),
	.w4(32'hbbbc6cbe),
	.w5(32'h38bfde0f),
	.w6(32'hbb0e5ad6),
	.w7(32'hbb3760ad),
	.w8(32'hbc1d5469),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb000f93),
	.w1(32'h3cb2e92d),
	.w2(32'h3cd8f63a),
	.w3(32'h3c12674f),
	.w4(32'h3ca9016e),
	.w5(32'hbadc7f5c),
	.w6(32'h3cada6fd),
	.w7(32'h3d1b02e4),
	.w8(32'h3bd408d9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcc933),
	.w1(32'h3b5139f1),
	.w2(32'hbbbfe72f),
	.w3(32'hbb179a8d),
	.w4(32'hbc0fddb4),
	.w5(32'h3b1a8075),
	.w6(32'h3b8ba2e6),
	.w7(32'hbb6e83f6),
	.w8(32'h3b71a906),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f39df),
	.w1(32'h3c2ce621),
	.w2(32'h3afe1ef2),
	.w3(32'h3baf05b7),
	.w4(32'h3b6e1a97),
	.w5(32'hb9977b37),
	.w6(32'h3b4317e4),
	.w7(32'hbb5bc890),
	.w8(32'h38615994),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1761ac),
	.w1(32'h3b8b8cb9),
	.w2(32'hbc163ef6),
	.w3(32'hba5d9e01),
	.w4(32'hbadddc41),
	.w5(32'h3bc31647),
	.w6(32'h3c85ec04),
	.w7(32'hbc2209b4),
	.w8(32'h3c5765e3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c032020),
	.w1(32'h3b7abe86),
	.w2(32'hbacabcdf),
	.w3(32'h38723af9),
	.w4(32'hbba00059),
	.w5(32'h3bc90574),
	.w6(32'h3c0df4f2),
	.w7(32'hbb57958e),
	.w8(32'h3bcbfd0a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bef70),
	.w1(32'h3b820641),
	.w2(32'h3ac5696b),
	.w3(32'h378cc92e),
	.w4(32'h39b7aae3),
	.w5(32'h3b08331d),
	.w6(32'hb985982b),
	.w7(32'hbae13bc4),
	.w8(32'h3bf3bf58),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2b719),
	.w1(32'h39e6d5f2),
	.w2(32'hbb0d3e2b),
	.w3(32'hbbc2b288),
	.w4(32'hbbafc5d7),
	.w5(32'h3bea0896),
	.w6(32'h3acb3c42),
	.w7(32'hba0fd650),
	.w8(32'h3bd8ef5f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26b831),
	.w1(32'h3b0e2764),
	.w2(32'h3b83116f),
	.w3(32'h3b3c0f30),
	.w4(32'h3b8d766e),
	.w5(32'h3b86e5f8),
	.w6(32'hbb1fe084),
	.w7(32'hba598784),
	.w8(32'h3b2c57a7),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fd3f5),
	.w1(32'h3a1d6f40),
	.w2(32'hba9114c0),
	.w3(32'h3acb94f8),
	.w4(32'h3b8a88ab),
	.w5(32'h3b4c00e3),
	.w6(32'hbb141889),
	.w7(32'hbb2126e5),
	.w8(32'h3b9b24c0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ef326),
	.w1(32'h3a7dee6f),
	.w2(32'hbad38a29),
	.w3(32'hba6fdcb8),
	.w4(32'hbb4cfcb6),
	.w5(32'h3bae30e2),
	.w6(32'hbac84af2),
	.w7(32'hbb0396e2),
	.w8(32'h3c14719f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be66768),
	.w1(32'h3b69c3b4),
	.w2(32'h3c8d0aa5),
	.w3(32'h3b0084fd),
	.w4(32'h3c3c885d),
	.w5(32'hba81ddf8),
	.w6(32'hbbae35f0),
	.w7(32'h3ca5e8f6),
	.w8(32'h3739a675),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81f9a3),
	.w1(32'h3a6a2ef0),
	.w2(32'hbc10f54e),
	.w3(32'hb879c9d9),
	.w4(32'h3c000ae0),
	.w5(32'hbc2feb80),
	.w6(32'hbae72ce9),
	.w7(32'hbb783a58),
	.w8(32'hbc02d661),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0f2b8),
	.w1(32'h3c39647f),
	.w2(32'h3a26e2e8),
	.w3(32'hbc0b2ebe),
	.w4(32'h3bf60964),
	.w5(32'hbbb96713),
	.w6(32'h3c0c1e8b),
	.w7(32'h3cad26b2),
	.w8(32'hbc0c4d75),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ab287),
	.w1(32'hbb8c46dd),
	.w2(32'h3bb95642),
	.w3(32'hbab6c389),
	.w4(32'h3b727f5d),
	.w5(32'hbb981365),
	.w6(32'hbaafe70a),
	.w7(32'h3c6ae5a5),
	.w8(32'hbbc17547),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10f1e4),
	.w1(32'hbc27abd0),
	.w2(32'hbb31dc9b),
	.w3(32'hbb81bb2e),
	.w4(32'h3c5b55c3),
	.w5(32'hbbacbb4f),
	.w6(32'hbc7db093),
	.w7(32'h3becd1e9),
	.w8(32'hbc4a57ae),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84e035),
	.w1(32'hbb785686),
	.w2(32'h3bdabfd2),
	.w3(32'h3c75260f),
	.w4(32'hbc0d5635),
	.w5(32'h3be1930a),
	.w6(32'h3cdc390c),
	.w7(32'h3b2ae804),
	.w8(32'h3a087221),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac74a21),
	.w1(32'h3c976cfe),
	.w2(32'h3cb70c74),
	.w3(32'h3cb96625),
	.w4(32'h3c74db7d),
	.w5(32'h3947fbd7),
	.w6(32'h3cf40a3b),
	.w7(32'h3cbd6c8d),
	.w8(32'hbaef4db1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda89b5),
	.w1(32'hbc633f08),
	.w2(32'hbbf923ac),
	.w3(32'hbba10eed),
	.w4(32'hbc4dc68a),
	.w5(32'h3a817851),
	.w6(32'h3a65817b),
	.w7(32'hbb8ca024),
	.w8(32'h3b09e23d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1de634),
	.w1(32'h3a658184),
	.w2(32'hbb70af55),
	.w3(32'hbb48a1a0),
	.w4(32'hbbec7c1f),
	.w5(32'hb98075eb),
	.w6(32'hba8fbcd3),
	.w7(32'hbb9e5249),
	.w8(32'h3ac4afa3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc074b87),
	.w1(32'h3bc34b41),
	.w2(32'h3a7ef0a2),
	.w3(32'hbb03bcde),
	.w4(32'h3a097da7),
	.w5(32'h3bb5e633),
	.w6(32'h3aafab3f),
	.w7(32'h3b70c15f),
	.w8(32'h3baa0e57),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca76e),
	.w1(32'h3b672fc3),
	.w2(32'hbab3d08c),
	.w3(32'h3ba84815),
	.w4(32'h3b13981e),
	.w5(32'h3b3ba078),
	.w6(32'h3c1fb759),
	.w7(32'h3b2096bb),
	.w8(32'hbb77a122),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7866),
	.w1(32'h3c229bb4),
	.w2(32'h3c1cb1d2),
	.w3(32'h3bcaeb5f),
	.w4(32'h3b8e00cb),
	.w5(32'hbc447af2),
	.w6(32'h3c4db822),
	.w7(32'h3bd8e6a3),
	.w8(32'hbc420e44),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f4c6),
	.w1(32'hbbda8a5f),
	.w2(32'hbbdba274),
	.w3(32'hbba307e8),
	.w4(32'hbbc7292e),
	.w5(32'hbb600c11),
	.w6(32'hbaf72ce0),
	.w7(32'hbb9eb2b6),
	.w8(32'hbc7cd8b7),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42ee45),
	.w1(32'h3c62e339),
	.w2(32'h3c8e25bb),
	.w3(32'h3cb8fabf),
	.w4(32'h3c0e3bfd),
	.w5(32'hbc433910),
	.w6(32'h3d125b2b),
	.w7(32'h3cb58f45),
	.w8(32'hbc7da644),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf50eb9),
	.w1(32'hbbda49b4),
	.w2(32'h3be37026),
	.w3(32'h3a285c84),
	.w4(32'h3b5131cb),
	.w5(32'hbb868116),
	.w6(32'h3c56ffcc),
	.w7(32'h3c627e6e),
	.w8(32'hbc1e0a48),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c038159),
	.w1(32'h3c40799c),
	.w2(32'hbbb94681),
	.w3(32'h3b923d32),
	.w4(32'h3ce1ead9),
	.w5(32'hba656c6f),
	.w6(32'hbac07a01),
	.w7(32'h3c8655f8),
	.w8(32'hbb8f338a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22b50b),
	.w1(32'hbb85e090),
	.w2(32'h39777283),
	.w3(32'hba8e2e0c),
	.w4(32'hba9787e4),
	.w5(32'hba4b0d4f),
	.w6(32'hbb4521bb),
	.w7(32'hba5ba1a0),
	.w8(32'hba76367f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aabcb),
	.w1(32'hb95fe1cb),
	.w2(32'hbbed4cf9),
	.w3(32'h3a0c170a),
	.w4(32'hb993f06e),
	.w5(32'hbbb66860),
	.w6(32'h3a34f1ec),
	.w7(32'hbc1075d9),
	.w8(32'hbc310ac1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c5e5f2),
	.w1(32'hbbea5f47),
	.w2(32'h3c4cc23d),
	.w3(32'hba767ba1),
	.w4(32'h3c1f5549),
	.w5(32'h3c2a13d9),
	.w6(32'hbae2cf0a),
	.w7(32'h3c16bc24),
	.w8(32'h3c217141),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7e6f2),
	.w1(32'h3b4aec7f),
	.w2(32'hbb16a8b6),
	.w3(32'hba4e7651),
	.w4(32'hbb88b139),
	.w5(32'h3bc792ad),
	.w6(32'hbacb0bd2),
	.w7(32'hbbf52adb),
	.w8(32'h3bd318fc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15a426),
	.w1(32'h3c18be32),
	.w2(32'h3b2f29b3),
	.w3(32'h3be9c8a7),
	.w4(32'h3b9fbaeb),
	.w5(32'h3ac1fd42),
	.w6(32'h3c2489e6),
	.w7(32'h3b40740a),
	.w8(32'h3a88c10d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b582a3a),
	.w1(32'h3b72c6c0),
	.w2(32'hbb59fe55),
	.w3(32'hba5fee69),
	.w4(32'hbb084773),
	.w5(32'hba1f7511),
	.w6(32'h3a36d50d),
	.w7(32'hbb94d604),
	.w8(32'h395ac069),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dd30d),
	.w1(32'hbb9d6454),
	.w2(32'h3b35a65d),
	.w3(32'hbafd2aba),
	.w4(32'hba1794a6),
	.w5(32'h3c007846),
	.w6(32'h3b182949),
	.w7(32'hba0a115a),
	.w8(32'hb91c4d9e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfeacf),
	.w1(32'hbbf683db),
	.w2(32'hbc283b35),
	.w3(32'hbb82315b),
	.w4(32'hbb7f4872),
	.w5(32'h3a2c0f71),
	.w6(32'hbbfc5ad1),
	.w7(32'hbb90b0a0),
	.w8(32'h3b1eb6fb),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dce56),
	.w1(32'hbabc3952),
	.w2(32'h3956f6d5),
	.w3(32'h3b45f98a),
	.w4(32'h3b98c5f0),
	.w5(32'hbb1b9ca3),
	.w6(32'h3b8a3b2c),
	.w7(32'h3bb91451),
	.w8(32'hbc021c4e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fd938),
	.w1(32'h3b78403f),
	.w2(32'h3a985bf3),
	.w3(32'h3b8366a8),
	.w4(32'h3ba5dbbe),
	.w5(32'hbb7c8a52),
	.w6(32'h3ab75616),
	.w7(32'h3bffbc18),
	.w8(32'hbc9386e5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7d97b),
	.w1(32'h3caf695b),
	.w2(32'h3ab85e7a),
	.w3(32'hbaa357e2),
	.w4(32'h3c9f5d89),
	.w5(32'hb879ec6c),
	.w6(32'h3c0fffb1),
	.w7(32'h3ca04545),
	.w8(32'h3ba1f03e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e8d38),
	.w1(32'h3afad0ac),
	.w2(32'hb7210998),
	.w3(32'h3b3af41a),
	.w4(32'h3ba51df0),
	.w5(32'hb933dddd),
	.w6(32'h3ba4a4e8),
	.w7(32'h3b9fb76d),
	.w8(32'hbb4d188e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf32608),
	.w1(32'h3b981d19),
	.w2(32'hbb444bd5),
	.w3(32'hbb7c3cea),
	.w4(32'h3b7b919b),
	.w5(32'h39e67954),
	.w6(32'hbaa17d10),
	.w7(32'h3b14364f),
	.w8(32'hbb892273),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8a15c),
	.w1(32'h3b47ec57),
	.w2(32'h3b8c4437),
	.w3(32'hb925bc0a),
	.w4(32'h3a1c595d),
	.w5(32'h3be5f51f),
	.w6(32'h39343c23),
	.w7(32'hba8b201f),
	.w8(32'hbb54f1f1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c894a4),
	.w1(32'h3c12dc18),
	.w2(32'h3a770541),
	.w3(32'h3c079578),
	.w4(32'h3c439ee8),
	.w5(32'h3bc7196e),
	.w6(32'h3b5773fd),
	.w7(32'h3c491a98),
	.w8(32'h3b3d634b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb037fd),
	.w1(32'h3a868796),
	.w2(32'hbbb1f73a),
	.w3(32'h3a996e92),
	.w4(32'hbb59f27c),
	.w5(32'hbba2893b),
	.w6(32'hbbe5217a),
	.w7(32'hbbdc18d9),
	.w8(32'hbc14fc56),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb98336),
	.w1(32'hbb115d31),
	.w2(32'h3c0387ac),
	.w3(32'hbc11a4fb),
	.w4(32'h3acbe9e6),
	.w5(32'hbbbc93a5),
	.w6(32'hbb6134b7),
	.w7(32'h3c3d490a),
	.w8(32'hbb811983),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf0240),
	.w1(32'hbc286f70),
	.w2(32'hbbcff88d),
	.w3(32'hbb6b1eb1),
	.w4(32'hbbdc3c0e),
	.w5(32'h3ba648df),
	.w6(32'h3aaffbc9),
	.w7(32'hbb28ff1b),
	.w8(32'h3b35b4df),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf554eb),
	.w1(32'hbb4cbe68),
	.w2(32'h3ba9f748),
	.w3(32'h38165701),
	.w4(32'h3bef8c31),
	.w5(32'h3a10eafc),
	.w6(32'hbbc514ec),
	.w7(32'h3c265b5c),
	.w8(32'h3bd8b5ab),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f48e9b),
	.w1(32'hbba3790c),
	.w2(32'hbbde59a6),
	.w3(32'h3af6b7ea),
	.w4(32'h3bc476dc),
	.w5(32'h3aa315d5),
	.w6(32'h3b26c496),
	.w7(32'hba7ff880),
	.w8(32'h3b839949),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b33e2),
	.w1(32'hbb853627),
	.w2(32'h3bb1f42f),
	.w3(32'hbc2cf059),
	.w4(32'hbb9ac353),
	.w5(32'hbb35dd35),
	.w6(32'h3a30a96e),
	.w7(32'h396ae551),
	.w8(32'hba947ee5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17f75f),
	.w1(32'hba530b25),
	.w2(32'hbc2e6583),
	.w3(32'hba86fd39),
	.w4(32'h3c4f9a01),
	.w5(32'h3abd9f65),
	.w6(32'hbbdc8c18),
	.w7(32'h3aad27b0),
	.w8(32'h3b582bac),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3fc99),
	.w1(32'h3ba5b576),
	.w2(32'h3ac2a23c),
	.w3(32'hba7953e2),
	.w4(32'hbb3830b4),
	.w5(32'h3c54920c),
	.w6(32'h3a83714c),
	.w7(32'hbb24e9fb),
	.w8(32'h3b3b5ecc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c6f96),
	.w1(32'h3c007701),
	.w2(32'h3c2203d8),
	.w3(32'h3b915c21),
	.w4(32'h3b5c3491),
	.w5(32'hb9d44027),
	.w6(32'h3c83c71f),
	.w7(32'h3c495469),
	.w8(32'hbb8fc517),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeae5ec),
	.w1(32'hbc2414c3),
	.w2(32'h3be79ad6),
	.w3(32'hbb0c6442),
	.w4(32'h3b52e25b),
	.w5(32'h3b6a2279),
	.w6(32'hbc505ef3),
	.w7(32'h3baefc12),
	.w8(32'h3baf5607),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc155bef),
	.w1(32'hbc615731),
	.w2(32'h3c044394),
	.w3(32'hbc5ee42d),
	.w4(32'h3b0512a3),
	.w5(32'h3af75207),
	.w6(32'hbb3a03e9),
	.w7(32'h3c179452),
	.w8(32'h3c862bc9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0068c6),
	.w1(32'h3b2efcbf),
	.w2(32'hbc0ee26b),
	.w3(32'h3bf9dd0c),
	.w4(32'hbaf2739a),
	.w5(32'hbb388ff1),
	.w6(32'h3ce769b0),
	.w7(32'hbbedf788),
	.w8(32'hbbab70ca),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3da65),
	.w1(32'hbc779781),
	.w2(32'hbc82b3b2),
	.w3(32'hbb8becf0),
	.w4(32'hbc99599e),
	.w5(32'hbb7ff2c8),
	.w6(32'hb9af46ac),
	.w7(32'hbc7f4e60),
	.w8(32'hbbd6ac9d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03d7fd),
	.w1(32'hb85fe61c),
	.w2(32'h3afce50c),
	.w3(32'hba017260),
	.w4(32'h3b05f72f),
	.w5(32'h3c0ff993),
	.w6(32'h3af59c96),
	.w7(32'hba8d6e8f),
	.w8(32'h3c0ea698),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d63a66),
	.w1(32'hb8bc1b30),
	.w2(32'hbb493d60),
	.w3(32'h3c4597b5),
	.w4(32'hbbe09a4d),
	.w5(32'h3b010c47),
	.w6(32'h3bec2008),
	.w7(32'hbc2db0d6),
	.w8(32'hbb8c5278),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4f7d0),
	.w1(32'h3bd71d22),
	.w2(32'hb95c2641),
	.w3(32'h3aac8598),
	.w4(32'h3b5fcfe2),
	.w5(32'h3a67d233),
	.w6(32'h3a6253a2),
	.w7(32'h3bfaf7d1),
	.w8(32'h3b220d70),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4574ca),
	.w1(32'h3c9a1191),
	.w2(32'h3bebd380),
	.w3(32'h3ba44de8),
	.w4(32'h3c179580),
	.w5(32'h3aebbc5f),
	.w6(32'h3d0a5ae7),
	.w7(32'h3c6992d1),
	.w8(32'hbada8863),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ae435),
	.w1(32'h39ee42e5),
	.w2(32'hbaaa82d0),
	.w3(32'h3b277565),
	.w4(32'h3b16b78e),
	.w5(32'h3bc557b5),
	.w6(32'hb9c1bbca),
	.w7(32'h3a9270cd),
	.w8(32'h3b11b8ca),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae204c2),
	.w1(32'h3a42a194),
	.w2(32'h3aa9ec5a),
	.w3(32'h3bf7e51a),
	.w4(32'h3beee0a9),
	.w5(32'h391c7b9c),
	.w6(32'h3a596e50),
	.w7(32'hbb7cbc91),
	.w8(32'h3bbd3b1a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8915ae),
	.w1(32'hb954b6b2),
	.w2(32'h3a89fffd),
	.w3(32'hbae729c7),
	.w4(32'hbb3f789b),
	.w5(32'h3939928c),
	.w6(32'hbaf8ac5e),
	.w7(32'hbb5e199c),
	.w8(32'hbb4fc9af),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399963b3),
	.w1(32'h3b658601),
	.w2(32'h3b1cbd04),
	.w3(32'hbb4f4aa9),
	.w4(32'hbae9b371),
	.w5(32'h39906daa),
	.w6(32'h3a281412),
	.w7(32'hbb4d1ea6),
	.w8(32'hbac36d42),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabccfc2),
	.w1(32'hbb849b86),
	.w2(32'h3c261828),
	.w3(32'hbac1b0fd),
	.w4(32'h3a799c3c),
	.w5(32'h3c1eb23e),
	.w6(32'hbb5bec50),
	.w7(32'h3b5fb8fd),
	.w8(32'h3c1777a9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c5a9),
	.w1(32'hbb0cc614),
	.w2(32'hbb74117a),
	.w3(32'h3bf42a02),
	.w4(32'h3b81ff5b),
	.w5(32'hbb03ea7d),
	.w6(32'hbb899e52),
	.w7(32'h3b438cf3),
	.w8(32'hb7804c16),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4cdb08),
	.w1(32'h3bfc7a47),
	.w2(32'h3a86a8ed),
	.w3(32'hb90475a2),
	.w4(32'h3c3e8f2c),
	.w5(32'hba967682),
	.w6(32'hbb4f36c0),
	.w7(32'h3b5e9223),
	.w8(32'h3c0a98d0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce2cdc),
	.w1(32'h398af41a),
	.w2(32'hbadf2768),
	.w3(32'h3ad1a897),
	.w4(32'h3b9791d5),
	.w5(32'h3b84a624),
	.w6(32'h3bb40de7),
	.w7(32'hb976ac3b),
	.w8(32'h3b4b3018),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae92280),
	.w1(32'hbc1a1e01),
	.w2(32'hbb3fc72b),
	.w3(32'hbabb28cb),
	.w4(32'h3b833314),
	.w5(32'h3b08903c),
	.w6(32'h3b636bda),
	.w7(32'h3bb29fd3),
	.w8(32'hb7d4c439),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb881ce89),
	.w1(32'h3a8aa6a6),
	.w2(32'h3ab23322),
	.w3(32'h3acc2747),
	.w4(32'h3ab1a6b3),
	.w5(32'hba22faa6),
	.w6(32'h3a0ea058),
	.w7(32'hb9213215),
	.w8(32'hbba9044c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d63ae),
	.w1(32'hbbba7574),
	.w2(32'hbb7d7fd1),
	.w3(32'hbb2f9ed3),
	.w4(32'hbb267ce6),
	.w5(32'hb9bc3412),
	.w6(32'hbbab5165),
	.w7(32'hbaafb5e0),
	.w8(32'h3a4200dc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e7a4d),
	.w1(32'hba80ae96),
	.w2(32'hbb150773),
	.w3(32'h3a116ce1),
	.w4(32'h39080103),
	.w5(32'hbaf6b328),
	.w6(32'h39b2a89d),
	.w7(32'hbabfc7c8),
	.w8(32'hbbae532d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f6274),
	.w1(32'hbb99cff0),
	.w2(32'hbac5799b),
	.w3(32'hbaaf57af),
	.w4(32'hba9e5f5b),
	.w5(32'h395b067c),
	.w6(32'hbafc9464),
	.w7(32'hba8aff94),
	.w8(32'h381809c1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba75233),
	.w1(32'h3af745b3),
	.w2(32'h3ba56d3c),
	.w3(32'hbad06ce3),
	.w4(32'h3b851118),
	.w5(32'hba6dda4c),
	.w6(32'hb9e60260),
	.w7(32'h3b2c8f28),
	.w8(32'hbaceaf36),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f8541),
	.w1(32'hbbadf4ac),
	.w2(32'h39818708),
	.w3(32'hbb325ec9),
	.w4(32'h3ad1a9e3),
	.w5(32'h3a9ccae7),
	.w6(32'hbaeabd17),
	.w7(32'h3b29ee30),
	.w8(32'h3b953409),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b671),
	.w1(32'h3ac50121),
	.w2(32'h3bb10131),
	.w3(32'hbb2fe45a),
	.w4(32'hba25f677),
	.w5(32'h3acafa5b),
	.w6(32'h3b8604be),
	.w7(32'h3b0a0b9d),
	.w8(32'h3c1b0025),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab86508),
	.w1(32'h3b16216c),
	.w2(32'hbb0a00df),
	.w3(32'h3b878c02),
	.w4(32'hbb02f537),
	.w5(32'h3afa8654),
	.w6(32'h3c164ae6),
	.w7(32'hbb77549a),
	.w8(32'hbac57129),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ace81),
	.w1(32'h3ababadb),
	.w2(32'h3b123a44),
	.w3(32'hbb655b17),
	.w4(32'hba6d8a2d),
	.w5(32'h3a889479),
	.w6(32'hbb4df18c),
	.w7(32'hbb946603),
	.w8(32'hba977ff6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a8720),
	.w1(32'hbab3843f),
	.w2(32'hbaaaef92),
	.w3(32'h3ae1af25),
	.w4(32'h3acab1e0),
	.w5(32'h3b92afcc),
	.w6(32'hba1de2c5),
	.w7(32'hba33a029),
	.w8(32'h3b2b1eb9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80af9d),
	.w1(32'h3b71dff8),
	.w2(32'hba81817e),
	.w3(32'h3bbad2f8),
	.w4(32'h3bbd772a),
	.w5(32'h3c067777),
	.w6(32'h3b8eb69e),
	.w7(32'h3a223819),
	.w8(32'h3b6e94bd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5a3ff),
	.w1(32'h3b4847cb),
	.w2(32'h3bae1581),
	.w3(32'h3c100498),
	.w4(32'h3bccf403),
	.w5(32'h3b72c534),
	.w6(32'h3be335b5),
	.w7(32'h3beb188b),
	.w8(32'h3b168ce1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b9ab4),
	.w1(32'h3a4ed8c3),
	.w2(32'hbaeb03e3),
	.w3(32'h3b9d46ed),
	.w4(32'h3acbaf61),
	.w5(32'h3b1e909c),
	.w6(32'hbb56d01f),
	.w7(32'h3b417d40),
	.w8(32'h3b741f53),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38575f53),
	.w1(32'h3b1a0ea6),
	.w2(32'h3ac72b04),
	.w3(32'hbac8401f),
	.w4(32'h3b13a964),
	.w5(32'hbad7ca53),
	.w6(32'hbafd4afa),
	.w7(32'h3b05143f),
	.w8(32'h38fbcdd7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3033de),
	.w1(32'hbb99fb50),
	.w2(32'hbb9f5ac7),
	.w3(32'hbb918f55),
	.w4(32'hbaeed373),
	.w5(32'hba2ef543),
	.w6(32'h39c45733),
	.w7(32'hbb467e25),
	.w8(32'h3c9a4017),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aede1),
	.w1(32'hbbd32737),
	.w2(32'hbaeb3c30),
	.w3(32'hbbde4dcc),
	.w4(32'hbbabffa7),
	.w5(32'hbbbd5759),
	.w6(32'h3c963237),
	.w7(32'h3c6c4819),
	.w8(32'hbb711f2f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f6dc1),
	.w1(32'h3a3819aa),
	.w2(32'hbb1357dc),
	.w3(32'hbb67b173),
	.w4(32'h3ad6cb8e),
	.w5(32'hbad3def5),
	.w6(32'hbb967763),
	.w7(32'hbb87cbde),
	.w8(32'h3c6fb53a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d97d68),
	.w1(32'h3ae493bd),
	.w2(32'h3b9f358b),
	.w3(32'hbc21c4b2),
	.w4(32'hbb8c6d1f),
	.w5(32'h3a3f05be),
	.w6(32'h3c3aa324),
	.w7(32'h3bb9ea15),
	.w8(32'hbb1187a0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dae1a2),
	.w1(32'h3b31fd26),
	.w2(32'h3c11803d),
	.w3(32'hb92239b7),
	.w4(32'h3a57c0bf),
	.w5(32'h3c03a0d6),
	.w6(32'h3aabd369),
	.w7(32'h3ae304bc),
	.w8(32'h3c1d4adc),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3d909),
	.w1(32'h3aa92b97),
	.w2(32'h3a0bcff9),
	.w3(32'h38975a75),
	.w4(32'h3a927258),
	.w5(32'h3af0e68e),
	.w6(32'h3b087541),
	.w7(32'h3a2faf29),
	.w8(32'h3b3d8ee3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c7a1b),
	.w1(32'h3ba23961),
	.w2(32'h3b8f6537),
	.w3(32'h3a5b2632),
	.w4(32'h3b991027),
	.w5(32'h3b2ee347),
	.w6(32'h3a1c0a48),
	.w7(32'h3b90a5ff),
	.w8(32'h3b8a0389),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule