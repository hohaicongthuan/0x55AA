module layer_10_featuremap_167(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35090368),
	.w1(32'hb607194a),
	.w2(32'hb50379ec),
	.w3(32'hb4de0e47),
	.w4(32'hb60da484),
	.w5(32'hb60435e1),
	.w6(32'h34953e00),
	.w7(32'h35395342),
	.w8(32'h35fba3a8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e65ca),
	.w1(32'h3964adb3),
	.w2(32'h385fc0c2),
	.w3(32'h38904972),
	.w4(32'h38e3bb82),
	.w5(32'h3894a052),
	.w6(32'hb8a50bad),
	.w7(32'h369d3a1a),
	.w8(32'h3841341d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35625c26),
	.w1(32'h355cb32b),
	.w2(32'h34c5dc70),
	.w3(32'hb3a04bd2),
	.w4(32'hb43daab0),
	.w5(32'hb5ab0f42),
	.w6(32'h3498a1a1),
	.w7(32'hb300388a),
	.w8(32'h34d2cec6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d3442d),
	.w1(32'h36369841),
	.w2(32'h386b2bcc),
	.w3(32'hb72f29cf),
	.w4(32'h364752ea),
	.w5(32'h366098a0),
	.w6(32'hb6baf6c7),
	.w7(32'hb73780ca),
	.w8(32'hb8ada04b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36407040),
	.w1(32'h36a24164),
	.w2(32'h368674bc),
	.w3(32'h3482108f),
	.w4(32'h368bec06),
	.w5(32'h3684cd50),
	.w6(32'hb648f213),
	.w7(32'h35c61285),
	.w8(32'h36559df8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ac90ca),
	.w1(32'h3613b6c2),
	.w2(32'h3556ceb9),
	.w3(32'hb4ccd5dc),
	.w4(32'h363b88e4),
	.w5(32'h34d50ad0),
	.w6(32'h35a1211d),
	.w7(32'h36969aaa),
	.w8(32'h3686eccf),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a82012),
	.w1(32'hb917b741),
	.w2(32'h38acac0a),
	.w3(32'hb9241caa),
	.w4(32'hb92f41ca),
	.w5(32'h38f38883),
	.w6(32'hb952a612),
	.w7(32'hb94858ec),
	.w8(32'h38018da8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60cc381),
	.w1(32'h38637c5f),
	.w2(32'h392ac318),
	.w3(32'h39e64689),
	.w4(32'h39a957cc),
	.w5(32'hb8ab34ea),
	.w6(32'h39c4e935),
	.w7(32'h39d057dc),
	.w8(32'h3987468d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3815c047),
	.w1(32'h3883c060),
	.w2(32'h3852fbf9),
	.w3(32'h36c523e2),
	.w4(32'h37864d03),
	.w5(32'h37d1a3ea),
	.w6(32'hb8c355be),
	.w7(32'h372ce949),
	.w8(32'h385871a5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9000bf7),
	.w1(32'hb7f45682),
	.w2(32'h3a1dd945),
	.w3(32'h39bd9322),
	.w4(32'h39d707e9),
	.w5(32'h39b1c684),
	.w6(32'h3a6f5402),
	.w7(32'h3a6882f0),
	.w8(32'h397399d5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79ad655),
	.w1(32'hb7381823),
	.w2(32'hb7826dbd),
	.w3(32'hb79cccf4),
	.w4(32'hb797e875),
	.w5(32'hb78ed924),
	.w6(32'hb7b24aed),
	.w7(32'hb6ca0faa),
	.w8(32'h37bc3bd7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb10b1),
	.w1(32'hb9d4ef7e),
	.w2(32'hb985d68a),
	.w3(32'hb8c4fb42),
	.w4(32'hb94c4073),
	.w5(32'h39006078),
	.w6(32'hb90b58f2),
	.w7(32'hb92faa1a),
	.w8(32'h38f1d044),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d51ce),
	.w1(32'hb9b92cc7),
	.w2(32'h39e0c118),
	.w3(32'h383c5146),
	.w4(32'h3a08e256),
	.w5(32'h3a11ad6d),
	.w6(32'h3a87bdce),
	.w7(32'h3ab82b7b),
	.w8(32'h3a30da98),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905c7c0),
	.w1(32'h37c37101),
	.w2(32'h38692644),
	.w3(32'h3911a2d4),
	.w4(32'h382a932f),
	.w5(32'hb8ff29c3),
	.w6(32'h38af0bb6),
	.w7(32'h39294f29),
	.w8(32'h38d0128b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db342a),
	.w1(32'hb901534b),
	.w2(32'hb9127af6),
	.w3(32'hb9232945),
	.w4(32'hb9606e0d),
	.w5(32'hb988ebbc),
	.w6(32'hb897a54b),
	.w7(32'hb8d882fd),
	.w8(32'hb94467f3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c66696),
	.w1(32'h391bb17b),
	.w2(32'h39ffa436),
	.w3(32'h38286cce),
	.w4(32'h3963c24a),
	.w5(32'h39c63fab),
	.w6(32'h3a1ab4af),
	.w7(32'h3a1edb4a),
	.w8(32'h39a6ddc1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368b5518),
	.w1(32'hb6164330),
	.w2(32'hb783a4cf),
	.w3(32'h36b8d0c4),
	.w4(32'hb7539a9f),
	.w5(32'h36061205),
	.w6(32'h377e4d1d),
	.w7(32'h346c518c),
	.w8(32'hb60bcd60),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25e5e0),
	.w1(32'hba05374a),
	.w2(32'h398311e8),
	.w3(32'hb8e7f0f7),
	.w4(32'hb8a0c1b7),
	.w5(32'hb7b0ac2c),
	.w6(32'h39c93a50),
	.w7(32'h38b66db3),
	.w8(32'hb8742ced),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984238a),
	.w1(32'hb80dd9dc),
	.w2(32'h39a99408),
	.w3(32'hb8a246a0),
	.w4(32'h3927ee23),
	.w5(32'h393e30ae),
	.w6(32'h39ee5573),
	.w7(32'h39ff9d1a),
	.w8(32'h398ccc17),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68f6006),
	.w1(32'hb5bb8ba5),
	.w2(32'hb73d3653),
	.w3(32'hb39389e2),
	.w4(32'h36014382),
	.w5(32'hb652bdd1),
	.w6(32'h367f4e37),
	.w7(32'h328dad46),
	.w8(32'hb5d791f8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb696530f),
	.w1(32'hb64eafee),
	.w2(32'hb63176bd),
	.w3(32'hb69bdb1f),
	.w4(32'hb6c95309),
	.w5(32'hb6aecc1d),
	.w6(32'hb589c7c7),
	.w7(32'hb60e1a79),
	.w8(32'hb6cf4db5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3640e413),
	.w1(32'hb83aa2c4),
	.w2(32'hb9262f5e),
	.w3(32'h381f10e0),
	.w4(32'hb70d1cbc),
	.w5(32'hb7c70980),
	.w6(32'h376fc79c),
	.w7(32'hb560eed4),
	.w8(32'h386ba422),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66d02f),
	.w1(32'hb9c9c1a4),
	.w2(32'h39f386c4),
	.w3(32'hba81a6e3),
	.w4(32'hb90dd3a2),
	.w5(32'h39bc4647),
	.w6(32'hb942bf1a),
	.w7(32'hba4aeff4),
	.w8(32'hba48055f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ad978c),
	.w1(32'h38996269),
	.w2(32'h39e1480e),
	.w3(32'h38ae7c5d),
	.w4(32'h3920ca8d),
	.w5(32'h390848d1),
	.w6(32'h39ccf761),
	.w7(32'h39b3e932),
	.w8(32'h387e3b3e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dcb53e),
	.w1(32'hb8a2a2f7),
	.w2(32'hb8b8c3f6),
	.w3(32'h3919b1ef),
	.w4(32'h3986c0d4),
	.w5(32'h3815ab8e),
	.w6(32'h3a0a2b8b),
	.w7(32'h3a071a63),
	.w8(32'h398d1ee3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cb9848),
	.w1(32'hb877513f),
	.w2(32'h382dd4e0),
	.w3(32'h37aeda43),
	.w4(32'hb86c4c6b),
	.w5(32'hb930ef3f),
	.w6(32'h36ca88b7),
	.w7(32'hb8259912),
	.w8(32'hb9a2095c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4ae4389),
	.w1(32'h3519b279),
	.w2(32'hb752c1d0),
	.w3(32'hb6a603e4),
	.w4(32'hb6346445),
	.w5(32'hb6b972d9),
	.w6(32'hb74e9046),
	.w7(32'hb73db060),
	.w8(32'hb6f812f4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8480d3e),
	.w1(32'h391fa539),
	.w2(32'h38d6bad8),
	.w3(32'h386a5212),
	.w4(32'h38e277d8),
	.w5(32'h3962ce38),
	.w6(32'h36e7cc93),
	.w7(32'h385e3961),
	.w8(32'h393eac2f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb771fea6),
	.w1(32'h36d2aed5),
	.w2(32'hb86c59fe),
	.w3(32'h368b0c82),
	.w4(32'hb7c1217b),
	.w5(32'h375088da),
	.w6(32'hb79f66f0),
	.w7(32'hb76657ea),
	.w8(32'h3899b7a2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85593ef),
	.w1(32'h38f40cee),
	.w2(32'h39e49b62),
	.w3(32'h393415e4),
	.w4(32'h39800cea),
	.w5(32'h3922a245),
	.w6(32'h39aca1f8),
	.w7(32'h399ec62b),
	.w8(32'hb8be1ba4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6620bfa),
	.w1(32'h33d1f741),
	.w2(32'hb5924e26),
	.w3(32'hb629befa),
	.w4(32'hb633b510),
	.w5(32'hb68df198),
	.w6(32'h3501c305),
	.w7(32'hb624e2d6),
	.w8(32'hb5e176e9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59c68cd),
	.w1(32'hb72d3602),
	.w2(32'hb6850e38),
	.w3(32'hb6932ce8),
	.w4(32'hb74e1e83),
	.w5(32'hb5cba1ca),
	.w6(32'hb487e418),
	.w7(32'hb6baf813),
	.w8(32'h36f6290e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c519bf),
	.w1(32'h3742fbc4),
	.w2(32'h3944153b),
	.w3(32'hb863b121),
	.w4(32'hb685f374),
	.w5(32'h382d8c74),
	.w6(32'h38d15811),
	.w7(32'h38698116),
	.w8(32'hb880ae5a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aadca9),
	.w1(32'hb7ee6fea),
	.w2(32'hb8c83fc4),
	.w3(32'h373f0476),
	.w4(32'hb7b58476),
	.w5(32'hb8d143be),
	.w6(32'h3768bb34),
	.w7(32'hb80620d2),
	.w8(32'hb8afc528),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c07e65),
	.w1(32'h35a03da7),
	.w2(32'h36ca1e79),
	.w3(32'hb7e92887),
	.w4(32'hb61155f9),
	.w5(32'h3787cc63),
	.w6(32'hb7452699),
	.w7(32'h37ef435d),
	.w8(32'h382a2c50),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb895efe8),
	.w1(32'hb8b949f3),
	.w2(32'h38869a61),
	.w3(32'hb87ad6fb),
	.w4(32'h36ea7248),
	.w5(32'h384c553b),
	.w6(32'h386b19c9),
	.w7(32'h38be124d),
	.w8(32'h38be49db),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2cc3b),
	.w1(32'hb9700069),
	.w2(32'h38c472a1),
	.w3(32'h3937c05d),
	.w4(32'hb8cd2efd),
	.w5(32'h378412bc),
	.w6(32'h39558192),
	.w7(32'h39178f58),
	.w8(32'hb877cef8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b8d4e),
	.w1(32'h38f68f2d),
	.w2(32'hba472f66),
	.w3(32'h386672ac),
	.w4(32'hb8cede17),
	.w5(32'hb980ab82),
	.w6(32'hb99d9bf0),
	.w7(32'hb99778d6),
	.w8(32'h38d08cd6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8800056),
	.w1(32'h38e621d7),
	.w2(32'hb8f0edb0),
	.w3(32'hb91f4e5d),
	.w4(32'hb8806a5a),
	.w5(32'h39613fc5),
	.w6(32'hba58e689),
	.w7(32'hba146029),
	.w8(32'h39072551),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380f976d),
	.w1(32'hb7bf42ea),
	.w2(32'hb8849f22),
	.w3(32'h39272aba),
	.w4(32'h39412a51),
	.w5(32'h38a26cf0),
	.w6(32'h39561b8c),
	.w7(32'h39b26985),
	.w8(32'h39884b0c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72db7c3),
	.w1(32'hb73afb30),
	.w2(32'h36765a8f),
	.w3(32'hb784a495),
	.w4(32'h35d7bd46),
	.w5(32'hb6579206),
	.w6(32'hb77aad61),
	.w7(32'hb68583bf),
	.w8(32'hb690ca02),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e7bbea),
	.w1(32'h3651d9ec),
	.w2(32'hb7e512e0),
	.w3(32'h36a68b00),
	.w4(32'h369b809a),
	.w5(32'hb7c93939),
	.w6(32'h3408eeff),
	.w7(32'hb67b9d97),
	.w8(32'hb7e71a3f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3808cf21),
	.w1(32'h39063c7f),
	.w2(32'hb8947e94),
	.w3(32'h38517b05),
	.w4(32'h39226755),
	.w5(32'h38faae1a),
	.w6(32'h38080d69),
	.w7(32'h391a0018),
	.w8(32'h390ab6ef),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898a686),
	.w1(32'h392e35ac),
	.w2(32'h3a45d377),
	.w3(32'h391a20a4),
	.w4(32'h3a224f85),
	.w5(32'h39fe9d90),
	.w6(32'h3a88adeb),
	.w7(32'h3a41ce5c),
	.w8(32'h3899e0b4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816abdd),
	.w1(32'h381f2866),
	.w2(32'h3953b154),
	.w3(32'hb6e48ac7),
	.w4(32'hb747895c),
	.w5(32'hb873b0b5),
	.w6(32'h3990a7b0),
	.w7(32'h392b1f60),
	.w8(32'hb90c8e8b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a20b1e),
	.w1(32'h38c73325),
	.w2(32'h3a1eaf4e),
	.w3(32'h38db0ef4),
	.w4(32'h395e4ad2),
	.w5(32'h392188e6),
	.w6(32'h3a18d9bf),
	.w7(32'h39fed3e7),
	.w8(32'h388798c3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382c76cd),
	.w1(32'hb88a0294),
	.w2(32'hb8c84029),
	.w3(32'h3899d5b7),
	.w4(32'h3884167e),
	.w5(32'h367a702e),
	.w6(32'h38eff2af),
	.w7(32'h38b4824f),
	.w8(32'h37d6e02c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1494b9),
	.w1(32'hb9d904a0),
	.w2(32'h39d33254),
	.w3(32'hb945601d),
	.w4(32'h397c1018),
	.w5(32'h39881a0d),
	.w6(32'h3a0dd6f7),
	.w7(32'h3a299a55),
	.w8(32'h390e18d3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da5c65),
	.w1(32'hb7f5a67f),
	.w2(32'h37949cbb),
	.w3(32'hb7c62ece),
	.w4(32'h3672ef6a),
	.w5(32'h3797a5f2),
	.w6(32'hb7064dfb),
	.w7(32'h36d3a2e5),
	.w8(32'hb650ee16),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d31a78),
	.w1(32'hb7b526bd),
	.w2(32'h37f71a33),
	.w3(32'h3585d30a),
	.w4(32'hb7db52a2),
	.w5(32'hb8c39bc1),
	.w6(32'hb7a08246),
	.w7(32'hb8fde3d8),
	.w8(32'hb92313fd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb747e472),
	.w1(32'hb816c4d7),
	.w2(32'hb7d83842),
	.w3(32'h378fdc07),
	.w4(32'hb7a32450),
	.w5(32'hb83c8623),
	.w6(32'h37f4070a),
	.w7(32'hb794fcf5),
	.w8(32'hb83c204b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b53dfa),
	.w1(32'hb58c4a10),
	.w2(32'h392ae879),
	.w3(32'h381e347c),
	.w4(32'h3854c6f9),
	.w5(32'h38c7dcf6),
	.w6(32'h398b60ca),
	.w7(32'h399f2508),
	.w8(32'hb85b696d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d2e977),
	.w1(32'hb74c6bdb),
	.w2(32'h37c2ad33),
	.w3(32'h368521ad),
	.w4(32'hb7935e65),
	.w5(32'hb7707321),
	.w6(32'h3797f66e),
	.w7(32'h357dc17c),
	.w8(32'hb6ea5c54),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cef22),
	.w1(32'hb9a99a6b),
	.w2(32'h39fd3fb9),
	.w3(32'hb91d5cb0),
	.w4(32'hb8659f0e),
	.w5(32'h3981e038),
	.w6(32'h3a08c280),
	.w7(32'h3861ba73),
	.w8(32'hb9c59f5b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35834387),
	.w1(32'hb805ecd4),
	.w2(32'hb8888674),
	.w3(32'hb61594d1),
	.w4(32'hb89eef65),
	.w5(32'hb883ccde),
	.w6(32'hb8350412),
	.w7(32'hb89e71fc),
	.w8(32'hb7b292c4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34271689),
	.w1(32'hb6016a63),
	.w2(32'h378eb229),
	.w3(32'h36a52d2a),
	.w4(32'hb649aa74),
	.w5(32'hb80749a9),
	.w6(32'h376b6607),
	.w7(32'hb8103fe1),
	.w8(32'hb8a4cf7c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb58f274b),
	.w1(32'h362e9d58),
	.w2(32'h362a6ec6),
	.w3(32'hb4313145),
	.w4(32'h3637cf82),
	.w5(32'h3559f1cf),
	.w6(32'h365a38ce),
	.w7(32'h364417b9),
	.w8(32'hb528d73f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bb1de4),
	.w1(32'h3723b8e6),
	.w2(32'h37c09570),
	.w3(32'hb65f62c8),
	.w4(32'h37b78bd8),
	.w5(32'h37b1243a),
	.w6(32'hb74ff1e8),
	.w7(32'h3704d16b),
	.w8(32'h37b8fd18),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375bfdbb),
	.w1(32'hb7263a9e),
	.w2(32'hb898e45d),
	.w3(32'h3749df01),
	.w4(32'hb7601fd0),
	.w5(32'hb71ef413),
	.w6(32'hb75ae30a),
	.w7(32'hb73758ef),
	.w8(32'h380a87f2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a2efc9),
	.w1(32'h368c7248),
	.w2(32'h3859a9da),
	.w3(32'h35e9a604),
	.w4(32'h37f41c38),
	.w5(32'h3892580b),
	.w6(32'hb7bb0a2a),
	.w7(32'h3723f791),
	.w8(32'h3862e12a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954b213),
	.w1(32'hb84f39c9),
	.w2(32'h397aa02b),
	.w3(32'h387996ba),
	.w4(32'h39941117),
	.w5(32'h3987cc8f),
	.w6(32'h39f93a4f),
	.w7(32'h39cfb683),
	.w8(32'h3938d468),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9238fe9),
	.w1(32'hb729462e),
	.w2(32'h38bd22e1),
	.w3(32'hb7e92783),
	.w4(32'h38325d58),
	.w5(32'h38931444),
	.w6(32'h39338a5e),
	.w7(32'hb823884f),
	.w8(32'hb9264357),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb665549d),
	.w1(32'hb46f9974),
	.w2(32'hb60f5048),
	.w3(32'h35e7c978),
	.w4(32'h37039fb6),
	.w5(32'h35698582),
	.w6(32'h36f0b5dd),
	.w7(32'h36806dd9),
	.w8(32'hb670e86e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6901d51),
	.w1(32'hb511aef1),
	.w2(32'h33349372),
	.w3(32'hb63122dd),
	.w4(32'hb6ad6de3),
	.w5(32'hb6f0d2a0),
	.w6(32'h352c9437),
	.w7(32'hb60d6ed8),
	.w8(32'hb70a1cf3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4ea19ed),
	.w1(32'h35fa73d5),
	.w2(32'h36ac16b0),
	.w3(32'hb6e7af34),
	.w4(32'hb6c65ece),
	.w5(32'hb50f40c3),
	.w6(32'hb61ebde0),
	.w7(32'h358df1ef),
	.w8(32'h362dba26),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5be1404),
	.w1(32'hb5222ed9),
	.w2(32'hb644aa3e),
	.w3(32'hb4b9864c),
	.w4(32'h360f5cdf),
	.w5(32'h35189f8d),
	.w6(32'hb61ad18f),
	.w7(32'h3616a021),
	.w8(32'h363fd07b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ae210),
	.w1(32'h38586832),
	.w2(32'h38341448),
	.w3(32'h39808754),
	.w4(32'h399f5970),
	.w5(32'h39a835af),
	.w6(32'h39df669a),
	.w7(32'h39c92c10),
	.w8(32'h39333b88),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f1fe4),
	.w1(32'h39bb57a2),
	.w2(32'h39b17ab1),
	.w3(32'h393a62dd),
	.w4(32'h37a4af94),
	.w5(32'hb7622582),
	.w6(32'h371c3ef5),
	.w7(32'hb8a94a22),
	.w8(32'hb7dca278),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e3dc83),
	.w1(32'hb89ce831),
	.w2(32'h37333548),
	.w3(32'hb93779b4),
	.w4(32'hb913a232),
	.w5(32'h3822f026),
	.w6(32'hb91a6a0f),
	.w7(32'hb91e7280),
	.w8(32'h39036038),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38af0356),
	.w1(32'hb893cc49),
	.w2(32'hb9401115),
	.w3(32'hb8936123),
	.w4(32'h39264541),
	.w5(32'h3846125b),
	.w6(32'h39d82fe5),
	.w7(32'h39e04a52),
	.w8(32'h39d95609),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65792b0),
	.w1(32'h34dc1157),
	.w2(32'hb42ad9c2),
	.w3(32'hb63b5f5e),
	.w4(32'h35d7b1cc),
	.w5(32'h348f1709),
	.w6(32'h34ee2458),
	.w7(32'h364cdcb0),
	.w8(32'h353e7da5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4a7952e),
	.w1(32'h35974d30),
	.w2(32'hb5d470ec),
	.w3(32'hb625ace1),
	.w4(32'hb5260f50),
	.w5(32'hb624586d),
	.w6(32'hb61c0bf3),
	.w7(32'hb4ae8815),
	.w8(32'hb485d18d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6087deb),
	.w1(32'h36a26516),
	.w2(32'h35d10d5f),
	.w3(32'h367acbe6),
	.w4(32'h3713e536),
	.w5(32'h36927519),
	.w6(32'h3730e4c3),
	.w7(32'h37085d5f),
	.w8(32'h35eaf737),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a12acf),
	.w1(32'hb80c20f1),
	.w2(32'hb69c9cc8),
	.w3(32'h374cb153),
	.w4(32'h38b0dd80),
	.w5(32'h38913a8c),
	.w6(32'h39020b31),
	.w7(32'h395afc96),
	.w8(32'h394159c2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb681bb8e),
	.w1(32'hb7120b7f),
	.w2(32'hb73b0b79),
	.w3(32'h377a2fbc),
	.w4(32'h37570d31),
	.w5(32'hb69d9743),
	.w6(32'h371fdeb0),
	.w7(32'h371819d0),
	.w8(32'hb765990f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a21d2a),
	.w1(32'hb9a97962),
	.w2(32'hb8c19b58),
	.w3(32'hb9278450),
	.w4(32'hb8a041b8),
	.w5(32'h3893a925),
	.w6(32'h375c7492),
	.w7(32'h38d0720b),
	.w8(32'hb7083712),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e05a20),
	.w1(32'h37475245),
	.w2(32'hb94e47fa),
	.w3(32'hb9242212),
	.w4(32'h39d51c46),
	.w5(32'h39bde0ee),
	.w6(32'h3a0dc998),
	.w7(32'h3a0b0dff),
	.w8(32'h39fad371),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9813d49),
	.w1(32'hb92a092a),
	.w2(32'h389523d3),
	.w3(32'hb8e2cdf7),
	.w4(32'h395e1a33),
	.w5(32'h394638b2),
	.w6(32'h39fb6f93),
	.w7(32'h3a457e9d),
	.w8(32'h39ee51f8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8261780),
	.w1(32'hb702e875),
	.w2(32'h38626ae9),
	.w3(32'hb8a380ff),
	.w4(32'hb887ec69),
	.w5(32'hb8c5a6d7),
	.w6(32'h3822267c),
	.w7(32'hb80c1557),
	.w8(32'hb91e729d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88eca3b),
	.w1(32'hb85626ba),
	.w2(32'h389d2c58),
	.w3(32'h3835ba79),
	.w4(32'h38804816),
	.w5(32'h39327097),
	.w6(32'h38e50d51),
	.w7(32'h39482924),
	.w8(32'h3911c43c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787ef65),
	.w1(32'h38056f92),
	.w2(32'h391a01d0),
	.w3(32'h374e89ff),
	.w4(32'hb7becea6),
	.w5(32'hb83b0a11),
	.w6(32'h391d84aa),
	.w7(32'h378c5f2f),
	.w8(32'hb9066888),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946340a),
	.w1(32'hb912021d),
	.w2(32'h39262177),
	.w3(32'hb927a7c0),
	.w4(32'h388efe9f),
	.w5(32'h39148113),
	.w6(32'h38f7e84c),
	.w7(32'h39c82f58),
	.w8(32'h39846e22),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ba49f2),
	.w1(32'h352f600a),
	.w2(32'hb5a8df15),
	.w3(32'h3512ca98),
	.w4(32'h34c6d468),
	.w5(32'hb53d8883),
	.w6(32'h3285a6e3),
	.w7(32'h34eb90a9),
	.w8(32'h34786f3f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d6692d),
	.w1(32'h3612bc72),
	.w2(32'h36267bb8),
	.w3(32'h353bc72d),
	.w4(32'hb4828573),
	.w5(32'h357ec33e),
	.w6(32'hb205e03a),
	.w7(32'h35e32b7b),
	.w8(32'h36470b68),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4e23f87),
	.w1(32'h3704f170),
	.w2(32'hb308f941),
	.w3(32'hb407f4d2),
	.w4(32'h371a6b22),
	.w5(32'hb3f859bb),
	.w6(32'h3732fe6e),
	.w7(32'h36613d7f),
	.w8(32'hb4fe1f04),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b22cca),
	.w1(32'h36dc656c),
	.w2(32'h3786c2c1),
	.w3(32'h37237224),
	.w4(32'h37fabe89),
	.w5(32'h3806ee45),
	.w6(32'h35d7b52a),
	.w7(32'h37767676),
	.w8(32'h376e37e7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f2b57),
	.w1(32'hb97577f2),
	.w2(32'hb9c61f14),
	.w3(32'hb90bc8d1),
	.w4(32'hb98b0b72),
	.w5(32'hb96c3e55),
	.w6(32'hb8c7e4b7),
	.w7(32'hb9785f63),
	.w8(32'hb9411437),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ef0634),
	.w1(32'hb8555762),
	.w2(32'hb8e4259d),
	.w3(32'hb7f9bb5b),
	.w4(32'hb77362bb),
	.w5(32'hb8759863),
	.w6(32'hb4d5cf37),
	.w7(32'h37284cc4),
	.w8(32'h382299ab),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382be7a1),
	.w1(32'h391a7d62),
	.w2(32'h39863a43),
	.w3(32'h3900e336),
	.w4(32'h39158a8b),
	.w5(32'hb844f5fb),
	.w6(32'h394a7c9b),
	.w7(32'h3934bda0),
	.w8(32'hb8e9b787),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddc91a),
	.w1(32'hba0ef31e),
	.w2(32'hb9a6496d),
	.w3(32'h38ca967f),
	.w4(32'h38613086),
	.w5(32'hb5801df6),
	.w6(32'h3a1ec83f),
	.w7(32'h39f97e91),
	.w8(32'h3906939f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a6dc26),
	.w1(32'hb8bcfded),
	.w2(32'hb923d9d8),
	.w3(32'hb8fa9a8e),
	.w4(32'hb91a229f),
	.w5(32'h375d4339),
	.w6(32'hb9a4f170),
	.w7(32'hb93032ee),
	.w8(32'h3809c798),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8d9a7),
	.w1(32'hb87700c6),
	.w2(32'h393f5f3a),
	.w3(32'h379e0f55),
	.w4(32'h399db683),
	.w5(32'h39dc7f2a),
	.w6(32'hb87f4bdc),
	.w7(32'hb83d530f),
	.w8(32'hb81c0354),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e36012),
	.w1(32'hb8c2ba1d),
	.w2(32'hb92ffd25),
	.w3(32'hb91e16ec),
	.w4(32'hb932c551),
	.w5(32'h3592ee52),
	.w6(32'hb9746123),
	.w7(32'hb8263f1c),
	.w8(32'h39151369),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c3cd4),
	.w1(32'hb95ad1c6),
	.w2(32'hb877e247),
	.w3(32'hb82e6ccd),
	.w4(32'hb93b2406),
	.w5(32'hb9de2c11),
	.w6(32'h390873bd),
	.w7(32'hb9b6055c),
	.w8(32'hba2817e6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b09213),
	.w1(32'h38edb34e),
	.w2(32'h39181347),
	.w3(32'h38af98de),
	.w4(32'h388515d6),
	.w5(32'h36b6dd73),
	.w6(32'hb785a165),
	.w7(32'hb8d2d337),
	.w8(32'hb8d36622),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9637f64),
	.w1(32'hb927eb57),
	.w2(32'hb8ad3e83),
	.w3(32'hb77952e0),
	.w4(32'h391c94fa),
	.w5(32'h38befcb6),
	.w6(32'h3848394e),
	.w7(32'h393bc123),
	.w8(32'hb6a5d22e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b68ac2),
	.w1(32'h377416aa),
	.w2(32'hb7c49714),
	.w3(32'h35b3b901),
	.w4(32'h37911545),
	.w5(32'hb819bb80),
	.w6(32'hb6fce9f0),
	.w7(32'hb7a5990f),
	.w8(32'hb81da11a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b853b),
	.w1(32'hb91ec839),
	.w2(32'h39875aa2),
	.w3(32'h38fdecca),
	.w4(32'h38ca58e3),
	.w5(32'hb8baf0b7),
	.w6(32'h39f8db44),
	.w7(32'h397e6628),
	.w8(32'hb970ccb1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39287753),
	.w1(32'h375d77b8),
	.w2(32'hb8d735bd),
	.w3(32'h37db0f47),
	.w4(32'h38a8a69c),
	.w5(32'h39503656),
	.w6(32'h35d20f95),
	.w7(32'h375757ec),
	.w8(32'h3955ccc8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9261f40),
	.w1(32'hb9c070f1),
	.w2(32'h3648ea16),
	.w3(32'hb9c88fb4),
	.w4(32'hb9b584c6),
	.w5(32'hb9b9da38),
	.w6(32'hb93a1523),
	.w7(32'hb9288c6b),
	.w8(32'hb9a89466),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f847c0),
	.w1(32'hb9ba82b2),
	.w2(32'hba904f6b),
	.w3(32'h370dd219),
	.w4(32'hb93959fd),
	.w5(32'hb9095151),
	.w6(32'hba2d7402),
	.w7(32'hba000df1),
	.w8(32'hb8823fed),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb851ed34),
	.w1(32'h3968993d),
	.w2(32'h3a1145a6),
	.w3(32'h3934d122),
	.w4(32'h3979c257),
	.w5(32'hb7813cf3),
	.w6(32'h3a079d04),
	.w7(32'h39eae83b),
	.w8(32'hb893d216),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912baa1),
	.w1(32'hb95c6279),
	.w2(32'h3992c18a),
	.w3(32'h38c86803),
	.w4(32'h37d397d5),
	.w5(32'h395a2a6d),
	.w6(32'h36cce7fa),
	.w7(32'hb75b7bbc),
	.w8(32'hb84f7b5c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897ee75),
	.w1(32'hb895ffb6),
	.w2(32'hb7fbf6c2),
	.w3(32'h3800350c),
	.w4(32'h362ef5f7),
	.w5(32'hb80adbd2),
	.w6(32'h3897a792),
	.w7(32'h3752b90a),
	.w8(32'hb78d338e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aaf385),
	.w1(32'hba0e0933),
	.w2(32'hba192e65),
	.w3(32'hb8e9daa5),
	.w4(32'hb9a87f1f),
	.w5(32'hba1fce0c),
	.w6(32'hb8e03c26),
	.w7(32'h39360e51),
	.w8(32'hb99f3408),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ec751),
	.w1(32'hb9b55888),
	.w2(32'hb9d99e11),
	.w3(32'hb92307da),
	.w4(32'hb9162a4f),
	.w5(32'hb64d7bb1),
	.w6(32'hb900fe9c),
	.w7(32'h3816a51d),
	.w8(32'h3960e8e8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ce9b7c),
	.w1(32'h37062fce),
	.w2(32'hb50e1567),
	.w3(32'h36bf220c),
	.w4(32'h3656c269),
	.w5(32'h365c0c45),
	.w6(32'h36ba4e3f),
	.w7(32'h368af364),
	.w8(32'h3608d8fd),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8237044),
	.w1(32'h380b7e60),
	.w2(32'h36e9e4a6),
	.w3(32'hb7434fe2),
	.w4(32'hb679e61d),
	.w5(32'hb79be9ae),
	.w6(32'h382a823f),
	.w7(32'h37531878),
	.w8(32'h37ce1655),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9521c90),
	.w1(32'hb762676e),
	.w2(32'h39f54377),
	.w3(32'hb824a39f),
	.w4(32'h39684f1e),
	.w5(32'h395d3455),
	.w6(32'h3a13f102),
	.w7(32'h3a131e94),
	.w8(32'h3908169e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a86d5),
	.w1(32'h3756ab72),
	.w2(32'h399e015d),
	.w3(32'hb73fde1b),
	.w4(32'h38eb558b),
	.w5(32'h3879186f),
	.w6(32'h39c950ba),
	.w7(32'h39bb994a),
	.w8(32'hb854d930),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365e91f4),
	.w1(32'h39155dd3),
	.w2(32'h37947890),
	.w3(32'h385ca9f2),
	.w4(32'h3a0e0603),
	.w5(32'h39e6a055),
	.w6(32'h393f51bb),
	.w7(32'h39ba626c),
	.w8(32'h3996c152),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39718bde),
	.w1(32'h399f25e0),
	.w2(32'h3974dd9a),
	.w3(32'hb69493ca),
	.w4(32'hb82de68a),
	.w5(32'h3880e70d),
	.w6(32'hb998c14c),
	.w7(32'hb981f51c),
	.w8(32'hb9065b55),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90968bf),
	.w1(32'hb90e7571),
	.w2(32'hb9215f1e),
	.w3(32'hb9284e02),
	.w4(32'hb9512b16),
	.w5(32'hb964431a),
	.w6(32'h372884d7),
	.w7(32'hb8814894),
	.w8(32'hb7ca22ea),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb790a59d),
	.w1(32'hb69bcd6c),
	.w2(32'h39261f02),
	.w3(32'h388f87ab),
	.w4(32'h39293506),
	.w5(32'h3805e87f),
	.w6(32'h39205a02),
	.w7(32'h391986e1),
	.w8(32'hb88837f7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb788042f),
	.w1(32'hb6bedd8a),
	.w2(32'h39502542),
	.w3(32'hb84f58f8),
	.w4(32'hb86474ad),
	.w5(32'hb8ce405f),
	.w6(32'h38e94173),
	.w7(32'hb6c7ccea),
	.w8(32'hb98fbca4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c0e3ac),
	.w1(32'h36685c2b),
	.w2(32'hb58e7fa4),
	.w3(32'h36a1fca5),
	.w4(32'h36666f76),
	.w5(32'h358f4cb2),
	.w6(32'h362b9037),
	.w7(32'hb546fdf3),
	.w8(32'hb59f32f3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ce807e),
	.w1(32'h361cb01e),
	.w2(32'hb6f61201),
	.w3(32'h37682dca),
	.w4(32'h36d267d1),
	.w5(32'hb7113a73),
	.w6(32'h37162ec6),
	.w7(32'hb58f66b6),
	.w8(32'hb5861caf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b3aa8b),
	.w1(32'hb67a34ad),
	.w2(32'hb53ad03f),
	.w3(32'hb72519db),
	.w4(32'hb700b116),
	.w5(32'hb532e86f),
	.w6(32'hb5cc680a),
	.w7(32'hb645a6d1),
	.w8(32'hb6c0b25d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb627ea65),
	.w1(32'h34e6f733),
	.w2(32'h34cee2b2),
	.w3(32'hb636d4be),
	.w4(32'hb50e284e),
	.w5(32'hb59baf06),
	.w6(32'hb5ab908d),
	.w7(32'h35822645),
	.w8(32'hb64af9d1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ec1701),
	.w1(32'h38cbd1fe),
	.w2(32'h39b30e0c),
	.w3(32'h38d64ff3),
	.w4(32'h392289b9),
	.w5(32'h38aedfcf),
	.w6(32'h39903623),
	.w7(32'h3993e0ef),
	.w8(32'h386c0e00),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70338bc),
	.w1(32'hb60f3da6),
	.w2(32'h37a8d8fb),
	.w3(32'hb6e3635d),
	.w4(32'hb30eb1d6),
	.w5(32'h379cadb5),
	.w6(32'hb68cf51d),
	.w7(32'h3688ac1f),
	.w8(32'h375987e5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f4e429),
	.w1(32'hb90a8d16),
	.w2(32'h390142d3),
	.w3(32'h37f7b5af),
	.w4(32'h3811ab0c),
	.w5(32'h38f65897),
	.w6(32'h393f682f),
	.w7(32'h3965b588),
	.w8(32'h39180732),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38920bb7),
	.w1(32'h3944046d),
	.w2(32'h392a1491),
	.w3(32'hb97a74b1),
	.w4(32'hb8e0193b),
	.w5(32'h38c731ff),
	.w6(32'hb98b84df),
	.w7(32'hb90988d4),
	.w8(32'h38b5183f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369879ce),
	.w1(32'h369d48b9),
	.w2(32'h3590a3ad),
	.w3(32'h351103fc),
	.w4(32'h35c18698),
	.w5(32'hb5c870c2),
	.w6(32'h35dc5e50),
	.w7(32'h3559672b),
	.w8(32'hb64a858a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79954b6),
	.w1(32'hb70a8614),
	.w2(32'hb8239377),
	.w3(32'h37a9497c),
	.w4(32'h372e429f),
	.w5(32'hb694470b),
	.w6(32'hb7019594),
	.w7(32'hb69bf91b),
	.w8(32'h37d42abd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365a1da5),
	.w1(32'h3595bf29),
	.w2(32'hb646b959),
	.w3(32'h355d4ac6),
	.w4(32'h3578e990),
	.w5(32'hb430283d),
	.w6(32'h35a8175e),
	.w7(32'hb417ed98),
	.w8(32'h36263013),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e9bf2),
	.w1(32'h387ef108),
	.w2(32'h38786511),
	.w3(32'h371a82cf),
	.w4(32'h38ddeeb1),
	.w5(32'h389a8693),
	.w6(32'h3889e832),
	.w7(32'h38d89d36),
	.w8(32'h38ae247b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38695db5),
	.w1(32'h3932215d),
	.w2(32'h39c2e414),
	.w3(32'h391aaf09),
	.w4(32'hb87fe0bf),
	.w5(32'h379e2bb1),
	.w6(32'h38211738),
	.w7(32'h37d6b9ba),
	.w8(32'h3639d873),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96eaaea),
	.w1(32'h37d5f287),
	.w2(32'h39f5a276),
	.w3(32'hb94f1b20),
	.w4(32'hb80e0986),
	.w5(32'h3690d0d3),
	.w6(32'h39288b4d),
	.w7(32'hb917c133),
	.w8(32'hb9a91515),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38070cf3),
	.w1(32'h366a9bd2),
	.w2(32'h3804837d),
	.w3(32'hb721af86),
	.w4(32'hb69a5768),
	.w5(32'h379c77a6),
	.w6(32'h370b21a7),
	.w7(32'h37447905),
	.w8(32'h36d30858),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385470bf),
	.w1(32'hb81c97a4),
	.w2(32'hb6f38b60),
	.w3(32'h373f65a6),
	.w4(32'hb89c0587),
	.w5(32'hb7372d32),
	.w6(32'hb78efd43),
	.w7(32'h38423365),
	.w8(32'h384f5c79),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ecddd),
	.w1(32'hb5b4ccfb),
	.w2(32'hb7c8cfb1),
	.w3(32'hb6c16c9f),
	.w4(32'h371fb8e3),
	.w5(32'h36ec2a65),
	.w6(32'hb819b8c9),
	.w7(32'hb75427bb),
	.w8(32'h3816ed3b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fac506),
	.w1(32'hb90116ba),
	.w2(32'h39083bd4),
	.w3(32'h39214a1e),
	.w4(32'hb61cbfed),
	.w5(32'h38a0ea74),
	.w6(32'h39826cbf),
	.w7(32'h37eec7b7),
	.w8(32'hb9081a13),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933e304),
	.w1(32'h39a07afe),
	.w2(32'h39428fa2),
	.w3(32'h38d94034),
	.w4(32'h38ac7ed5),
	.w5(32'h383bff7f),
	.w6(32'hb7046b1d),
	.w7(32'h37cb246f),
	.w8(32'h388258c4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1120d3),
	.w1(32'hb9e9521e),
	.w2(32'h39cec578),
	.w3(32'hb994a74b),
	.w4(32'hb8df5c39),
	.w5(32'h39847db3),
	.w6(32'h389810bf),
	.w7(32'h389f51ee),
	.w8(32'hb9004fc8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389cf4e6),
	.w1(32'h38d6dace),
	.w2(32'hb7b1d101),
	.w3(32'h3787c9fb),
	.w4(32'h3854d1e0),
	.w5(32'hb82bfa17),
	.w6(32'hb8ab6e05),
	.w7(32'hb83ad37d),
	.w8(32'hb96002a8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81eb1a2),
	.w1(32'hb8bd929e),
	.w2(32'hb700fc49),
	.w3(32'h3877f919),
	.w4(32'h3981d9e5),
	.w5(32'h3943b64d),
	.w6(32'h395738fe),
	.w7(32'h383baa8b),
	.w8(32'h38ce8a48),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6748e),
	.w1(32'hb8f14c82),
	.w2(32'h3902d525),
	.w3(32'hb91e0e64),
	.w4(32'hb91ab6d2),
	.w5(32'hb866fa50),
	.w6(32'hb84a831c),
	.w7(32'hb92e8a61),
	.w8(32'hb98727fb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88579a1),
	.w1(32'hb8e76fe6),
	.w2(32'hb88f1488),
	.w3(32'hb8c9b555),
	.w4(32'hb92ae1a5),
	.w5(32'hb96b3c89),
	.w6(32'hb909da95),
	.w7(32'hb907d134),
	.w8(32'hb90e29fa),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8904218),
	.w1(32'h37cee377),
	.w2(32'h3954aaa9),
	.w3(32'hb8c6a58c),
	.w4(32'h38a1bade),
	.w5(32'h3802c639),
	.w6(32'h388413ce),
	.w7(32'hb883f801),
	.w8(32'hb93f7837),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375ac435),
	.w1(32'h386774ce),
	.w2(32'h392323a9),
	.w3(32'h3800b589),
	.w4(32'h3826857d),
	.w5(32'h383885cb),
	.w6(32'h390d8d9a),
	.w7(32'h390a9f81),
	.w8(32'hb66f1bdc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a6de8),
	.w1(32'h373d3923),
	.w2(32'h39d3ee52),
	.w3(32'hb9a0a4f9),
	.w4(32'hb7db914b),
	.w5(32'h3a01cde7),
	.w6(32'hb9c465a8),
	.w7(32'hb91e9928),
	.w8(32'h387d2593),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e4da3),
	.w1(32'hb94749f9),
	.w2(32'hb9674d92),
	.w3(32'hb994a05b),
	.w4(32'hb9d200f8),
	.w5(32'hb9ac25a7),
	.w6(32'hb9bf13fc),
	.w7(32'hb9e4f386),
	.w8(32'hb9cb2f0f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381af693),
	.w1(32'h37627da1),
	.w2(32'h37160cd6),
	.w3(32'h383f2071),
	.w4(32'h37508a4f),
	.w5(32'h36112744),
	.w6(32'h3782626a),
	.w7(32'h366f1667),
	.w8(32'hb6a2516d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d594a8),
	.w1(32'hb857436c),
	.w2(32'hb7d3be25),
	.w3(32'hb6cae04a),
	.w4(32'hb7efe2da),
	.w5(32'hb782e3a5),
	.w6(32'hb802c2ba),
	.w7(32'hb70f793d),
	.w8(32'h3777a68b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8323ae9),
	.w1(32'hb82d2115),
	.w2(32'h3835ef72),
	.w3(32'hb8bab9a0),
	.w4(32'h3750a032),
	.w5(32'h383c027a),
	.w6(32'hb82af76c),
	.w7(32'h3836b49f),
	.w8(32'h38a5b74e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f3877),
	.w1(32'hb9597d47),
	.w2(32'hb7f6c92d),
	.w3(32'hb8b9a21c),
	.w4(32'hb9104ee1),
	.w5(32'h38a47937),
	.w6(32'hb7ed5347),
	.w7(32'h38d303d8),
	.w8(32'hb6b63f64),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a8965),
	.w1(32'h39006541),
	.w2(32'h3a1cded4),
	.w3(32'h38985b6f),
	.w4(32'h39e76460),
	.w5(32'h39f7cf29),
	.w6(32'h3a538b7c),
	.w7(32'h3a804f0b),
	.w8(32'h3a1021b4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72cac04),
	.w1(32'h3719e254),
	.w2(32'hb49ebfdd),
	.w3(32'hb73a1f30),
	.w4(32'h3652f774),
	.w5(32'hb6f5ebbb),
	.w6(32'h37cd63a1),
	.w7(32'h37029a47),
	.w8(32'hb7449297),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90634e4),
	.w1(32'h3867c775),
	.w2(32'h39c1dd28),
	.w3(32'h37bacd7c),
	.w4(32'h3865ecc0),
	.w5(32'h393127a3),
	.w6(32'h39ae8c95),
	.w7(32'h39ed690d),
	.w8(32'h394c00e7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888c07f),
	.w1(32'hb8c81ede),
	.w2(32'h395e9995),
	.w3(32'hb85c2ed5),
	.w4(32'hb83b0e29),
	.w5(32'hb91bf39e),
	.w6(32'h38ecaab4),
	.w7(32'hb7585a8b),
	.w8(32'hb99a0e16),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992cb0f),
	.w1(32'hb984415e),
	.w2(32'h392c5a04),
	.w3(32'hb85af374),
	.w4(32'h390926a0),
	.w5(32'h397dff44),
	.w6(32'h398a3941),
	.w7(32'h39c1c7f9),
	.w8(32'h392e1d52),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374d28ed),
	.w1(32'h393b884d),
	.w2(32'h38977ff1),
	.w3(32'h38bd4dcf),
	.w4(32'h39551d53),
	.w5(32'h399d4c35),
	.w6(32'hb6c95f33),
	.w7(32'h3912bae2),
	.w8(32'h39682a04),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927e697),
	.w1(32'hb97b828e),
	.w2(32'hb9886ae6),
	.w3(32'hb97cec1a),
	.w4(32'hb9604c2a),
	.w5(32'hb9372457),
	.w6(32'hb9c0522e),
	.w7(32'hb9be00a7),
	.w8(32'hb99d9ebd),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b20312),
	.w1(32'hb86f3475),
	.w2(32'hb826dab4),
	.w3(32'hb64b952d),
	.w4(32'h37e3f9a7),
	.w5(32'h36782cff),
	.w6(32'h37d2adc1),
	.w7(32'h35dfd425),
	.w8(32'h37062301),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abf174),
	.w1(32'hb908d3fb),
	.w2(32'hb88a35b0),
	.w3(32'h38b50c57),
	.w4(32'h37df99eb),
	.w5(32'hb8b5cd58),
	.w6(32'h392fa177),
	.w7(32'h3823cdc1),
	.w8(32'hb8fe5c86),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381c5a73),
	.w1(32'hb9025bd0),
	.w2(32'hb9af7bd0),
	.w3(32'hb8de6e6a),
	.w4(32'hb9a336fc),
	.w5(32'hb960707a),
	.w6(32'hb8e5559c),
	.w7(32'hb9b02d46),
	.w8(32'hb8efce99),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f3ba88),
	.w1(32'hb8540f75),
	.w2(32'hb91c2bf7),
	.w3(32'hb8043eb1),
	.w4(32'hb8929067),
	.w5(32'hb8b45f08),
	.w6(32'hb80e5bb7),
	.w7(32'hb887737f),
	.w8(32'h379c30b2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c5cd3d),
	.w1(32'hb84a735b),
	.w2(32'h36544f95),
	.w3(32'hb8248703),
	.w4(32'hb7cdd912),
	.w5(32'hb4c9defd),
	.w6(32'hb6a78b13),
	.w7(32'hb78da5dd),
	.w8(32'hb7beac9e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb667a63c),
	.w1(32'hb7396bdd),
	.w2(32'hb7b6cc8a),
	.w3(32'hb755577c),
	.w4(32'hb7b95a55),
	.w5(32'hb79d03ff),
	.w6(32'hb740c53c),
	.w7(32'hb79fac21),
	.w8(32'hb8181785),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376af2ce),
	.w1(32'h38c8e258),
	.w2(32'h3938b73a),
	.w3(32'h37b4f4e9),
	.w4(32'h38c2219a),
	.w5(32'h38d3561b),
	.w6(32'h39015b43),
	.w7(32'h388cb064),
	.w8(32'h38a3b65c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fef9e6),
	.w1(32'hb79fb80c),
	.w2(32'h37d06743),
	.w3(32'hb7ca6151),
	.w4(32'hb7b0018a),
	.w5(32'h380e7595),
	.w6(32'hb6f5677d),
	.w7(32'h37c763a3),
	.w8(32'h371df3df),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b6d78f),
	.w1(32'h3727ce68),
	.w2(32'h3857e542),
	.w3(32'h36ecfbfa),
	.w4(32'h372e49e3),
	.w5(32'hb707f976),
	.w6(32'h3885a161),
	.w7(32'h389d214d),
	.w8(32'hb8ad2426),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c922de),
	.w1(32'hb772d739),
	.w2(32'hb7be46eb),
	.w3(32'hb838e74d),
	.w4(32'hb7496dca),
	.w5(32'h3743823a),
	.w6(32'hb6f240fa),
	.w7(32'h3665ddb7),
	.w8(32'h379edd47),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1b37d),
	.w1(32'h3822137d),
	.w2(32'h39bbf44a),
	.w3(32'hb9104263),
	.w4(32'h39933ab5),
	.w5(32'h39f516e2),
	.w6(32'h398f424e),
	.w7(32'h39a4d825),
	.w8(32'h396dc8bb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6594179),
	.w1(32'h375a5b27),
	.w2(32'h38275c12),
	.w3(32'hb73e7102),
	.w4(32'hb6ed85e3),
	.w5(32'h379450ed),
	.w6(32'h36ce4024),
	.w7(32'h37ebd2bc),
	.w8(32'h373eb94f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38079409),
	.w1(32'h3706a1d2),
	.w2(32'hb673da87),
	.w3(32'h37b06990),
	.w4(32'hb70af2ae),
	.w5(32'hb706e998),
	.w6(32'h37502a8c),
	.w7(32'hb78b7467),
	.w8(32'hb7c1770c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f9bd1),
	.w1(32'h36b55302),
	.w2(32'hb8150454),
	.w3(32'hb7d75a1f),
	.w4(32'hb8f2dec8),
	.w5(32'hb9887afe),
	.w6(32'hb8fc11ab),
	.w7(32'hb94e0826),
	.w8(32'hb9d91769),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924cd49),
	.w1(32'h3855bb18),
	.w2(32'h39f8c366),
	.w3(32'h38ad7063),
	.w4(32'hb826d5a6),
	.w5(32'hb85686d7),
	.w6(32'h38cd1bed),
	.w7(32'hb979c395),
	.w8(32'hb9afb314),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a5a693),
	.w1(32'hb76db3a6),
	.w2(32'hb7b331ea),
	.w3(32'hb6f1b0d9),
	.w4(32'hb83cbaaf),
	.w5(32'hb76d000c),
	.w6(32'hb6c48191),
	.w7(32'hb7f00ba9),
	.w8(32'h3788b740),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37da3e7e),
	.w1(32'hb7d54995),
	.w2(32'h3944e1ec),
	.w3(32'h38139af7),
	.w4(32'h389b4bca),
	.w5(32'hb90d251f),
	.w6(32'h397de24d),
	.w7(32'h396491bd),
	.w8(32'hb98c7de8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7353c2a),
	.w1(32'h3892c19b),
	.w2(32'h393a7575),
	.w3(32'h389be740),
	.w4(32'h38d68083),
	.w5(32'h38e381f9),
	.w6(32'h3888f8ec),
	.w7(32'h389a8b27),
	.w8(32'h3805e0c1),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98155fd),
	.w1(32'hb8f69e44),
	.w2(32'h39220aa1),
	.w3(32'h3928412a),
	.w4(32'h39dc2e54),
	.w5(32'h39bb0b0c),
	.w6(32'h3a789e14),
	.w7(32'h3a6ff73b),
	.w8(32'h3a0e398e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c5539b),
	.w1(32'hb892f5a6),
	.w2(32'hb8278fbe),
	.w3(32'hb88d64cd),
	.w4(32'hb9117447),
	.w5(32'hb8cb503c),
	.w6(32'hb8e1ba92),
	.w7(32'hb8c304b4),
	.w8(32'hb8472201),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93955fa),
	.w1(32'h3861aa39),
	.w2(32'h3a2a7dd2),
	.w3(32'hb896aa28),
	.w4(32'h38ca8a98),
	.w5(32'h388bfa44),
	.w6(32'h39cdad8f),
	.w7(32'h37a21066),
	.w8(32'hb9e8685d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38570279),
	.w1(32'hb887466a),
	.w2(32'hb79a7e18),
	.w3(32'h38872540),
	.w4(32'hb85dec7c),
	.w5(32'hb79b0228),
	.w6(32'hb6018754),
	.w7(32'h37781110),
	.w8(32'h379c534b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8278c99),
	.w1(32'hb8cd83e5),
	.w2(32'h3926511e),
	.w3(32'hb8515be5),
	.w4(32'hb8c69430),
	.w5(32'hb9280282),
	.w6(32'h388cc831),
	.w7(32'hb969ae27),
	.w8(32'hb9c1595c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb745fe5f),
	.w1(32'h373c0eac),
	.w2(32'hb6c60641),
	.w3(32'hb768509b),
	.w4(32'h37057928),
	.w5(32'hb6be1cca),
	.w6(32'h37c0d9c3),
	.w7(32'h372c7316),
	.w8(32'hb5faa23b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e7cfee),
	.w1(32'h39340f48),
	.w2(32'h39454222),
	.w3(32'h37d7c9de),
	.w4(32'h38de67e1),
	.w5(32'h390cf400),
	.w6(32'h381d6c2d),
	.w7(32'h383d1d5c),
	.w8(32'h38a3f4f1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e62661),
	.w1(32'hb7e5f557),
	.w2(32'hb934caf5),
	.w3(32'hb84bf4a1),
	.w4(32'h38039279),
	.w5(32'hb873429f),
	.w6(32'h379bbeb5),
	.w7(32'hb7c438cd),
	.w8(32'hb7a015f5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901f768),
	.w1(32'h37b0315f),
	.w2(32'h38325291),
	.w3(32'hb87a3753),
	.w4(32'h38b0a4ae),
	.w5(32'h3938ccd6),
	.w6(32'h3918c8ab),
	.w7(32'h393c3ede),
	.w8(32'h394c4013),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382c0a79),
	.w1(32'hb7f6da0b),
	.w2(32'hb6a79fb9),
	.w3(32'h3847a75f),
	.w4(32'hb7e2e50c),
	.w5(32'h37d5cff5),
	.w6(32'hb815ea73),
	.w7(32'h3756c989),
	.w8(32'h37935d8e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c86f14),
	.w1(32'hb804d983),
	.w2(32'hb7b74a01),
	.w3(32'h380fb16e),
	.w4(32'hb7e1569e),
	.w5(32'hb7a02852),
	.w6(32'hb7d8d787),
	.w7(32'hb7c55952),
	.w8(32'hb7bd40cb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e85158),
	.w1(32'h388fda4e),
	.w2(32'h37c257ce),
	.w3(32'hb80fae9d),
	.w4(32'hb7c713d5),
	.w5(32'hb86c12a9),
	.w6(32'h383c7f0f),
	.w7(32'h372f46f2),
	.w8(32'h37fc2bb6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d784a),
	.w1(32'h38ff31b3),
	.w2(32'h3903ea0a),
	.w3(32'h37d9581f),
	.w4(32'h38321ba9),
	.w5(32'h390e930e),
	.w6(32'h38a35d1e),
	.w7(32'h38a5ee73),
	.w8(32'h3909bc56),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39063688),
	.w1(32'hb8b2ba6d),
	.w2(32'hb8ec0b68),
	.w3(32'h388c49a9),
	.w4(32'hb885ad14),
	.w5(32'h3581a3c0),
	.w6(32'hb6d2cd54),
	.w7(32'h37fd82ed),
	.w8(32'hb886bdca),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33219dee),
	.w1(32'h37e3f4f1),
	.w2(32'h38545cfc),
	.w3(32'hb853c134),
	.w4(32'h37cef641),
	.w5(32'h37fa2655),
	.w6(32'hb6cecea2),
	.w7(32'h35cbf511),
	.w8(32'h371d49ea),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27ccf8),
	.w1(32'hba25dcf3),
	.w2(32'h39df8c63),
	.w3(32'hb78a57f1),
	.w4(32'h3a4bf10b),
	.w5(32'h3a69bde6),
	.w6(32'h3afc016f),
	.w7(32'h3b00e1eb),
	.w8(32'h3a980ae2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c09354),
	.w1(32'h391e146c),
	.w2(32'hb922bf48),
	.w3(32'h39b8f481),
	.w4(32'h383fc3a2),
	.w5(32'hb9c013ef),
	.w6(32'h391a890d),
	.w7(32'h37a8fc31),
	.w8(32'hb6ce1058),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d1cfc),
	.w1(32'hb716f3db),
	.w2(32'h3714a186),
	.w3(32'hb7614eb2),
	.w4(32'hb5c67c36),
	.w5(32'h386d5f76),
	.w6(32'hb6b95bec),
	.w7(32'h36bc6ff2),
	.w8(32'h36dc64f3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb728dc2f),
	.w1(32'h38b3f1e6),
	.w2(32'h375dc16a),
	.w3(32'hb78888c0),
	.w4(32'h389a7095),
	.w5(32'hb70cbde3),
	.w6(32'h3864c7fe),
	.w7(32'hb7bed65a),
	.w8(32'hb412e962),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b7dc65),
	.w1(32'hb5e54d3a),
	.w2(32'h37c4c61c),
	.w3(32'h381cff00),
	.w4(32'h38238781),
	.w5(32'h383648da),
	.w6(32'h3739c8c9),
	.w7(32'h38731b29),
	.w8(32'h383e1883),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38025ed3),
	.w1(32'hb75337fe),
	.w2(32'hb7a70d34),
	.w3(32'h37f7d292),
	.w4(32'hb7f477b9),
	.w5(32'hb7eb6f79),
	.w6(32'hb7eaf0b4),
	.w7(32'hb816531c),
	.w8(32'hb844d079),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82717ec),
	.w1(32'hb80b74b8),
	.w2(32'h38114023),
	.w3(32'h38498abb),
	.w4(32'h3881154d),
	.w5(32'h386e1377),
	.w6(32'h389c3ab2),
	.w7(32'h389652f6),
	.w8(32'hb88a3f5f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78b0487),
	.w1(32'hb97afbf4),
	.w2(32'hb951b1c8),
	.w3(32'hb8a2890b),
	.w4(32'hb9639150),
	.w5(32'hb9bc84c5),
	.w6(32'hb816413f),
	.w7(32'hb90d9449),
	.w8(32'hb8a164c9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c8579),
	.w1(32'hb8d86430),
	.w2(32'hb839b7b8),
	.w3(32'h38a8b180),
	.w4(32'h395e5353),
	.w5(32'hb93473d4),
	.w6(32'h3a6c5407),
	.w7(32'h3a2f193a),
	.w8(32'h38299b0a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d2cef8),
	.w1(32'h38f0755a),
	.w2(32'h38abb764),
	.w3(32'hb8be8ee4),
	.w4(32'h38e68a51),
	.w5(32'h38e46f8f),
	.w6(32'hb7d49736),
	.w7(32'hb7250d22),
	.w8(32'hb842037d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d5d03),
	.w1(32'hb9074ef6),
	.w2(32'h39878270),
	.w3(32'h387b5c82),
	.w4(32'h3969be2a),
	.w5(32'h3980cf81),
	.w6(32'h3a1d018e),
	.w7(32'h3a1a8e85),
	.w8(32'h3989a657),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3651d8a6),
	.w1(32'hb83a9048),
	.w2(32'h378af2c4),
	.w3(32'hb80d921e),
	.w4(32'hb85e454c),
	.w5(32'hb83e8e62),
	.w6(32'h37a04b92),
	.w7(32'h3767531e),
	.w8(32'h36f71202),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37252da7),
	.w1(32'h354a3ae4),
	.w2(32'hb73806b3),
	.w3(32'hb66109a6),
	.w4(32'hb7654ff0),
	.w5(32'hb74458d3),
	.w6(32'h35f2a837),
	.w7(32'hb663af18),
	.w8(32'hb77aff43),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369c12ec),
	.w1(32'h382812e8),
	.w2(32'hb7ebf605),
	.w3(32'h37870c09),
	.w4(32'h380db3f3),
	.w5(32'hb8101093),
	.w6(32'h3810ec3d),
	.w7(32'h37d75169),
	.w8(32'hb7e67561),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7014f70),
	.w1(32'h359814b4),
	.w2(32'hb6f30331),
	.w3(32'hb7103807),
	.w4(32'hb7068efd),
	.w5(32'hb728d1fe),
	.w6(32'hb673e407),
	.w7(32'h35f8fd74),
	.w8(32'hb74bff6c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ff6d8),
	.w1(32'hb8b51dc5),
	.w2(32'h38dbac53),
	.w3(32'h388c44df),
	.w4(32'h398beb4b),
	.w5(32'h386bcc14),
	.w6(32'h397e20c2),
	.w7(32'h39bebff0),
	.w8(32'h38e98203),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9e757),
	.w1(32'hb898c751),
	.w2(32'hb9ae5105),
	.w3(32'hb99481ce),
	.w4(32'hb984ea5e),
	.w5(32'hb8d5d76d),
	.w6(32'hb9905fed),
	.w7(32'hb99eef92),
	.w8(32'h3886246b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6eb66),
	.w1(32'h387fa9a8),
	.w2(32'h386e3b59),
	.w3(32'h379ec0f2),
	.w4(32'hb8408541),
	.w5(32'hb8ca782f),
	.w6(32'h35168527),
	.w7(32'hb88dff3d),
	.w8(32'hb90c393d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f1fe7b),
	.w1(32'hb842f646),
	.w2(32'hb879a325),
	.w3(32'hb7b15fa2),
	.w4(32'hb84129d8),
	.w5(32'hb80af48d),
	.w6(32'hb83865d9),
	.w7(32'hb8741f36),
	.w8(32'h35b237b2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ee6e7),
	.w1(32'h36153f37),
	.w2(32'hb92521b8),
	.w3(32'hb7857232),
	.w4(32'hb8d16e6d),
	.w5(32'hb97fc477),
	.w6(32'hb8910e25),
	.w7(32'hb8a5733e),
	.w8(32'hb98741b1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e707ce),
	.w1(32'hb82cc755),
	.w2(32'h397d773f),
	.w3(32'h37c0fbe7),
	.w4(32'h3881ddaf),
	.w5(32'h372c9deb),
	.w6(32'h39c49bcb),
	.w7(32'h392c3814),
	.w8(32'hb94b06a3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0938d),
	.w1(32'hb99a60a3),
	.w2(32'h39e18be3),
	.w3(32'hb8f4bfb1),
	.w4(32'h39e9b05b),
	.w5(32'h3a09db4d),
	.w6(32'h3a5d7331),
	.w7(32'h3a8aca77),
	.w8(32'h3a437694),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83c6704),
	.w1(32'hb6e4118b),
	.w2(32'hb5fe9003),
	.w3(32'hb7f8149a),
	.w4(32'hb789ccb1),
	.w5(32'hb7004425),
	.w6(32'h3545a57f),
	.w7(32'h36ce1885),
	.w8(32'h366592fc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81cae98),
	.w1(32'hb8290b58),
	.w2(32'hb795c9bc),
	.w3(32'hb818894d),
	.w4(32'hb7a47ed1),
	.w5(32'hb6f4e725),
	.w6(32'h3650de14),
	.w7(32'hb7a69d85),
	.w8(32'hb72e607a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909eb60),
	.w1(32'h38886d6c),
	.w2(32'h3926bd0a),
	.w3(32'h36d6fcd1),
	.w4(32'hb88c80ae),
	.w5(32'h380d7764),
	.w6(32'hb7ee1091),
	.w7(32'h37c64a59),
	.w8(32'h39224dae),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2d79f),
	.w1(32'hb896cc08),
	.w2(32'h3987eac2),
	.w3(32'hb84e859d),
	.w4(32'hb92e5e99),
	.w5(32'hb928a11e),
	.w6(32'hb82d28a2),
	.w7(32'hb944144e),
	.w8(32'hb9c787a8),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88201ac),
	.w1(32'h37b4105c),
	.w2(32'h3959a234),
	.w3(32'hb930cd31),
	.w4(32'hb8e6fbee),
	.w5(32'hb92bfce0),
	.w6(32'h39491c07),
	.w7(32'h37bcd3fa),
	.w8(32'hb922f710),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377ae295),
	.w1(32'hb95006a7),
	.w2(32'hb88412af),
	.w3(32'h3682c993),
	.w4(32'hb88cfe51),
	.w5(32'h38d2c6a2),
	.w6(32'h383bdfc8),
	.w7(32'hb8a81e37),
	.w8(32'hb80f142f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375f92d9),
	.w1(32'h37b32565),
	.w2(32'h3556387f),
	.w3(32'h3684566d),
	.w4(32'hb5b271d4),
	.w5(32'hb6918603),
	.w6(32'h378b955f),
	.w7(32'h3590c98b),
	.w8(32'hb6d4c16a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ff4776),
	.w1(32'h344356ea),
	.w2(32'h32923c82),
	.w3(32'hb6bc5d5a),
	.w4(32'hb81930a5),
	.w5(32'hb81dc117),
	.w6(32'hb79590d4),
	.w7(32'hb7d14da1),
	.w8(32'hb7f2d4f5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377957ee),
	.w1(32'hb92e0de4),
	.w2(32'h390c174a),
	.w3(32'h37cfe78d),
	.w4(32'hb72e94a1),
	.w5(32'h39485c58),
	.w6(32'h384ef8eb),
	.w7(32'h38060c2e),
	.w8(32'h387f6c9a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71dce5),
	.w1(32'hba23197a),
	.w2(32'h379429bd),
	.w3(32'hb842a51d),
	.w4(32'h39c1e192),
	.w5(32'h3a0033c1),
	.w6(32'h3a8b6816),
	.w7(32'h3aa5bc49),
	.w8(32'h3a7a5fac),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e751b),
	.w1(32'h37d6b6c9),
	.w2(32'h39297b4b),
	.w3(32'hb811a6cb),
	.w4(32'h384a597e),
	.w5(32'h390cdc9d),
	.w6(32'hb7872930),
	.w7(32'h391d9f9d),
	.w8(32'h37eb1922),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389689a9),
	.w1(32'hb788ef87),
	.w2(32'hb9716085),
	.w3(32'h38f48ff6),
	.w4(32'h32ead862),
	.w5(32'hb8a4c92a),
	.w6(32'hb8036e1e),
	.w7(32'hb69e8c62),
	.w8(32'h38851e3e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bbdff3),
	.w1(32'hb93b0626),
	.w2(32'hb93f08be),
	.w3(32'hb68c1a52),
	.w4(32'hb89136c7),
	.w5(32'hb96bb5cb),
	.w6(32'h39268f3c),
	.w7(32'hb6eb122c),
	.w8(32'hb944de83),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb850049f),
	.w1(32'hb7c3c0d5),
	.w2(32'hb4f635fc),
	.w3(32'hb82590d7),
	.w4(32'hb80ca89a),
	.w5(32'hb7c3fee3),
	.w6(32'hb7c48416),
	.w7(32'hb719eb1e),
	.w8(32'hb7c807a1),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb774b3ef),
	.w1(32'hb74ff318),
	.w2(32'hb731ff9e),
	.w3(32'hb7f8be1b),
	.w4(32'hb7c20263),
	.w5(32'hb70e059d),
	.w6(32'h34071354),
	.w7(32'h370cc33d),
	.w8(32'h37178368),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38259f27),
	.w1(32'hb7077093),
	.w2(32'hb7c27a7a),
	.w3(32'hb7a9c032),
	.w4(32'hb765c1f8),
	.w5(32'hb53d9ece),
	.w6(32'h355d67ca),
	.w7(32'hb6f9badd),
	.w8(32'hb76189be),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81370f1),
	.w1(32'h373aa43a),
	.w2(32'hb84957f2),
	.w3(32'hb7e44d41),
	.w4(32'h37659cee),
	.w5(32'hb8067cee),
	.w6(32'h3738e7d2),
	.w7(32'hb80655d1),
	.w8(32'hb621c8b7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37402585),
	.w1(32'h364abf10),
	.w2(32'h37a73832),
	.w3(32'h38223a1f),
	.w4(32'hb7690f44),
	.w5(32'h389e89d4),
	.w6(32'hb84cd94b),
	.w7(32'hb60247cd),
	.w8(32'h3841f7b2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0fb9a),
	.w1(32'hb8a2de8d),
	.w2(32'h36c488b9),
	.w3(32'hb889e41f),
	.w4(32'hb88bee84),
	.w5(32'hb8828851),
	.w6(32'h3948f64e),
	.w7(32'h359fa20e),
	.w8(32'hb904679f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bb11ae),
	.w1(32'hb8dcb761),
	.w2(32'h3711373e),
	.w3(32'hb8c6d4fc),
	.w4(32'hb9130c95),
	.w5(32'hb8a9dfa7),
	.w6(32'hb91cd6c0),
	.w7(32'hb8f043fc),
	.w8(32'hb8980f83),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377811a2),
	.w1(32'hb883709d),
	.w2(32'hb93e1167),
	.w3(32'hb83e07b1),
	.w4(32'hb8808436),
	.w5(32'hb820296f),
	.w6(32'hb7f6566a),
	.w7(32'hb7f14134),
	.w8(32'h36c81d63),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94edf68),
	.w1(32'hb9abcc73),
	.w2(32'h384dda8a),
	.w3(32'hb90d72e3),
	.w4(32'hb82c6af4),
	.w5(32'h3920a3d5),
	.w6(32'h38a1937d),
	.w7(32'h39a0b874),
	.w8(32'h39087e3e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935f45e),
	.w1(32'hb874ef2a),
	.w2(32'h3961ff93),
	.w3(32'hb9544d9b),
	.w4(32'hb886da35),
	.w5(32'hb82f0616),
	.w6(32'h38a50055),
	.w7(32'hb83ccc8a),
	.w8(32'hb946da3f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ba5a10),
	.w1(32'h378e53e1),
	.w2(32'h375507a3),
	.w3(32'hb81c99d8),
	.w4(32'hb656baa0),
	.w5(32'hb6ce0d45),
	.w6(32'hb836c0af),
	.w7(32'hb7cfa616),
	.w8(32'hb7fab0dd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a46638),
	.w1(32'hb783e0d8),
	.w2(32'h394a6cda),
	.w3(32'h384c9a02),
	.w4(32'h38abe260),
	.w5(32'h38fdf373),
	.w6(32'h395f2be4),
	.w7(32'h39311d75),
	.w8(32'h3884d629),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b4ed7d),
	.w1(32'hb757f3cc),
	.w2(32'hb6959a7e),
	.w3(32'hb657cfd1),
	.w4(32'hb7c99eae),
	.w5(32'hb7dab6e2),
	.w6(32'hb80c86c6),
	.w7(32'hb75f105b),
	.w8(32'hb808b3a0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bd3226),
	.w1(32'hb72327fc),
	.w2(32'hb482a774),
	.w3(32'hb829c2fe),
	.w4(32'hb72669e3),
	.w5(32'hb6dc58db),
	.w6(32'h37c00fae),
	.w7(32'h3743481f),
	.w8(32'hb5b611f1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7af2182),
	.w1(32'h370291fd),
	.w2(32'hb729ea19),
	.w3(32'hb7bfa3ec),
	.w4(32'h36b66007),
	.w5(32'hb69cb49f),
	.w6(32'h376f9587),
	.w7(32'h361ec0ff),
	.w8(32'h3552febe),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb703860c),
	.w1(32'hb609eb98),
	.w2(32'hb82ceef2),
	.w3(32'hb71d18ab),
	.w4(32'hb7a0c3bf),
	.w5(32'hb80a59ad),
	.w6(32'hb75a8247),
	.w7(32'hb813d3e3),
	.w8(32'hb81acf83),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ad46e),
	.w1(32'hb99e670d),
	.w2(32'hb9e79bea),
	.w3(32'hb92e1f89),
	.w4(32'hb95f7654),
	.w5(32'hb9644d9d),
	.w6(32'hb919d234),
	.w7(32'hb8fcb775),
	.w8(32'hb9147903),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957f654),
	.w1(32'h3781b4e1),
	.w2(32'h39fa50a2),
	.w3(32'hb9133916),
	.w4(32'hb78e1b08),
	.w5(32'h38196f56),
	.w6(32'h38f5e428),
	.w7(32'hb8f4bca3),
	.w8(32'hb95942e9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c2f3f9),
	.w1(32'hb874db87),
	.w2(32'h399f77c8),
	.w3(32'h386a7df5),
	.w4(32'hb8cad8e4),
	.w5(32'hb843bda3),
	.w6(32'h395363fb),
	.w7(32'hb91b1c3e),
	.w8(32'hb9cc19a9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb2c02),
	.w1(32'hb9532ee7),
	.w2(32'h39c5e95f),
	.w3(32'h3971ff35),
	.w4(32'h39cfff30),
	.w5(32'h39b202e5),
	.w6(32'h3a4565ca),
	.w7(32'h39f6347e),
	.w8(32'h38923a79),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78bd928),
	.w1(32'h379f4c0e),
	.w2(32'h37bc8d15),
	.w3(32'hb80a7905),
	.w4(32'h36093689),
	.w5(32'h36bae6d6),
	.w6(32'h381c745d),
	.w7(32'hb6c54f61),
	.w8(32'hb7d3085a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372589bd),
	.w1(32'h37ae68ea),
	.w2(32'hb60858d4),
	.w3(32'h3798c341),
	.w4(32'h37221102),
	.w5(32'hb6831662),
	.w6(32'h3792f3c3),
	.w7(32'h366fee43),
	.w8(32'h36bc630a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79264b1),
	.w1(32'hb6cdbfe6),
	.w2(32'hb79615d3),
	.w3(32'hb7467ab1),
	.w4(32'hb6e42473),
	.w5(32'hb70f1870),
	.w6(32'hb51c1492),
	.w7(32'hb72373d6),
	.w8(32'hb72fbb33),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77577ad),
	.w1(32'h3423c681),
	.w2(32'hb780f654),
	.w3(32'hb726e9db),
	.w4(32'h36652d38),
	.w5(32'hb6818f4d),
	.w6(32'h37265e46),
	.w7(32'hb43e700d),
	.w8(32'hb52c3a47),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958bf73),
	.w1(32'hb948f82f),
	.w2(32'hb8f1ca99),
	.w3(32'hb96a0599),
	.w4(32'hb9961616),
	.w5(32'hb97edb06),
	.w6(32'hb8d43072),
	.w7(32'hb97f77c0),
	.w8(32'hb93652c6),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7061d37),
	.w1(32'h35022514),
	.w2(32'h37929d9a),
	.w3(32'hb716e4c4),
	.w4(32'hb637e967),
	.w5(32'h37e5b202),
	.w6(32'h378e37d7),
	.w7(32'h385a04b8),
	.w8(32'hb689d3df),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e8cff),
	.w1(32'hb871e08d),
	.w2(32'hb7eade76),
	.w3(32'hb85ac086),
	.w4(32'hb8869826),
	.w5(32'hb74577ce),
	.w6(32'hb8a1f35e),
	.w7(32'hb8492474),
	.w8(32'h36a1dfab),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37390276),
	.w1(32'h38066a92),
	.w2(32'hb80c8c62),
	.w3(32'h3627aee9),
	.w4(32'h3739dfd0),
	.w5(32'hb7ca799b),
	.w6(32'h38768852),
	.w7(32'h371fe11f),
	.w8(32'hb8336595),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb640e573),
	.w1(32'h3804b412),
	.w2(32'h3771d831),
	.w3(32'h36909add),
	.w4(32'h37fa24b1),
	.w5(32'h3770e36c),
	.w6(32'h378c11bb),
	.w7(32'h37bb177a),
	.w8(32'h36ea5133),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8570b23),
	.w1(32'h385318ae),
	.w2(32'h38e77d6f),
	.w3(32'hb825be6a),
	.w4(32'h389c3c58),
	.w5(32'h38edfe6a),
	.w6(32'h394eb357),
	.w7(32'h3989e162),
	.w8(32'h3944dd01),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387ee7c7),
	.w1(32'h384a6f9c),
	.w2(32'h3816dcf5),
	.w3(32'hb71329f4),
	.w4(32'h37feab3c),
	.w5(32'h381058a6),
	.w6(32'h381b2e8a),
	.w7(32'h3819db91),
	.w8(32'h37f7ed36),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f805bc),
	.w1(32'h3818dcae),
	.w2(32'h39718995),
	.w3(32'h3828876f),
	.w4(32'h38fca343),
	.w5(32'h393c7d77),
	.w6(32'h38d3ebb1),
	.w7(32'hb91b4d56),
	.w8(32'hb926d71a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71a5159),
	.w1(32'h36f262fa),
	.w2(32'hb6dc1377),
	.w3(32'hb767bab8),
	.w4(32'h369a203f),
	.w5(32'hb6707fa3),
	.w6(32'hb690600f),
	.w7(32'hb6443335),
	.w8(32'hb5f78a1d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17051d),
	.w1(32'h3a0ef2e8),
	.w2(32'h39448ced),
	.w3(32'h39144a22),
	.w4(32'h39bd6fab),
	.w5(32'hb8d7b1cf),
	.w6(32'hb9e07d01),
	.w7(32'hb9e81e82),
	.w8(32'hba47a091),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule