module layer_10_featuremap_492(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fab3f),
	.w1(32'h3bcd0a51),
	.w2(32'h3aca027b),
	.w3(32'hb8ff5589),
	.w4(32'h3c2ae96b),
	.w5(32'h3b06deb7),
	.w6(32'h3b9f6127),
	.w7(32'h3a878bdf),
	.w8(32'hbb090aa2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8732eb),
	.w1(32'h3bad75b8),
	.w2(32'hbaf70f6b),
	.w3(32'h3b47b5f6),
	.w4(32'h3abab34b),
	.w5(32'hbbd8fe39),
	.w6(32'hbacb4788),
	.w7(32'hbabf17c3),
	.w8(32'hbbccc0cc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb258114),
	.w1(32'hbabd2c33),
	.w2(32'hbb7083dd),
	.w3(32'hba9615ad),
	.w4(32'hbb52a5ed),
	.w5(32'h39b49116),
	.w6(32'hbaa37c67),
	.w7(32'hbbb58fc6),
	.w8(32'h3a82afdd),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8227),
	.w1(32'hbb7fbc5b),
	.w2(32'hbb783e04),
	.w3(32'hbbc30393),
	.w4(32'hbb9f1be6),
	.w5(32'hbc00d7bd),
	.w6(32'hba1aeb51),
	.w7(32'h3b0f78ae),
	.w8(32'h3a8dddc9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d9c16),
	.w1(32'h3b078058),
	.w2(32'h3aa949fa),
	.w3(32'hba343cf6),
	.w4(32'hba47c33c),
	.w5(32'h3a37964d),
	.w6(32'h3a3ed3c0),
	.w7(32'hbb193257),
	.w8(32'hba9f58a0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87f64e),
	.w1(32'h3944e1b6),
	.w2(32'hbaac291a),
	.w3(32'h3ac1407f),
	.w4(32'hbaffb5dc),
	.w5(32'hbb42b627),
	.w6(32'hb738ed6c),
	.w7(32'hbaf4be93),
	.w8(32'hb9ffb868),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d4cf2),
	.w1(32'hba51212a),
	.w2(32'h3bfc7fc8),
	.w3(32'hbb412f20),
	.w4(32'hbb882f48),
	.w5(32'hbbd21b7e),
	.w6(32'hbb25e10d),
	.w7(32'h37e8ff4f),
	.w8(32'hbbbf96e0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01f9f0),
	.w1(32'hbc002cee),
	.w2(32'h3bf878d6),
	.w3(32'hbc4c93ad),
	.w4(32'hb94de0c5),
	.w5(32'h3c1cfeae),
	.w6(32'hbc3bf530),
	.w7(32'hbbc0d9e7),
	.w8(32'hbb8ebc33),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ada54),
	.w1(32'h38e6160d),
	.w2(32'h38baf895),
	.w3(32'hbb1b938a),
	.w4(32'h3b0e1090),
	.w5(32'hbbc4386b),
	.w6(32'hbc0a5b6a),
	.w7(32'h3b9cf26d),
	.w8(32'h3b0cf503),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb153c7c),
	.w1(32'h3ba592f7),
	.w2(32'h3b0d08ce),
	.w3(32'hbb682e02),
	.w4(32'hbb3b72c4),
	.w5(32'hb9b9035c),
	.w6(32'hbb1fd24b),
	.w7(32'hbb1e1b70),
	.w8(32'hbb976e89),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f252b),
	.w1(32'h3aecfcb0),
	.w2(32'h3a403ef6),
	.w3(32'hba5b04ac),
	.w4(32'hb9ac52ef),
	.w5(32'h3a22eb36),
	.w6(32'hbadb3ad3),
	.w7(32'hbb1e0fc2),
	.w8(32'hbb13af48),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81baf7),
	.w1(32'h3b133246),
	.w2(32'h3be201cf),
	.w3(32'hbb8fda13),
	.w4(32'h3bb70697),
	.w5(32'h3c19d7a3),
	.w6(32'hbbeae09e),
	.w7(32'h3b58362a),
	.w8(32'hbaa328d3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af444da),
	.w1(32'h39876815),
	.w2(32'h3b3b5379),
	.w3(32'hbaaff99e),
	.w4(32'h3aa8e329),
	.w5(32'h3b11a8f8),
	.w6(32'hbbbc9931),
	.w7(32'h3ba5abcb),
	.w8(32'h3b5a0c9a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3475e7),
	.w1(32'hba9a1cc8),
	.w2(32'hbb755d49),
	.w3(32'h3b76e2c0),
	.w4(32'h3aaf7e8f),
	.w5(32'h3afe2133),
	.w6(32'h3b8d64e1),
	.w7(32'hbac808ca),
	.w8(32'h3afd55d6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c5b92),
	.w1(32'h3b3619be),
	.w2(32'hb943e86b),
	.w3(32'hb8aeead9),
	.w4(32'hbafb00cc),
	.w5(32'h3b605ea3),
	.w6(32'h3b4476d5),
	.w7(32'hbb46cc69),
	.w8(32'hbb866802),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbacb3e),
	.w1(32'h3c04f429),
	.w2(32'h3c2fe0c8),
	.w3(32'hbae4432d),
	.w4(32'h3bc3068c),
	.w5(32'h3c9967b7),
	.w6(32'hbba911a1),
	.w7(32'h3bf39f90),
	.w8(32'h3aac12c3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b412e34),
	.w1(32'h39b7b06c),
	.w2(32'h3a8f2071),
	.w3(32'h3b9082f1),
	.w4(32'hbb24bd02),
	.w5(32'hbb79f848),
	.w6(32'h3a47ce32),
	.w7(32'hbaa7e4af),
	.w8(32'hbb333bd3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5070d7),
	.w1(32'h3b2182d9),
	.w2(32'h3c04e2c7),
	.w3(32'hbc4609aa),
	.w4(32'h3bc23a4a),
	.w5(32'h3b65927a),
	.w6(32'hbc301411),
	.w7(32'h3b120622),
	.w8(32'hbba20a5e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16b0bb),
	.w1(32'h3acd6461),
	.w2(32'h3b81cc9c),
	.w3(32'hbb9fa1e2),
	.w4(32'h380c6c0c),
	.w5(32'h3af81f24),
	.w6(32'hbbc4b714),
	.w7(32'h3a9cf78e),
	.w8(32'h3bb0bca6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccbfe5),
	.w1(32'hba3cfa46),
	.w2(32'h3b60c134),
	.w3(32'hbae33c69),
	.w4(32'hbb862be3),
	.w5(32'hbc05d770),
	.w6(32'h39791673),
	.w7(32'hbbc33a35),
	.w8(32'hbc0fd95e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c090e),
	.w1(32'hbb53607f),
	.w2(32'hbbc2bb55),
	.w3(32'hba92e694),
	.w4(32'hbb44b4ab),
	.w5(32'hbab37808),
	.w6(32'hbb5b11a1),
	.w7(32'hbb689a3e),
	.w8(32'h3a3c4840),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7b26),
	.w1(32'hbb5e707f),
	.w2(32'hbb0948cf),
	.w3(32'hba1abe05),
	.w4(32'hbafc51b4),
	.w5(32'hbb9cdfcc),
	.w6(32'h3a539211),
	.w7(32'hbaa4f62c),
	.w8(32'hbaa6d574),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f76e4),
	.w1(32'hbb08c49c),
	.w2(32'h3b5227ae),
	.w3(32'hbc32ca13),
	.w4(32'h3ae4a748),
	.w5(32'h3b97f48a),
	.w6(32'hbcb85f7e),
	.w7(32'h3a6f772b),
	.w8(32'hbc21ae42),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399168e1),
	.w1(32'h3886d973),
	.w2(32'hbb107821),
	.w3(32'hba8477c5),
	.w4(32'hba40e567),
	.w5(32'hbb1ff87a),
	.w6(32'hbb93f505),
	.w7(32'hb9327084),
	.w8(32'hbbb63edb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfef1ef),
	.w1(32'h3b23116e),
	.w2(32'hbbb59bc9),
	.w3(32'hbafb2b9a),
	.w4(32'hbb277ce9),
	.w5(32'hbbd2bc05),
	.w6(32'h3b75a221),
	.w7(32'hbad9b23b),
	.w8(32'hbbf1a90f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30cfc8),
	.w1(32'hbaf408c0),
	.w2(32'hbb593885),
	.w3(32'hbb82cf19),
	.w4(32'hbb8ca84e),
	.w5(32'hbb4dbf37),
	.w6(32'hbb146e5b),
	.w7(32'hbb489272),
	.w8(32'hbb9f28f7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfccf6),
	.w1(32'h3be4d1ba),
	.w2(32'hba806bfb),
	.w3(32'hbb0ef085),
	.w4(32'h3be9ae11),
	.w5(32'hbac05d66),
	.w6(32'hbaccc08a),
	.w7(32'h3c53f680),
	.w8(32'h3c2aaec8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ba05d),
	.w1(32'hbb2a7808),
	.w2(32'hbc106c53),
	.w3(32'h3ca35ff9),
	.w4(32'hbb974046),
	.w5(32'hbbab74ea),
	.w6(32'h3cc48fb6),
	.w7(32'h3b1a46f0),
	.w8(32'h3b605a3b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e86c),
	.w1(32'h3b0025ff),
	.w2(32'h3ac13abf),
	.w3(32'h3962b607),
	.w4(32'h3b5b7709),
	.w5(32'hbb21bd92),
	.w6(32'hb9983edc),
	.w7(32'h3ba90613),
	.w8(32'hb9979622),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7258ea),
	.w1(32'h3b3df043),
	.w2(32'hbbfe1a7a),
	.w3(32'h3b384edd),
	.w4(32'hb9b9f351),
	.w5(32'hbbfbd7ce),
	.w6(32'h3c49ff60),
	.w7(32'h3b71a6ad),
	.w8(32'hbc530a5a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb158458),
	.w1(32'h3b7fad2b),
	.w2(32'h3c2ba6b8),
	.w3(32'hbb15df83),
	.w4(32'h3b927386),
	.w5(32'h3bb24da7),
	.w6(32'hbb9eb685),
	.w7(32'h3a87cabe),
	.w8(32'hbb9cc99f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30bce3),
	.w1(32'h39d5348b),
	.w2(32'hb878d1c8),
	.w3(32'h3b8e422a),
	.w4(32'hbabf45c6),
	.w5(32'h3b0f5c51),
	.w6(32'hbb39ae2a),
	.w7(32'h3a8f72d5),
	.w8(32'h3af6f54b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8caef4d),
	.w1(32'h3b8ed5a4),
	.w2(32'h3bce6b56),
	.w3(32'h3a76fca4),
	.w4(32'h3c073443),
	.w5(32'hba87da3a),
	.w6(32'h3a539904),
	.w7(32'hbb245fba),
	.w8(32'hba046a42),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b67a8),
	.w1(32'h3aa523b9),
	.w2(32'hb792155f),
	.w3(32'hbb41d4f3),
	.w4(32'hbbb0cd50),
	.w5(32'hbbcb916f),
	.w6(32'hb9c3bc13),
	.w7(32'hbbca1303),
	.w8(32'hbbab43e2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e55e3),
	.w1(32'hbabb5eb9),
	.w2(32'hba94168d),
	.w3(32'h3b30a144),
	.w4(32'hbb81d86d),
	.w5(32'h3b3ebe95),
	.w6(32'h3a472a67),
	.w7(32'hbb826b8f),
	.w8(32'hba932c72),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24366f),
	.w1(32'hbb1e82cb),
	.w2(32'h3b0eb4d8),
	.w3(32'hbbc1f62a),
	.w4(32'hba9e481c),
	.w5(32'hbb575007),
	.w6(32'hbc05674a),
	.w7(32'hb89a18ea),
	.w8(32'hbb5786a8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13b98b),
	.w1(32'hbb351c9f),
	.w2(32'hbc0c2186),
	.w3(32'hbb5d20ed),
	.w4(32'h3b9c4bdb),
	.w5(32'h3b0978a4),
	.w6(32'hbbe14317),
	.w7(32'h3c096f21),
	.w8(32'hbc1ada3e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4328ce),
	.w1(32'h3b841930),
	.w2(32'hbc0521fa),
	.w3(32'h3bd83229),
	.w4(32'hbb59eed6),
	.w5(32'hbc836a48),
	.w6(32'h3aa3ba37),
	.w7(32'hbbbf788b),
	.w8(32'hbcaad4ec),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d2fdc),
	.w1(32'hbaaa666b),
	.w2(32'hbcafb136),
	.w3(32'h3c594589),
	.w4(32'hbab38472),
	.w5(32'hbcb8037c),
	.w6(32'h3c686429),
	.w7(32'hbbbe8fd2),
	.w8(32'hbc9d7548),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac51076),
	.w1(32'hbada3068),
	.w2(32'hbb74550a),
	.w3(32'hbaac3980),
	.w4(32'hbb093e9e),
	.w5(32'hbb885e80),
	.w6(32'hbb02beb9),
	.w7(32'hbac3fc7d),
	.w8(32'hbb6b9e17),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b65b02),
	.w1(32'h3b0e2359),
	.w2(32'h3aaf3c61),
	.w3(32'h39ba60a4),
	.w4(32'h3b952826),
	.w5(32'hbb04e9b2),
	.w6(32'hba9f4fbb),
	.w7(32'h3b50c891),
	.w8(32'hbae7d641),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec8d69),
	.w1(32'h3b5331f4),
	.w2(32'h3b2d5900),
	.w3(32'hb69c3e10),
	.w4(32'h39d76148),
	.w5(32'hbadd8901),
	.w6(32'h3b2a6d69),
	.w7(32'h3b119c96),
	.w8(32'h3b0f184c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c571e),
	.w1(32'hbaa941ca),
	.w2(32'hbb28d16b),
	.w3(32'hb885cb04),
	.w4(32'hb996829a),
	.w5(32'hb9338132),
	.w6(32'hba944195),
	.w7(32'h3b3e9c23),
	.w8(32'h39a7e179),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1734d2),
	.w1(32'h3c26f0a6),
	.w2(32'hba37dea6),
	.w3(32'hbc236b98),
	.w4(32'h3c3365c4),
	.w5(32'h3b6dff37),
	.w6(32'hbbcbeb8d),
	.w7(32'h3c01f91e),
	.w8(32'hb63e8e10),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe25d7),
	.w1(32'h3baaa6b6),
	.w2(32'hba04ab73),
	.w3(32'h3ac0f1e8),
	.w4(32'h3a230776),
	.w5(32'hbab1fcdc),
	.w6(32'h378995f6),
	.w7(32'hb9b0b977),
	.w8(32'hbac505c6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c009170),
	.w1(32'h3c105304),
	.w2(32'h3c2ae99d),
	.w3(32'hbb1bf549),
	.w4(32'h3b354c5d),
	.w5(32'h3ccabec7),
	.w6(32'hbbba7fc5),
	.w7(32'h3b59f1ae),
	.w8(32'hbb7b1ec1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc084fd),
	.w1(32'h3b8b8c69),
	.w2(32'hba77cc23),
	.w3(32'h39a3c4e3),
	.w4(32'h3aefff46),
	.w5(32'hbb88b726),
	.w6(32'h3b1f3f5d),
	.w7(32'h3b864e2f),
	.w8(32'h3bdc0402),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23751a),
	.w1(32'hb9f7d02a),
	.w2(32'h3b574e4f),
	.w3(32'hbb65eb8c),
	.w4(32'hbb37a040),
	.w5(32'hba8bee6e),
	.w6(32'hbbaad51d),
	.w7(32'h3ab136b0),
	.w8(32'hba286064),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21418d),
	.w1(32'h39d048fd),
	.w2(32'hba539e36),
	.w3(32'hbb7ef366),
	.w4(32'h3b994da6),
	.w5(32'hb971fd45),
	.w6(32'hbaa7c798),
	.w7(32'h3b675ef4),
	.w8(32'h3bcc09dc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f79c8),
	.w1(32'h3a015ff2),
	.w2(32'hb9a16a20),
	.w3(32'h3a9b555e),
	.w4(32'h389b25d4),
	.w5(32'h3b8915bd),
	.w6(32'h3b963501),
	.w7(32'h3a92c6a1),
	.w8(32'h3bd3e838),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a39a8),
	.w1(32'hbaff62d5),
	.w2(32'hbb4a8a1f),
	.w3(32'h3bcd10ee),
	.w4(32'hba0eda6d),
	.w5(32'hbacb7e73),
	.w6(32'h3bab80b3),
	.w7(32'h3b2a17d9),
	.w8(32'h3a7cee4a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc121ed5),
	.w1(32'h3bd1d372),
	.w2(32'hbb159e4b),
	.w3(32'hbab2ee60),
	.w4(32'h3c0ad401),
	.w5(32'hbb9ff04d),
	.w6(32'hbaa636f6),
	.w7(32'h3b74caa9),
	.w8(32'hbbc5e431),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3790ad),
	.w1(32'hba70256d),
	.w2(32'h38bbc7c3),
	.w3(32'hbb91d232),
	.w4(32'hba1ea53b),
	.w5(32'hbb4e6990),
	.w6(32'hbbcf712e),
	.w7(32'hbb3e3059),
	.w8(32'hbb45eaf3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc379bb8),
	.w1(32'hb92b1e19),
	.w2(32'hbb1136a7),
	.w3(32'hbc41c14b),
	.w4(32'h3bbde4d3),
	.w5(32'h3ae7ec06),
	.w6(32'hbc1be6d1),
	.w7(32'h3b8753cd),
	.w8(32'h3abb991a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50c849),
	.w1(32'hbbaea28c),
	.w2(32'h3b92a194),
	.w3(32'hbb9f0d67),
	.w4(32'hbbaadfd3),
	.w5(32'hbb02d7de),
	.w6(32'hba1e93ca),
	.w7(32'h3b2f3058),
	.w8(32'h3aa6ded4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6a4bd),
	.w1(32'h3a39b4d2),
	.w2(32'h3b5ef890),
	.w3(32'h3aa189c0),
	.w4(32'h3b8f17ae),
	.w5(32'h3b262797),
	.w6(32'h3af5a9b9),
	.w7(32'h3a39bd8e),
	.w8(32'hbb0e805f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb625699),
	.w1(32'h3b18e6c7),
	.w2(32'h3950a5e3),
	.w3(32'hba923d54),
	.w4(32'h3b5eb38f),
	.w5(32'h3aef28a6),
	.w6(32'h3a99704f),
	.w7(32'h3b49a0fd),
	.w8(32'h3b1dfddb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf1efd),
	.w1(32'h3a8ddbea),
	.w2(32'h3b16c424),
	.w3(32'h3b896d66),
	.w4(32'hbb848b46),
	.w5(32'h3aec9af3),
	.w6(32'h3bada2cc),
	.w7(32'hbb1af64d),
	.w8(32'hba92c365),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb127ca0),
	.w1(32'hbb4a708c),
	.w2(32'hba3fd29b),
	.w3(32'hb9c14e47),
	.w4(32'hba94f82b),
	.w5(32'hb99d45c8),
	.w6(32'hbb26c70a),
	.w7(32'hba963e72),
	.w8(32'hba7bdb1d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6e7e2),
	.w1(32'hbba949e8),
	.w2(32'hbb3464ac),
	.w3(32'h3b05d1e8),
	.w4(32'hbbb5fb82),
	.w5(32'hbb8d99bc),
	.w6(32'h3b743e8f),
	.w7(32'hbb9f6f71),
	.w8(32'hbb2aadb3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb174301),
	.w1(32'hbab819cb),
	.w2(32'hbb9e2195),
	.w3(32'hbb4fbc80),
	.w4(32'hbb0fe0fc),
	.w5(32'hbaacde8a),
	.w6(32'h3b45c6f2),
	.w7(32'h3bd7ee1f),
	.w8(32'h3c0b632a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79fd32),
	.w1(32'h3b0f78d1),
	.w2(32'h3881a607),
	.w3(32'hb9ef039a),
	.w4(32'h3b57d803),
	.w5(32'hba61ced6),
	.w6(32'h3c72f17a),
	.w7(32'h3c01df78),
	.w8(32'h3bca2e5c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b702115),
	.w1(32'hbbf2fad6),
	.w2(32'hbbc0f0b3),
	.w3(32'hb88f6485),
	.w4(32'hbb9128d5),
	.w5(32'hbb811bfc),
	.w6(32'hbb125f66),
	.w7(32'h38b591c6),
	.w8(32'hb867602d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b148bfe),
	.w1(32'h3b8af599),
	.w2(32'h3b3af2e7),
	.w3(32'hbb3cf314),
	.w4(32'h3b8f54dd),
	.w5(32'h3c114fff),
	.w6(32'h3b1d14c4),
	.w7(32'h3b8789a3),
	.w8(32'h3b11875f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82ae9b),
	.w1(32'h3ba71983),
	.w2(32'h3a2a7dbd),
	.w3(32'h3bc5721f),
	.w4(32'h3b9d19d3),
	.w5(32'hba87eda2),
	.w6(32'h3b23eb05),
	.w7(32'h3bae1bcd),
	.w8(32'h3b0969c7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77ed28),
	.w1(32'h3ad1a2d0),
	.w2(32'h3b4f641d),
	.w3(32'h3b8b9c09),
	.w4(32'h3b841bd3),
	.w5(32'hbaabbb75),
	.w6(32'h3b2a9011),
	.w7(32'h3b1e81c2),
	.w8(32'h39c44e75),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3044bd),
	.w1(32'hbb90c15f),
	.w2(32'hbbbdd902),
	.w3(32'hbbfc6d02),
	.w4(32'h3be507e5),
	.w5(32'h3c074286),
	.w6(32'hbc16b5a1),
	.w7(32'h3b27c01d),
	.w8(32'h3bf19d16),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb64cb),
	.w1(32'h3ba2a561),
	.w2(32'h3b0797b7),
	.w3(32'hbbe1f8c8),
	.w4(32'hbbca1b08),
	.w5(32'hbc345260),
	.w6(32'hbbe4240d),
	.w7(32'hbb607f3f),
	.w8(32'hbb601336),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a48e16),
	.w1(32'h3bcdcdfb),
	.w2(32'hbaacc171),
	.w3(32'hbb1b2ed4),
	.w4(32'h3bc78da5),
	.w5(32'hbb8a6653),
	.w6(32'hb5360e6c),
	.w7(32'h3be28e04),
	.w8(32'h39e9ef90),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c407463),
	.w1(32'h3bfc5ca4),
	.w2(32'hbb964473),
	.w3(32'hbaa21ed0),
	.w4(32'hbbaf61d8),
	.w5(32'hbc74cff2),
	.w6(32'h3b3c8ec7),
	.w7(32'hbc5b35d1),
	.w8(32'hbcf1135c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd22e72),
	.w1(32'hbb563983),
	.w2(32'hbb93cdf7),
	.w3(32'hbbee8029),
	.w4(32'hbb7e887c),
	.w5(32'hbb127168),
	.w6(32'hbc020406),
	.w7(32'hbaba72e7),
	.w8(32'hbb23fbde),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba980244),
	.w1(32'hba922e7f),
	.w2(32'h386b033d),
	.w3(32'hbb1a41cc),
	.w4(32'hbb670a00),
	.w5(32'h3a0a75fd),
	.w6(32'hbabab73f),
	.w7(32'hbb577b4d),
	.w8(32'hbb558766),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba387e06),
	.w1(32'hba9569a7),
	.w2(32'hbb04993c),
	.w3(32'hb9dd9384),
	.w4(32'hbb86ed8b),
	.w5(32'hbb9237bb),
	.w6(32'hbaf65fdb),
	.w7(32'hbb8587d3),
	.w8(32'hbbc44cfc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba36d97),
	.w1(32'hbb5b6408),
	.w2(32'hbb6d21a0),
	.w3(32'hbbe8c593),
	.w4(32'h3a5a53ea),
	.w5(32'h3ac0a891),
	.w6(32'hbc09e09b),
	.w7(32'hbaef777c),
	.w8(32'hba9270a7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0c10),
	.w1(32'hbbb6fb15),
	.w2(32'hbb33b99f),
	.w3(32'hbaa301da),
	.w4(32'hbb4e3e6c),
	.w5(32'hbb8653f9),
	.w6(32'hbace4a53),
	.w7(32'h3b6c87b0),
	.w8(32'h3b52e1a1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6e531),
	.w1(32'hbb9a1368),
	.w2(32'hbbabef09),
	.w3(32'hbbd63892),
	.w4(32'hbb5859c0),
	.w5(32'h3b3cd4d2),
	.w6(32'hba1b5f37),
	.w7(32'hbb504efe),
	.w8(32'hba864339),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cb35c),
	.w1(32'hbc029a0a),
	.w2(32'hbae277a4),
	.w3(32'hbb9ecbb2),
	.w4(32'hbc01a3cd),
	.w5(32'hbb4b7932),
	.w6(32'hbc02f321),
	.w7(32'hbbb81b33),
	.w8(32'hba06b849),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e7222),
	.w1(32'hba67ede1),
	.w2(32'hbbde3643),
	.w3(32'hbbdc75d8),
	.w4(32'h3b176d9d),
	.w5(32'h3bb194da),
	.w6(32'hbb345127),
	.w7(32'hbb84e14f),
	.w8(32'hbc33fa6f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc183cdd),
	.w1(32'h3a7ef44e),
	.w2(32'hba1d4e2c),
	.w3(32'hbbceb040),
	.w4(32'h3b3c7a3b),
	.w5(32'hb97176a4),
	.w6(32'hbc2527af),
	.w7(32'h3b57ca83),
	.w8(32'h3ab5b3ae),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43d7f7),
	.w1(32'hbb897a8b),
	.w2(32'hbb9ce45e),
	.w3(32'hbbd3c111),
	.w4(32'hbb34fb2c),
	.w5(32'h3b48e0fc),
	.w6(32'hbb9f232e),
	.w7(32'hbad27e20),
	.w8(32'hbadaba8d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e293b),
	.w1(32'h3bf4b29b),
	.w2(32'hbb225850),
	.w3(32'hbbb88724),
	.w4(32'h3c20a117),
	.w5(32'h3b735f1f),
	.w6(32'hbb3a4cc1),
	.w7(32'h3b979578),
	.w8(32'h3bb99308),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce552b),
	.w1(32'h3b217063),
	.w2(32'h3b260734),
	.w3(32'h3b0247a3),
	.w4(32'h3b4b1cd8),
	.w5(32'h3b24b39d),
	.w6(32'h3b1249a4),
	.w7(32'h3b83dbc6),
	.w8(32'h3b08541c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39826c46),
	.w1(32'hba7de07c),
	.w2(32'hbaed2276),
	.w3(32'h39956807),
	.w4(32'h3a021db9),
	.w5(32'hbaf32b27),
	.w6(32'hbb0ba5be),
	.w7(32'hbace2df8),
	.w8(32'h399e1522),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1fedc),
	.w1(32'hbbd85c78),
	.w2(32'hbc2b19d6),
	.w3(32'hbacbb511),
	.w4(32'hba5fc378),
	.w5(32'hbaee2025),
	.w6(32'h3b13fb3b),
	.w7(32'hbba23f4d),
	.w8(32'hbb714f9e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71a472),
	.w1(32'hba2c9770),
	.w2(32'h3a1228e0),
	.w3(32'hba6c439d),
	.w4(32'hb9aedef0),
	.w5(32'hbadf6a42),
	.w6(32'hbbc2f251),
	.w7(32'h3ad74f48),
	.w8(32'hbaad82c2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1f306),
	.w1(32'hbb4dbe7e),
	.w2(32'hbbf4cd4c),
	.w3(32'h3b86fe2b),
	.w4(32'hbb955ec1),
	.w5(32'hbbbf1cad),
	.w6(32'h3a5719d9),
	.w7(32'hbbbb7dba),
	.w8(32'hbbbd9c58),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d8d2b),
	.w1(32'hb83fbcdc),
	.w2(32'hbb86be0b),
	.w3(32'hbbaf761e),
	.w4(32'hb9f15f42),
	.w5(32'hbb22310e),
	.w6(32'hbb9c6205),
	.w7(32'hbb60ec56),
	.w8(32'hbb978e4b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a517000),
	.w1(32'h39839af6),
	.w2(32'hbb690f82),
	.w3(32'h3916b90b),
	.w4(32'h3b390ec6),
	.w5(32'h3b3119ef),
	.w6(32'hbb8ba29b),
	.w7(32'h3b11236e),
	.w8(32'h3bc4b1fd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03a35a),
	.w1(32'h3adafa82),
	.w2(32'hbb1b2ddd),
	.w3(32'hb99add4c),
	.w4(32'hbb2cf473),
	.w5(32'hbb96ec3f),
	.w6(32'hbbaa9589),
	.w7(32'hbbc082d6),
	.w8(32'hbbe24acf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd01afc),
	.w1(32'h3a9ca505),
	.w2(32'h3ba0d8b4),
	.w3(32'hbc0a0b02),
	.w4(32'h3a2cb04c),
	.w5(32'h3bb0c551),
	.w6(32'hbc7ab777),
	.w7(32'hbb38898c),
	.w8(32'hbace3c34),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c033f62),
	.w1(32'h3a15e012),
	.w2(32'hbbdb2e47),
	.w3(32'h3be051e7),
	.w4(32'hbb8c96b8),
	.w5(32'hbc461da8),
	.w6(32'h3baf90a4),
	.w7(32'hbb401706),
	.w8(32'hbc4b83d9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04336c),
	.w1(32'hbbec0b3f),
	.w2(32'hbb75a3b0),
	.w3(32'hbc22ec19),
	.w4(32'hbb1434e4),
	.w5(32'h3b9fed44),
	.w6(32'hbc87e1c1),
	.w7(32'hb89dd30c),
	.w8(32'h3ac9795f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab5e17),
	.w1(32'h3bbb0a22),
	.w2(32'h3bc38d7d),
	.w3(32'hb83bc5b8),
	.w4(32'h3aed3bc7),
	.w5(32'hbabaed69),
	.w6(32'h3b45d31f),
	.w7(32'hba84ddd1),
	.w8(32'hbb8cc215),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01125e),
	.w1(32'h3bb52792),
	.w2(32'h3aac3c1d),
	.w3(32'h3ab99f2d),
	.w4(32'h3c037f3f),
	.w5(32'h3beefce0),
	.w6(32'hbbc742ec),
	.w7(32'hbb629554),
	.w8(32'hbb4b121e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75fdae),
	.w1(32'hb890a199),
	.w2(32'hbb92b066),
	.w3(32'h3a61beb2),
	.w4(32'h3ba3af04),
	.w5(32'h3c3fd86c),
	.w6(32'hbb3d031c),
	.w7(32'hbab4ddaf),
	.w8(32'hbbaf643a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efed61),
	.w1(32'hbb95eb4f),
	.w2(32'hbc1ee5ff),
	.w3(32'h3b26169d),
	.w4(32'hbb9a3e2d),
	.w5(32'hbbec3178),
	.w6(32'h3b52ac40),
	.w7(32'hbbdad120),
	.w8(32'hbc192f57),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf53a2d),
	.w1(32'hba698b73),
	.w2(32'hbb6d814a),
	.w3(32'h3a06f0e9),
	.w4(32'hba829c21),
	.w5(32'hbb606e7d),
	.w6(32'h397c93e3),
	.w7(32'h3a3ad690),
	.w8(32'hbb6c34e3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bd4de),
	.w1(32'h3befde73),
	.w2(32'h3aaa10a5),
	.w3(32'hbc059bce),
	.w4(32'h3b8d76b4),
	.w5(32'h39f197f8),
	.w6(32'hbc33996c),
	.w7(32'h3b5a7698),
	.w8(32'h39667068),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf76859),
	.w1(32'hbb09f1cf),
	.w2(32'hba8895a2),
	.w3(32'hbbdfd828),
	.w4(32'hba8cf7de),
	.w5(32'h3ab9227e),
	.w6(32'hba83279b),
	.w7(32'h3b8f77ed),
	.w8(32'h39e58262),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e57d5),
	.w1(32'hbc2e5f47),
	.w2(32'hbb529364),
	.w3(32'hbbedb3be),
	.w4(32'hbbd627cc),
	.w5(32'h3b9685b6),
	.w6(32'hbc748ab3),
	.w7(32'hbb0bf187),
	.w8(32'hbbda95d6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28d30a),
	.w1(32'hbbb5a29b),
	.w2(32'hbc37751f),
	.w3(32'hbbd35802),
	.w4(32'hbb886a51),
	.w5(32'hbb8f7779),
	.w6(32'hbc06682a),
	.w7(32'hbc208e09),
	.w8(32'hbc42e7f4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfee4b7),
	.w1(32'h3c277797),
	.w2(32'h3a3734b3),
	.w3(32'h3b63ce1c),
	.w4(32'h3b74d0b0),
	.w5(32'hba54399b),
	.w6(32'hb908bb50),
	.w7(32'h3b8305ab),
	.w8(32'hbb85adea),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed4963),
	.w1(32'hbbbda2be),
	.w2(32'hba61c323),
	.w3(32'hba475e36),
	.w4(32'hba9fa7f0),
	.w5(32'h3bbf16f0),
	.w6(32'hbaed00ea),
	.w7(32'h395cfb00),
	.w8(32'h3b16c349),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819fd5),
	.w1(32'hbaf03661),
	.w2(32'h3a88c355),
	.w3(32'hba5f9a8a),
	.w4(32'h3a96fff9),
	.w5(32'h3a6047bb),
	.w6(32'hbbb6c9fe),
	.w7(32'h3bb9d631),
	.w8(32'hba479d21),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c2aad),
	.w1(32'h3ac5a8a5),
	.w2(32'hbbf617fe),
	.w3(32'hbb9b534e),
	.w4(32'h3ba32350),
	.w5(32'h3bae476f),
	.w6(32'hbc211ada),
	.w7(32'h3b8883ca),
	.w8(32'hbb9d5949),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac548e1),
	.w1(32'h3b47608e),
	.w2(32'hb9f0ec5b),
	.w3(32'hbb6f32f4),
	.w4(32'h3b8bbb73),
	.w5(32'hbb242b77),
	.w6(32'hbafcf3c7),
	.w7(32'h3add8b29),
	.w8(32'hb95f8cb5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bae8e),
	.w1(32'hba9475d0),
	.w2(32'hba8285f4),
	.w3(32'h3b028fc3),
	.w4(32'h3b3b88e6),
	.w5(32'h3a9480f4),
	.w6(32'h39c1d27a),
	.w7(32'h3b4a35d0),
	.w8(32'h3b7c4596),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb842811),
	.w1(32'hbac25a8f),
	.w2(32'hb7df2139),
	.w3(32'hbac7b644),
	.w4(32'hbb3366ee),
	.w5(32'hb9468978),
	.w6(32'hb92aba42),
	.w7(32'hbbb9d5b4),
	.w8(32'hbbcf76a9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f59bf),
	.w1(32'h3bb5462e),
	.w2(32'h3b109bb5),
	.w3(32'hbbe382a0),
	.w4(32'h3b4f31e1),
	.w5(32'h3a99baf7),
	.w6(32'hbc0c1610),
	.w7(32'h3b4b5cd1),
	.w8(32'hb9f9f5f3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be774e1),
	.w1(32'h39065907),
	.w2(32'hbbdc570f),
	.w3(32'h3a98c7d9),
	.w4(32'hbb60b1b8),
	.w5(32'hbba7cf64),
	.w6(32'h3b9a90e8),
	.w7(32'h3a35cdf1),
	.w8(32'hbba42432),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0349a),
	.w1(32'hbb8f8243),
	.w2(32'hbb9deaf3),
	.w3(32'hbb48cc4f),
	.w4(32'hbb37f021),
	.w5(32'hbab8fbfe),
	.w6(32'h3b208543),
	.w7(32'hbb74507a),
	.w8(32'hbc2f6561),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a974912),
	.w1(32'h38ab1506),
	.w2(32'hbbac64ac),
	.w3(32'h3b4796f8),
	.w4(32'hbb318ad9),
	.w5(32'hba628fb6),
	.w6(32'hbb3ad984),
	.w7(32'hbbfc3bc2),
	.w8(32'hbc1e0aae),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc047206),
	.w1(32'h3a5b864d),
	.w2(32'hbad85216),
	.w3(32'hbc476251),
	.w4(32'hbb9b2e0b),
	.w5(32'hb984d5f7),
	.w6(32'hbc36e4d3),
	.w7(32'hbae5afed),
	.w8(32'h3acf53d1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64689a),
	.w1(32'hbac00d25),
	.w2(32'hbbaada20),
	.w3(32'h3a250d24),
	.w4(32'h3bf8091d),
	.w5(32'h3b9b6f13),
	.w6(32'hbb663e3b),
	.w7(32'h3ab02f80),
	.w8(32'hba88c4dc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a2c8e),
	.w1(32'h3a8d5597),
	.w2(32'hba900bd0),
	.w3(32'hbb8afe63),
	.w4(32'hb9ec542a),
	.w5(32'hbb9970a6),
	.w6(32'hbb7ea680),
	.w7(32'hbbb93c12),
	.w8(32'hbc15edde),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae351c8),
	.w1(32'hbbbb7fe8),
	.w2(32'hbba9455e),
	.w3(32'h3b8c5e05),
	.w4(32'hbb728122),
	.w5(32'hbb3a4117),
	.w6(32'hbb2933cb),
	.w7(32'hbb88e403),
	.w8(32'hbb5dc7d6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd50ac),
	.w1(32'h3b16738a),
	.w2(32'hbaacd89b),
	.w3(32'hbbb841cd),
	.w4(32'h3b7fbdbe),
	.w5(32'hba6c451c),
	.w6(32'hbb853c2f),
	.w7(32'h3b85c34f),
	.w8(32'h3b01cf90),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e83f4a),
	.w1(32'h3a99e5c4),
	.w2(32'h3b12a38a),
	.w3(32'h3b02c4df),
	.w4(32'h3b7bb45f),
	.w5(32'hba049da1),
	.w6(32'h3a9a0d88),
	.w7(32'h3a021eb6),
	.w8(32'hbb3f0520),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc0e20),
	.w1(32'hbb26c767),
	.w2(32'hbb3d46a9),
	.w3(32'h39516d48),
	.w4(32'hbba7ef52),
	.w5(32'hbb2917ed),
	.w6(32'hb8b9a702),
	.w7(32'hbad38da9),
	.w8(32'hbb10b3ab),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58469d),
	.w1(32'h3b13d643),
	.w2(32'hbb69f71d),
	.w3(32'hbb34a4bd),
	.w4(32'h3b222409),
	.w5(32'h3aae9251),
	.w6(32'hba65048c),
	.w7(32'h3a5fe6fb),
	.w8(32'h37d2f29e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fc6b5),
	.w1(32'hbb817083),
	.w2(32'hbb138abf),
	.w3(32'h3ad9a6dd),
	.w4(32'hbb903302),
	.w5(32'hbbae1140),
	.w6(32'h3b9a60e0),
	.w7(32'hbb48249c),
	.w8(32'h3b2664a8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb633b1),
	.w1(32'h3b1814e0),
	.w2(32'hba1b107e),
	.w3(32'hbc2e50c6),
	.w4(32'hbbb8813d),
	.w5(32'hbb8aff13),
	.w6(32'hbc1fb01d),
	.w7(32'hbbafcd71),
	.w8(32'hbbd59476),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeb18c),
	.w1(32'h3a0fb90d),
	.w2(32'hbc421cb4),
	.w3(32'h3aec4759),
	.w4(32'h3aa4161b),
	.w5(32'hbbc40dee),
	.w6(32'hba23712a),
	.w7(32'hbb1323f2),
	.w8(32'hbc2e20d3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d3178),
	.w1(32'h3b8e64f1),
	.w2(32'hba42ebef),
	.w3(32'hbb0f9763),
	.w4(32'h3a975bc4),
	.w5(32'h3baec19d),
	.w6(32'hbb0d1324),
	.w7(32'h3b8a8046),
	.w8(32'h3ac8228d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef8da2),
	.w1(32'h3aa379c9),
	.w2(32'h3b4625fb),
	.w3(32'h3baadd2c),
	.w4(32'h3b50140d),
	.w5(32'h3b3df5be),
	.w6(32'h3bf85a28),
	.w7(32'h3b9bfdae),
	.w8(32'hba80dfae),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ead0c9),
	.w1(32'hbb87f99b),
	.w2(32'hba03e588),
	.w3(32'h396ad032),
	.w4(32'hbba617a2),
	.w5(32'hbafb79d6),
	.w6(32'h3af9685b),
	.w7(32'hbb859ccd),
	.w8(32'hbb4a4ece),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abad3c8),
	.w1(32'hbabc512e),
	.w2(32'hba1ea2d0),
	.w3(32'hbb2eb9f7),
	.w4(32'hbb10ff89),
	.w5(32'hbb8e602f),
	.w6(32'hbb97993a),
	.w7(32'h3ae7e669),
	.w8(32'hbbb1a215),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add089b),
	.w1(32'hbba8c896),
	.w2(32'h37b826b6),
	.w3(32'hbc08fb8f),
	.w4(32'hbc2520a2),
	.w5(32'hbbb545a8),
	.w6(32'hbc77d43a),
	.w7(32'hbbc0dae1),
	.w8(32'hbc2b2de0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd21a07),
	.w1(32'hbb087b17),
	.w2(32'hbb170757),
	.w3(32'hbbbc4469),
	.w4(32'hbac549db),
	.w5(32'h3b2bb6b8),
	.w6(32'hbbb02d43),
	.w7(32'h389ad665),
	.w8(32'h3b5b6df9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84d588),
	.w1(32'hbbafde7f),
	.w2(32'hbb25c9db),
	.w3(32'hb98d34e9),
	.w4(32'hbbd9a46d),
	.w5(32'h3946b00c),
	.w6(32'h3b492318),
	.w7(32'hbba77876),
	.w8(32'hbb093a4d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba63867),
	.w1(32'h3a9cbd9e),
	.w2(32'hbb952365),
	.w3(32'hbba64981),
	.w4(32'h3b40813d),
	.w5(32'h39f8a62b),
	.w6(32'hbb2b282e),
	.w7(32'hbad448db),
	.w8(32'h3a6fb2bc),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39708072),
	.w1(32'hb8b9d920),
	.w2(32'h3b4417c6),
	.w3(32'h3b1a81e6),
	.w4(32'h3b11491f),
	.w5(32'h3b753751),
	.w6(32'h3b467519),
	.w7(32'hba7aed5c),
	.w8(32'hba563b8e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e2d6d),
	.w1(32'hbb45065e),
	.w2(32'hbb3d88f8),
	.w3(32'hbb602f6b),
	.w4(32'hbb1ba05f),
	.w5(32'h39d3ba77),
	.w6(32'hbb815185),
	.w7(32'hbad8c6d8),
	.w8(32'hba10a066),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccb9d2),
	.w1(32'h3bafb1df),
	.w2(32'hbb0ee206),
	.w3(32'hbb3f91ae),
	.w4(32'h3bf3185d),
	.w5(32'h3bf93b9b),
	.w6(32'h3b0bacfb),
	.w7(32'h3b33bc10),
	.w8(32'hbbec4eaa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f9d0a),
	.w1(32'hbbb50261),
	.w2(32'hbb052fbf),
	.w3(32'hbb8269b1),
	.w4(32'h3afe9c3a),
	.w5(32'h3c0e70d6),
	.w6(32'hbbd3a403),
	.w7(32'h3a0b1f81),
	.w8(32'h3ad123bb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01a42a),
	.w1(32'h3ac1e827),
	.w2(32'hbb8bc399),
	.w3(32'h3be99d86),
	.w4(32'h3a8a7820),
	.w5(32'hbafcb5ae),
	.w6(32'h3ba1d4b8),
	.w7(32'hbbc47e2c),
	.w8(32'hbc0ba213),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab58c5),
	.w1(32'hbaa164e4),
	.w2(32'h3b2eee9f),
	.w3(32'hbaffb0d7),
	.w4(32'h3bc46b08),
	.w5(32'h3b8c790e),
	.w6(32'hbc13115a),
	.w7(32'h3bbf3d84),
	.w8(32'h3aa8276f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb838363),
	.w1(32'hbbcf1be5),
	.w2(32'h3a5f274a),
	.w3(32'hbbb1d0c7),
	.w4(32'hba912578),
	.w5(32'h3a7a243c),
	.w6(32'hbbe99928),
	.w7(32'h3ad9f66d),
	.w8(32'h3a5d3fad),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c37614),
	.w1(32'h3a75e919),
	.w2(32'hb9dd39b1),
	.w3(32'hbb36c6fe),
	.w4(32'hbada5153),
	.w5(32'h3a9cd2e3),
	.w6(32'hbb523307),
	.w7(32'hbb313704),
	.w8(32'hbb8de184),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3908a8),
	.w1(32'hbb633814),
	.w2(32'hbb850881),
	.w3(32'hbac82028),
	.w4(32'hba343867),
	.w5(32'hbad1c6f1),
	.w6(32'hbb78ecbe),
	.w7(32'h3a7d860b),
	.w8(32'hb9f89f3d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9210a5),
	.w1(32'hbb385c4e),
	.w2(32'h3a9a1831),
	.w3(32'hbba2ad18),
	.w4(32'h3b5c785b),
	.w5(32'hba808f99),
	.w6(32'hbb6615b8),
	.w7(32'hba8bb478),
	.w8(32'hba7b381c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74e62b),
	.w1(32'h3b2c6671),
	.w2(32'hbba12db2),
	.w3(32'h3bdf6416),
	.w4(32'hbb4dc84c),
	.w5(32'hbc403ee5),
	.w6(32'h3c3fc123),
	.w7(32'hbbc8e2f4),
	.w8(32'hbc878ca4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79e39f),
	.w1(32'hbb064283),
	.w2(32'hbb524c91),
	.w3(32'h3ad513dc),
	.w4(32'hbb2721c0),
	.w5(32'hbb9da11a),
	.w6(32'hbacbb9e4),
	.w7(32'hb9a2e64c),
	.w8(32'hbbbeb96f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11bf67),
	.w1(32'h3988a6aa),
	.w2(32'hba856373),
	.w3(32'hba86c166),
	.w4(32'h3b7765e7),
	.w5(32'h3ad6145f),
	.w6(32'hbb2d1381),
	.w7(32'h3b1fa05a),
	.w8(32'h39b77097),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2966da),
	.w1(32'hbc0cdf2b),
	.w2(32'hbc1bff1a),
	.w3(32'h3a8ef877),
	.w4(32'hbbd4ed50),
	.w5(32'hbba89962),
	.w6(32'hbb293bc7),
	.w7(32'hbb26d657),
	.w8(32'hbab83512),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbca128),
	.w1(32'hbb2300ec),
	.w2(32'hbb41f690),
	.w3(32'hbbfd6215),
	.w4(32'h3b001957),
	.w5(32'hba8f066a),
	.w6(32'hbb93f943),
	.w7(32'hba0dc6f2),
	.w8(32'h3ab063ae),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc55781),
	.w1(32'h3b472190),
	.w2(32'hbb3c32cc),
	.w3(32'h3b9e413a),
	.w4(32'h3af9b09d),
	.w5(32'hbb361f6a),
	.w6(32'h3ae86a27),
	.w7(32'h3b03a6d5),
	.w8(32'hbbb23d3a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cc188),
	.w1(32'hb9ef423e),
	.w2(32'h3a71faa4),
	.w3(32'hbaea669f),
	.w4(32'hbb7eeb91),
	.w5(32'hbacddb67),
	.w6(32'h3ab8b762),
	.w7(32'hb9c0626c),
	.w8(32'hbb1835dc),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8db49),
	.w1(32'hba926159),
	.w2(32'hbaac786b),
	.w3(32'hb84c7772),
	.w4(32'hba51cca8),
	.w5(32'hbb624968),
	.w6(32'hbbc23b90),
	.w7(32'hbaffb4c6),
	.w8(32'hbb95e826),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73b0ff),
	.w1(32'hbac11ab4),
	.w2(32'hbb825661),
	.w3(32'hbb8f2832),
	.w4(32'hbad5214e),
	.w5(32'hbbaca756),
	.w6(32'hbbc5aa13),
	.w7(32'hba1f78bb),
	.w8(32'hbc27846a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bc035),
	.w1(32'hbab61f25),
	.w2(32'hbb831975),
	.w3(32'hbbdb320f),
	.w4(32'hbac57f87),
	.w5(32'hbb5413c1),
	.w6(32'hbc0e4785),
	.w7(32'hbb544ac9),
	.w8(32'hbb5e934c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a7eeb),
	.w1(32'hbbbc5c7c),
	.w2(32'h3a7b88a5),
	.w3(32'hbc14d2cc),
	.w4(32'hbbaa5606),
	.w5(32'h3abcaa5e),
	.w6(32'hbbefe19d),
	.w7(32'hbba0a975),
	.w8(32'hbb833ca6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a7960),
	.w1(32'h3b0a731d),
	.w2(32'hbc15d224),
	.w3(32'h3c07474d),
	.w4(32'h37fdf474),
	.w5(32'hbbe2559e),
	.w6(32'h3c202b1c),
	.w7(32'hba980573),
	.w8(32'hbc3aed73),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aee3c),
	.w1(32'h3a3b1088),
	.w2(32'hbb4c9329),
	.w3(32'h3ab91fe7),
	.w4(32'hbaea17bf),
	.w5(32'hbc0034a9),
	.w6(32'hbb9e0895),
	.w7(32'hbbdc7081),
	.w8(32'hbc3031a0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa73463),
	.w1(32'h3b95d4cd),
	.w2(32'hbaf35aea),
	.w3(32'hba6f603a),
	.w4(32'h3b0fd6a4),
	.w5(32'hbb6483a7),
	.w6(32'hbbe986ae),
	.w7(32'hbb8ff125),
	.w8(32'hbc0126a9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8135f5),
	.w1(32'h3b82e557),
	.w2(32'h3ae07726),
	.w3(32'h3a2008c2),
	.w4(32'h3956299d),
	.w5(32'hbb9a9c3a),
	.w6(32'hbc0def14),
	.w7(32'hbb682cb1),
	.w8(32'hbbdef248),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b6fe5),
	.w1(32'hbaefd4ed),
	.w2(32'hbbdb32a8),
	.w3(32'hba23083c),
	.w4(32'hba4c75e0),
	.w5(32'hbb88f108),
	.w6(32'hbb05dd60),
	.w7(32'h3a46cd08),
	.w8(32'hbb35d322),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9843c50),
	.w1(32'h3be3d148),
	.w2(32'h3a8ac6a8),
	.w3(32'hba9f78ad),
	.w4(32'h3b53e0ae),
	.w5(32'hbaa3dbe4),
	.w6(32'h3b864558),
	.w7(32'h3ac73e32),
	.w8(32'hbadea26b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa52702),
	.w1(32'hbbaae16f),
	.w2(32'hbae69a59),
	.w3(32'h37ef5f3f),
	.w4(32'hbbfcc96d),
	.w5(32'hbae704a7),
	.w6(32'hbb81c7fb),
	.w7(32'h3afb79e8),
	.w8(32'h3b5de171),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66e2ca),
	.w1(32'h39879ab9),
	.w2(32'hbb812377),
	.w3(32'hbacd3bfb),
	.w4(32'h3bc2bbef),
	.w5(32'h3b590177),
	.w6(32'h3b316392),
	.w7(32'h3ae90de3),
	.w8(32'h3b6812dc),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe344),
	.w1(32'hbb023f4a),
	.w2(32'hbb8c4fd4),
	.w3(32'hbb37f89a),
	.w4(32'hb9ef9057),
	.w5(32'h3a16c6a4),
	.w6(32'hbad4d0cf),
	.w7(32'hbb5f5460),
	.w8(32'hbb1c13aa),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4405f1),
	.w1(32'hbab9a651),
	.w2(32'hbb413be7),
	.w3(32'hbb31854d),
	.w4(32'h3b743384),
	.w5(32'h3b7f590f),
	.w6(32'hbbac5519),
	.w7(32'hbb3a3d98),
	.w8(32'hbb40132f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6d7e7),
	.w1(32'h3babf565),
	.w2(32'h3a5f8db9),
	.w3(32'h3b31a3e5),
	.w4(32'hb9c2098b),
	.w5(32'hbbdcf72f),
	.w6(32'hbab9884a),
	.w7(32'hbbacce82),
	.w8(32'hbbfda995),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043082),
	.w1(32'hbaa15602),
	.w2(32'hbab09f1c),
	.w3(32'h3b3e402a),
	.w4(32'h38f406da),
	.w5(32'hb95475e7),
	.w6(32'hbacda2e2),
	.w7(32'hbb2e30a1),
	.w8(32'hbb2f7189),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9171e),
	.w1(32'hbb112152),
	.w2(32'hba9a4b7a),
	.w3(32'hbade52df),
	.w4(32'hbb647573),
	.w5(32'hbaa2d4a0),
	.w6(32'hbba3e3cd),
	.w7(32'hbb25917c),
	.w8(32'hbb6b94b9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb426ad8),
	.w1(32'hbb69d971),
	.w2(32'hbb368385),
	.w3(32'hb9bec10c),
	.w4(32'h3b8398c6),
	.w5(32'h3b18b3c9),
	.w6(32'h385e48b4),
	.w7(32'h3a445a34),
	.w8(32'h3b1f1155),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe65e0a),
	.w1(32'hb8cb697a),
	.w2(32'h3a95958b),
	.w3(32'hb7ae7d81),
	.w4(32'hb981138a),
	.w5(32'h3ab8ecdc),
	.w6(32'h3a716c1b),
	.w7(32'h3b3873cb),
	.w8(32'h3b650e18),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba76fa3),
	.w1(32'hba73972d),
	.w2(32'hbb764c42),
	.w3(32'h3b69340c),
	.w4(32'h37d550a7),
	.w5(32'hbb49b1c5),
	.w6(32'h3be06ae8),
	.w7(32'hbb8fb541),
	.w8(32'hbbc63610),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d9210),
	.w1(32'hbad41f9b),
	.w2(32'h3b083401),
	.w3(32'hbbfa339b),
	.w4(32'hbc1d27d7),
	.w5(32'hbc29a4ad),
	.w6(32'hbc711f5a),
	.w7(32'hbc0178fa),
	.w8(32'hbc22a9b3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0d436),
	.w1(32'h3b4a55f2),
	.w2(32'hba03a741),
	.w3(32'hbb9c1a28),
	.w4(32'hba877421),
	.w5(32'hbb317153),
	.w6(32'hbc25884b),
	.w7(32'hb930d637),
	.w8(32'hbb685ce4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9addc9),
	.w1(32'h3b991a93),
	.w2(32'hb91b37ca),
	.w3(32'h3b3243ef),
	.w4(32'h3bce6225),
	.w5(32'h3aa4281c),
	.w6(32'h3b5b0970),
	.w7(32'h3b064d78),
	.w8(32'hba5b77de),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a360bf0),
	.w1(32'hba063235),
	.w2(32'h3909939d),
	.w3(32'h3b31022a),
	.w4(32'h3acf854f),
	.w5(32'h3aabb3fc),
	.w6(32'h3ab32ca2),
	.w7(32'hba55b4d9),
	.w8(32'h39b17358),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f808d),
	.w1(32'h3bcedf42),
	.w2(32'h3964cee1),
	.w3(32'hbbb2df28),
	.w4(32'h3bdc5bc6),
	.w5(32'h3abe4eab),
	.w6(32'hbb73ede8),
	.w7(32'h3be9d8dc),
	.w8(32'hbad434a8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29e756),
	.w1(32'h3af8076d),
	.w2(32'hbb5b1e5a),
	.w3(32'hbb7e1b07),
	.w4(32'h3b897d0a),
	.w5(32'h3b85c317),
	.w6(32'hbbd4b79c),
	.w7(32'h3b669dac),
	.w8(32'h3a1871df),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc653),
	.w1(32'hbb34f6dd),
	.w2(32'hbb39c016),
	.w3(32'hbb8b21fa),
	.w4(32'hb9604134),
	.w5(32'hbaad438a),
	.w6(32'hbbb3ede6),
	.w7(32'hb9e639ab),
	.w8(32'hbb4c7eee),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a411e1e),
	.w1(32'h3b30c4dd),
	.w2(32'h3acd77d0),
	.w3(32'hbb101104),
	.w4(32'h3a7b90bc),
	.w5(32'h3ae434ad),
	.w6(32'hbb3b657f),
	.w7(32'hb9860a32),
	.w8(32'hbad20ded),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0dcf2),
	.w1(32'h3a827e57),
	.w2(32'hba9d5965),
	.w3(32'h3a5a9285),
	.w4(32'h3a47a135),
	.w5(32'hbb029e8b),
	.w6(32'h3ab281e5),
	.w7(32'h3be2759a),
	.w8(32'h3a5dcc63),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27ce96),
	.w1(32'h3b11e17a),
	.w2(32'hbb793d29),
	.w3(32'h3a1be580),
	.w4(32'hbaccd535),
	.w5(32'hbb8b6b99),
	.w6(32'hba78f9f9),
	.w7(32'hbb265b48),
	.w8(32'hba903fed),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab527ad),
	.w1(32'hbb298d7a),
	.w2(32'hba462b75),
	.w3(32'h3ae40743),
	.w4(32'hbbdf39bc),
	.w5(32'hbb740401),
	.w6(32'hbb3aa033),
	.w7(32'hbbe6a0d0),
	.w8(32'hbbd04e31),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd32b35),
	.w1(32'hba26ebc5),
	.w2(32'hbb473d9f),
	.w3(32'hbbe30eb0),
	.w4(32'hbafe91ed),
	.w5(32'hbb4f0fb6),
	.w6(32'hbb90b8ce),
	.w7(32'hbb6596fe),
	.w8(32'hbba61981),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd148d5),
	.w1(32'h3c14e7ad),
	.w2(32'h3c027122),
	.w3(32'hbc0b6ead),
	.w4(32'h3c11e3c7),
	.w5(32'h3bf06d5f),
	.w6(32'hbbcaa3b6),
	.w7(32'h3a7ded9e),
	.w8(32'h36f46f5c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb141d8),
	.w1(32'hbb461745),
	.w2(32'hbb00b7b9),
	.w3(32'h3bbecdf5),
	.w4(32'h3b1be10d),
	.w5(32'h3ac5284f),
	.w6(32'hbb0ffc58),
	.w7(32'hbb204d37),
	.w8(32'hbaa83ea4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b3ed8),
	.w1(32'hbb046e68),
	.w2(32'h3a6de264),
	.w3(32'h3bac800b),
	.w4(32'hbb3edf29),
	.w5(32'hba6a8db0),
	.w6(32'hbb8d6f68),
	.w7(32'hbbada920),
	.w8(32'hbb4862cf),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948eb9),
	.w1(32'hb9f7e40f),
	.w2(32'h393df634),
	.w3(32'hbb213249),
	.w4(32'h3b9686f3),
	.w5(32'h3bb316ae),
	.w6(32'hbb4181ee),
	.w7(32'h3a9b8c0e),
	.w8(32'h3b500d2d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb607a00),
	.w1(32'h3ba8a1a6),
	.w2(32'hbb0b1c63),
	.w3(32'h3a09fdf3),
	.w4(32'h3b95c130),
	.w5(32'h3ba79522),
	.w6(32'hbb04b883),
	.w7(32'h3bfbe1fc),
	.w8(32'h3b20587d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc211183),
	.w1(32'hbbb6b708),
	.w2(32'h39412cff),
	.w3(32'hbb8498a0),
	.w4(32'hbb012621),
	.w5(32'hbb605762),
	.w6(32'h3b6c1e8f),
	.w7(32'hbb97faa4),
	.w8(32'hbc3c1f86),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c7d1f),
	.w1(32'hba4b0e80),
	.w2(32'h392a01c8),
	.w3(32'hbba17fe1),
	.w4(32'hbad7729a),
	.w5(32'hbb4cb2a6),
	.w6(32'hbbc8aebf),
	.w7(32'hba681a36),
	.w8(32'hbb782bc8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d567f),
	.w1(32'h39c70df5),
	.w2(32'h3b0131c7),
	.w3(32'hbc591b2a),
	.w4(32'h3b84792a),
	.w5(32'hba26c054),
	.w6(32'hbc5e67b3),
	.w7(32'h39aa3662),
	.w8(32'hbb10b969),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeefdad),
	.w1(32'h3bf0b5a6),
	.w2(32'hbbd2a137),
	.w3(32'h3b01622c),
	.w4(32'h39ab3cc4),
	.w5(32'h3a1a1e4e),
	.w6(32'h3a4836b6),
	.w7(32'hbba02621),
	.w8(32'hbc64dfec),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecca46),
	.w1(32'hba37a470),
	.w2(32'hbb5033e9),
	.w3(32'hbbbe766a),
	.w4(32'hb7e91b4d),
	.w5(32'h3acfd23b),
	.w6(32'hbc237fbe),
	.w7(32'hbb1c453f),
	.w8(32'hbad426de),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecc9e5),
	.w1(32'hbb713975),
	.w2(32'hbb0be596),
	.w3(32'h3ab05c1f),
	.w4(32'hbae37f9b),
	.w5(32'hba6c61f5),
	.w6(32'hbb00e0e4),
	.w7(32'h3b147e77),
	.w8(32'h3b4e44a6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d4160),
	.w1(32'hbbc7ed4d),
	.w2(32'hbb6a120b),
	.w3(32'h3993ebee),
	.w4(32'hbb205bbe),
	.w5(32'hba205674),
	.w6(32'h3ad7f021),
	.w7(32'h3ae2ec6d),
	.w8(32'h3b58f29f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb8b16),
	.w1(32'h3b17a96e),
	.w2(32'hb9819103),
	.w3(32'hbbb0083f),
	.w4(32'h3bd7dcfe),
	.w5(32'h3b8e83d2),
	.w6(32'hbacdb271),
	.w7(32'h3bd97ba8),
	.w8(32'h3bf42ae8),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c8f46),
	.w1(32'hbbd4e29b),
	.w2(32'hbb6fcf94),
	.w3(32'h3b18d271),
	.w4(32'hbb0a044e),
	.w5(32'h3abf5ecd),
	.w6(32'h3b5cea56),
	.w7(32'hbac900d1),
	.w8(32'hbb616abf),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899c267),
	.w1(32'h3bba91cd),
	.w2(32'h3bb87661),
	.w3(32'h3c09e2bc),
	.w4(32'h3b776afb),
	.w5(32'hbadfc849),
	.w6(32'hba3e3f7c),
	.w7(32'h3b27c6d9),
	.w8(32'hbaa4a606),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0de294),
	.w1(32'h3ba75fa4),
	.w2(32'hbb92c71a),
	.w3(32'h3b18e287),
	.w4(32'h3b77566d),
	.w5(32'h3a468a27),
	.w6(32'h3acf4aa7),
	.w7(32'hbaaa7e3b),
	.w8(32'hbb999226),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbce2a),
	.w1(32'hbaaa71a9),
	.w2(32'hbaf660f7),
	.w3(32'h3bb50a46),
	.w4(32'hbb8f8ee9),
	.w5(32'hbb729798),
	.w6(32'hbb0a8d91),
	.w7(32'hbb80c28e),
	.w8(32'hbb814f45),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2c84e),
	.w1(32'h3b820f47),
	.w2(32'h3bf94557),
	.w3(32'hbbf3816a),
	.w4(32'h3b03b15f),
	.w5(32'h393fa886),
	.w6(32'hbbe1aab4),
	.w7(32'h3b091e1c),
	.w8(32'h3b75e55c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00e30b),
	.w1(32'hbac19b6b),
	.w2(32'h3b3f0d41),
	.w3(32'hba890b6e),
	.w4(32'hba930dff),
	.w5(32'hbb36aac4),
	.w6(32'hbb26e285),
	.w7(32'h3a311f98),
	.w8(32'hbb41337f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d66325),
	.w1(32'hbadc8173),
	.w2(32'h3b2aaaac),
	.w3(32'hbc3f8416),
	.w4(32'hbc34c30c),
	.w5(32'hbb702816),
	.w6(32'hbacf4fc3),
	.w7(32'hbc16f434),
	.w8(32'hbc14b6fd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c2693),
	.w1(32'h3b93fe0f),
	.w2(32'h3b5b9711),
	.w3(32'hbb9373ae),
	.w4(32'h39dc7edc),
	.w5(32'h3bd6b522),
	.w6(32'hbb5722af),
	.w7(32'h3c2b9366),
	.w8(32'h3bd0c138),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d90c),
	.w1(32'hbbccf132),
	.w2(32'hbb7c1ee0),
	.w3(32'hba170194),
	.w4(32'h3c17d4bb),
	.w5(32'h3c74f4cf),
	.w6(32'hb98771a9),
	.w7(32'h3a9fa419),
	.w8(32'h3c1e7b4b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38abc001),
	.w1(32'h39e042ba),
	.w2(32'h3afab9e8),
	.w3(32'h3c18b84c),
	.w4(32'hbc956b09),
	.w5(32'hbcd963ef),
	.w6(32'h3b05403c),
	.w7(32'hbbc0c5fb),
	.w8(32'hbcac613a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a9470),
	.w1(32'h3bea6369),
	.w2(32'hbc2be17f),
	.w3(32'hbc5ecb92),
	.w4(32'h3c8d5719),
	.w5(32'h3cb52c69),
	.w6(32'hbcaa6bb1),
	.w7(32'hbb077f00),
	.w8(32'h3bf48d7d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcda51b),
	.w1(32'h3b138562),
	.w2(32'hbb959bc4),
	.w3(32'hba2b7ff8),
	.w4(32'h3a600f10),
	.w5(32'hbbdbfd32),
	.w6(32'hba3ecdba),
	.w7(32'h3b5df541),
	.w8(32'h39f81dc4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcde1bb),
	.w1(32'hbc387a84),
	.w2(32'hbb7e46f7),
	.w3(32'hbb7d0783),
	.w4(32'h3b73296e),
	.w5(32'h3d19db19),
	.w6(32'h3a8c9039),
	.w7(32'hbb1f9df8),
	.w8(32'h3c4b4a14),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92ce51),
	.w1(32'h3b9e1baf),
	.w2(32'h3bc7dc45),
	.w3(32'hb9b8402f),
	.w4(32'h3b5fafcf),
	.w5(32'h3a1fa4ec),
	.w6(32'hbadac390),
	.w7(32'h3bb99145),
	.w8(32'hbbaa3e66),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997a823),
	.w1(32'h3b3a58c0),
	.w2(32'hbbaa4876),
	.w3(32'h3bae8319),
	.w4(32'hb9948480),
	.w5(32'hba3fe803),
	.w6(32'hbb1128f0),
	.w7(32'h3b8d6fe8),
	.w8(32'h3b8974cf),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8526),
	.w1(32'h3c73a796),
	.w2(32'h3c8f5375),
	.w3(32'hbb951b4a),
	.w4(32'h3b9f77a9),
	.w5(32'h3b07bd2d),
	.w6(32'hbbe3015f),
	.w7(32'h3c16ce07),
	.w8(32'hbadc15d9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34b368),
	.w1(32'h3932931c),
	.w2(32'h39812f31),
	.w3(32'h3c64d4c1),
	.w4(32'h3a17f831),
	.w5(32'h3b48b1d6),
	.w6(32'h3c7eb5a8),
	.w7(32'hbac1e04f),
	.w8(32'h3b5d9673),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4253aa),
	.w1(32'hbc6c26c4),
	.w2(32'hbc3e6fc4),
	.w3(32'hba47fe80),
	.w4(32'hbc7f93e9),
	.w5(32'hbcc57c44),
	.w6(32'hbb147e43),
	.w7(32'hbc678dd6),
	.w8(32'hbcb464ba),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5189f8),
	.w1(32'h3b85896d),
	.w2(32'h3b266fb6),
	.w3(32'hbccf98bc),
	.w4(32'h3b0cd94a),
	.w5(32'hbbcb7a72),
	.w6(32'hbc9e4e88),
	.w7(32'h3a6356c2),
	.w8(32'hbb7048b0),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40a575),
	.w1(32'hbb983b69),
	.w2(32'hbb96155e),
	.w3(32'hbb44d20d),
	.w4(32'hbbe33558),
	.w5(32'hbc3009db),
	.w6(32'hbc58a98b),
	.w7(32'hbb2a34ee),
	.w8(32'hbc5105fb),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd17701),
	.w1(32'h3b9f9d60),
	.w2(32'hba7b4984),
	.w3(32'hbafa5dd1),
	.w4(32'h3a88cd9c),
	.w5(32'h3b699578),
	.w6(32'hbc017cfc),
	.w7(32'hbbecdaa6),
	.w8(32'hbbc93c65),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda1c43),
	.w1(32'hbc5f5c93),
	.w2(32'hba3918a0),
	.w3(32'hbb219d78),
	.w4(32'hba712ca6),
	.w5(32'h3cd8cb1f),
	.w6(32'hbae86f04),
	.w7(32'hbb2026cc),
	.w8(32'h3c13c565),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bc8ee),
	.w1(32'hbb434db7),
	.w2(32'hbc0d283a),
	.w3(32'h3b8ac918),
	.w4(32'h3b441080),
	.w5(32'h3d04cb11),
	.w6(32'h39830fe6),
	.w7(32'h3b43d009),
	.w8(32'h3ba4ec4e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b8958),
	.w1(32'hbb32d83c),
	.w2(32'h3b020c7d),
	.w3(32'h3b559172),
	.w4(32'h3bc46352),
	.w5(32'hbbd4f45b),
	.w6(32'h38a3b2e4),
	.w7(32'h3b51f9d3),
	.w8(32'h3ac39fe8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfde24f),
	.w1(32'hbadd62c3),
	.w2(32'hba868f5f),
	.w3(32'hbbf4d1e0),
	.w4(32'hb828fd5f),
	.w5(32'h3c3e335a),
	.w6(32'hbc1fd13b),
	.w7(32'h3abf9392),
	.w8(32'h3c13e5d6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81bce2),
	.w1(32'hbaec364e),
	.w2(32'h3b83657d),
	.w3(32'hbbd86ed7),
	.w4(32'hba9b63dd),
	.w5(32'hba1d23c5),
	.w6(32'hbc225fd4),
	.w7(32'hbb6bd562),
	.w8(32'hba3f044b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90d48a),
	.w1(32'hbc2598f1),
	.w2(32'h3a9a848c),
	.w3(32'hbc0b601d),
	.w4(32'hbc04d384),
	.w5(32'hbb338fec),
	.w6(32'hbbd8756e),
	.w7(32'hbbae4f24),
	.w8(32'hbbc44561),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ab0b),
	.w1(32'hbc075328),
	.w2(32'hbc9431c0),
	.w3(32'h39d17c01),
	.w4(32'hbc6963a8),
	.w5(32'hbc9b4f13),
	.w6(32'hba78a66d),
	.w7(32'hbc5a9a92),
	.w8(32'hbccebd89),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec4863),
	.w1(32'h3c8d4292),
	.w2(32'h3c9d5293),
	.w3(32'hbbdf96fd),
	.w4(32'h3c7db37b),
	.w5(32'h3cbfed24),
	.w6(32'hbb2547b8),
	.w7(32'h3b24c1c1),
	.w8(32'h3bb0dbfa),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c364c80),
	.w1(32'h3b2448da),
	.w2(32'h3aafb6fb),
	.w3(32'h3c6ab4b7),
	.w4(32'h3af5e92d),
	.w5(32'hb9cf36a0),
	.w6(32'h3c0b4f25),
	.w7(32'h3bc89599),
	.w8(32'h3b0830e7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69e7f5),
	.w1(32'hbb6fd761),
	.w2(32'hbc712545),
	.w3(32'hbad8f3f4),
	.w4(32'h3b8c75df),
	.w5(32'hbc27403b),
	.w6(32'h3b9978a8),
	.w7(32'h3c4d686c),
	.w8(32'hba5d63b8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0befe6),
	.w1(32'hbb8e9e53),
	.w2(32'hbbc10615),
	.w3(32'hbb759192),
	.w4(32'hbb98cff7),
	.w5(32'hbbab12a8),
	.w6(32'hbb6f726d),
	.w7(32'h3c09cef1),
	.w8(32'hbb4d7a31),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ebb0a),
	.w1(32'h3bd15df4),
	.w2(32'h3b9940d7),
	.w3(32'hb9e9fb05),
	.w4(32'hbc273e26),
	.w5(32'h3c0eb6cc),
	.w6(32'hbb7c54f8),
	.w7(32'hbc4e2d77),
	.w8(32'hba0b2bcf),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa52c2a),
	.w1(32'hb7e26b79),
	.w2(32'hbbe3356d),
	.w3(32'hbb8a50e3),
	.w4(32'hba771e54),
	.w5(32'hbb4f4a6d),
	.w6(32'hbbc25581),
	.w7(32'hbbbbf3b0),
	.w8(32'h39140d2c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb965641),
	.w1(32'h3b697e90),
	.w2(32'h3aefd187),
	.w3(32'hbc1974ef),
	.w4(32'h3c437dad),
	.w5(32'h3c8b3c0b),
	.w6(32'hbb9ae5c9),
	.w7(32'h3b82f366),
	.w8(32'h3c01215d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f8696),
	.w1(32'h3c1ea45b),
	.w2(32'h37ce3f3b),
	.w3(32'h3aaf9852),
	.w4(32'h3c2f0e36),
	.w5(32'h3c8764c5),
	.w6(32'h3b80bd8f),
	.w7(32'h3aa9ec51),
	.w8(32'h3c160d47),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c2ef3),
	.w1(32'hbc2e32c3),
	.w2(32'hbc363aa8),
	.w3(32'h3c3c5f27),
	.w4(32'hbbb83534),
	.w5(32'hbbb23048),
	.w6(32'h3b72939a),
	.w7(32'hbc1f4743),
	.w8(32'hbca08224),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74f032),
	.w1(32'hbc299802),
	.w2(32'h3c56843d),
	.w3(32'hbc3953d6),
	.w4(32'hbc762dfd),
	.w5(32'hbbd2694b),
	.w6(32'hbcbe06f8),
	.w7(32'hbc541048),
	.w8(32'hbb54c529),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fb49b),
	.w1(32'hbbdd7ea0),
	.w2(32'hbc2b99f7),
	.w3(32'hbcac897e),
	.w4(32'hbc045bae),
	.w5(32'hbc549906),
	.w6(32'hbc0cb7ed),
	.w7(32'hbb411d26),
	.w8(32'hbcaab0a0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0faf54),
	.w1(32'hbb9cef04),
	.w2(32'hbc64ef66),
	.w3(32'h3ad914c8),
	.w4(32'hbb2ea04c),
	.w5(32'hbbcb2b63),
	.w6(32'hbc3a3758),
	.w7(32'h3b1e7dd8),
	.w8(32'hbc5c7754),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85d43d),
	.w1(32'hbb7d5fcb),
	.w2(32'hbb6bae4e),
	.w3(32'hbc4ef754),
	.w4(32'hbb9ef2d0),
	.w5(32'hb96c71a8),
	.w6(32'hbb8e650f),
	.w7(32'hbae1a9df),
	.w8(32'hbb4086ef),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61f03e),
	.w1(32'h3b9a9ecf),
	.w2(32'hbbc3e864),
	.w3(32'hbb562842),
	.w4(32'h3be2c6d5),
	.w5(32'hba5953eb),
	.w6(32'h3ac56f04),
	.w7(32'h3b10d77c),
	.w8(32'h3c297c72),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29e489),
	.w1(32'hbb368dca),
	.w2(32'h3b7dc089),
	.w3(32'hbbe82197),
	.w4(32'hbae64376),
	.w5(32'h3c0ea33d),
	.w6(32'h39d2af48),
	.w7(32'h3a80b5f2),
	.w8(32'h3aec00f3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a7bdf),
	.w1(32'h3b68dc72),
	.w2(32'hbad6ec57),
	.w3(32'h3a33b5fb),
	.w4(32'h3a50be9f),
	.w5(32'h3a76e869),
	.w6(32'h3b45617c),
	.w7(32'h3b8845ce),
	.w8(32'hbc0a29e7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a35825),
	.w1(32'h3a085dfa),
	.w2(32'hbb71627f),
	.w3(32'hbb5c44e5),
	.w4(32'h3b8653b8),
	.w5(32'h3c5d11fd),
	.w6(32'hbad7053e),
	.w7(32'h3c0cc137),
	.w8(32'hbc155a46),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977006),
	.w1(32'h3c052c97),
	.w2(32'h3b309dcf),
	.w3(32'hbba33b62),
	.w4(32'hbaa851c8),
	.w5(32'hbc008750),
	.w6(32'hbb7184a0),
	.w7(32'h3a89487f),
	.w8(32'h3a237601),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee7ad2),
	.w1(32'h3c3e3827),
	.w2(32'hbb1897f7),
	.w3(32'hbbd841ea),
	.w4(32'h3be6942d),
	.w5(32'h3990e55a),
	.w6(32'hba804263),
	.w7(32'h3c1f8eac),
	.w8(32'h3c01ce44),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3824a),
	.w1(32'hbb88b273),
	.w2(32'hba4f9ad5),
	.w3(32'hbbae55ae),
	.w4(32'hbbe4645e),
	.w5(32'hbba776f9),
	.w6(32'hbabbdf43),
	.w7(32'h39e55497),
	.w8(32'hb959eb1f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa8f97),
	.w1(32'hbbf6d07a),
	.w2(32'hbceadea4),
	.w3(32'hbb3ce3b5),
	.w4(32'h3c1299df),
	.w5(32'hbc6a77a2),
	.w6(32'hbbfa799a),
	.w7(32'h3c0d37f0),
	.w8(32'h3c198d2d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5aafde),
	.w1(32'h3c332c1d),
	.w2(32'h3b137c85),
	.w3(32'hbbdd958f),
	.w4(32'h3b7edab0),
	.w5(32'h3b2da7f0),
	.w6(32'hbb1841a3),
	.w7(32'h3aac962d),
	.w8(32'hba026e9c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c71c45),
	.w1(32'hba430fdd),
	.w2(32'h3bccb3f3),
	.w3(32'hb9b8dde7),
	.w4(32'hbb2914a9),
	.w5(32'h3b9f4dcd),
	.w6(32'h3abaaf31),
	.w7(32'hbacdc0ba),
	.w8(32'hbb16e2bb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f2d68),
	.w1(32'h39e27533),
	.w2(32'hbb993fce),
	.w3(32'hbb42389f),
	.w4(32'h3b90249e),
	.w5(32'h3bbed026),
	.w6(32'h3bba71ce),
	.w7(32'h3ba4ab96),
	.w8(32'h3b57c2ac),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cd0f4),
	.w1(32'h3bb1abe6),
	.w2(32'h3b9b2c10),
	.w3(32'h3a727957),
	.w4(32'hbb459fe0),
	.w5(32'hbb459b43),
	.w6(32'h3b9b8f68),
	.w7(32'h3ac221fc),
	.w8(32'h3a118f4a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0fe3f),
	.w1(32'h3b8371c4),
	.w2(32'h3bd042f1),
	.w3(32'hbbb9902b),
	.w4(32'h3c6df0a6),
	.w5(32'h3cc9ed13),
	.w6(32'hbbf8a228),
	.w7(32'h3c1504cb),
	.w8(32'h3b95561e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c001792),
	.w1(32'hba2d408c),
	.w2(32'h3b937458),
	.w3(32'h3c4338b9),
	.w4(32'h3a2b1aa8),
	.w5(32'h3c93e963),
	.w6(32'hbaab98a3),
	.w7(32'hbcc0c940),
	.w8(32'hbc79eff8),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc955fde),
	.w1(32'hba8d019c),
	.w2(32'h39311e3c),
	.w3(32'h37d0c9dc),
	.w4(32'h3bc732c5),
	.w5(32'hba4d2723),
	.w6(32'h3b22f217),
	.w7(32'h3b196e8d),
	.w8(32'h3aabe1f5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb957916),
	.w1(32'h3a033f0e),
	.w2(32'hbba03545),
	.w3(32'h392c6542),
	.w4(32'h3a02daa8),
	.w5(32'hbc195f72),
	.w6(32'h3bec4004),
	.w7(32'h3be13e99),
	.w8(32'h3c352a18),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ca146),
	.w1(32'hbb9710cd),
	.w2(32'h3b175207),
	.w3(32'h39dd7ce3),
	.w4(32'hbbbf8fa1),
	.w5(32'hbaf5d93e),
	.w6(32'h3c149eb7),
	.w7(32'hbb367294),
	.w8(32'hbb706722),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9d7d5),
	.w1(32'h3b7386ba),
	.w2(32'h3b8338ec),
	.w3(32'hbc13b7ad),
	.w4(32'hbb216c73),
	.w5(32'hbbb10fab),
	.w6(32'hbb403c65),
	.w7(32'h3ae48acc),
	.w8(32'hbba30261),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b415a),
	.w1(32'h3c0bdab9),
	.w2(32'hb9dde1e2),
	.w3(32'h3ba7ae98),
	.w4(32'hb9699539),
	.w5(32'h3c82d624),
	.w6(32'h3ab72304),
	.w7(32'h3b8ef576),
	.w8(32'h3b2371fb),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81ec4e),
	.w1(32'h3c014bfc),
	.w2(32'hbb7c8a7a),
	.w3(32'hbb034292),
	.w4(32'h3c55f58c),
	.w5(32'h3b8b2b94),
	.w6(32'hbb877097),
	.w7(32'h3c085cc8),
	.w8(32'hbb7a5c00),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa8809),
	.w1(32'hbbd72ace),
	.w2(32'hbc13b770),
	.w3(32'hba95582d),
	.w4(32'hbac3e98d),
	.w5(32'hbc055956),
	.w6(32'hbb1a6753),
	.w7(32'hbb786204),
	.w8(32'h3bd2d112),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0334e),
	.w1(32'h3c579b7c),
	.w2(32'h3c638f66),
	.w3(32'hbb04a86d),
	.w4(32'h3ba977b8),
	.w5(32'hbabd4206),
	.w6(32'hbbea5357),
	.w7(32'hbb34e019),
	.w8(32'h3a21a078),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule