module layer_10_featuremap_6(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb906684),
	.w1(32'h3b5ddcc5),
	.w2(32'h3c6c7cef),
	.w3(32'hbcbb31e7),
	.w4(32'h3b1a771f),
	.w5(32'h3c984302),
	.w6(32'hbb86eb40),
	.w7(32'h3996a266),
	.w8(32'hbc4b9e3d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c958192),
	.w1(32'hbc97bff3),
	.w2(32'h3af5b256),
	.w3(32'h3cb452ba),
	.w4(32'hbc806834),
	.w5(32'hbb7fcdab),
	.w6(32'h3ca71255),
	.w7(32'hbb993792),
	.w8(32'hb985cef0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26ca50),
	.w1(32'hbcd39e29),
	.w2(32'hbb11e3d5),
	.w3(32'h3ca4943e),
	.w4(32'hbc6c0c53),
	.w5(32'hbad2313a),
	.w6(32'h3c2f0716),
	.w7(32'h3b943138),
	.w8(32'h3ba9946d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba732c2),
	.w1(32'hbbc855ed),
	.w2(32'h3b98a68b),
	.w3(32'hbc267ad6),
	.w4(32'hbc9fa167),
	.w5(32'hbc44fb86),
	.w6(32'hbb30a370),
	.w7(32'hbc4e95cf),
	.w8(32'hbc86a343),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42345b),
	.w1(32'hbc202f2c),
	.w2(32'h3cdbbd82),
	.w3(32'h3c9abb88),
	.w4(32'h3bdc8cf9),
	.w5(32'hbca46c47),
	.w6(32'hbb12d706),
	.w7(32'hbaaf52ff),
	.w8(32'h3c2aeca3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9e8fb),
	.w1(32'h3ba1b26b),
	.w2(32'h3a80df55),
	.w3(32'h39e11a6b),
	.w4(32'h3c2447b3),
	.w5(32'hbb60a976),
	.w6(32'hbbf6239f),
	.w7(32'hba0a0f2b),
	.w8(32'hbb8e18b4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9900a52),
	.w1(32'hbad9533a),
	.w2(32'h3b2c2b48),
	.w3(32'hbb667f85),
	.w4(32'h3b30fab2),
	.w5(32'hba22fa21),
	.w6(32'hbba2a9f6),
	.w7(32'hb9754c01),
	.w8(32'hbc195782),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b059e35),
	.w1(32'hbb23bc09),
	.w2(32'h3b3d1178),
	.w3(32'h3bd9cf84),
	.w4(32'h3b2ef0c6),
	.w5(32'hbbef755d),
	.w6(32'hba7e2221),
	.w7(32'h3c01845a),
	.w8(32'h3beb4f4a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b930c45),
	.w1(32'h3a1cf9eb),
	.w2(32'hbaaf3d26),
	.w3(32'hbc5c1b07),
	.w4(32'h3aa123fc),
	.w5(32'h3bbb1a9e),
	.w6(32'h395e0bdf),
	.w7(32'hbb17c8e3),
	.w8(32'h3bd2963a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5387a),
	.w1(32'hbb89da69),
	.w2(32'h3b0a5d9d),
	.w3(32'hbb66bfc3),
	.w4(32'hbc6b7fc0),
	.w5(32'hbb0717e4),
	.w6(32'h39ba0525),
	.w7(32'hbbfaef06),
	.w8(32'h3b15f434),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0be5),
	.w1(32'h3ad39146),
	.w2(32'hbb036c0f),
	.w3(32'hba76c565),
	.w4(32'hbac0179e),
	.w5(32'h3b86ec93),
	.w6(32'hb9ff3aea),
	.w7(32'hbb02898c),
	.w8(32'h3c22fa29),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b8b2f),
	.w1(32'h3b519702),
	.w2(32'hbb0b9067),
	.w3(32'hbc4e3949),
	.w4(32'hbcc40d91),
	.w5(32'h3a8ab6a7),
	.w6(32'h3c0a486b),
	.w7(32'hbcbd71b4),
	.w8(32'h38fafd8f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959d3ec),
	.w1(32'h3b5cef97),
	.w2(32'hbae9a5f5),
	.w3(32'h39edf80d),
	.w4(32'h3b4aba57),
	.w5(32'hba27a637),
	.w6(32'hba286d8e),
	.w7(32'h3b057c36),
	.w8(32'h3b9f3812),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b080c63),
	.w1(32'h3ba6fc23),
	.w2(32'h39781cf6),
	.w3(32'hba67047f),
	.w4(32'h3c1a3096),
	.w5(32'hbbe48715),
	.w6(32'h3af38274),
	.w7(32'hb940b8b5),
	.w8(32'hbb7c2a44),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45ad3),
	.w1(32'hbca333a9),
	.w2(32'hbb336540),
	.w3(32'h3cacb9e4),
	.w4(32'h3c5da85e),
	.w5(32'hbba477c3),
	.w6(32'h3c40b02d),
	.w7(32'h3c36244e),
	.w8(32'h3a968b10),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86f5ad),
	.w1(32'hbb5dd43c),
	.w2(32'h3b10f38c),
	.w3(32'hbbce0bd1),
	.w4(32'hbbb5f5f6),
	.w5(32'hba093961),
	.w6(32'hbb04e97b),
	.w7(32'hbb8854fc),
	.w8(32'h3b7e498b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add7ff3),
	.w1(32'h3a9f491b),
	.w2(32'hbb2ab9ea),
	.w3(32'hba7a8018),
	.w4(32'hb8ab0fa1),
	.w5(32'hbbafd383),
	.w6(32'hb9698077),
	.w7(32'hbaf1008c),
	.w8(32'hb9c3a11b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c95a3),
	.w1(32'h3b8de218),
	.w2(32'hbb1703c8),
	.w3(32'h3b09e14b),
	.w4(32'h3c31ed7e),
	.w5(32'h3a50e2c5),
	.w6(32'h3b00b470),
	.w7(32'h3c4af636),
	.w8(32'h3b65ff9a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997945c),
	.w1(32'hbb13a8cb),
	.w2(32'h3ad8cbf8),
	.w3(32'hbb9730cf),
	.w4(32'h3b828b08),
	.w5(32'h3a9e829f),
	.w6(32'hbadde8f1),
	.w7(32'h3bce7bfd),
	.w8(32'hb95263d8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d6837),
	.w1(32'h3a5a0583),
	.w2(32'hb833800b),
	.w3(32'hbba4fb11),
	.w4(32'hbc4166be),
	.w5(32'h3ad5c255),
	.w6(32'hbadf7e83),
	.w7(32'hbc120eec),
	.w8(32'h3bcd8120),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa30cd9),
	.w1(32'hbb5789b4),
	.w2(32'h3ab3b22c),
	.w3(32'h3be0a9d2),
	.w4(32'hba979214),
	.w5(32'h3c38323f),
	.w6(32'h3bf31f7d),
	.w7(32'h3b19bb29),
	.w8(32'hbbc68d91),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77ca2b),
	.w1(32'h3b809d53),
	.w2(32'hb9eab60e),
	.w3(32'hbbdde96d),
	.w4(32'hba8f06bd),
	.w5(32'hbb18d325),
	.w6(32'hbb0d8304),
	.w7(32'h3b579b9a),
	.w8(32'hbae4ad30),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37842b),
	.w1(32'hbac24460),
	.w2(32'h3b0c926c),
	.w3(32'hbb9c2fc2),
	.w4(32'hbc27ab84),
	.w5(32'h3a15ef99),
	.w6(32'hbb8741ed),
	.w7(32'h3a886c6c),
	.w8(32'h3b452daa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39b4b2),
	.w1(32'hbb761d21),
	.w2(32'hbb17035b),
	.w3(32'hbb1a9a85),
	.w4(32'hbb5e8679),
	.w5(32'hbc0ce2f8),
	.w6(32'h3b9f0e58),
	.w7(32'h3b19cca7),
	.w8(32'hbb3a9146),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77dda8),
	.w1(32'h3c021d62),
	.w2(32'h3b07fac2),
	.w3(32'h3aa34318),
	.w4(32'h3beab681),
	.w5(32'hba7d77af),
	.w6(32'hbbfc4357),
	.w7(32'h3b7cf616),
	.w8(32'h3a1074a9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd70c6c),
	.w1(32'hbc9a235e),
	.w2(32'h3bf44215),
	.w3(32'h3be57e2a),
	.w4(32'hbc29d936),
	.w5(32'hbc528dc9),
	.w6(32'hbc7ed2ee),
	.w7(32'hbc8992d5),
	.w8(32'hbcf6e596),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b437c),
	.w1(32'h38665fc4),
	.w2(32'h39a61b76),
	.w3(32'h3cabe196),
	.w4(32'h3d05f4e1),
	.w5(32'hb8cebc60),
	.w6(32'hbc86258d),
	.w7(32'h3c6345b6),
	.w8(32'h39944b0a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bde57),
	.w1(32'h39b8066a),
	.w2(32'h3b7a77c7),
	.w3(32'h3b4cddb2),
	.w4(32'h39bc8a62),
	.w5(32'h3a6ec2a9),
	.w6(32'h3b915a4d),
	.w7(32'h3b921d3a),
	.w8(32'hbac60866),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7985c),
	.w1(32'hbbf92ac0),
	.w2(32'h3ba571e3),
	.w3(32'hbb24b4dc),
	.w4(32'hbbb8281d),
	.w5(32'hbcc73d0c),
	.w6(32'hbb703e7a),
	.w7(32'hbb8c2139),
	.w8(32'h3b48915e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b96dc),
	.w1(32'h3c936c30),
	.w2(32'hbb8b59ca),
	.w3(32'hbcbe7851),
	.w4(32'hbb6b329d),
	.w5(32'h3a96019f),
	.w6(32'hbb89e481),
	.w7(32'hbbd37ecd),
	.w8(32'h39f7128b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3464f4),
	.w1(32'hb9e6f51d),
	.w2(32'hba1fc570),
	.w3(32'hb95a56ce),
	.w4(32'h3a0c9af6),
	.w5(32'hbb2b1d11),
	.w6(32'hbb3609cb),
	.w7(32'hba9d42dd),
	.w8(32'hbb05adb1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8529bd),
	.w1(32'h3c33ff13),
	.w2(32'hba4bf251),
	.w3(32'hbc2b9bb7),
	.w4(32'hbc0e5c04),
	.w5(32'hbc66edf0),
	.w6(32'h3ab55835),
	.w7(32'hbbb5e913),
	.w8(32'hbb1962cb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b851858),
	.w1(32'hbb22172c),
	.w2(32'h3a7b1a01),
	.w3(32'hbbfe0e26),
	.w4(32'hbc058ccf),
	.w5(32'h3b233bca),
	.w6(32'hbbb44ef5),
	.w7(32'hbc260ce7),
	.w8(32'h3a582885),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8d8ee),
	.w1(32'hbb155e4c),
	.w2(32'hb922e958),
	.w3(32'hbab5eb1e),
	.w4(32'hbb0c777e),
	.w5(32'hbb1f7870),
	.w6(32'hbab8444d),
	.w7(32'hbaf18974),
	.w8(32'hbc477018),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0034c5),
	.w1(32'h3bdbac23),
	.w2(32'hbb128999),
	.w3(32'h3ad45a33),
	.w4(32'h3bbeb6d4),
	.w5(32'hbb3de773),
	.w6(32'hbc98601d),
	.w7(32'hbc336d81),
	.w8(32'hbb511200),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3e762),
	.w1(32'hbb4a6881),
	.w2(32'h3cfe7f28),
	.w3(32'hba39d4dc),
	.w4(32'h38942f3e),
	.w5(32'hbb157e7b),
	.w6(32'hbba86094),
	.w7(32'hbb4b2d7a),
	.w8(32'hbd0e7282),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce54481),
	.w1(32'h3cb37721),
	.w2(32'hba23c663),
	.w3(32'h3be76fb5),
	.w4(32'h3d070f25),
	.w5(32'h3841d3ca),
	.w6(32'hbd86426b),
	.w7(32'hbcc8a16d),
	.w8(32'h3a4344e9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f521f4),
	.w1(32'h398f67e9),
	.w2(32'hbc149627),
	.w3(32'hb8b0683c),
	.w4(32'hbb370431),
	.w5(32'h3ba7f26e),
	.w6(32'h3c069cb2),
	.w7(32'h3b43ffba),
	.w8(32'hb88ee2c1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b326),
	.w1(32'hbc3bce67),
	.w2(32'h3bb3e8bd),
	.w3(32'h3caf47ee),
	.w4(32'h3c68481b),
	.w5(32'hbb94dccd),
	.w6(32'h3c622de5),
	.w7(32'h3ba967ea),
	.w8(32'h3ba2e2ef),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96499b),
	.w1(32'h3bf9bf53),
	.w2(32'hbaf3caab),
	.w3(32'hbc965711),
	.w4(32'hbc18688c),
	.w5(32'hba84971b),
	.w6(32'h3b3970de),
	.w7(32'hbbd3bb36),
	.w8(32'hbc020a53),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02765c),
	.w1(32'hbbee7f27),
	.w2(32'h3a65ac94),
	.w3(32'hbb6babb0),
	.w4(32'h392d27c3),
	.w5(32'h3ba0f384),
	.w6(32'hbc31273b),
	.w7(32'h3a1b311a),
	.w8(32'hbbc0763d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b288f34),
	.w1(32'hbb0c556f),
	.w2(32'hbb714cc8),
	.w3(32'h3c807f91),
	.w4(32'h3c7bb50a),
	.w5(32'hb91dcd5e),
	.w6(32'hbbd9bb77),
	.w7(32'hbc0808ab),
	.w8(32'hbb882647),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8cab1),
	.w1(32'hbacc2b6c),
	.w2(32'h3b2ca324),
	.w3(32'hbc128883),
	.w4(32'hbbfe3457),
	.w5(32'hba767ce5),
	.w6(32'hbb3ed3ab),
	.w7(32'h3bc22be4),
	.w8(32'h3b2d8791),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08d021),
	.w1(32'h3b4f6fdb),
	.w2(32'h3bb8c5fc),
	.w3(32'h3b971530),
	.w4(32'h3ab9e54a),
	.w5(32'h3b81e898),
	.w6(32'h3b86f9f4),
	.w7(32'h3b24d34f),
	.w8(32'h3c38e966),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8de035),
	.w1(32'h3b125f9f),
	.w2(32'hbb749427),
	.w3(32'hbb1fb3b0),
	.w4(32'hbd0c2972),
	.w5(32'hbcd668c3),
	.w6(32'h3ce210d2),
	.w7(32'h3c67cac8),
	.w8(32'h3bcfd2d8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbcc1ab),
	.w1(32'h3bf20813),
	.w2(32'hbb89b1cf),
	.w3(32'hbd124a54),
	.w4(32'hbc6155c7),
	.w5(32'h3c156b0d),
	.w6(32'hbabb2f0d),
	.w7(32'hbbcadc73),
	.w8(32'h3b85fe43),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c255e),
	.w1(32'hbcb4f07e),
	.w2(32'hbbce96b4),
	.w3(32'h3cb30c15),
	.w4(32'h3c040e36),
	.w5(32'h3bf1060a),
	.w6(32'h3bf17a03),
	.w7(32'h3c95dde8),
	.w8(32'hb8d5f932),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ac3b),
	.w1(32'h3beaab8a),
	.w2(32'h3a2a97ac),
	.w3(32'h3c8aabd9),
	.w4(32'h3c9a33f8),
	.w5(32'hbbb81c78),
	.w6(32'hbc85c0bf),
	.w7(32'hbbc44e86),
	.w8(32'hbb2cc0de),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a2566),
	.w1(32'hba944eb8),
	.w2(32'hbc074aa6),
	.w3(32'hbb0c3e5b),
	.w4(32'hbb184a11),
	.w5(32'h3a0bef03),
	.w6(32'hba08ec2a),
	.w7(32'hbb62fa21),
	.w8(32'hbb729fac),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba820db),
	.w1(32'hbb8b3c5e),
	.w2(32'h3ba6a8c8),
	.w3(32'hbb82ba50),
	.w4(32'hbbee7bcc),
	.w5(32'hbc7410fe),
	.w6(32'h3c702da2),
	.w7(32'h3c02c01d),
	.w8(32'hbc528236),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c36db),
	.w1(32'h3ca5f968),
	.w2(32'hbb81862c),
	.w3(32'hbc86c1b5),
	.w4(32'h3b6e4889),
	.w5(32'hbc3b19a5),
	.w6(32'hbcfc3ec9),
	.w7(32'hbcb5c387),
	.w8(32'hbb9dd6ca),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c792a0a),
	.w1(32'hb95ac371),
	.w2(32'h3b85d696),
	.w3(32'hbc88b065),
	.w4(32'hbbc397b5),
	.w5(32'hbc8a330e),
	.w6(32'h3b2c91d4),
	.w7(32'hbab40f21),
	.w8(32'hbc89944e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c65e0),
	.w1(32'h3c96ae41),
	.w2(32'hbb875254),
	.w3(32'hbc583818),
	.w4(32'h3c030684),
	.w5(32'hbb1fdddb),
	.w6(32'hbce397f8),
	.w7(32'hbc7cea91),
	.w8(32'h3b448dc0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca682e),
	.w1(32'hbbcd8086),
	.w2(32'h3bc12caa),
	.w3(32'hbac8edcc),
	.w4(32'h3b06efe4),
	.w5(32'hbba4a2a2),
	.w6(32'hbbcc1c8f),
	.w7(32'hbc09ed96),
	.w8(32'hba721e31),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8075f0),
	.w1(32'h3c73007f),
	.w2(32'h3bf6462e),
	.w3(32'hbc1bde95),
	.w4(32'h3c286386),
	.w5(32'hbbbd3490),
	.w6(32'hbc084634),
	.w7(32'hbbebbfc5),
	.w8(32'hbc501416),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d2ba5),
	.w1(32'h3bd0e0ef),
	.w2(32'hbb757538),
	.w3(32'h3bbf6b0d),
	.w4(32'h3be8fad7),
	.w5(32'h3b069a51),
	.w6(32'hbc83d11e),
	.w7(32'hbbbb8563),
	.w8(32'h3c277fbc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc505ac2),
	.w1(32'hbbdedf4a),
	.w2(32'h37ef3cc6),
	.w3(32'hbc3f9efe),
	.w4(32'hbc6676bb),
	.w5(32'hbb1f55be),
	.w6(32'h3c38d025),
	.w7(32'hbb4c2b7d),
	.w8(32'h3a88fb24),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6752d),
	.w1(32'hbad8abb5),
	.w2(32'hbb93819b),
	.w3(32'h3ba5ac3c),
	.w4(32'hbb2f6eec),
	.w5(32'hbba50486),
	.w6(32'h3c07f701),
	.w7(32'hbb3f1b54),
	.w8(32'h3baf110c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6476c5),
	.w1(32'hbc03ca0b),
	.w2(32'hbb62a58e),
	.w3(32'hbb0868c4),
	.w4(32'hbbdea1cd),
	.w5(32'h39bcc973),
	.w6(32'h3c1f1f30),
	.w7(32'h3a803e55),
	.w8(32'h3c189b69),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4783d),
	.w1(32'h3ad1efd8),
	.w2(32'hbbcd0f08),
	.w3(32'hb972f2d3),
	.w4(32'h3b68a708),
	.w5(32'hbbe98d17),
	.w6(32'h3bc7f256),
	.w7(32'hbc099588),
	.w8(32'h3bc2e068),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8881d5),
	.w1(32'hba71eb67),
	.w2(32'hbc061deb),
	.w3(32'hbba22878),
	.w4(32'hbb44ffa3),
	.w5(32'h3bcc6738),
	.w6(32'hbbb52bd8),
	.w7(32'hbb9b48b5),
	.w8(32'h3b619468),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfc613),
	.w1(32'hbc38dc29),
	.w2(32'hbc251237),
	.w3(32'h3b247074),
	.w4(32'h3b39a4c2),
	.w5(32'h3c4e4535),
	.w6(32'h3c4a2562),
	.w7(32'h3bb90a75),
	.w8(32'h3a89c021),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4daae),
	.w1(32'hbb658a3b),
	.w2(32'h3b11839d),
	.w3(32'hbc051ccc),
	.w4(32'hbbb472c0),
	.w5(32'hba6ba694),
	.w6(32'h3ca42f56),
	.w7(32'h3c807c07),
	.w8(32'h3a4bcc98),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac0c66),
	.w1(32'h397db2da),
	.w2(32'h3b3b3b7c),
	.w3(32'h3a37882c),
	.w4(32'hbbb6d761),
	.w5(32'h3b7c1af8),
	.w6(32'h3b019e46),
	.w7(32'hbb2f79b1),
	.w8(32'h3c2dc1e3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7d79b),
	.w1(32'h3bf7da5d),
	.w2(32'h3a6e01ef),
	.w3(32'hba9804a2),
	.w4(32'h3b3323ad),
	.w5(32'hbae7016e),
	.w6(32'h3b37adce),
	.w7(32'hbb828d56),
	.w8(32'hbb67c8d8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f07c2),
	.w1(32'h3ae74375),
	.w2(32'h3b85c351),
	.w3(32'hbb083bfd),
	.w4(32'h3938e272),
	.w5(32'h3b4b3313),
	.w6(32'hbbdc4313),
	.w7(32'hbba9555d),
	.w8(32'h3b627851),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fc700),
	.w1(32'hbb2f6bc6),
	.w2(32'h3c20cff1),
	.w3(32'h399e017f),
	.w4(32'hbba693bd),
	.w5(32'hbaac5b49),
	.w6(32'h3b01ed80),
	.w7(32'hbaff33a8),
	.w8(32'hbc253095),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc48670),
	.w1(32'h3c82b72c),
	.w2(32'h3bde835e),
	.w3(32'h3c2eae68),
	.w4(32'h3c39ff5d),
	.w5(32'h3b80e1e6),
	.w6(32'hbd1fc769),
	.w7(32'hbca9ea42),
	.w8(32'h3b0d4205),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fa633),
	.w1(32'h3bfa868d),
	.w2(32'h3aab072a),
	.w3(32'hbc59cbda),
	.w4(32'h3b51dace),
	.w5(32'h3a4972a5),
	.w6(32'hbc36d0a8),
	.w7(32'hbc2c2a01),
	.w8(32'hbb65cf55),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c17004),
	.w1(32'hbadae9df),
	.w2(32'h3a1a998f),
	.w3(32'hb89f3c73),
	.w4(32'hbadaa5e8),
	.w5(32'h3c505806),
	.w6(32'hb9e2d9f7),
	.w7(32'hbab80b28),
	.w8(32'h3b5ca1dd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2421df),
	.w1(32'hbc044042),
	.w2(32'hbae5a98c),
	.w3(32'h3b500508),
	.w4(32'h3af80fb8),
	.w5(32'h3be2d39e),
	.w6(32'hbb3e8966),
	.w7(32'hb9c57e16),
	.w8(32'hbb6820bf),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89840d),
	.w1(32'hba0314f6),
	.w2(32'hb8cb046d),
	.w3(32'hbb5fd19a),
	.w4(32'h3b4ba687),
	.w5(32'h3c57f03c),
	.w6(32'hbb9923fe),
	.w7(32'hbb1519a7),
	.w8(32'hbc010a44),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f233c),
	.w1(32'hbca39801),
	.w2(32'hb9d5e5eb),
	.w3(32'h3cc494b4),
	.w4(32'h3ca197aa),
	.w5(32'hbc5aeb93),
	.w6(32'hbbd56647),
	.w7(32'h3c926eb5),
	.w8(32'h3c9ae5b6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36c570),
	.w1(32'h3c2a8f63),
	.w2(32'hbb1d3090),
	.w3(32'hbcef0bae),
	.w4(32'hbcd7f7ed),
	.w5(32'hbb2ded91),
	.w6(32'h3cca56b9),
	.w7(32'h3b9a2f10),
	.w8(32'h3ac7f475),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ac763),
	.w1(32'hbbaa3e8f),
	.w2(32'hbb9ea33a),
	.w3(32'hba0e11d6),
	.w4(32'hbb0c7cc9),
	.w5(32'hbbae6690),
	.w6(32'hba012d91),
	.w7(32'hbb4ce9bd),
	.w8(32'hbb057cb1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14a19e),
	.w1(32'hbba3e2d0),
	.w2(32'hbb852bf5),
	.w3(32'hbb312d40),
	.w4(32'hb9854bed),
	.w5(32'hbb37987c),
	.w6(32'hbb92bc75),
	.w7(32'h3a629770),
	.w8(32'h3be390d5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c038354),
	.w1(32'h3c3c8bf3),
	.w2(32'hba8bf5a5),
	.w3(32'hbc6c0ea2),
	.w4(32'hbc07a1c4),
	.w5(32'hbc8795ed),
	.w6(32'hbbfb6542),
	.w7(32'hbcb2dc35),
	.w8(32'h3c308a3d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f995c),
	.w1(32'h3b1010d7),
	.w2(32'hbb352b79),
	.w3(32'hbca3a8a3),
	.w4(32'hbc8cd61b),
	.w5(32'h3c11caae),
	.w6(32'hbbe92507),
	.w7(32'hbc9476cd),
	.w8(32'h3ba73c36),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8d492),
	.w1(32'hbc1315ae),
	.w2(32'h3a82caaa),
	.w3(32'h3c1f62ae),
	.w4(32'hbb8685c6),
	.w5(32'h3b187b8a),
	.w6(32'h3be7c6aa),
	.w7(32'h3c2483cf),
	.w8(32'h38b5a78e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036f58),
	.w1(32'hba03faa2),
	.w2(32'hbb8702b9),
	.w3(32'hbba6478f),
	.w4(32'h3a65ed27),
	.w5(32'hbae7889a),
	.w6(32'hbc22c8e1),
	.w7(32'h3a4efd14),
	.w8(32'hbbd55e71),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b03c0),
	.w1(32'hbac76089),
	.w2(32'hbb0c978e),
	.w3(32'hbacbc0dc),
	.w4(32'h3b906c33),
	.w5(32'h37a273de),
	.w6(32'hbc6174df),
	.w7(32'hbb9537bc),
	.w8(32'h3a2ef79a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de6b16),
	.w1(32'h3a1d56ff),
	.w2(32'h3b0c3a8a),
	.w3(32'h3aa22b6d),
	.w4(32'h3a83f34c),
	.w5(32'h3b38ea76),
	.w6(32'hbaa1b3aa),
	.w7(32'hba1c8323),
	.w8(32'h39d1a531),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a023f1),
	.w1(32'hbc559ffb),
	.w2(32'h3b0c5636),
	.w3(32'h3caa6f68),
	.w4(32'h3c697c98),
	.w5(32'h3af6b397),
	.w6(32'hbc2cc873),
	.w7(32'hbb9a90d2),
	.w8(32'h3b0a6a80),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d3b1f),
	.w1(32'hbb7f5dea),
	.w2(32'hbbf17fbb),
	.w3(32'h3ba9cd48),
	.w4(32'h3ad5085f),
	.w5(32'h3bdc43b0),
	.w6(32'hbbec3e74),
	.w7(32'hbb8355ee),
	.w8(32'h3b806d7d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd075378),
	.w1(32'hbd22b336),
	.w2(32'h3bab7b18),
	.w3(32'h3bf17931),
	.w4(32'hbbecd6c8),
	.w5(32'h3c18c960),
	.w6(32'h3c5b14f5),
	.w7(32'h3cc1507a),
	.w8(32'hbcb00e1d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc26c2),
	.w1(32'h3ab9801e),
	.w2(32'hbb2b1a48),
	.w3(32'h3c688561),
	.w4(32'hbaeacc95),
	.w5(32'hbbad55ed),
	.w6(32'hbc111cc8),
	.w7(32'hbb841fca),
	.w8(32'hbbdef025),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92ad6a),
	.w1(32'hba4b58f4),
	.w2(32'h3acedffe),
	.w3(32'h39b7ceae),
	.w4(32'h3a9b4077),
	.w5(32'h3943f906),
	.w6(32'hbb33e3df),
	.w7(32'hbb96af1c),
	.w8(32'hbaac9655),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc9acb),
	.w1(32'hba1c0c99),
	.w2(32'h39e615cc),
	.w3(32'h39dc7275),
	.w4(32'hba96e051),
	.w5(32'hbc6d7a95),
	.w6(32'hbb0948e4),
	.w7(32'hbb70569b),
	.w8(32'hbcd0748e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f0376),
	.w1(32'h3c9491e4),
	.w2(32'h3b74ac77),
	.w3(32'hbb9beafd),
	.w4(32'h3a9509b9),
	.w5(32'h3ae5f965),
	.w6(32'hbd17483b),
	.w7(32'hbcac9088),
	.w8(32'hbc1d3bed),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf48ee),
	.w1(32'h3bc0c793),
	.w2(32'hbbbcd96c),
	.w3(32'h3be87ee5),
	.w4(32'h3c716b44),
	.w5(32'hbc077e1a),
	.w6(32'hbc48a568),
	.w7(32'hbc18ffb7),
	.w8(32'h398d9995),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb186b1e),
	.w1(32'hbb61e952),
	.w2(32'h3bb883a1),
	.w3(32'hbb9cccee),
	.w4(32'h3750a3c2),
	.w5(32'h3bceec0b),
	.w6(32'h3b827e87),
	.w7(32'h398a28ff),
	.w8(32'h3c3f0ec1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11044d),
	.w1(32'hbb9a87d7),
	.w2(32'hbb2177d3),
	.w3(32'hbb432988),
	.w4(32'hbbcb2165),
	.w5(32'hbb8080f9),
	.w6(32'h3c4cd7ff),
	.w7(32'h3bd6211a),
	.w8(32'hbbd42893),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16dc7c),
	.w1(32'hbb042a35),
	.w2(32'h3974e0d9),
	.w3(32'hbae50a2a),
	.w4(32'hbae69bae),
	.w5(32'h38610d11),
	.w6(32'hbbc9b29b),
	.w7(32'hbacd413f),
	.w8(32'hb90f9ce4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d17435),
	.w1(32'h3b357826),
	.w2(32'h3c011b29),
	.w3(32'h3a6c26e7),
	.w4(32'h3a9030c7),
	.w5(32'hbb2259e5),
	.w6(32'hbb4858d3),
	.w7(32'hba2413a6),
	.w8(32'h3b177b1f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf657df),
	.w1(32'h3bd80466),
	.w2(32'hbc4450e9),
	.w3(32'hbc0b1675),
	.w4(32'h3bf70be5),
	.w5(32'h3c04350c),
	.w6(32'hbc3091a0),
	.w7(32'hbbbe26cd),
	.w8(32'h3c5a9a67),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82fcf3),
	.w1(32'hbc32763d),
	.w2(32'hbb8323a2),
	.w3(32'hbbd19ca2),
	.w4(32'hbc42e9a2),
	.w5(32'hbc10fa80),
	.w6(32'h3cfdbb17),
	.w7(32'h3c51c0c2),
	.w8(32'hb921a9f3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e609f),
	.w1(32'hbb51a167),
	.w2(32'hbc8755b7),
	.w3(32'hbbdcb081),
	.w4(32'h3ae4dead),
	.w5(32'h3b44aeeb),
	.w6(32'hbc49b1bc),
	.w7(32'hbafacc0f),
	.w8(32'h3b112432),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfd65cc),
	.w1(32'hbc5ab6e4),
	.w2(32'hbc2189f7),
	.w3(32'hbbb9e065),
	.w4(32'hbc02988b),
	.w5(32'hbc813f1a),
	.w6(32'h3c2a5623),
	.w7(32'h3b9c12dd),
	.w8(32'h3bbc6f5f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab15079),
	.w1(32'h3aa9a685),
	.w2(32'h3a95418f),
	.w3(32'hbc64c5f2),
	.w4(32'hbbc989ff),
	.w5(32'hbb7955b6),
	.w6(32'hbbd9fb5b),
	.w7(32'hbc580f58),
	.w8(32'hbac25632),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a434de4),
	.w1(32'h3b3ba7a2),
	.w2(32'h3b278440),
	.w3(32'hbb0a033d),
	.w4(32'h3b80f6d7),
	.w5(32'h3afecc21),
	.w6(32'hbbba366d),
	.w7(32'hb7b86a8d),
	.w8(32'hbc0efe0d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2cd24),
	.w1(32'h3b6ee32e),
	.w2(32'hbb38a6b0),
	.w3(32'hbb9eebfa),
	.w4(32'hbb8f3fe1),
	.w5(32'hb960c107),
	.w6(32'h3bd8a9d3),
	.w7(32'h3bf8f464),
	.w8(32'h3a19bc6f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9edcd),
	.w1(32'h3c11d124),
	.w2(32'hbb33d6b7),
	.w3(32'hbae4deb1),
	.w4(32'hbb592c83),
	.w5(32'hbb08aa80),
	.w6(32'hbb90d924),
	.w7(32'hbbe0e480),
	.w8(32'h3b94314f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb01bd6),
	.w1(32'h3b45f158),
	.w2(32'hbb488e63),
	.w3(32'h3c3bbb5c),
	.w4(32'h3c492027),
	.w5(32'h3adabac3),
	.w6(32'h3c416cd1),
	.w7(32'h3c45771b),
	.w8(32'h3b90a72d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6788d1),
	.w1(32'hbb1457f5),
	.w2(32'h3af26407),
	.w3(32'h3b7e5626),
	.w4(32'h3ba6e240),
	.w5(32'h3b5d243a),
	.w6(32'h3ac0ff3d),
	.w7(32'hbade6b19),
	.w8(32'hbcb1cbc5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19d4eb),
	.w1(32'h3bd41526),
	.w2(32'h3a01e04e),
	.w3(32'h3c87a51a),
	.w4(32'h3bc09deb),
	.w5(32'hb9df23f5),
	.w6(32'hbc3516aa),
	.w7(32'hbbd02758),
	.w8(32'hbbe8eb73),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabebbe5),
	.w1(32'hbb97b023),
	.w2(32'hb97f30c4),
	.w3(32'h3afc3f44),
	.w4(32'hba81f5a0),
	.w5(32'h3b0b3b5c),
	.w6(32'h3b039443),
	.w7(32'hb9e11f3d),
	.w8(32'hbc1d5f78),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb258b76),
	.w1(32'hbbaf2293),
	.w2(32'hbc0eac8f),
	.w3(32'hb935d7ab),
	.w4(32'hbb5bc043),
	.w5(32'hbb10ae5c),
	.w6(32'hbbee9f70),
	.w7(32'hbc119711),
	.w8(32'h3ad7208c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d0871),
	.w1(32'hbb0ee3f8),
	.w2(32'hbc72f2b5),
	.w3(32'hbbd60ae2),
	.w4(32'hbc103e6b),
	.w5(32'h3c341663),
	.w6(32'hbbc27e7b),
	.w7(32'hbaf6b363),
	.w8(32'hbae10bb3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd052df6),
	.w1(32'hbcd775c1),
	.w2(32'h3b121dab),
	.w3(32'h3bc086e9),
	.w4(32'hbc0a06f6),
	.w5(32'hbc04ddb6),
	.w6(32'h3c9d8b0a),
	.w7(32'h3c8ec67d),
	.w8(32'h3b6d25bb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b912fe0),
	.w1(32'h3bcb229f),
	.w2(32'hbc803605),
	.w3(32'hbbded56e),
	.w4(32'hbc0f53c7),
	.w5(32'h3bd5960d),
	.w6(32'h3b5d2c3e),
	.w7(32'hbc12ecb4),
	.w8(32'h3a84930d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93b32f),
	.w1(32'hbc0442a5),
	.w2(32'h3bc306eb),
	.w3(32'hbb3da10b),
	.w4(32'hbbc4032c),
	.w5(32'h3c1165e4),
	.w6(32'h3c4c4675),
	.w7(32'h39bee019),
	.w8(32'hbb685a0d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ef95e),
	.w1(32'h3a552d1e),
	.w2(32'h3af77b8f),
	.w3(32'h3c8e0ee1),
	.w4(32'h3c4bc191),
	.w5(32'h3b785ba2),
	.w6(32'hbbbe398b),
	.w7(32'h3bf17c6c),
	.w8(32'hbbcad661),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dce0f6),
	.w1(32'hbb892365),
	.w2(32'hbc557567),
	.w3(32'h3c628972),
	.w4(32'h3b93ab60),
	.w5(32'hbb881fca),
	.w6(32'hbc860786),
	.w7(32'hbc205e90),
	.w8(32'h3b130a23),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c84c),
	.w1(32'hbb71895f),
	.w2(32'h3bb38740),
	.w3(32'hbc9d13ef),
	.w4(32'hbc8eb391),
	.w5(32'hbb6f68d8),
	.w6(32'h3bc3f392),
	.w7(32'hbb4e0f3f),
	.w8(32'h3b4e5206),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b779ce6),
	.w1(32'h3b944610),
	.w2(32'h3b8ec6db),
	.w3(32'hbc18bad3),
	.w4(32'h3b426a7c),
	.w5(32'h3b5fbbe6),
	.w6(32'hbbaa18af),
	.w7(32'hbc7471b3),
	.w8(32'h3b236efa),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f16ea),
	.w1(32'hba8f48c7),
	.w2(32'h3bb734bc),
	.w3(32'hbaddb3b9),
	.w4(32'h3a9e0075),
	.w5(32'hbafc0b7f),
	.w6(32'hbb8a1109),
	.w7(32'hbbd9c040),
	.w8(32'hbbfef695),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba089fd),
	.w1(32'hba97106e),
	.w2(32'h3aba310e),
	.w3(32'hba84ae53),
	.w4(32'h3badb28a),
	.w5(32'h3a0db3c7),
	.w6(32'hbc5859c2),
	.w7(32'h3b0456e5),
	.w8(32'h3bd4070e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec4e92),
	.w1(32'h3af5ca67),
	.w2(32'hbbcd96b3),
	.w3(32'h3a717a76),
	.w4(32'h3a3cb97c),
	.w5(32'hbc75dd44),
	.w6(32'h3b5ff1d0),
	.w7(32'hba071b8a),
	.w8(32'hbaa15384),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f604),
	.w1(32'hbb5e1c14),
	.w2(32'hba358785),
	.w3(32'hbc588ebd),
	.w4(32'hbbc7d4ad),
	.w5(32'hbb467c39),
	.w6(32'hbb854562),
	.w7(32'hbc6eb039),
	.w8(32'hba4adbc3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ecd1c),
	.w1(32'h3bb987ab),
	.w2(32'hbbd4e0a1),
	.w3(32'hbc12c174),
	.w4(32'hbc2c5e9a),
	.w5(32'hbb885da9),
	.w6(32'h3b18733b),
	.w7(32'h3a5664e8),
	.w8(32'h3b8840c0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfba239),
	.w1(32'hbc049917),
	.w2(32'hb98d85cb),
	.w3(32'hbc006b85),
	.w4(32'hbb683417),
	.w5(32'h39e4b727),
	.w6(32'h3c4b4471),
	.w7(32'h3c1e8799),
	.w8(32'h3ae8487a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7eecf3),
	.w1(32'hb97f9a44),
	.w2(32'hbb047191),
	.w3(32'h3abf4941),
	.w4(32'h3a77807b),
	.w5(32'hbae0d6c7),
	.w6(32'h3a576d78),
	.w7(32'h3a458e42),
	.w8(32'hbb971e43),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ced11),
	.w1(32'hbb40a6e6),
	.w2(32'hbba07dba),
	.w3(32'h3a45e4c8),
	.w4(32'hba80718d),
	.w5(32'hb6ed6c74),
	.w6(32'hbb97703f),
	.w7(32'hbaff9c67),
	.w8(32'hbb9eaa69),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2c777),
	.w1(32'h3bafdf58),
	.w2(32'h3b5e3852),
	.w3(32'hbab45c59),
	.w4(32'h3c13a239),
	.w5(32'h3bc46aa1),
	.w6(32'hbc238618),
	.w7(32'hbc1cc5e7),
	.w8(32'h3be0bfc8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32d8ec),
	.w1(32'hbb25e5e8),
	.w2(32'hba8688c0),
	.w3(32'h3b53bbc3),
	.w4(32'hb9d01f2f),
	.w5(32'hbc03ff39),
	.w6(32'h3bdb7706),
	.w7(32'h3b04a054),
	.w8(32'hbc2f30f7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f5c6),
	.w1(32'h3b9f2bea),
	.w2(32'h3bdee48d),
	.w3(32'hbb3238b0),
	.w4(32'hbb0e581d),
	.w5(32'h3c1612f3),
	.w6(32'hbc82e484),
	.w7(32'hbbcfff49),
	.w8(32'hbcac7866),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25332f),
	.w1(32'h3c6bc0ca),
	.w2(32'h3be27557),
	.w3(32'h3cc01de5),
	.w4(32'h3ca262e1),
	.w5(32'h3c335ef6),
	.w6(32'hbcd61627),
	.w7(32'hbba82ffb),
	.w8(32'hbca27dde),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97db17),
	.w1(32'h3bd8790d),
	.w2(32'hbb2685f9),
	.w3(32'h3cf4bf4d),
	.w4(32'h3c9b8234),
	.w5(32'h3bf91432),
	.w6(32'hbcd50bc2),
	.w7(32'hbc18633a),
	.w8(32'hba6de48b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e3d81),
	.w1(32'h3b984273),
	.w2(32'h3b64c741),
	.w3(32'hbba57e8b),
	.w4(32'h3add5681),
	.w5(32'h3c47c9af),
	.w6(32'hbb0b9ecd),
	.w7(32'hbc02db9a),
	.w8(32'hbba9e322),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeefc80),
	.w1(32'hbc080605),
	.w2(32'hbb28c948),
	.w3(32'h3cabc780),
	.w4(32'h3c50926a),
	.w5(32'h3a831297),
	.w6(32'h3b55c2dc),
	.w7(32'h3b7914fc),
	.w8(32'h3c06b3e0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10d23c),
	.w1(32'hbb6e2126),
	.w2(32'hbb4c1462),
	.w3(32'hbc2d9994),
	.w4(32'hbb94070b),
	.w5(32'hbacbab26),
	.w6(32'hb9f69625),
	.w7(32'hbb3db74c),
	.w8(32'h3c09938b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52d079),
	.w1(32'hbb2ea961),
	.w2(32'hbc2f091e),
	.w3(32'hbbf59afe),
	.w4(32'hbc5cd026),
	.w5(32'hbc50d39c),
	.w6(32'h3ae99345),
	.w7(32'h3c3eedc8),
	.w8(32'h3c9fdfba),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc069fe9),
	.w1(32'hbb53060f),
	.w2(32'h3c116722),
	.w3(32'hbcbbba99),
	.w4(32'hbc10c32b),
	.w5(32'h3cea8364),
	.w6(32'h3c278d42),
	.w7(32'hbc03236a),
	.w8(32'hbc9be69c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55c714),
	.w1(32'hbb0bd980),
	.w2(32'h3a134212),
	.w3(32'h3cdb29ae),
	.w4(32'h385fbc45),
	.w5(32'hb977b342),
	.w6(32'h3b7d2adb),
	.w7(32'h3b4963af),
	.w8(32'h3b4cb0b4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bc0a1),
	.w1(32'h3ad8f50f),
	.w2(32'h3accb4a3),
	.w3(32'h3a32b61c),
	.w4(32'h3b36ba31),
	.w5(32'hbc328808),
	.w6(32'h3a89c3cd),
	.w7(32'h3b38efde),
	.w8(32'h3ba022fa),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11166d),
	.w1(32'h3b76d494),
	.w2(32'hbc067f10),
	.w3(32'hbc6b9aa3),
	.w4(32'hbb899e6b),
	.w5(32'h3b162f89),
	.w6(32'h3ab59e26),
	.w7(32'hbb24c8b1),
	.w8(32'h3a53367a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd89239),
	.w1(32'hba00fa0d),
	.w2(32'h3b3123a1),
	.w3(32'hbb98a9b8),
	.w4(32'h3b1f7a7a),
	.w5(32'h3bb65371),
	.w6(32'hbb2c3769),
	.w7(32'h3b97758a),
	.w8(32'h3be3a620),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2083f),
	.w1(32'hbb179edb),
	.w2(32'hbac1eb72),
	.w3(32'hbb95d6c3),
	.w4(32'hbb757029),
	.w5(32'hba91b16e),
	.w6(32'hbad4b931),
	.w7(32'hbae17af4),
	.w8(32'hbb4ae268),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff7229),
	.w1(32'hbaa97e62),
	.w2(32'h3b7543fe),
	.w3(32'hbb036bb0),
	.w4(32'h3a6cf7e6),
	.w5(32'hbc261fca),
	.w6(32'hbb7944bd),
	.w7(32'hbb0f16de),
	.w8(32'hbb292538),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0f0d0),
	.w1(32'h3aa1daca),
	.w2(32'hba9b30e8),
	.w3(32'hbc0fbfc1),
	.w4(32'hbb945c5c),
	.w5(32'hba719d95),
	.w6(32'h3bfe2e5d),
	.w7(32'h3c10edd2),
	.w8(32'h3b14ba7f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58a920),
	.w1(32'hbb40b81a),
	.w2(32'h3ac7b4cf),
	.w3(32'hbab71261),
	.w4(32'hbb8dbc2c),
	.w5(32'h3920d7c7),
	.w6(32'h3a6fc7d1),
	.w7(32'hb9a05b3a),
	.w8(32'h3ac92646),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ab247),
	.w1(32'h3b7d9bc3),
	.w2(32'hbb2fcba1),
	.w3(32'hbb531405),
	.w4(32'h3ac64b77),
	.w5(32'h3c900427),
	.w6(32'hba4dc273),
	.w7(32'h3b399815),
	.w8(32'h3c886cd9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01721b),
	.w1(32'h3afedac5),
	.w2(32'h39266171),
	.w3(32'h3c58f97e),
	.w4(32'hbb830b60),
	.w5(32'h3a531ba6),
	.w6(32'h3cd6dd54),
	.w7(32'h3c1e9bed),
	.w8(32'h3b814dfb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e48698),
	.w1(32'hbb841db7),
	.w2(32'hbb6a59b4),
	.w3(32'hbbdbecaf),
	.w4(32'hbb21cd4e),
	.w5(32'hba2be998),
	.w6(32'hbb55970b),
	.w7(32'h3a4cadc7),
	.w8(32'hbb5494fe),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed58a6),
	.w1(32'hba060082),
	.w2(32'hbbdbbe74),
	.w3(32'h3acfe679),
	.w4(32'h3b3df3e2),
	.w5(32'hbb76dbf5),
	.w6(32'hbaee4e0b),
	.w7(32'h3aa67597),
	.w8(32'h3bc9a6f2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cff75),
	.w1(32'hbbc64018),
	.w2(32'h3ae843f0),
	.w3(32'hbb4bad84),
	.w4(32'hbbc2db58),
	.w5(32'h3b2abb2f),
	.w6(32'h3bc85cf7),
	.w7(32'h3b30a18b),
	.w8(32'h3bdc61ec),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55243e),
	.w1(32'hbbd1980b),
	.w2(32'hbba33fd7),
	.w3(32'hbb4edc52),
	.w4(32'h3b5094a0),
	.w5(32'h3b0db47e),
	.w6(32'h3bdff109),
	.w7(32'hba126e92),
	.w8(32'hbb8b5599),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7277ed),
	.w1(32'hbc81be30),
	.w2(32'hbac5cfcf),
	.w3(32'h3b84366c),
	.w4(32'hba8ac14d),
	.w5(32'hbad7c7e1),
	.w6(32'h3bb1c94d),
	.w7(32'h3bdbbc8f),
	.w8(32'hba42ce67),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a5e6),
	.w1(32'hba8876ea),
	.w2(32'hbc5d1f2a),
	.w3(32'hba81e885),
	.w4(32'hbb541e9b),
	.w5(32'h3b4d4064),
	.w6(32'hb9dcae92),
	.w7(32'hbb78a4b1),
	.w8(32'h3c1b27bb),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05aa4d),
	.w1(32'hbc871325),
	.w2(32'h3b1b0eaa),
	.w3(32'hbb81d03a),
	.w4(32'hbc025651),
	.w5(32'h3b59f630),
	.w6(32'h3c6ce00b),
	.w7(32'h3c3bad7f),
	.w8(32'hbb658de1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b380a5b),
	.w1(32'h3be9b9b2),
	.w2(32'h3a8e438c),
	.w3(32'hbb5228de),
	.w4(32'hbb8654e0),
	.w5(32'h3abf01e4),
	.w6(32'hbb53599f),
	.w7(32'hbb3584ee),
	.w8(32'hba9acff3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ec92),
	.w1(32'hb94db4fc),
	.w2(32'h3ba0e2fd),
	.w3(32'hbadcfaa2),
	.w4(32'hbb86194c),
	.w5(32'hb9297d11),
	.w6(32'hbb96fa26),
	.w7(32'h3abe4b26),
	.w8(32'hb9a1e447),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15cebd),
	.w1(32'h3aa6404b),
	.w2(32'hbb86a4bd),
	.w3(32'hbbc69a34),
	.w4(32'h3bb8c9a5),
	.w5(32'h3c7d7169),
	.w6(32'hb991adea),
	.w7(32'hbc475bff),
	.w8(32'hbaa458ba),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e023f),
	.w1(32'hbc06936e),
	.w2(32'hbbdbcaa8),
	.w3(32'h3d10e7ae),
	.w4(32'h3c84131a),
	.w5(32'hbbf5db7a),
	.w6(32'h3c49613e),
	.w7(32'h3cb11d9f),
	.w8(32'h3bd7437d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfbb51),
	.w1(32'h3c28ec9c),
	.w2(32'hbb900224),
	.w3(32'hbccc962c),
	.w4(32'hbbe287ce),
	.w5(32'hbbf24579),
	.w6(32'hbbbcb2b7),
	.w7(32'hbc84de72),
	.w8(32'hbad797ad),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc351384),
	.w1(32'hbbdb1778),
	.w2(32'h3a73d94f),
	.w3(32'hbcd3cff4),
	.w4(32'hbc4de2ff),
	.w5(32'h3b2ee007),
	.w6(32'hbc19a7d3),
	.w7(32'hbb880bf6),
	.w8(32'h3c502ba5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88fd39),
	.w1(32'hb9bc4797),
	.w2(32'h3afe8658),
	.w3(32'h3ab82ae0),
	.w4(32'h3b3aea59),
	.w5(32'h3b3deecc),
	.w6(32'h3c21a17d),
	.w7(32'h3c1e5553),
	.w8(32'h3b6e0eed),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50d625),
	.w1(32'hbac52ba7),
	.w2(32'h3bb53383),
	.w3(32'h3b546a9a),
	.w4(32'h3b8740cc),
	.w5(32'hbba71713),
	.w6(32'h3b8b8c3a),
	.w7(32'hb9ee78c3),
	.w8(32'hbae611aa),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93b9b8),
	.w1(32'hb98dc7cf),
	.w2(32'hbaa3785e),
	.w3(32'hbcfd4326),
	.w4(32'hbcb7a986),
	.w5(32'h3a808e01),
	.w6(32'hbcf303ff),
	.w7(32'hbc8a5969),
	.w8(32'h3b299883),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaade57),
	.w1(32'h3aa1cac5),
	.w2(32'h3b0a646e),
	.w3(32'hb9ed69c6),
	.w4(32'hbb17120e),
	.w5(32'h3ba4bdf2),
	.w6(32'hb926e74a),
	.w7(32'hb9e33600),
	.w8(32'hba9e6dba),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e113e),
	.w1(32'h3acb663a),
	.w2(32'h3c96f03c),
	.w3(32'h3bf94fce),
	.w4(32'h3c0bf72f),
	.w5(32'h3acdba66),
	.w6(32'hbbb07ff1),
	.w7(32'hbbbf42ec),
	.w8(32'hbb99c494),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c946c75),
	.w1(32'h3c6d4565),
	.w2(32'h3ad7773a),
	.w3(32'hbb94f13c),
	.w4(32'hbb980fd4),
	.w5(32'h39f1c4a4),
	.w6(32'hbcba07e0),
	.w7(32'hbc85e06b),
	.w8(32'hba98e002),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd7905),
	.w1(32'hbb845ffe),
	.w2(32'h3aa7bb56),
	.w3(32'hbbab157e),
	.w4(32'hbb75ef15),
	.w5(32'h3c356c93),
	.w6(32'hbc2b3f8b),
	.w7(32'hbb6f01f2),
	.w8(32'h3bcc7bb2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c338afc),
	.w1(32'h3bc7cef8),
	.w2(32'h3bb92619),
	.w3(32'h3d059232),
	.w4(32'h3cbdf104),
	.w5(32'h379b537c),
	.w6(32'h3cd52604),
	.w7(32'h3c922a58),
	.w8(32'h3aaaed07),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933f23),
	.w1(32'h3b2dfbb4),
	.w2(32'h3c5e6067),
	.w3(32'hbb84da81),
	.w4(32'hbb1bda9b),
	.w5(32'h3c220d6a),
	.w6(32'hbb380a19),
	.w7(32'hbc5e2bac),
	.w8(32'hbb8e852c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2ea9c),
	.w1(32'h3ca1f254),
	.w2(32'h3b86af8d),
	.w3(32'h3c347b76),
	.w4(32'h3c23723c),
	.w5(32'h3bb8cbc6),
	.w6(32'hbc481abd),
	.w7(32'hbbc838ac),
	.w8(32'h3bf992fb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b084556),
	.w1(32'h37a412dd),
	.w2(32'h3b8b6ca2),
	.w3(32'hbb1c4278),
	.w4(32'h3a13f016),
	.w5(32'h3a8ef632),
	.w6(32'h3b9af5f4),
	.w7(32'h3adf2523),
	.w8(32'hbacb09d8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948b7e4),
	.w1(32'hbc074ddc),
	.w2(32'hbb2ada44),
	.w3(32'hbbc0f549),
	.w4(32'hbbe60b48),
	.w5(32'hbb9e2781),
	.w6(32'hbbcbfda2),
	.w7(32'hbc131db7),
	.w8(32'hb934b5f9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67d76f),
	.w1(32'hbb7d007d),
	.w2(32'h3bddd80f),
	.w3(32'hbc04bcb7),
	.w4(32'hbc226eb9),
	.w5(32'hb9fb51a3),
	.w6(32'hbc0e25be),
	.w7(32'hbbe4725e),
	.w8(32'hbbb5284f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ff0e2),
	.w1(32'h3b25dd55),
	.w2(32'hbacb600b),
	.w3(32'hb9ac7330),
	.w4(32'h3b117748),
	.w5(32'hba1e2345),
	.w6(32'hbb915b0f),
	.w7(32'hbb8b3a23),
	.w8(32'h3aaf1774),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedb287),
	.w1(32'hbb2688da),
	.w2(32'hbd000189),
	.w3(32'hbaa92eba),
	.w4(32'hbb07fd26),
	.w5(32'hbc99121c),
	.w6(32'hbac26450),
	.w7(32'h3a9cc19c),
	.w8(32'h3ba76651),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2998f6),
	.w1(32'hbd0946b6),
	.w2(32'h3afdbdb4),
	.w3(32'hbce6ba14),
	.w4(32'hbcacea65),
	.w5(32'hba08f44e),
	.w6(32'h3b9afeba),
	.w7(32'h3b7e27a4),
	.w8(32'h3b8339e0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a069c7e),
	.w1(32'hbc161fc1),
	.w2(32'h3b25953b),
	.w3(32'hbb072ca2),
	.w4(32'hbb24bbc6),
	.w5(32'hbb83e78b),
	.w6(32'hbb78340f),
	.w7(32'hbabf3fe3),
	.w8(32'hbb18ec3f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1182f4),
	.w1(32'hbb1d1084),
	.w2(32'h3aeae3b5),
	.w3(32'h3a53bfc4),
	.w4(32'h3ad61b9f),
	.w5(32'hba81f525),
	.w6(32'hba6bd980),
	.w7(32'h3bd1f272),
	.w8(32'hbb00a3ef),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393acc4e),
	.w1(32'h3abc70a4),
	.w2(32'hbae8950d),
	.w3(32'h3bb92741),
	.w4(32'h3adc1612),
	.w5(32'hbbd31f21),
	.w6(32'h3acc78bc),
	.w7(32'h3b1aa2cc),
	.w8(32'hbb55e208),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a83c4),
	.w1(32'h3ab9e45d),
	.w2(32'hbc0f23c9),
	.w3(32'hbc42eb09),
	.w4(32'hbaecd400),
	.w5(32'h3c40e1c8),
	.w6(32'hbc38039e),
	.w7(32'hbc051b38),
	.w8(32'h3b50af24),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba53c02),
	.w1(32'hba9fb177),
	.w2(32'h3bdbe58d),
	.w3(32'h3d2f14b6),
	.w4(32'h3cfb33a2),
	.w5(32'h3be275c9),
	.w6(32'h3d1a3ef0),
	.w7(32'h3cbe50cd),
	.w8(32'h3b21114b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba67119),
	.w1(32'h3acba722),
	.w2(32'h39e7f071),
	.w3(32'h3b1dc326),
	.w4(32'h3b8f660f),
	.w5(32'h3aba5fc0),
	.w6(32'h3b9c4a4c),
	.w7(32'h3bc1ab93),
	.w8(32'h3a054263),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba085feb),
	.w1(32'hbb1ca978),
	.w2(32'h3b83c5ec),
	.w3(32'h3a837bc4),
	.w4(32'hbb29e701),
	.w5(32'hbaae2c68),
	.w6(32'h3a2acf24),
	.w7(32'h39eeb351),
	.w8(32'h3a056c21),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2314),
	.w1(32'h39103dda),
	.w2(32'h3b1f8d2d),
	.w3(32'hbb3eaec5),
	.w4(32'hbb975c6e),
	.w5(32'h3aebbacc),
	.w6(32'hbb6aa902),
	.w7(32'hbbe5b8e5),
	.w8(32'h3b840132),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af750bc),
	.w1(32'h3b75c47b),
	.w2(32'h3bbaf253),
	.w3(32'h3aa93e3c),
	.w4(32'h3bce01f9),
	.w5(32'hbad32edd),
	.w6(32'h3bc814f9),
	.w7(32'h3b2f6e82),
	.w8(32'hbb2a99b9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9322da),
	.w1(32'h3b9a8371),
	.w2(32'h3c1ce3b0),
	.w3(32'hbb597561),
	.w4(32'hbb0f40e8),
	.w5(32'h3bb399df),
	.w6(32'hbb33f87e),
	.w7(32'hbb24d3aa),
	.w8(32'hb98e6369),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e8b3f),
	.w1(32'h3b60ea0a),
	.w2(32'h3b73f610),
	.w3(32'h3b462d04),
	.w4(32'hbb78810b),
	.w5(32'h3b734465),
	.w6(32'h3a801fa7),
	.w7(32'hbb0c1119),
	.w8(32'h3946475e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88f5af),
	.w1(32'h383294ff),
	.w2(32'h3ae207ef),
	.w3(32'hbb8d948e),
	.w4(32'hbb88156d),
	.w5(32'hba87db94),
	.w6(32'hbbca3c74),
	.w7(32'hbc016529),
	.w8(32'hbb969bc7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab72e5d),
	.w1(32'h3aa4378c),
	.w2(32'h3ad86641),
	.w3(32'hbb5d7902),
	.w4(32'h3bc81823),
	.w5(32'h3b55713d),
	.w6(32'hba4d64a2),
	.w7(32'hba0026de),
	.w8(32'h3ad278a5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73380b),
	.w1(32'h3b96227c),
	.w2(32'hbaa72cab),
	.w3(32'hbb7025d9),
	.w4(32'h3bbde08a),
	.w5(32'h3aa11995),
	.w6(32'hbb3a8087),
	.w7(32'h3b6fa2d8),
	.w8(32'h3c52c9a1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bf249),
	.w1(32'hbbeeed41),
	.w2(32'h3c177c64),
	.w3(32'hbbf5cb30),
	.w4(32'hbc90f02a),
	.w5(32'hba2e4134),
	.w6(32'hb9b6d11a),
	.w7(32'hbc88899a),
	.w8(32'h3a6344aa),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed2783),
	.w1(32'h3bcae0ff),
	.w2(32'h3bbac1fd),
	.w3(32'h3b39d362),
	.w4(32'h3aa41e34),
	.w5(32'h3bdb99b2),
	.w6(32'hb9364fc1),
	.w7(32'h3b22887e),
	.w8(32'h3b89d7aa),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc1888),
	.w1(32'hbb783318),
	.w2(32'h3afb03b8),
	.w3(32'h3bb7fe36),
	.w4(32'hba7f0b07),
	.w5(32'h3baabe7c),
	.w6(32'h3be076a9),
	.w7(32'h3bb79592),
	.w8(32'h3bb72b14),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb50207),
	.w1(32'hba10166f),
	.w2(32'h3a960493),
	.w3(32'h3a5f742c),
	.w4(32'h39ec5a94),
	.w5(32'h3b93e287),
	.w6(32'hbb2f972c),
	.w7(32'hb9b53531),
	.w8(32'h3b867d7a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b657e1e),
	.w1(32'h3bf3e3f1),
	.w2(32'h3a529120),
	.w3(32'hbb33e4da),
	.w4(32'h3ab299b8),
	.w5(32'h3b1f3bff),
	.w6(32'h3b5a8309),
	.w7(32'h3b3ae5db),
	.w8(32'h3b208bb5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b896bac),
	.w1(32'h3a7c4675),
	.w2(32'h3aa63e34),
	.w3(32'h3b8e26a1),
	.w4(32'h3b3c5414),
	.w5(32'hbb6e5d8f),
	.w6(32'h3b2fb8aa),
	.w7(32'hbad4157b),
	.w8(32'h3b3ccbe2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ff12b),
	.w1(32'hbb0e26d6),
	.w2(32'hb729fef7),
	.w3(32'hb9620827),
	.w4(32'h39e49a73),
	.w5(32'hbb9260b3),
	.w6(32'hb9e9c8c0),
	.w7(32'h3aefe65f),
	.w8(32'hbb628814),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a959e8),
	.w1(32'hba1e127f),
	.w2(32'hbcd16378),
	.w3(32'hbb1c47ca),
	.w4(32'hb9b1377c),
	.w5(32'hbd06f002),
	.w6(32'hbbbaff27),
	.w7(32'hbb104034),
	.w8(32'hbb3eb992),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4c9579),
	.w1(32'hbd0b6127),
	.w2(32'h3994d93d),
	.w3(32'hbd9807f6),
	.w4(32'hbd4b2f49),
	.w5(32'h3aad0cb1),
	.w6(32'hbd0c7b87),
	.w7(32'hbc97ca64),
	.w8(32'h3b76e8ce),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bea6b),
	.w1(32'hbb3e825c),
	.w2(32'h3af0f41a),
	.w3(32'hbbb668a3),
	.w4(32'hb997679a),
	.w5(32'h3b95eb29),
	.w6(32'hbb2ce324),
	.w7(32'h3a9a1339),
	.w8(32'h3b15cfc1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b304fc8),
	.w1(32'h3a2e9422),
	.w2(32'h3a3990f3),
	.w3(32'h3aa197f8),
	.w4(32'h3a6023a4),
	.w5(32'hbb3e9a8a),
	.w6(32'hb805167a),
	.w7(32'hbac9729a),
	.w8(32'hbb326e24),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05010d),
	.w1(32'h39c798de),
	.w2(32'h3bd9d1ad),
	.w3(32'hbb9b442d),
	.w4(32'hbba50446),
	.w5(32'h3bf51151),
	.w6(32'hbba5febe),
	.w7(32'hbb477117),
	.w8(32'hb9f95ad2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be87155),
	.w1(32'hbab5f95e),
	.w2(32'h3b0f78c7),
	.w3(32'h3bc3074c),
	.w4(32'h3a58b536),
	.w5(32'h3a6371f0),
	.w6(32'h3b117a2f),
	.w7(32'hbb22c78c),
	.w8(32'h3b27c435),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53a585),
	.w1(32'h3b076aa2),
	.w2(32'h3b12bf8c),
	.w3(32'hb8e7e7bf),
	.w4(32'h3b5b9b1b),
	.w5(32'h3abea224),
	.w6(32'hbb26b15f),
	.w7(32'h3a8372c0),
	.w8(32'h3a37d566),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd18211),
	.w1(32'hba9874e4),
	.w2(32'h3b96a169),
	.w3(32'hbc0503c3),
	.w4(32'hba174980),
	.w5(32'h3b5961bf),
	.w6(32'hbb13a997),
	.w7(32'h3a87bbf0),
	.w8(32'hb9788a01),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb831b5f),
	.w1(32'hbae0d0af),
	.w2(32'hbc871a4d),
	.w3(32'hbb20d595),
	.w4(32'hbb295ee0),
	.w5(32'hb9c62c50),
	.w6(32'hbbb25e09),
	.w7(32'h3af19b03),
	.w8(32'h3b547399),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32164b),
	.w1(32'hbc44559c),
	.w2(32'hbb0dccf4),
	.w3(32'h3c4ee440),
	.w4(32'h3c103015),
	.w5(32'hbbca0a72),
	.w6(32'h3c9efbd6),
	.w7(32'h3c6ed1d2),
	.w8(32'hbb79be3e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba965b0),
	.w1(32'hbb182a97),
	.w2(32'h39ddd7fb),
	.w3(32'hbb9ed3f7),
	.w4(32'hbb849eaf),
	.w5(32'h3befaa62),
	.w6(32'hbb815f0d),
	.w7(32'hbb6dea89),
	.w8(32'h3ac1be4c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b032553),
	.w1(32'h3ae0b210),
	.w2(32'h3bc2e51b),
	.w3(32'h3ae5f866),
	.w4(32'h3b514a08),
	.w5(32'h3a85dff2),
	.w6(32'h3c0d43cf),
	.w7(32'h3b8a22da),
	.w8(32'h3ae534f1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1d889),
	.w1(32'h3a682a8c),
	.w2(32'hba8996fc),
	.w3(32'hbb37368d),
	.w4(32'hbb280d8e),
	.w5(32'hb9ab64f9),
	.w6(32'h3a752942),
	.w7(32'hb76e8a2e),
	.w8(32'h3abfc20d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac366e7),
	.w1(32'hb86e9d3c),
	.w2(32'hbba7422f),
	.w3(32'hbbe8e838),
	.w4(32'hbb7b2370),
	.w5(32'hbbf7680a),
	.w6(32'hbc13c52e),
	.w7(32'h3a7adc4d),
	.w8(32'hba263972),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71f2e),
	.w1(32'hbbf58024),
	.w2(32'h3a12a334),
	.w3(32'hbce9d4ac),
	.w4(32'hbc899089),
	.w5(32'hbb805209),
	.w6(32'hbc3d0a7a),
	.w7(32'hbbac127a),
	.w8(32'hbacd3b3e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e274c),
	.w1(32'h3ad3c91e),
	.w2(32'hbcda273f),
	.w3(32'hbae8fd1f),
	.w4(32'hbb191ddb),
	.w5(32'hbd1a2ebe),
	.w6(32'hbb9eccb0),
	.w7(32'hbab8bb2a),
	.w8(32'hbc575d16),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6cc05b),
	.w1(32'hbd274865),
	.w2(32'h3a1cc7a5),
	.w3(32'hbdc50704),
	.w4(32'hbd8bf13b),
	.w5(32'hbb2fbaf0),
	.w6(32'hbd78953a),
	.w7(32'hbd0ec75b),
	.w8(32'h3b30f965),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05f781),
	.w1(32'h3b05db54),
	.w2(32'h3b66eba7),
	.w3(32'hbaa22139),
	.w4(32'h3978f8d5),
	.w5(32'h3b99e162),
	.w6(32'hb80f9aa3),
	.w7(32'h3a48e0af),
	.w8(32'h3b11249b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcac1ee),
	.w1(32'h39bc9133),
	.w2(32'hbac5a818),
	.w3(32'h3b14e27c),
	.w4(32'hbb46335b),
	.w5(32'h3b172f50),
	.w6(32'hbaf40e0c),
	.w7(32'hbbc92a5f),
	.w8(32'hb9a8e9a2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a036ae),
	.w1(32'h3a9b6379),
	.w2(32'h3a39e5d2),
	.w3(32'hbb4b06c6),
	.w4(32'h3ab3594b),
	.w5(32'hbb90b623),
	.w6(32'hbb43c474),
	.w7(32'h3b1df0e2),
	.w8(32'hbadd1099),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb943cff),
	.w1(32'h3be8ec37),
	.w2(32'hbb8c09b8),
	.w3(32'hbc3a870c),
	.w4(32'h3bb0ce22),
	.w5(32'hbbe549c6),
	.w6(32'hbad4a0dd),
	.w7(32'h3b63aa33),
	.w8(32'hbb987713),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ee7c8),
	.w1(32'h3aa8d657),
	.w2(32'hbbd48c2a),
	.w3(32'hbba0196c),
	.w4(32'hbac75af5),
	.w5(32'hbc5df5fc),
	.w6(32'hbc0a62bd),
	.w7(32'hbb5c015c),
	.w8(32'hbaa7ad36),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9250b5),
	.w1(32'hbc58249c),
	.w2(32'h3b0649a6),
	.w3(32'hbcb2914d),
	.w4(32'hbc7f64c2),
	.w5(32'h3b8884e4),
	.w6(32'hbc085efd),
	.w7(32'hbae46972),
	.w8(32'h3a88ff1b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d62f4),
	.w1(32'h3a4d2ff7),
	.w2(32'h3bc35318),
	.w3(32'hbac9e9c9),
	.w4(32'h3b7bec32),
	.w5(32'h3b827ac8),
	.w6(32'hbabd3b1f),
	.w7(32'h3ae62e4a),
	.w8(32'h3b08ea83),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d3936),
	.w1(32'h3b177c6e),
	.w2(32'h3bf00001),
	.w3(32'hbb85a9d6),
	.w4(32'hbb8a34fd),
	.w5(32'h3b8c86cc),
	.w6(32'hbb9aab1a),
	.w7(32'hbb2f6c10),
	.w8(32'hbb9fee12),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b912c3b),
	.w1(32'hb721ca68),
	.w2(32'h3ba0465f),
	.w3(32'hba26cd90),
	.w4(32'hbab67561),
	.w5(32'h3c764eb7),
	.w6(32'hbbcb88ae),
	.w7(32'hbb30dcf1),
	.w8(32'h3beb70e5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec3218),
	.w1(32'h3b09492b),
	.w2(32'h3ac1bc8f),
	.w3(32'h3c998884),
	.w4(32'h3bdbeefa),
	.w5(32'hbb6f3a8a),
	.w6(32'h3c26c6ac),
	.w7(32'h3ac33cdf),
	.w8(32'hbaf84090),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e9a1c),
	.w1(32'h3b821f38),
	.w2(32'hbccbb18c),
	.w3(32'hbb301934),
	.w4(32'hbb3a9654),
	.w5(32'hbcb8982f),
	.w6(32'h3a9cf88d),
	.w7(32'h3b2d22b8),
	.w8(32'h3a9a9925),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2da373),
	.w1(32'hbcf951db),
	.w2(32'h3b36cecf),
	.w3(32'hbd510299),
	.w4(32'hbd10e794),
	.w5(32'h3b0e96af),
	.w6(32'hbc73b82b),
	.w7(32'hbbbd4746),
	.w8(32'h3b8a1143),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a445c0c),
	.w1(32'hbb382488),
	.w2(32'h3b43010d),
	.w3(32'h3af2c314),
	.w4(32'hbac45b02),
	.w5(32'hbb3b2250),
	.w6(32'h3b8590a6),
	.w7(32'h3b54f968),
	.w8(32'hba9ccb72),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b902fb5),
	.w1(32'hbaf4602d),
	.w2(32'h3b876449),
	.w3(32'hbb34a13c),
	.w4(32'h3911c152),
	.w5(32'hba88ebb4),
	.w6(32'hbb0c5569),
	.w7(32'hba12d009),
	.w8(32'h3b67a2e9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95bcee),
	.w1(32'hba4721a5),
	.w2(32'h3b846296),
	.w3(32'hbbc77d5a),
	.w4(32'hbbc4694d),
	.w5(32'h3af2c3f5),
	.w6(32'hba8f53fc),
	.w7(32'hba25be40),
	.w8(32'hbb3e58d7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac3787),
	.w1(32'hbac33779),
	.w2(32'h38c9fc81),
	.w3(32'h3a6f462b),
	.w4(32'h3b0186b6),
	.w5(32'hb9a8fe76),
	.w6(32'hbb8939dd),
	.w7(32'hbb2abec2),
	.w8(32'h3b2dc91a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8429dd),
	.w1(32'h3ab9ddd4),
	.w2(32'h3b30723e),
	.w3(32'hbb6766a9),
	.w4(32'h3b8c0fc0),
	.w5(32'h3a85f013),
	.w6(32'hbab96bf3),
	.w7(32'hbb38f4c3),
	.w8(32'h3b6d56b4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa61461),
	.w1(32'h3ab84bed),
	.w2(32'hbb72477b),
	.w3(32'hbb76c529),
	.w4(32'hbb97aea6),
	.w5(32'hbabff984),
	.w6(32'hbb5e419c),
	.w7(32'hb9b694d0),
	.w8(32'h3ac803cc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5ad18),
	.w1(32'h3900a749),
	.w2(32'h3a5b49b3),
	.w3(32'hbbe5ab53),
	.w4(32'h39386bb1),
	.w5(32'hbb023d48),
	.w6(32'h3ab7bbb5),
	.w7(32'h3b1bd70d),
	.w8(32'h38949a3d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82eba2),
	.w1(32'hba0d72e6),
	.w2(32'h393751d0),
	.w3(32'hb9a4c963),
	.w4(32'hb9a45ab2),
	.w5(32'hbb736b43),
	.w6(32'hbb143ad4),
	.w7(32'h38f5ff22),
	.w8(32'hbb2465de),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9542b),
	.w1(32'h3b91be20),
	.w2(32'h3bed00e9),
	.w3(32'h393209d9),
	.w4(32'h3b4a20ee),
	.w5(32'hba0f93cd),
	.w6(32'hbb80f440),
	.w7(32'hba5b7b98),
	.w8(32'hbb9fc89a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932c8f),
	.w1(32'h3ba63ca6),
	.w2(32'h3b88f512),
	.w3(32'hbb24e8d0),
	.w4(32'hbaa0fe71),
	.w5(32'hbaf05244),
	.w6(32'hbbf6d68b),
	.w7(32'hbb9475c5),
	.w8(32'hbaa2ab79),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b610a13),
	.w1(32'hba4524a5),
	.w2(32'h3a9c57cd),
	.w3(32'h3ae9ce85),
	.w4(32'h39ba82dc),
	.w5(32'hbaf7a415),
	.w6(32'h3b496163),
	.w7(32'h3a8b7046),
	.w8(32'hbb1a3513),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca3c33),
	.w1(32'h3bd30782),
	.w2(32'hb8e6e36f),
	.w3(32'hb9da615d),
	.w4(32'h3aa8321e),
	.w5(32'hbb9489ed),
	.w6(32'hbb7dd5f6),
	.w7(32'h399c8e9a),
	.w8(32'hbb5171ca),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8211aa),
	.w1(32'h3ba79042),
	.w2(32'hba43cfa3),
	.w3(32'hbb6c5b01),
	.w4(32'h3b51cd9c),
	.w5(32'hbc013bb4),
	.w6(32'hbbd75cce),
	.w7(32'h3a3c1d12),
	.w8(32'hbb1f60f4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19e91c),
	.w1(32'h3aba5061),
	.w2(32'h3b4b670f),
	.w3(32'hbb4963ec),
	.w4(32'hbb9d6121),
	.w5(32'h3b146dc8),
	.w6(32'hbb132e05),
	.w7(32'hbb0f9c89),
	.w8(32'h3b4360a1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10263f),
	.w1(32'h3b034be6),
	.w2(32'hb907129a),
	.w3(32'h3bb559a5),
	.w4(32'h3bd784b4),
	.w5(32'h3b28a7d2),
	.w6(32'h3a8ed5fe),
	.w7(32'hba731589),
	.w8(32'hbbbf2509),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ad2b5),
	.w1(32'hba94d290),
	.w2(32'hbb85192b),
	.w3(32'hba20a32f),
	.w4(32'h3b54e64e),
	.w5(32'hbacc856c),
	.w6(32'hbbb07223),
	.w7(32'hbba30a35),
	.w8(32'hba92ec95),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4eb847),
	.w1(32'hb9d186f3),
	.w2(32'h3b16c216),
	.w3(32'hbbaaedd9),
	.w4(32'hbad615bd),
	.w5(32'hbab4605e),
	.w6(32'h3a6ce0be),
	.w7(32'hbb722cd7),
	.w8(32'h39946db4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42ff06),
	.w1(32'hb91ec3ec),
	.w2(32'h3bc36db8),
	.w3(32'hba94af2e),
	.w4(32'h390fcd69),
	.w5(32'hb9405ad4),
	.w6(32'h3b3078f4),
	.w7(32'h3b4a572f),
	.w8(32'h3b8e42ed),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e868c),
	.w1(32'h3b7108fe),
	.w2(32'h3ba14cc2),
	.w3(32'hbb85ddad),
	.w4(32'hbb93bb60),
	.w5(32'hbad089a7),
	.w6(32'hbbd7e1cf),
	.w7(32'hbb6991bb),
	.w8(32'h3a972da3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fb1f3),
	.w1(32'hbbaeb009),
	.w2(32'h3b227da5),
	.w3(32'h3ab51fb2),
	.w4(32'hbb5940d6),
	.w5(32'h3bb1ee93),
	.w6(32'hba900c45),
	.w7(32'hbb3f9da4),
	.w8(32'h3b9068c2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03f06d),
	.w1(32'h3b1b654c),
	.w2(32'hbb1f2b42),
	.w3(32'h3a1f23da),
	.w4(32'hbb23b02e),
	.w5(32'hb9584bb6),
	.w6(32'hbb079e30),
	.w7(32'hbb8904e2),
	.w8(32'h3c05e270),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa95460),
	.w1(32'hb9adf5b1),
	.w2(32'h3b5170b8),
	.w3(32'h3a2fca1d),
	.w4(32'hb9078f69),
	.w5(32'h3b536217),
	.w6(32'h3c02c314),
	.w7(32'h3bbd3bf3),
	.w8(32'hba2f4f39),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a220969),
	.w1(32'hbaad79cd),
	.w2(32'hba482850),
	.w3(32'hbb793cfc),
	.w4(32'hbb319991),
	.w5(32'hbaf4282a),
	.w6(32'hbbd159b0),
	.w7(32'hbbe1f836),
	.w8(32'h3bc897ae),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3dbc40),
	.w1(32'h3b227024),
	.w2(32'h38a2f621),
	.w3(32'hbb3bd24b),
	.w4(32'hb938cd59),
	.w5(32'h39bc68f3),
	.w6(32'h3ba07ac7),
	.w7(32'h3b41b444),
	.w8(32'hba94c53d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45f94f),
	.w1(32'hb9b4eb14),
	.w2(32'h399e6bf2),
	.w3(32'hbb04912c),
	.w4(32'hba24d37f),
	.w5(32'h3a0bcbaa),
	.w6(32'hbb77ba92),
	.w7(32'hbac98ae6),
	.w8(32'h3b5f85d4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b142a13),
	.w1(32'h3ab3f490),
	.w2(32'hb93bbff6),
	.w3(32'h3a8c279a),
	.w4(32'h3a4539f4),
	.w5(32'h3b664407),
	.w6(32'h3bcf5a65),
	.w7(32'h3ba985a2),
	.w8(32'h38b089cb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3348e5),
	.w1(32'h3ac3a3b0),
	.w2(32'h3b879f3f),
	.w3(32'h3b892ac1),
	.w4(32'h3a90efd1),
	.w5(32'h3bdd90a9),
	.w6(32'h3b9508fe),
	.w7(32'h3b2faa73),
	.w8(32'hb9825823),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c142887),
	.w1(32'h3c106659),
	.w2(32'h3bb516a4),
	.w3(32'h3c8341e4),
	.w4(32'h3c650351),
	.w5(32'h3adb2425),
	.w6(32'h3c0ef6ad),
	.w7(32'h3be4d785),
	.w8(32'hbb12b6b8),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94651f),
	.w1(32'h3bca0018),
	.w2(32'h39a502d6),
	.w3(32'hbb7caf2c),
	.w4(32'hbadf1503),
	.w5(32'hbaf531c6),
	.w6(32'hbc05280b),
	.w7(32'hbb62713a),
	.w8(32'hb9b5040f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c0fbc),
	.w1(32'hbb0bad06),
	.w2(32'hbaf6a47e),
	.w3(32'hbbee20e1),
	.w4(32'hbc085e72),
	.w5(32'hba9c5219),
	.w6(32'hbb37d820),
	.w7(32'hbb58df63),
	.w8(32'h3a37e234),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac44e6),
	.w1(32'h398524be),
	.w2(32'h3b907726),
	.w3(32'h398a5002),
	.w4(32'h3b5a5e9e),
	.w5(32'h3b14c64b),
	.w6(32'h3b12bae6),
	.w7(32'h3b3c4a24),
	.w8(32'h3b616c28),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4bde7),
	.w1(32'h3b62a646),
	.w2(32'h3b99c04e),
	.w3(32'h3b81f854),
	.w4(32'hba96cff5),
	.w5(32'h3ac5f827),
	.w6(32'h3b608243),
	.w7(32'h3b8d66f2),
	.w8(32'h3bd1c4c0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbada140),
	.w1(32'hb9e98f4a),
	.w2(32'hbb854006),
	.w3(32'hbba6a659),
	.w4(32'hba8fd959),
	.w5(32'hbb757d19),
	.w6(32'hba9f4697),
	.w7(32'hbb1ef7b8),
	.w8(32'h39ceb1db),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b3393),
	.w1(32'h3b16c64a),
	.w2(32'h3aa478c4),
	.w3(32'hbb3e34b1),
	.w4(32'h3ae8b4bb),
	.w5(32'hbb39407c),
	.w6(32'hbb801f95),
	.w7(32'h3a5c2e86),
	.w8(32'h3acb11fc),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule