module layer_8_featuremap_231(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c3ce2),
	.w1(32'h3c5f10b0),
	.w2(32'h3c9494f9),
	.w3(32'h3bcf4afc),
	.w4(32'hbb751785),
	.w5(32'h3c49d73c),
	.w6(32'h3b30bd06),
	.w7(32'h3c2616d1),
	.w8(32'h3bae0df2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ac18),
	.w1(32'hbc05caf9),
	.w2(32'hbc3c0bf3),
	.w3(32'h3bbc590f),
	.w4(32'hbc2a5834),
	.w5(32'hbc4a1e51),
	.w6(32'hbc2e6d60),
	.w7(32'hbc3789ab),
	.w8(32'hbc330fb5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ab44),
	.w1(32'hbc44dc65),
	.w2(32'hbcd7d2d7),
	.w3(32'hbc0bed59),
	.w4(32'hbc356583),
	.w5(32'hbc8f0125),
	.w6(32'hbc866c25),
	.w7(32'hbc397f8a),
	.w8(32'hbc2860ff),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1c153),
	.w1(32'h3b1ebef5),
	.w2(32'hbb57a45c),
	.w3(32'hbcd107ab),
	.w4(32'hbbb839e3),
	.w5(32'hba94a516),
	.w6(32'hbb773244),
	.w7(32'h38a406e6),
	.w8(32'h3b7a8cd3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386c06e7),
	.w1(32'h3bbc4558),
	.w2(32'h3c621033),
	.w3(32'hbb3845aa),
	.w4(32'h3b3cf51a),
	.w5(32'h3c44576d),
	.w6(32'h3a1b68db),
	.w7(32'h3bad3a51),
	.w8(32'h3a0eb498),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5df8ec),
	.w1(32'h3ca39340),
	.w2(32'h3c4b70be),
	.w3(32'h3c6eb480),
	.w4(32'h3c584e9e),
	.w5(32'h3bb7b65e),
	.w6(32'h3cb177fd),
	.w7(32'h3cabd8da),
	.w8(32'h3c4b5e19),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1154c1),
	.w1(32'h3c28c6c1),
	.w2(32'h3c937725),
	.w3(32'h3bcfa326),
	.w4(32'h3c120b65),
	.w5(32'h3c8256fe),
	.w6(32'hba073ae4),
	.w7(32'h3c0b6907),
	.w8(32'h3bfb0105),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c951c68),
	.w1(32'h3be29d28),
	.w2(32'h3c14bf1a),
	.w3(32'h3c31ff0d),
	.w4(32'hbc3b428c),
	.w5(32'hbc81847a),
	.w6(32'hbb9b3144),
	.w7(32'h3c2b50be),
	.w8(32'h3c26b3be),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b5155),
	.w1(32'hbb6e447d),
	.w2(32'hbbdbcad2),
	.w3(32'hbc2dbc53),
	.w4(32'hbaf84288),
	.w5(32'hbb7e34bc),
	.w6(32'hbc056d84),
	.w7(32'hbc4b591d),
	.w8(32'hbc12611e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2b001),
	.w1(32'hbba15ae1),
	.w2(32'h3bea0dfa),
	.w3(32'hbb4886c2),
	.w4(32'hbb235113),
	.w5(32'h3c1ab3c3),
	.w6(32'hbb77880f),
	.w7(32'h3b9a2bfd),
	.w8(32'h3bc51c77),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92122d),
	.w1(32'h3c11aa30),
	.w2(32'h3c03d27e),
	.w3(32'h3b53681a),
	.w4(32'h3ba9eca9),
	.w5(32'h3cae7e3c),
	.w6(32'h3af31dd3),
	.w7(32'h3a163551),
	.w8(32'hb8dcbd0c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a8b65),
	.w1(32'h3c1ee7f9),
	.w2(32'h3cc5c698),
	.w3(32'h3c12f5ac),
	.w4(32'h3bded5cf),
	.w5(32'h3c24be9d),
	.w6(32'h3c0416d1),
	.w7(32'h3c412bd0),
	.w8(32'h385078d3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14072d),
	.w1(32'h3af40455),
	.w2(32'hba948e5a),
	.w3(32'h3b277d4a),
	.w4(32'h3a575d08),
	.w5(32'hb93efcc6),
	.w6(32'hbb381204),
	.w7(32'h3999ef8d),
	.w8(32'hbafec79a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf21c8),
	.w1(32'hbc0406ba),
	.w2(32'hbcda014c),
	.w3(32'hbb8afc61),
	.w4(32'hbc23b519),
	.w5(32'hbc4eda8d),
	.w6(32'hbc805f90),
	.w7(32'hbc772932),
	.w8(32'hbbbfee31),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5cdfe),
	.w1(32'h3bc7b9a4),
	.w2(32'h3bc0f111),
	.w3(32'hbc9713a7),
	.w4(32'h3be2589b),
	.w5(32'h3ba28759),
	.w6(32'h3b1c730f),
	.w7(32'h3a5d746c),
	.w8(32'h3bca9a59),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed2f41),
	.w1(32'h3c06111f),
	.w2(32'hbbd3d7a7),
	.w3(32'h3b97c3c1),
	.w4(32'h3c0b819e),
	.w5(32'hbacf7af4),
	.w6(32'h3c05228b),
	.w7(32'hbc83f952),
	.w8(32'hbc5e7781),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97a51b),
	.w1(32'h3c899478),
	.w2(32'h3c3c7752),
	.w3(32'h3bfb5a87),
	.w4(32'h3cbdfc29),
	.w5(32'h3cb75d65),
	.w6(32'h3c144da2),
	.w7(32'h3b579573),
	.w8(32'h3c4f9944),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c574477),
	.w1(32'hbce1b555),
	.w2(32'hbd0a2eb3),
	.w3(32'h3a439c95),
	.w4(32'hbc71b47b),
	.w5(32'hbd03dcad),
	.w6(32'hbc8ce44a),
	.w7(32'hbcb473f7),
	.w8(32'hbc701307),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5ca46),
	.w1(32'hba57fae4),
	.w2(32'h3c30b1d5),
	.w3(32'hbd0f2580),
	.w4(32'hbc0493ef),
	.w5(32'hbaf749ed),
	.w6(32'h3bfc4fbe),
	.w7(32'h3b8f0e1b),
	.w8(32'h3c34feaa),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15fcd1),
	.w1(32'hbc24e1f0),
	.w2(32'hbc5b2cd8),
	.w3(32'h3b0b0612),
	.w4(32'hbb4710c5),
	.w5(32'hbc1f3dee),
	.w6(32'hbb8ed574),
	.w7(32'hbbdc0a66),
	.w8(32'hba8d79b9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf165d),
	.w1(32'hbc60257e),
	.w2(32'hbca90278),
	.w3(32'hba94ceee),
	.w4(32'hbbcb15c8),
	.w5(32'hbc50b78d),
	.w6(32'hbbc30728),
	.w7(32'hbc581594),
	.w8(32'hbc389570),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc592baf),
	.w1(32'hbbb75263),
	.w2(32'hbc96bc6f),
	.w3(32'hbbe26cb6),
	.w4(32'hb94b5b67),
	.w5(32'hbc44efb7),
	.w6(32'hbb8dd79a),
	.w7(32'hbc19ee28),
	.w8(32'hbb9655fc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e8365),
	.w1(32'h3a3ea6d5),
	.w2(32'h3c8667fc),
	.w3(32'hbc8d5e37),
	.w4(32'hbc3bb36c),
	.w5(32'h3c0ee676),
	.w6(32'h3b28f700),
	.w7(32'h3c15afb9),
	.w8(32'h3c72f792),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c058f46),
	.w1(32'hbb8d38a2),
	.w2(32'hbc968e8e),
	.w3(32'h3bfd350f),
	.w4(32'hbc000571),
	.w5(32'hbc176642),
	.w6(32'hbae97ee1),
	.w7(32'hbc2e0735),
	.w8(32'hbc3ec7b6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67fef0),
	.w1(32'h3bde1fb7),
	.w2(32'h3c359b7c),
	.w3(32'hbc31c200),
	.w4(32'h3b0590f0),
	.w5(32'h3ba4dd1d),
	.w6(32'h3bbefb80),
	.w7(32'h3c431367),
	.w8(32'h3bdadb39),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c397d13),
	.w1(32'h3c848c26),
	.w2(32'h3c5c762d),
	.w3(32'h3a964d2e),
	.w4(32'h3b5dfcde),
	.w5(32'h3b8137cf),
	.w6(32'h3c7e7b46),
	.w7(32'h3c40157e),
	.w8(32'hbbc3307b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86d28c),
	.w1(32'h3ba900b0),
	.w2(32'h3c4ece82),
	.w3(32'h3b8e5d6d),
	.w4(32'h39aa4035),
	.w5(32'h3ac3ba67),
	.w6(32'h3bdbf536),
	.w7(32'h3c0a61ae),
	.w8(32'h3c6173c3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b330481),
	.w1(32'hbc0ab582),
	.w2(32'hbbd2b95b),
	.w3(32'hba0d5b16),
	.w4(32'hbce3f372),
	.w5(32'hbcda0c69),
	.w6(32'hbc7cbd49),
	.w7(32'hbbc6010d),
	.w8(32'hbc8ad6b9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd72ac),
	.w1(32'h38bab758),
	.w2(32'h3b81d8c2),
	.w3(32'hbc274cbd),
	.w4(32'hbbd1743d),
	.w5(32'hba38001b),
	.w6(32'h3a61093d),
	.w7(32'h3aa59160),
	.w8(32'h3b84dda7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03e2a0),
	.w1(32'h3c23ec2b),
	.w2(32'h3c6610bb),
	.w3(32'h3bc801c4),
	.w4(32'h3c778774),
	.w5(32'h3c9be4f0),
	.w6(32'h3bdfaac0),
	.w7(32'h3c3a0b39),
	.w8(32'h3c1ae9e2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c250cd6),
	.w1(32'h3c268980),
	.w2(32'h3be2dcd0),
	.w3(32'h3c7f86f9),
	.w4(32'h3b93e0ec),
	.w5(32'h3c23e804),
	.w6(32'h3b65e2a7),
	.w7(32'h3aac26dc),
	.w8(32'hbb74c6ce),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb51551),
	.w1(32'hba03317b),
	.w2(32'hbb97cb89),
	.w3(32'h3bd9915e),
	.w4(32'h3bbdac9c),
	.w5(32'hbb09edd7),
	.w6(32'hbb8037e4),
	.w7(32'hbb9c0a96),
	.w8(32'hbc252c66),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58bb81),
	.w1(32'hbc8c26b7),
	.w2(32'hbd1a438c),
	.w3(32'hbb0e68e4),
	.w4(32'hbb99c5be),
	.w5(32'hbcbd9555),
	.w6(32'hbc313d3b),
	.w7(32'hbcbe098a),
	.w8(32'hbc7fc6ed),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb7cf3),
	.w1(32'h3d1cea27),
	.w2(32'h3d8678a0),
	.w3(32'hbcc67970),
	.w4(32'h3cd819e8),
	.w5(32'h3d527216),
	.w6(32'h3cbe5394),
	.w7(32'h3d2e4c47),
	.w8(32'h3c99d5db),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d449a6d),
	.w1(32'h3b9b17ec),
	.w2(32'hbc20f096),
	.w3(32'h3d2d1aec),
	.w4(32'hbb6b9341),
	.w5(32'hbc84ef10),
	.w6(32'h3618bffe),
	.w7(32'hbb8c566b),
	.w8(32'hbb8f982c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1c072),
	.w1(32'h3c65c93e),
	.w2(32'h3cc8bf88),
	.w3(32'hbc938dc6),
	.w4(32'h3a6f7228),
	.w5(32'h3c136b53),
	.w6(32'hba84503f),
	.w7(32'h3c07d1ff),
	.w8(32'h3c21595e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50f08d),
	.w1(32'h3a3f903a),
	.w2(32'hbbbedea7),
	.w3(32'h3bda637c),
	.w4(32'h3ac359ef),
	.w5(32'hbb287c36),
	.w6(32'h396b8852),
	.w7(32'hbbbe658e),
	.w8(32'hbb748252),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42efe3),
	.w1(32'hb8c5589d),
	.w2(32'hbbca6775),
	.w3(32'hba3f166d),
	.w4(32'h3a99d379),
	.w5(32'hbb46b6d6),
	.w6(32'hbaa09856),
	.w7(32'hbc246a36),
	.w8(32'hbae4ab4d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90cfda),
	.w1(32'hbc000de9),
	.w2(32'hbb7ccd6f),
	.w3(32'hbb41a934),
	.w4(32'hbc0ea6d8),
	.w5(32'hbb6f58b9),
	.w6(32'hbc5fc1c4),
	.w7(32'hbc027aa5),
	.w8(32'hbc0f6326),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb35052),
	.w1(32'h3c94e416),
	.w2(32'h3cbea779),
	.w3(32'hbc28cdc8),
	.w4(32'h3c935774),
	.w5(32'h3cbc1b5e),
	.w6(32'h3c30d85b),
	.w7(32'h3ca639e2),
	.w8(32'h3c5cb433),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3554e2),
	.w1(32'hbc97f033),
	.w2(32'hbd0b0b1c),
	.w3(32'h3bcb29f0),
	.w4(32'hbcb981f9),
	.w5(32'hbd188950),
	.w6(32'hbc63de43),
	.w7(32'hbcc66e0a),
	.w8(32'hbc8b760a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc8398),
	.w1(32'h3c75fcc1),
	.w2(32'h3bfbbcf6),
	.w3(32'hbcc4cdb0),
	.w4(32'h3c3106a9),
	.w5(32'h3befa77b),
	.w6(32'h3b0f409f),
	.w7(32'h3a329189),
	.w8(32'hbc55c459),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdcd4d),
	.w1(32'h3b82e034),
	.w2(32'h3c12ba1b),
	.w3(32'hbba36305),
	.w4(32'hba22ab94),
	.w5(32'h3c086a17),
	.w6(32'h3bc192a1),
	.w7(32'h3c21dab3),
	.w8(32'h3ba20b27),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0599f2),
	.w1(32'h3a8847b0),
	.w2(32'h3c7da90c),
	.w3(32'h3bb80e49),
	.w4(32'hbbbfc68d),
	.w5(32'h3a91fe14),
	.w6(32'hba61dc7f),
	.w7(32'hb97f2b5c),
	.w8(32'hba48e521),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbac0a),
	.w1(32'hbc8436ef),
	.w2(32'hbd3384f9),
	.w3(32'hbb966164),
	.w4(32'hbc79213b),
	.w5(32'hbcfe150d),
	.w6(32'hbc102722),
	.w7(32'hbcaf725f),
	.w8(32'hbc27162f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd120cd4),
	.w1(32'hbbcbbb37),
	.w2(32'hbb480586),
	.w3(32'hbd057c98),
	.w4(32'hbb6941dd),
	.w5(32'hbab5df34),
	.w6(32'hbc0a86cd),
	.w7(32'hbb68c248),
	.w8(32'h3bdb727f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfab5b2),
	.w1(32'h3d131b16),
	.w2(32'h3d70af75),
	.w3(32'h3c0b73e9),
	.w4(32'h3cc4a0a5),
	.w5(32'h3d4201e1),
	.w6(32'h3c98c16e),
	.w7(32'h3d04ef16),
	.w8(32'h3cc18026),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3da56e),
	.w1(32'hbc4b93f0),
	.w2(32'hbc830f57),
	.w3(32'h3d0b2803),
	.w4(32'hbc51ae52),
	.w5(32'hbc7279f4),
	.w6(32'hb7c92373),
	.w7(32'hbb803105),
	.w8(32'h3a962c27),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc161c83),
	.w1(32'hbc18b258),
	.w2(32'hbcc33ada),
	.w3(32'hbc383e34),
	.w4(32'hbc3e0a6a),
	.w5(32'hbca152ab),
	.w6(32'hbb44e87b),
	.w7(32'hbb8e8b57),
	.w8(32'h3a9b8fb2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc955eaf),
	.w1(32'hbc234365),
	.w2(32'hbbde09d6),
	.w3(32'hbc8dd498),
	.w4(32'hbb67bcdd),
	.w5(32'hbc1308b9),
	.w6(32'hbb1b06fe),
	.w7(32'hbb9d2496),
	.w8(32'hbc45180e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf7b44),
	.w1(32'h3b16e038),
	.w2(32'h3983c3e4),
	.w3(32'hbbc98be3),
	.w4(32'h3ba90fd4),
	.w5(32'h3b3d0c41),
	.w6(32'h3b9e0250),
	.w7(32'h3bc03d52),
	.w8(32'h3b17d7d5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f6700),
	.w1(32'h3c3fb25e),
	.w2(32'h3b752695),
	.w3(32'hbc116845),
	.w4(32'hbbd4a5ae),
	.w5(32'hbbc69ff4),
	.w6(32'hbbcad551),
	.w7(32'hbc2b31bc),
	.w8(32'h3ba52c5d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae201b),
	.w1(32'h3c02aa24),
	.w2(32'h3c028236),
	.w3(32'h3bb2d2cb),
	.w4(32'h3b5f33a1),
	.w5(32'h3be39984),
	.w6(32'h3b05018d),
	.w7(32'h39c6914a),
	.w8(32'h3bdee3fd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be78264),
	.w1(32'h3aa15d29),
	.w2(32'h3a780cf2),
	.w3(32'h3c0e89cf),
	.w4(32'hbb2b8559),
	.w5(32'hbacf6e45),
	.w6(32'h39cafe7f),
	.w7(32'h3bf4e675),
	.w8(32'h3c509a77),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04448b),
	.w1(32'hbbaa7fed),
	.w2(32'hbb2acd70),
	.w3(32'h3bf13a5b),
	.w4(32'hbaaec333),
	.w5(32'hbbf6e18d),
	.w6(32'hbbd750fd),
	.w7(32'hbb5aae3b),
	.w8(32'h3af0eb18),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52c205),
	.w1(32'hbbc9d34e),
	.w2(32'h3bc162c9),
	.w3(32'hbc15e768),
	.w4(32'hbc9c75e9),
	.w5(32'hbb77fd2a),
	.w6(32'hbc09cbe8),
	.w7(32'hbb7b10a1),
	.w8(32'hbb559f8b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54383),
	.w1(32'h3c0bc9f5),
	.w2(32'h3c39bfb7),
	.w3(32'hbb505907),
	.w4(32'h3ba7dfe6),
	.w5(32'h3c06175c),
	.w6(32'h3bea402d),
	.w7(32'h3c2cbe92),
	.w8(32'h3c0e4d87),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f308f),
	.w1(32'h3b688012),
	.w2(32'h3c81c608),
	.w3(32'hbb8c46cc),
	.w4(32'hbb71f030),
	.w5(32'h3c0276a5),
	.w6(32'hbb8468b6),
	.w7(32'h3b4dd2a0),
	.w8(32'h3b9c5b93),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfde5ae),
	.w1(32'hb9de5bdf),
	.w2(32'h3b24db00),
	.w3(32'h3bc5bac5),
	.w4(32'hbbace94d),
	.w5(32'hba9a9eeb),
	.w6(32'hba5db158),
	.w7(32'hbb8417de),
	.w8(32'hbb21338a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4de93a),
	.w1(32'hbbb847cb),
	.w2(32'hbcb30184),
	.w3(32'hbb0d20c5),
	.w4(32'hbbdc4d7c),
	.w5(32'hbc9b7920),
	.w6(32'hbc69fdeb),
	.w7(32'hbc829ce5),
	.w8(32'hbbb50232),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69eb46),
	.w1(32'h3b36e805),
	.w2(32'h3bbdd103),
	.w3(32'hbbb60414),
	.w4(32'hbb9a8251),
	.w5(32'h3b93d29f),
	.w6(32'hbb8c0342),
	.w7(32'h3b5e51c9),
	.w8(32'h3a9347f9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ef5aa),
	.w1(32'h3c6d3a4c),
	.w2(32'h3c81ea10),
	.w3(32'h39441d55),
	.w4(32'h3c4f379b),
	.w5(32'h3c5d1e49),
	.w6(32'hbc00b12f),
	.w7(32'hbbd6675b),
	.w8(32'hbb391344),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2be06e),
	.w1(32'hba9ca19b),
	.w2(32'h39993489),
	.w3(32'h3b9431fb),
	.w4(32'h3b1f0de1),
	.w5(32'h3b859b45),
	.w6(32'h3b01312e),
	.w7(32'h3aeec6dd),
	.w8(32'h3a97e19c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3521ba),
	.w1(32'h3c16e1c7),
	.w2(32'h3c131568),
	.w3(32'h3be091cf),
	.w4(32'h3c02ea21),
	.w5(32'h3c0c5d16),
	.w6(32'h3c183e57),
	.w7(32'h3c2a906f),
	.w8(32'h3c13b16a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19b0a9),
	.w1(32'hb95866f2),
	.w2(32'hbaf3a2c8),
	.w3(32'h3c00f1c4),
	.w4(32'hbabb49c0),
	.w5(32'hbac7fe7a),
	.w6(32'hb9da5c17),
	.w7(32'hbac6a679),
	.w8(32'hbb39ce9d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6654db),
	.w1(32'h3c60476b),
	.w2(32'h3cb1d09b),
	.w3(32'hbba099d8),
	.w4(32'h3c2d7772),
	.w5(32'h3ca31002),
	.w6(32'h3bedbf2d),
	.w7(32'h3c4de805),
	.w8(32'h3c133948),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb04056),
	.w1(32'h3c078946),
	.w2(32'h3be8ec9f),
	.w3(32'h3c4d3260),
	.w4(32'h3c12501f),
	.w5(32'h3bcb23ae),
	.w6(32'h3a68ff70),
	.w7(32'h3909a64c),
	.w8(32'h3bc5c29e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04bebb),
	.w1(32'h3c553fb0),
	.w2(32'h3d09b518),
	.w3(32'h3b34065b),
	.w4(32'h3b592f9d),
	.w5(32'h3c953b93),
	.w6(32'h3b737ba2),
	.w7(32'h3c382c90),
	.w8(32'h3b303052),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90dee8),
	.w1(32'hbc52ddbc),
	.w2(32'hbbe0520b),
	.w3(32'h3c159209),
	.w4(32'hbc2c75a7),
	.w5(32'hbc6c5220),
	.w6(32'hbc719778),
	.w7(32'hbc4cb4ce),
	.w8(32'hbc0ce57a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01eecf),
	.w1(32'hbcb1db4d),
	.w2(32'hbceacb01),
	.w3(32'hbc8e4255),
	.w4(32'hbc24caa3),
	.w5(32'hbce44a3f),
	.w6(32'hbb98c28a),
	.w7(32'hbc55fe60),
	.w8(32'hbc2599bc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc817eb5),
	.w1(32'hba8b40dc),
	.w2(32'h3c137288),
	.w3(32'hbc83cf57),
	.w4(32'hbb1697dd),
	.w5(32'h3bcfa7ce),
	.w6(32'hbbbf6498),
	.w7(32'h3b90df3d),
	.w8(32'h3ba0a105),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d06fd),
	.w1(32'h3c6525cc),
	.w2(32'h3cc6cf17),
	.w3(32'h3c3d7574),
	.w4(32'h3c51c42d),
	.w5(32'h3c21ef77),
	.w6(32'h3b98ce87),
	.w7(32'h3c4de5ac),
	.w8(32'h3ba53890),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e7d28),
	.w1(32'h3c3ead89),
	.w2(32'h3c6afc7c),
	.w3(32'h3b780095),
	.w4(32'h3c2408fe),
	.w5(32'h3c59331e),
	.w6(32'h3b79ab53),
	.w7(32'h3c51d4b6),
	.w8(32'h3c2d93c8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c9f1b),
	.w1(32'hbbdfc64b),
	.w2(32'h3a56ab66),
	.w3(32'h3aa9b01e),
	.w4(32'hbadb4c9f),
	.w5(32'h3c1074ec),
	.w6(32'hbbe0e93b),
	.w7(32'h3b92ef65),
	.w8(32'h3bb20fe2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba918312),
	.w1(32'h3bff9329),
	.w2(32'h3c40b2df),
	.w3(32'h3b6c3067),
	.w4(32'hbada134c),
	.w5(32'h3ab1471d),
	.w6(32'hbb0aa85e),
	.w7(32'h3c09fd7e),
	.w8(32'h3b8104c0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be51188),
	.w1(32'hbc894429),
	.w2(32'hbcd5c413),
	.w3(32'hbb95ed00),
	.w4(32'hbc4a9513),
	.w5(32'hbcc5fbb9),
	.w6(32'hbc3d45ef),
	.w7(32'hbc9bc01f),
	.w8(32'hbc033cc6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99b82e),
	.w1(32'h3b45f44b),
	.w2(32'h3bb374df),
	.w3(32'hbc911a8a),
	.w4(32'hb90bdbcd),
	.w5(32'h3b7bd356),
	.w6(32'hba34ca97),
	.w7(32'h3b1802a0),
	.w8(32'h3ba6b2a8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe4f83),
	.w1(32'hb9bd31ce),
	.w2(32'h3b98759c),
	.w3(32'hb9ae7069),
	.w4(32'hbc00353d),
	.w5(32'hba8255aa),
	.w6(32'h36073660),
	.w7(32'hbac6cd4a),
	.w8(32'h3bb9b280),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f6944),
	.w1(32'hbb3bdf18),
	.w2(32'h3bf3558b),
	.w3(32'h3b8bf6f7),
	.w4(32'hbb7bb20e),
	.w5(32'h3bd0ea3f),
	.w6(32'hba5fdf34),
	.w7(32'h3a35a9c4),
	.w8(32'h37af9206),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa300b2),
	.w1(32'h3b9c8ff3),
	.w2(32'h3bd9c8dd),
	.w3(32'h3bfa05d9),
	.w4(32'hbb58c470),
	.w5(32'h3a84ca86),
	.w6(32'hbb46b94c),
	.w7(32'hba62541a),
	.w8(32'hbb2c428e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62ef0f),
	.w1(32'hbc6ffe49),
	.w2(32'hbcc55a9a),
	.w3(32'hbb8ae14a),
	.w4(32'hbc2482cb),
	.w5(32'hbc8e383b),
	.w6(32'hbc5fcc6a),
	.w7(32'hbc9036db),
	.w8(32'hbc6df19f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84d6eb),
	.w1(32'hbc8b192e),
	.w2(32'hbbbcdb5c),
	.w3(32'hbcb1dc19),
	.w4(32'hbc24090a),
	.w5(32'hbc78a6a9),
	.w6(32'hbc483943),
	.w7(32'hbc0a37c3),
	.w8(32'hbc6aac25),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55ba6c),
	.w1(32'hbc8170bd),
	.w2(32'hbd0e9dfc),
	.w3(32'hbc9f137a),
	.w4(32'hbcb01b93),
	.w5(32'hbd027539),
	.w6(32'hbc662305),
	.w7(32'hbca00aab),
	.w8(32'hbc4a6386),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7b03d),
	.w1(32'h3c428723),
	.w2(32'h3c9703c9),
	.w3(32'hbcfbeffb),
	.w4(32'h3c2e9b25),
	.w5(32'h3c446ecd),
	.w6(32'h3c50edd5),
	.w7(32'h3cbb89cc),
	.w8(32'h3c985e5b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdec9ac),
	.w1(32'hbcb52a21),
	.w2(32'hbd070d88),
	.w3(32'hbbe5ccff),
	.w4(32'hbcd98869),
	.w5(32'hbd11bb65),
	.w6(32'hbc9aa166),
	.w7(32'hbcc7b312),
	.w8(32'hbc30d801),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee0693),
	.w1(32'h3c5c6b34),
	.w2(32'h3c38421a),
	.w3(32'hbce736c5),
	.w4(32'h3be92629),
	.w5(32'h3c212b8b),
	.w6(32'h3c69fcb0),
	.w7(32'h3ba82457),
	.w8(32'h3c0749f0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c190292),
	.w1(32'hba0aac43),
	.w2(32'h3b200cbb),
	.w3(32'h3bbc67dd),
	.w4(32'hbb70e66d),
	.w5(32'h39399685),
	.w6(32'h3b3c14c7),
	.w7(32'h3ab69c9a),
	.w8(32'h3ae8c065),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdc9b1),
	.w1(32'h3bade579),
	.w2(32'h3b85547e),
	.w3(32'h3af02682),
	.w4(32'h3b907619),
	.w5(32'h3b4e9557),
	.w6(32'h3b136ad5),
	.w7(32'h3ba62ccf),
	.w8(32'h3ba78704),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a067762),
	.w1(32'h3b7b0dd6),
	.w2(32'h3bebdbc5),
	.w3(32'hba7577fb),
	.w4(32'h3b7acc17),
	.w5(32'h3bb279c3),
	.w6(32'h3ae81d04),
	.w7(32'h3ae82fed),
	.w8(32'h3ab4adf5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99d897),
	.w1(32'hbc63db2f),
	.w2(32'hbca2b0ef),
	.w3(32'h3b578867),
	.w4(32'hbbee80a7),
	.w5(32'hbc66c07f),
	.w6(32'hbbba670c),
	.w7(32'hbbbc6bfe),
	.w8(32'hbbf16be7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f7a3c),
	.w1(32'h3cafdc0c),
	.w2(32'h3d04ad74),
	.w3(32'hbc5ee7b5),
	.w4(32'h3c89901f),
	.w5(32'h3ca6eab1),
	.w6(32'h3c44514c),
	.w7(32'h3c8bddf5),
	.w8(32'h3c75d3bf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd25d24),
	.w1(32'h3d1b9861),
	.w2(32'h3d9c0e2d),
	.w3(32'h3c5d7a70),
	.w4(32'h3c6b4444),
	.w5(32'h3d5687c6),
	.w6(32'h3c8ded54),
	.w7(32'h3ce06f85),
	.w8(32'h3c8859a5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d49380c),
	.w1(32'hb8fb7b07),
	.w2(32'hba526fca),
	.w3(32'h3d23910c),
	.w4(32'h3b2287d8),
	.w5(32'h3a5e4a58),
	.w6(32'hba85d959),
	.w7(32'h39b2248f),
	.w8(32'h39d1bd7a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab955c4),
	.w1(32'h3ad7f3d2),
	.w2(32'h3bae418a),
	.w3(32'h3aab2194),
	.w4(32'hbb828592),
	.w5(32'hb95b58d4),
	.w6(32'hbb46fdf7),
	.w7(32'h3a68b450),
	.w8(32'h3987a682),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5e264),
	.w1(32'h3c97fcd5),
	.w2(32'h3ca49cc9),
	.w3(32'h3b88943c),
	.w4(32'h3c74d398),
	.w5(32'h3c2f6f71),
	.w6(32'h3ca022ab),
	.w7(32'h3c0215c6),
	.w8(32'h3a657327),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f802d),
	.w1(32'h3ac32ff3),
	.w2(32'hb989b80a),
	.w3(32'h3bdb52cb),
	.w4(32'h376a17c1),
	.w5(32'hbab4c51b),
	.w6(32'h3ab40631),
	.w7(32'hbab68496),
	.w8(32'h3b0ec17d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b105c60),
	.w1(32'hbc23e6c7),
	.w2(32'hbcac1cbd),
	.w3(32'hbb83d2f8),
	.w4(32'hbc279a69),
	.w5(32'hbc1c3e67),
	.w6(32'hbc194058),
	.w7(32'hbbeb2df0),
	.w8(32'hbad09394),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50dc1c),
	.w1(32'hbc36031b),
	.w2(32'hbc99ae77),
	.w3(32'hbc0cda29),
	.w4(32'hbc2607ca),
	.w5(32'hbc9a3289),
	.w6(32'hbc31b3ea),
	.w7(32'hbc88b30b),
	.w8(32'hbbb0f0f2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5de867),
	.w1(32'hbb86f637),
	.w2(32'h3bbc552e),
	.w3(32'hbc91a9b5),
	.w4(32'hbbcdc91c),
	.w5(32'h3a13fbe9),
	.w6(32'hbc4e39fc),
	.w7(32'h3b3e0927),
	.w8(32'h3978532b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b957ed1),
	.w1(32'h3bbdf402),
	.w2(32'h3c142d8d),
	.w3(32'h3ae41ffb),
	.w4(32'hba91f68f),
	.w5(32'h3bf95831),
	.w6(32'hbabea8ad),
	.w7(32'h3bd856d8),
	.w8(32'h3a24f360),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b6e78),
	.w1(32'h3bcce091),
	.w2(32'h3b42e82f),
	.w3(32'hbb9a94a1),
	.w4(32'h3bb688e2),
	.w5(32'h3b6f985a),
	.w6(32'h3bae5a37),
	.w7(32'h3c95b43d),
	.w8(32'h3cc8ec49),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c719e),
	.w1(32'hbae6faca),
	.w2(32'hbbd1e21b),
	.w3(32'h3c09368f),
	.w4(32'h3c304faa),
	.w5(32'h3c10499f),
	.w6(32'h3be703fe),
	.w7(32'h3b4013e1),
	.w8(32'h3b439ee3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea84d6),
	.w1(32'h3c06019e),
	.w2(32'h3cc42933),
	.w3(32'h3b963639),
	.w4(32'h3bf7c5f4),
	.w5(32'h3c475683),
	.w6(32'h385623e8),
	.w7(32'h3c2d70a0),
	.w8(32'hbacf61ca),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e307f),
	.w1(32'h3b1147f7),
	.w2(32'h3b8e6b99),
	.w3(32'h3c5285a4),
	.w4(32'h3b8d676c),
	.w5(32'h3c1b1019),
	.w6(32'hbc37d4d9),
	.w7(32'hbacc5ebc),
	.w8(32'h3bdf1a38),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ce9da),
	.w1(32'h3c1a969f),
	.w2(32'h3c6162f0),
	.w3(32'h3c4acd67),
	.w4(32'h3bd3be83),
	.w5(32'h3c66635a),
	.w6(32'hb9ebadcb),
	.w7(32'h3c2d45ce),
	.w8(32'h3c688292),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c824f09),
	.w1(32'h3a85595a),
	.w2(32'h3bb3c88c),
	.w3(32'h3c0dc77f),
	.w4(32'hbbc612e0),
	.w5(32'hba28877e),
	.w6(32'hbc2f22e4),
	.w7(32'hbbfad613),
	.w8(32'h3a4dd4e3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bd992),
	.w1(32'hba999573),
	.w2(32'hbb29f4e5),
	.w3(32'h3bea932d),
	.w4(32'hbb389075),
	.w5(32'h3b2eddb1),
	.w6(32'h39de38c5),
	.w7(32'h3b210c7e),
	.w8(32'h3bbd10d5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e9b43),
	.w1(32'hba860ee7),
	.w2(32'h3b65cba9),
	.w3(32'h3bb4de80),
	.w4(32'hbbc66109),
	.w5(32'hbb3ec3d8),
	.w6(32'hb9dffe39),
	.w7(32'h3b09a770),
	.w8(32'h3b9a2a5a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be997ef),
	.w1(32'h3cce26a6),
	.w2(32'h3d570740),
	.w3(32'h3baddb76),
	.w4(32'h3c8653c3),
	.w5(32'h3d101f6d),
	.w6(32'h3bf04585),
	.w7(32'h3cb1a186),
	.w8(32'h3bcc2ab3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1430b1),
	.w1(32'h3b6e2dec),
	.w2(32'h3bdbece8),
	.w3(32'h3ce00d6d),
	.w4(32'hba29cb7e),
	.w5(32'h3be890e4),
	.w6(32'hb8ad0717),
	.w7(32'h3aae398e),
	.w8(32'h3a911d7c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cb3a6),
	.w1(32'h3b4551ae),
	.w2(32'h3c9c85ae),
	.w3(32'h3b0bf4aa),
	.w4(32'h3c05569a),
	.w5(32'h3c452991),
	.w6(32'h3b8ecbfb),
	.w7(32'h3bdbce7d),
	.w8(32'h3ba25f03),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47f9d3),
	.w1(32'h3c78f026),
	.w2(32'h3c4d40bb),
	.w3(32'h3c44342f),
	.w4(32'h3c549ade),
	.w5(32'h3c3e3d24),
	.w6(32'h3c672524),
	.w7(32'h3c64dca3),
	.w8(32'h3c240232),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ac07d),
	.w1(32'h3cd51a7b),
	.w2(32'h3d3b3c12),
	.w3(32'h3c85cf07),
	.w4(32'h3c502709),
	.w5(32'h3d252635),
	.w6(32'h3c6ce187),
	.w7(32'h3cc90f90),
	.w8(32'h3c27f747),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd47ff6),
	.w1(32'hbacac91f),
	.w2(32'hbaa50d6a),
	.w3(32'h3b85a47e),
	.w4(32'h3bb8d030),
	.w5(32'h3b1fd0dd),
	.w6(32'h3af1acb2),
	.w7(32'h3bc11aa7),
	.w8(32'h3a0e9548),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da9b42),
	.w1(32'h3bd12ee9),
	.w2(32'h3c0be540),
	.w3(32'h3abd900b),
	.w4(32'h3bbeefb0),
	.w5(32'h3c0b1a84),
	.w6(32'h3bb81bd8),
	.w7(32'h3ae3297e),
	.w8(32'hbba56af6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85cdc6),
	.w1(32'hbb0af6c7),
	.w2(32'hbb904e12),
	.w3(32'h3c0bdcee),
	.w4(32'hbb394403),
	.w5(32'hbb11d2a9),
	.w6(32'hba29a0d7),
	.w7(32'hbb0e8b69),
	.w8(32'hbaaf0e1f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57ca75),
	.w1(32'hbc1e8d61),
	.w2(32'hbc8d8276),
	.w3(32'hbb76b56d),
	.w4(32'hbbad2469),
	.w5(32'hbc115391),
	.w6(32'hbc2f764a),
	.w7(32'hbc5cac9b),
	.w8(32'hbb862b06),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb47048),
	.w1(32'h3c95d1fb),
	.w2(32'h3d14b76e),
	.w3(32'h3ae41da1),
	.w4(32'h3c18df4a),
	.w5(32'h3cc2d57a),
	.w6(32'h3c06ce67),
	.w7(32'h3c9c923d),
	.w8(32'h3c3d5f96),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d5d97),
	.w1(32'h3b825279),
	.w2(32'h3c2a1cfe),
	.w3(32'h3c487629),
	.w4(32'h3b55621d),
	.w5(32'h3b602a7b),
	.w6(32'h3bbd7de3),
	.w7(32'h3ba06266),
	.w8(32'hbb4b6418),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9e989),
	.w1(32'hb7ca46ca),
	.w2(32'h3acdaec5),
	.w3(32'h3b19cd1e),
	.w4(32'hb9f0516a),
	.w5(32'h39ce44be),
	.w6(32'hbb1fe56e),
	.w7(32'h39358e3f),
	.w8(32'h3ba28592),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b844fad),
	.w1(32'hbbf7eee6),
	.w2(32'h3acc14dc),
	.w3(32'h3becd3ae),
	.w4(32'hbbed936b),
	.w5(32'hbbf3d906),
	.w6(32'hbc795a62),
	.w7(32'hbc841cba),
	.w8(32'hbc551e50),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc129803),
	.w1(32'hbc01e00f),
	.w2(32'hbc761df1),
	.w3(32'hbc20ac77),
	.w4(32'hbc4c6b9d),
	.w5(32'hbc0a0763),
	.w6(32'hbc387490),
	.w7(32'hbc4a1d51),
	.w8(32'hbc06f566),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f12b4),
	.w1(32'h3adb9d81),
	.w2(32'h3c193172),
	.w3(32'hbc462760),
	.w4(32'hbb0db95c),
	.w5(32'h3b6b8cfc),
	.w6(32'hbb020343),
	.w7(32'h3b89c461),
	.w8(32'hbb0b82eb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1d2e0),
	.w1(32'h3c8d851b),
	.w2(32'h3cdddd73),
	.w3(32'h3b8acccd),
	.w4(32'h3c08be1c),
	.w5(32'h3c52e551),
	.w6(32'h3b9ec69e),
	.w7(32'h3c848687),
	.w8(32'hb9b00189),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d51f),
	.w1(32'h3b2009da),
	.w2(32'h3b8d5709),
	.w3(32'hbc086b52),
	.w4(32'h3ad10d99),
	.w5(32'h3aa7e982),
	.w6(32'h3b68c163),
	.w7(32'h3c065a74),
	.w8(32'h3b7ea5dd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81a0c3),
	.w1(32'hbbff6863),
	.w2(32'hbb9ccdf0),
	.w3(32'hb714b71c),
	.w4(32'hbb1c04b6),
	.w5(32'hbc3c83d0),
	.w6(32'hbbdbae6e),
	.w7(32'h3b953bae),
	.w8(32'hbb0f3cb6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc237564),
	.w1(32'h3aa6a812),
	.w2(32'h39a5cc5e),
	.w3(32'hbb3eeea8),
	.w4(32'hb92744ae),
	.w5(32'hbb0debfe),
	.w6(32'h3a2bd90e),
	.w7(32'hba8228fe),
	.w8(32'hb902c7a2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbdcca),
	.w1(32'hbcc8950e),
	.w2(32'hbd1431f8),
	.w3(32'hbac2b78a),
	.w4(32'hbccf01b9),
	.w5(32'hbceaaefe),
	.w6(32'hbc39c7d7),
	.w7(32'hbce6f5e8),
	.w8(32'h3b5e6091),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule