module layer_9 (
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 2048;
	parameter IMG_SIZE = 26;

	wire	valid_out_0,
		valid_out_1,
		valid_out_2,
		valid_out_3,
		valid_out_4,
		valid_out_5,
		valid_out_6,
		valid_out_7,
		valid_out_8,
		valid_out_9,
		valid_out_10,
		valid_out_11,
		valid_out_12,
		valid_out_13,
		valid_out_14,
		valid_out_15,
		valid_out_16,
		valid_out_17,
		valid_out_18,
		valid_out_19,
		valid_out_20,
		valid_out_21,
		valid_out_22,
		valid_out_23,
		valid_out_24,
		valid_out_25,
		valid_out_26,
		valid_out_27,
		valid_out_28,
		valid_out_29,
		valid_out_30,
		valid_out_31,
		valid_out_32,
		valid_out_33,
		valid_out_34,
		valid_out_35,
		valid_out_36,
		valid_out_37,
		valid_out_38,
		valid_out_39,
		valid_out_40,
		valid_out_41,
		valid_out_42,
		valid_out_43,
		valid_out_44,
		valid_out_45,
		valid_out_46,
		valid_out_47,
		valid_out_48,
		valid_out_49,
		valid_out_50,
		valid_out_51,
		valid_out_52,
		valid_out_53,
		valid_out_54,
		valid_out_55,
		valid_out_56,
		valid_out_57,
		valid_out_58,
		valid_out_59,
		valid_out_60,
		valid_out_61,
		valid_out_62,
		valid_out_63,
		valid_out_64,
		valid_out_65,
		valid_out_66,
		valid_out_67,
		valid_out_68,
		valid_out_69,
		valid_out_70,
		valid_out_71,
		valid_out_72,
		valid_out_73,
		valid_out_74,
		valid_out_75,
		valid_out_76,
		valid_out_77,
		valid_out_78,
		valid_out_79,
		valid_out_80,
		valid_out_81,
		valid_out_82,
		valid_out_83,
		valid_out_84,
		valid_out_85,
		valid_out_86,
		valid_out_87,
		valid_out_88,
		valid_out_89,
		valid_out_90,
		valid_out_91,
		valid_out_92,
		valid_out_93,
		valid_out_94,
		valid_out_95,
		valid_out_96,
		valid_out_97,
		valid_out_98,
		valid_out_99,
		valid_out_100,
		valid_out_101,
		valid_out_102,
		valid_out_103,
		valid_out_104,
		valid_out_105,
		valid_out_106,
		valid_out_107,
		valid_out_108,
		valid_out_109,
		valid_out_110,
		valid_out_111,
		valid_out_112,
		valid_out_113,
		valid_out_114,
		valid_out_115,
		valid_out_116,
		valid_out_117,
		valid_out_118,
		valid_out_119,
		valid_out_120,
		valid_out_121,
		valid_out_122,
		valid_out_123,
		valid_out_124,
		valid_out_125,
		valid_out_126,
		valid_out_127,
		valid_out_128,
		valid_out_129,
		valid_out_130,
		valid_out_131,
		valid_out_132,
		valid_out_133,
		valid_out_134,
		valid_out_135,
		valid_out_136,
		valid_out_137,
		valid_out_138,
		valid_out_139,
		valid_out_140,
		valid_out_141,
		valid_out_142,
		valid_out_143,
		valid_out_144,
		valid_out_145,
		valid_out_146,
		valid_out_147,
		valid_out_148,
		valid_out_149,
		valid_out_150,
		valid_out_151,
		valid_out_152,
		valid_out_153,
		valid_out_154,
		valid_out_155,
		valid_out_156,
		valid_out_157,
		valid_out_158,
		valid_out_159,
		valid_out_160,
		valid_out_161,
		valid_out_162,
		valid_out_163,
		valid_out_164,
		valid_out_165,
		valid_out_166,
		valid_out_167,
		valid_out_168,
		valid_out_169,
		valid_out_170,
		valid_out_171,
		valid_out_172,
		valid_out_173,
		valid_out_174,
		valid_out_175,
		valid_out_176,
		valid_out_177,
		valid_out_178,
		valid_out_179,
		valid_out_180,
		valid_out_181,
		valid_out_182,
		valid_out_183,
		valid_out_184,
		valid_out_185,
		valid_out_186,
		valid_out_187,
		valid_out_188,
		valid_out_189,
		valid_out_190,
		valid_out_191,
		valid_out_192,
		valid_out_193,
		valid_out_194,
		valid_out_195,
		valid_out_196,
		valid_out_197,
		valid_out_198,
		valid_out_199,
		valid_out_200,
		valid_out_201,
		valid_out_202,
		valid_out_203,
		valid_out_204,
		valid_out_205,
		valid_out_206,
		valid_out_207,
		valid_out_208,
		valid_out_209,
		valid_out_210,
		valid_out_211,
		valid_out_212,
		valid_out_213,
		valid_out_214,
		valid_out_215,
		valid_out_216,
		valid_out_217,
		valid_out_218,
		valid_out_219,
		valid_out_220,
		valid_out_221,
		valid_out_222,
		valid_out_223,
		valid_out_224,
		valid_out_225,
		valid_out_226,
		valid_out_227,
		valid_out_228,
		valid_out_229,
		valid_out_230,
		valid_out_231,
		valid_out_232,
		valid_out_233,
		valid_out_234,
		valid_out_235,
		valid_out_236,
		valid_out_237,
		valid_out_238,
		valid_out_239,
		valid_out_240,
		valid_out_241,
		valid_out_242,
		valid_out_243,
		valid_out_244,
		valid_out_245,
		valid_out_246,
		valid_out_247,
		valid_out_248,
		valid_out_249,
		valid_out_250,
		valid_out_251,
		valid_out_252,
		valid_out_253,
		valid_out_254,
		valid_out_255;
Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7:0]),
	.valid_in(valid_in),
	.data_out(data_out[7:0]),
	.valid_out(valid_out_0)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15:8]),
	.valid_in(valid_in),
	.data_out(data_out[15:8]),
	.valid_out(valid_out_1)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[23:16]),
	.valid_in(valid_in),
	.data_out(data_out[23:16]),
	.valid_out(valid_out_2)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:24]),
	.valid_in(valid_in),
	.data_out(data_out[31:24]),
	.valid_out(valid_out_3)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[39:32]),
	.valid_in(valid_in),
	.data_out(data_out[39:32]),
	.valid_out(valid_out_4)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[47:40]),
	.valid_in(valid_in),
	.data_out(data_out[47:40]),
	.valid_out(valid_out_5)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[55:48]),
	.valid_in(valid_in),
	.data_out(data_out[55:48]),
	.valid_out(valid_out_6)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:56]),
	.valid_in(valid_in),
	.data_out(data_out[63:56]),
	.valid_out(valid_out_7)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[71:64]),
	.valid_in(valid_in),
	.data_out(data_out[71:64]),
	.valid_out(valid_out_8)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[79:72]),
	.valid_in(valid_in),
	.data_out(data_out[79:72]),
	.valid_out(valid_out_9)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[87:80]),
	.valid_in(valid_in),
	.data_out(data_out[87:80]),
	.valid_out(valid_out_10)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:88]),
	.valid_in(valid_in),
	.data_out(data_out[95:88]),
	.valid_out(valid_out_11)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[103:96]),
	.valid_in(valid_in),
	.data_out(data_out[103:96]),
	.valid_out(valid_out_12)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[111:104]),
	.valid_in(valid_in),
	.data_out(data_out[111:104]),
	.valid_out(valid_out_13)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[119:112]),
	.valid_in(valid_in),
	.data_out(data_out[119:112]),
	.valid_out(valid_out_14)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:120]),
	.valid_in(valid_in),
	.data_out(data_out[127:120]),
	.valid_out(valid_out_15)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[135:128]),
	.valid_in(valid_in),
	.data_out(data_out[135:128]),
	.valid_out(valid_out_16)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[143:136]),
	.valid_in(valid_in),
	.data_out(data_out[143:136]),
	.valid_out(valid_out_17)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[151:144]),
	.valid_in(valid_in),
	.data_out(data_out[151:144]),
	.valid_out(valid_out_18)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:152]),
	.valid_in(valid_in),
	.data_out(data_out[159:152]),
	.valid_out(valid_out_19)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[167:160]),
	.valid_in(valid_in),
	.data_out(data_out[167:160]),
	.valid_out(valid_out_20)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[175:168]),
	.valid_in(valid_in),
	.data_out(data_out[175:168]),
	.valid_out(valid_out_21)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[183:176]),
	.valid_in(valid_in),
	.data_out(data_out[183:176]),
	.valid_out(valid_out_22)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:184]),
	.valid_in(valid_in),
	.data_out(data_out[191:184]),
	.valid_out(valid_out_23)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[199:192]),
	.valid_in(valid_in),
	.data_out(data_out[199:192]),
	.valid_out(valid_out_24)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[207:200]),
	.valid_in(valid_in),
	.data_out(data_out[207:200]),
	.valid_out(valid_out_25)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[215:208]),
	.valid_in(valid_in),
	.data_out(data_out[215:208]),
	.valid_out(valid_out_26)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:216]),
	.valid_in(valid_in),
	.data_out(data_out[223:216]),
	.valid_out(valid_out_27)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[231:224]),
	.valid_in(valid_in),
	.data_out(data_out[231:224]),
	.valid_out(valid_out_28)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[239:232]),
	.valid_in(valid_in),
	.data_out(data_out[239:232]),
	.valid_out(valid_out_29)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[247:240]),
	.valid_in(valid_in),
	.data_out(data_out[247:240]),
	.valid_out(valid_out_30)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:248]),
	.valid_in(valid_in),
	.data_out(data_out[255:248]),
	.valid_out(valid_out_31)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[263:256]),
	.valid_in(valid_in),
	.data_out(data_out[263:256]),
	.valid_out(valid_out_32)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[271:264]),
	.valid_in(valid_in),
	.data_out(data_out[271:264]),
	.valid_out(valid_out_33)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[279:272]),
	.valid_in(valid_in),
	.data_out(data_out[279:272]),
	.valid_out(valid_out_34)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:280]),
	.valid_in(valid_in),
	.data_out(data_out[287:280]),
	.valid_out(valid_out_35)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[295:288]),
	.valid_in(valid_in),
	.data_out(data_out[295:288]),
	.valid_out(valid_out_36)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[303:296]),
	.valid_in(valid_in),
	.data_out(data_out[303:296]),
	.valid_out(valid_out_37)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[311:304]),
	.valid_in(valid_in),
	.data_out(data_out[311:304]),
	.valid_out(valid_out_38)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:312]),
	.valid_in(valid_in),
	.data_out(data_out[319:312]),
	.valid_out(valid_out_39)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[327:320]),
	.valid_in(valid_in),
	.data_out(data_out[327:320]),
	.valid_out(valid_out_40)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[335:328]),
	.valid_in(valid_in),
	.data_out(data_out[335:328]),
	.valid_out(valid_out_41)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[343:336]),
	.valid_in(valid_in),
	.data_out(data_out[343:336]),
	.valid_out(valid_out_42)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:344]),
	.valid_in(valid_in),
	.data_out(data_out[351:344]),
	.valid_out(valid_out_43)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[359:352]),
	.valid_in(valid_in),
	.data_out(data_out[359:352]),
	.valid_out(valid_out_44)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[367:360]),
	.valid_in(valid_in),
	.data_out(data_out[367:360]),
	.valid_out(valid_out_45)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[375:368]),
	.valid_in(valid_in),
	.data_out(data_out[375:368]),
	.valid_out(valid_out_46)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:376]),
	.valid_in(valid_in),
	.data_out(data_out[383:376]),
	.valid_out(valid_out_47)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[391:384]),
	.valid_in(valid_in),
	.data_out(data_out[391:384]),
	.valid_out(valid_out_48)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[399:392]),
	.valid_in(valid_in),
	.data_out(data_out[399:392]),
	.valid_out(valid_out_49)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[407:400]),
	.valid_in(valid_in),
	.data_out(data_out[407:400]),
	.valid_out(valid_out_50)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:408]),
	.valid_in(valid_in),
	.data_out(data_out[415:408]),
	.valid_out(valid_out_51)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[423:416]),
	.valid_in(valid_in),
	.data_out(data_out[423:416]),
	.valid_out(valid_out_52)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[431:424]),
	.valid_in(valid_in),
	.data_out(data_out[431:424]),
	.valid_out(valid_out_53)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[439:432]),
	.valid_in(valid_in),
	.data_out(data_out[439:432]),
	.valid_out(valid_out_54)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:440]),
	.valid_in(valid_in),
	.data_out(data_out[447:440]),
	.valid_out(valid_out_55)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[455:448]),
	.valid_in(valid_in),
	.data_out(data_out[455:448]),
	.valid_out(valid_out_56)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[463:456]),
	.valid_in(valid_in),
	.data_out(data_out[463:456]),
	.valid_out(valid_out_57)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[471:464]),
	.valid_in(valid_in),
	.data_out(data_out[471:464]),
	.valid_out(valid_out_58)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:472]),
	.valid_in(valid_in),
	.data_out(data_out[479:472]),
	.valid_out(valid_out_59)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[487:480]),
	.valid_in(valid_in),
	.data_out(data_out[487:480]),
	.valid_out(valid_out_60)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[495:488]),
	.valid_in(valid_in),
	.data_out(data_out[495:488]),
	.valid_out(valid_out_61)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[503:496]),
	.valid_in(valid_in),
	.data_out(data_out[503:496]),
	.valid_out(valid_out_62)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:504]),
	.valid_in(valid_in),
	.data_out(data_out[511:504]),
	.valid_out(valid_out_63)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[519:512]),
	.valid_in(valid_in),
	.data_out(data_out[519:512]),
	.valid_out(valid_out_64)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[527:520]),
	.valid_in(valid_in),
	.data_out(data_out[527:520]),
	.valid_out(valid_out_65)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[535:528]),
	.valid_in(valid_in),
	.data_out(data_out[535:528]),
	.valid_out(valid_out_66)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:536]),
	.valid_in(valid_in),
	.data_out(data_out[543:536]),
	.valid_out(valid_out_67)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[551:544]),
	.valid_in(valid_in),
	.data_out(data_out[551:544]),
	.valid_out(valid_out_68)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[559:552]),
	.valid_in(valid_in),
	.data_out(data_out[559:552]),
	.valid_out(valid_out_69)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[567:560]),
	.valid_in(valid_in),
	.data_out(data_out[567:560]),
	.valid_out(valid_out_70)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:568]),
	.valid_in(valid_in),
	.data_out(data_out[575:568]),
	.valid_out(valid_out_71)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[583:576]),
	.valid_in(valid_in),
	.data_out(data_out[583:576]),
	.valid_out(valid_out_72)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[591:584]),
	.valid_in(valid_in),
	.data_out(data_out[591:584]),
	.valid_out(valid_out_73)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[599:592]),
	.valid_in(valid_in),
	.data_out(data_out[599:592]),
	.valid_out(valid_out_74)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:600]),
	.valid_in(valid_in),
	.data_out(data_out[607:600]),
	.valid_out(valid_out_75)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[615:608]),
	.valid_in(valid_in),
	.data_out(data_out[615:608]),
	.valid_out(valid_out_76)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[623:616]),
	.valid_in(valid_in),
	.data_out(data_out[623:616]),
	.valid_out(valid_out_77)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[631:624]),
	.valid_in(valid_in),
	.data_out(data_out[631:624]),
	.valid_out(valid_out_78)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:632]),
	.valid_in(valid_in),
	.data_out(data_out[639:632]),
	.valid_out(valid_out_79)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[647:640]),
	.valid_in(valid_in),
	.data_out(data_out[647:640]),
	.valid_out(valid_out_80)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[655:648]),
	.valid_in(valid_in),
	.data_out(data_out[655:648]),
	.valid_out(valid_out_81)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[663:656]),
	.valid_in(valid_in),
	.data_out(data_out[663:656]),
	.valid_out(valid_out_82)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:664]),
	.valid_in(valid_in),
	.data_out(data_out[671:664]),
	.valid_out(valid_out_83)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[679:672]),
	.valid_in(valid_in),
	.data_out(data_out[679:672]),
	.valid_out(valid_out_84)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[687:680]),
	.valid_in(valid_in),
	.data_out(data_out[687:680]),
	.valid_out(valid_out_85)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[695:688]),
	.valid_in(valid_in),
	.data_out(data_out[695:688]),
	.valid_out(valid_out_86)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:696]),
	.valid_in(valid_in),
	.data_out(data_out[703:696]),
	.valid_out(valid_out_87)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[711:704]),
	.valid_in(valid_in),
	.data_out(data_out[711:704]),
	.valid_out(valid_out_88)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[719:712]),
	.valid_in(valid_in),
	.data_out(data_out[719:712]),
	.valid_out(valid_out_89)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[727:720]),
	.valid_in(valid_in),
	.data_out(data_out[727:720]),
	.valid_out(valid_out_90)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:728]),
	.valid_in(valid_in),
	.data_out(data_out[735:728]),
	.valid_out(valid_out_91)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[743:736]),
	.valid_in(valid_in),
	.data_out(data_out[743:736]),
	.valid_out(valid_out_92)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[751:744]),
	.valid_in(valid_in),
	.data_out(data_out[751:744]),
	.valid_out(valid_out_93)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[759:752]),
	.valid_in(valid_in),
	.data_out(data_out[759:752]),
	.valid_out(valid_out_94)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:760]),
	.valid_in(valid_in),
	.data_out(data_out[767:760]),
	.valid_out(valid_out_95)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[775:768]),
	.valid_in(valid_in),
	.data_out(data_out[775:768]),
	.valid_out(valid_out_96)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[783:776]),
	.valid_in(valid_in),
	.data_out(data_out[783:776]),
	.valid_out(valid_out_97)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[791:784]),
	.valid_in(valid_in),
	.data_out(data_out[791:784]),
	.valid_out(valid_out_98)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:792]),
	.valid_in(valid_in),
	.data_out(data_out[799:792]),
	.valid_out(valid_out_99)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[807:800]),
	.valid_in(valid_in),
	.data_out(data_out[807:800]),
	.valid_out(valid_out_100)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[815:808]),
	.valid_in(valid_in),
	.data_out(data_out[815:808]),
	.valid_out(valid_out_101)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[823:816]),
	.valid_in(valid_in),
	.data_out(data_out[823:816]),
	.valid_out(valid_out_102)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:824]),
	.valid_in(valid_in),
	.data_out(data_out[831:824]),
	.valid_out(valid_out_103)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[839:832]),
	.valid_in(valid_in),
	.data_out(data_out[839:832]),
	.valid_out(valid_out_104)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[847:840]),
	.valid_in(valid_in),
	.data_out(data_out[847:840]),
	.valid_out(valid_out_105)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[855:848]),
	.valid_in(valid_in),
	.data_out(data_out[855:848]),
	.valid_out(valid_out_106)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:856]),
	.valid_in(valid_in),
	.data_out(data_out[863:856]),
	.valid_out(valid_out_107)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[871:864]),
	.valid_in(valid_in),
	.data_out(data_out[871:864]),
	.valid_out(valid_out_108)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[879:872]),
	.valid_in(valid_in),
	.data_out(data_out[879:872]),
	.valid_out(valid_out_109)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[887:880]),
	.valid_in(valid_in),
	.data_out(data_out[887:880]),
	.valid_out(valid_out_110)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:888]),
	.valid_in(valid_in),
	.data_out(data_out[895:888]),
	.valid_out(valid_out_111)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[903:896]),
	.valid_in(valid_in),
	.data_out(data_out[903:896]),
	.valid_out(valid_out_112)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[911:904]),
	.valid_in(valid_in),
	.data_out(data_out[911:904]),
	.valid_out(valid_out_113)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[919:912]),
	.valid_in(valid_in),
	.data_out(data_out[919:912]),
	.valid_out(valid_out_114)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:920]),
	.valid_in(valid_in),
	.data_out(data_out[927:920]),
	.valid_out(valid_out_115)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[935:928]),
	.valid_in(valid_in),
	.data_out(data_out[935:928]),
	.valid_out(valid_out_116)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[943:936]),
	.valid_in(valid_in),
	.data_out(data_out[943:936]),
	.valid_out(valid_out_117)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[951:944]),
	.valid_in(valid_in),
	.data_out(data_out[951:944]),
	.valid_out(valid_out_118)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:952]),
	.valid_in(valid_in),
	.data_out(data_out[959:952]),
	.valid_out(valid_out_119)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[967:960]),
	.valid_in(valid_in),
	.data_out(data_out[967:960]),
	.valid_out(valid_out_120)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[975:968]),
	.valid_in(valid_in),
	.data_out(data_out[975:968]),
	.valid_out(valid_out_121)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[983:976]),
	.valid_in(valid_in),
	.data_out(data_out[983:976]),
	.valid_out(valid_out_122)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:984]),
	.valid_in(valid_in),
	.data_out(data_out[991:984]),
	.valid_out(valid_out_123)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[999:992]),
	.valid_in(valid_in),
	.data_out(data_out[999:992]),
	.valid_out(valid_out_124)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1007:1000]),
	.valid_in(valid_in),
	.data_out(data_out[1007:1000]),
	.valid_out(valid_out_125)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1015:1008]),
	.valid_in(valid_in),
	.data_out(data_out[1015:1008]),
	.valid_out(valid_out_126)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:1016]),
	.valid_in(valid_in),
	.data_out(data_out[1023:1016]),
	.valid_out(valid_out_127)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1031:1024]),
	.valid_in(valid_in),
	.data_out(data_out[1031:1024]),
	.valid_out(valid_out_128)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1039:1032]),
	.valid_in(valid_in),
	.data_out(data_out[1039:1032]),
	.valid_out(valid_out_129)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1047:1040]),
	.valid_in(valid_in),
	.data_out(data_out[1047:1040]),
	.valid_out(valid_out_130)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1048]),
	.valid_in(valid_in),
	.data_out(data_out[1055:1048]),
	.valid_out(valid_out_131)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1063:1056]),
	.valid_in(valid_in),
	.data_out(data_out[1063:1056]),
	.valid_out(valid_out_132)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1071:1064]),
	.valid_in(valid_in),
	.data_out(data_out[1071:1064]),
	.valid_out(valid_out_133)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1079:1072]),
	.valid_in(valid_in),
	.data_out(data_out[1079:1072]),
	.valid_out(valid_out_134)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1080]),
	.valid_in(valid_in),
	.data_out(data_out[1087:1080]),
	.valid_out(valid_out_135)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1095:1088]),
	.valid_in(valid_in),
	.data_out(data_out[1095:1088]),
	.valid_out(valid_out_136)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1103:1096]),
	.valid_in(valid_in),
	.data_out(data_out[1103:1096]),
	.valid_out(valid_out_137)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1111:1104]),
	.valid_in(valid_in),
	.data_out(data_out[1111:1104]),
	.valid_out(valid_out_138)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1112]),
	.valid_in(valid_in),
	.data_out(data_out[1119:1112]),
	.valid_out(valid_out_139)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1127:1120]),
	.valid_in(valid_in),
	.data_out(data_out[1127:1120]),
	.valid_out(valid_out_140)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1135:1128]),
	.valid_in(valid_in),
	.data_out(data_out[1135:1128]),
	.valid_out(valid_out_141)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1143:1136]),
	.valid_in(valid_in),
	.data_out(data_out[1143:1136]),
	.valid_out(valid_out_142)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1144]),
	.valid_in(valid_in),
	.data_out(data_out[1151:1144]),
	.valid_out(valid_out_143)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1159:1152]),
	.valid_in(valid_in),
	.data_out(data_out[1159:1152]),
	.valid_out(valid_out_144)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1167:1160]),
	.valid_in(valid_in),
	.data_out(data_out[1167:1160]),
	.valid_out(valid_out_145)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1175:1168]),
	.valid_in(valid_in),
	.data_out(data_out[1175:1168]),
	.valid_out(valid_out_146)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1176]),
	.valid_in(valid_in),
	.data_out(data_out[1183:1176]),
	.valid_out(valid_out_147)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1191:1184]),
	.valid_in(valid_in),
	.data_out(data_out[1191:1184]),
	.valid_out(valid_out_148)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1199:1192]),
	.valid_in(valid_in),
	.data_out(data_out[1199:1192]),
	.valid_out(valid_out_149)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1207:1200]),
	.valid_in(valid_in),
	.data_out(data_out[1207:1200]),
	.valid_out(valid_out_150)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1208]),
	.valid_in(valid_in),
	.data_out(data_out[1215:1208]),
	.valid_out(valid_out_151)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1223:1216]),
	.valid_in(valid_in),
	.data_out(data_out[1223:1216]),
	.valid_out(valid_out_152)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1231:1224]),
	.valid_in(valid_in),
	.data_out(data_out[1231:1224]),
	.valid_out(valid_out_153)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1239:1232]),
	.valid_in(valid_in),
	.data_out(data_out[1239:1232]),
	.valid_out(valid_out_154)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1240]),
	.valid_in(valid_in),
	.data_out(data_out[1247:1240]),
	.valid_out(valid_out_155)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1255:1248]),
	.valid_in(valid_in),
	.data_out(data_out[1255:1248]),
	.valid_out(valid_out_156)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1263:1256]),
	.valid_in(valid_in),
	.data_out(data_out[1263:1256]),
	.valid_out(valid_out_157)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1271:1264]),
	.valid_in(valid_in),
	.data_out(data_out[1271:1264]),
	.valid_out(valid_out_158)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1272]),
	.valid_in(valid_in),
	.data_out(data_out[1279:1272]),
	.valid_out(valid_out_159)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1287:1280]),
	.valid_in(valid_in),
	.data_out(data_out[1287:1280]),
	.valid_out(valid_out_160)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1295:1288]),
	.valid_in(valid_in),
	.data_out(data_out[1295:1288]),
	.valid_out(valid_out_161)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1303:1296]),
	.valid_in(valid_in),
	.data_out(data_out[1303:1296]),
	.valid_out(valid_out_162)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1304]),
	.valid_in(valid_in),
	.data_out(data_out[1311:1304]),
	.valid_out(valid_out_163)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1319:1312]),
	.valid_in(valid_in),
	.data_out(data_out[1319:1312]),
	.valid_out(valid_out_164)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1327:1320]),
	.valid_in(valid_in),
	.data_out(data_out[1327:1320]),
	.valid_out(valid_out_165)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1335:1328]),
	.valid_in(valid_in),
	.data_out(data_out[1335:1328]),
	.valid_out(valid_out_166)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1336]),
	.valid_in(valid_in),
	.data_out(data_out[1343:1336]),
	.valid_out(valid_out_167)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1351:1344]),
	.valid_in(valid_in),
	.data_out(data_out[1351:1344]),
	.valid_out(valid_out_168)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1359:1352]),
	.valid_in(valid_in),
	.data_out(data_out[1359:1352]),
	.valid_out(valid_out_169)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1367:1360]),
	.valid_in(valid_in),
	.data_out(data_out[1367:1360]),
	.valid_out(valid_out_170)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1368]),
	.valid_in(valid_in),
	.data_out(data_out[1375:1368]),
	.valid_out(valid_out_171)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1383:1376]),
	.valid_in(valid_in),
	.data_out(data_out[1383:1376]),
	.valid_out(valid_out_172)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1391:1384]),
	.valid_in(valid_in),
	.data_out(data_out[1391:1384]),
	.valid_out(valid_out_173)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1399:1392]),
	.valid_in(valid_in),
	.data_out(data_out[1399:1392]),
	.valid_out(valid_out_174)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1400]),
	.valid_in(valid_in),
	.data_out(data_out[1407:1400]),
	.valid_out(valid_out_175)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1415:1408]),
	.valid_in(valid_in),
	.data_out(data_out[1415:1408]),
	.valid_out(valid_out_176)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1423:1416]),
	.valid_in(valid_in),
	.data_out(data_out[1423:1416]),
	.valid_out(valid_out_177)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1431:1424]),
	.valid_in(valid_in),
	.data_out(data_out[1431:1424]),
	.valid_out(valid_out_178)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1432]),
	.valid_in(valid_in),
	.data_out(data_out[1439:1432]),
	.valid_out(valid_out_179)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1447:1440]),
	.valid_in(valid_in),
	.data_out(data_out[1447:1440]),
	.valid_out(valid_out_180)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1455:1448]),
	.valid_in(valid_in),
	.data_out(data_out[1455:1448]),
	.valid_out(valid_out_181)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1463:1456]),
	.valid_in(valid_in),
	.data_out(data_out[1463:1456]),
	.valid_out(valid_out_182)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1464]),
	.valid_in(valid_in),
	.data_out(data_out[1471:1464]),
	.valid_out(valid_out_183)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1479:1472]),
	.valid_in(valid_in),
	.data_out(data_out[1479:1472]),
	.valid_out(valid_out_184)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1487:1480]),
	.valid_in(valid_in),
	.data_out(data_out[1487:1480]),
	.valid_out(valid_out_185)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1495:1488]),
	.valid_in(valid_in),
	.data_out(data_out[1495:1488]),
	.valid_out(valid_out_186)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1496]),
	.valid_in(valid_in),
	.data_out(data_out[1503:1496]),
	.valid_out(valid_out_187)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1511:1504]),
	.valid_in(valid_in),
	.data_out(data_out[1511:1504]),
	.valid_out(valid_out_188)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1519:1512]),
	.valid_in(valid_in),
	.data_out(data_out[1519:1512]),
	.valid_out(valid_out_189)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1527:1520]),
	.valid_in(valid_in),
	.data_out(data_out[1527:1520]),
	.valid_out(valid_out_190)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1528]),
	.valid_in(valid_in),
	.data_out(data_out[1535:1528]),
	.valid_out(valid_out_191)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1543:1536]),
	.valid_in(valid_in),
	.data_out(data_out[1543:1536]),
	.valid_out(valid_out_192)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1551:1544]),
	.valid_in(valid_in),
	.data_out(data_out[1551:1544]),
	.valid_out(valid_out_193)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1559:1552]),
	.valid_in(valid_in),
	.data_out(data_out[1559:1552]),
	.valid_out(valid_out_194)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1560]),
	.valid_in(valid_in),
	.data_out(data_out[1567:1560]),
	.valid_out(valid_out_195)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1575:1568]),
	.valid_in(valid_in),
	.data_out(data_out[1575:1568]),
	.valid_out(valid_out_196)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1583:1576]),
	.valid_in(valid_in),
	.data_out(data_out[1583:1576]),
	.valid_out(valid_out_197)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1591:1584]),
	.valid_in(valid_in),
	.data_out(data_out[1591:1584]),
	.valid_out(valid_out_198)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1592]),
	.valid_in(valid_in),
	.data_out(data_out[1599:1592]),
	.valid_out(valid_out_199)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1607:1600]),
	.valid_in(valid_in),
	.data_out(data_out[1607:1600]),
	.valid_out(valid_out_200)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1615:1608]),
	.valid_in(valid_in),
	.data_out(data_out[1615:1608]),
	.valid_out(valid_out_201)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1623:1616]),
	.valid_in(valid_in),
	.data_out(data_out[1623:1616]),
	.valid_out(valid_out_202)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1624]),
	.valid_in(valid_in),
	.data_out(data_out[1631:1624]),
	.valid_out(valid_out_203)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1639:1632]),
	.valid_in(valid_in),
	.data_out(data_out[1639:1632]),
	.valid_out(valid_out_204)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1647:1640]),
	.valid_in(valid_in),
	.data_out(data_out[1647:1640]),
	.valid_out(valid_out_205)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1655:1648]),
	.valid_in(valid_in),
	.data_out(data_out[1655:1648]),
	.valid_out(valid_out_206)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1656]),
	.valid_in(valid_in),
	.data_out(data_out[1663:1656]),
	.valid_out(valid_out_207)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1671:1664]),
	.valid_in(valid_in),
	.data_out(data_out[1671:1664]),
	.valid_out(valid_out_208)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1679:1672]),
	.valid_in(valid_in),
	.data_out(data_out[1679:1672]),
	.valid_out(valid_out_209)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1687:1680]),
	.valid_in(valid_in),
	.data_out(data_out[1687:1680]),
	.valid_out(valid_out_210)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1688]),
	.valid_in(valid_in),
	.data_out(data_out[1695:1688]),
	.valid_out(valid_out_211)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1703:1696]),
	.valid_in(valid_in),
	.data_out(data_out[1703:1696]),
	.valid_out(valid_out_212)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1711:1704]),
	.valid_in(valid_in),
	.data_out(data_out[1711:1704]),
	.valid_out(valid_out_213)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1719:1712]),
	.valid_in(valid_in),
	.data_out(data_out[1719:1712]),
	.valid_out(valid_out_214)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1720]),
	.valid_in(valid_in),
	.data_out(data_out[1727:1720]),
	.valid_out(valid_out_215)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1735:1728]),
	.valid_in(valid_in),
	.data_out(data_out[1735:1728]),
	.valid_out(valid_out_216)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1743:1736]),
	.valid_in(valid_in),
	.data_out(data_out[1743:1736]),
	.valid_out(valid_out_217)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1751:1744]),
	.valid_in(valid_in),
	.data_out(data_out[1751:1744]),
	.valid_out(valid_out_218)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1752]),
	.valid_in(valid_in),
	.data_out(data_out[1759:1752]),
	.valid_out(valid_out_219)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1767:1760]),
	.valid_in(valid_in),
	.data_out(data_out[1767:1760]),
	.valid_out(valid_out_220)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1775:1768]),
	.valid_in(valid_in),
	.data_out(data_out[1775:1768]),
	.valid_out(valid_out_221)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1783:1776]),
	.valid_in(valid_in),
	.data_out(data_out[1783:1776]),
	.valid_out(valid_out_222)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1784]),
	.valid_in(valid_in),
	.data_out(data_out[1791:1784]),
	.valid_out(valid_out_223)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1799:1792]),
	.valid_in(valid_in),
	.data_out(data_out[1799:1792]),
	.valid_out(valid_out_224)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1807:1800]),
	.valid_in(valid_in),
	.data_out(data_out[1807:1800]),
	.valid_out(valid_out_225)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1815:1808]),
	.valid_in(valid_in),
	.data_out(data_out[1815:1808]),
	.valid_out(valid_out_226)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1816]),
	.valid_in(valid_in),
	.data_out(data_out[1823:1816]),
	.valid_out(valid_out_227)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1831:1824]),
	.valid_in(valid_in),
	.data_out(data_out[1831:1824]),
	.valid_out(valid_out_228)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1839:1832]),
	.valid_in(valid_in),
	.data_out(data_out[1839:1832]),
	.valid_out(valid_out_229)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1847:1840]),
	.valid_in(valid_in),
	.data_out(data_out[1847:1840]),
	.valid_out(valid_out_230)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1848]),
	.valid_in(valid_in),
	.data_out(data_out[1855:1848]),
	.valid_out(valid_out_231)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1863:1856]),
	.valid_in(valid_in),
	.data_out(data_out[1863:1856]),
	.valid_out(valid_out_232)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1871:1864]),
	.valid_in(valid_in),
	.data_out(data_out[1871:1864]),
	.valid_out(valid_out_233)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1879:1872]),
	.valid_in(valid_in),
	.data_out(data_out[1879:1872]),
	.valid_out(valid_out_234)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1880]),
	.valid_in(valid_in),
	.data_out(data_out[1887:1880]),
	.valid_out(valid_out_235)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1895:1888]),
	.valid_in(valid_in),
	.data_out(data_out[1895:1888]),
	.valid_out(valid_out_236)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1903:1896]),
	.valid_in(valid_in),
	.data_out(data_out[1903:1896]),
	.valid_out(valid_out_237)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1911:1904]),
	.valid_in(valid_in),
	.data_out(data_out[1911:1904]),
	.valid_out(valid_out_238)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1912]),
	.valid_in(valid_in),
	.data_out(data_out[1919:1912]),
	.valid_out(valid_out_239)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1927:1920]),
	.valid_in(valid_in),
	.data_out(data_out[1927:1920]),
	.valid_out(valid_out_240)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1935:1928]),
	.valid_in(valid_in),
	.data_out(data_out[1935:1928]),
	.valid_out(valid_out_241)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1943:1936]),
	.valid_in(valid_in),
	.data_out(data_out[1943:1936]),
	.valid_out(valid_out_242)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1944]),
	.valid_in(valid_in),
	.data_out(data_out[1951:1944]),
	.valid_out(valid_out_243)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1959:1952]),
	.valid_in(valid_in),
	.data_out(data_out[1959:1952]),
	.valid_out(valid_out_244)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1967:1960]),
	.valid_in(valid_in),
	.data_out(data_out[1967:1960]),
	.valid_out(valid_out_245)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1975:1968]),
	.valid_in(valid_in),
	.data_out(data_out[1975:1968]),
	.valid_out(valid_out_246)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1976]),
	.valid_in(valid_in),
	.data_out(data_out[1983:1976]),
	.valid_out(valid_out_247)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1991:1984]),
	.valid_in(valid_in),
	.data_out(data_out[1991:1984]),
	.valid_out(valid_out_248)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1999:1992]),
	.valid_in(valid_in),
	.data_out(data_out[1999:1992]),
	.valid_out(valid_out_249)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2007:2000]),
	.valid_in(valid_in),
	.data_out(data_out[2007:2000]),
	.valid_out(valid_out_250)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:2008]),
	.valid_in(valid_in),
	.data_out(data_out[2015:2008]),
	.valid_out(valid_out_251)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2023:2016]),
	.valid_in(valid_in),
	.data_out(data_out[2023:2016]),
	.valid_out(valid_out_252)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2031:2024]),
	.valid_in(valid_in),
	.data_out(data_out[2031:2024]),
	.valid_out(valid_out_253)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2039:2032]),
	.valid_in(valid_in),
	.data_out(data_out[2039:2032]),
	.valid_out(valid_out_254)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2040]),
	.valid_in(valid_in),
	.data_out(data_out[2047:2040]),
	.valid_out(valid_out_255)
);

	assign valid_out = valid_out_0 & valid_out_1 & valid_out_2 & valid_out_3 & valid_out_4 & valid_out_5 & valid_out_6 & valid_out_7 & valid_out_8 & valid_out_9 & valid_out_10 & valid_out_11 & valid_out_12 & valid_out_13 & valid_out_14 & valid_out_15 & valid_out_16 & valid_out_17 & valid_out_18 & valid_out_19 & valid_out_20 & valid_out_21 & valid_out_22 & valid_out_23 & valid_out_24 & valid_out_25 & valid_out_26 & valid_out_27 & valid_out_28 & valid_out_29 & valid_out_30 & valid_out_31 & valid_out_32 & valid_out_33 & valid_out_34 & valid_out_35 & valid_out_36 & valid_out_37 & valid_out_38 & valid_out_39 & valid_out_40 & valid_out_41 & valid_out_42 & valid_out_43 & valid_out_44 & valid_out_45 & valid_out_46 & valid_out_47 & valid_out_48 & valid_out_49 & valid_out_50 & valid_out_51 & valid_out_52 & valid_out_53 & valid_out_54 & valid_out_55 & valid_out_56 & valid_out_57 & valid_out_58 & valid_out_59 & valid_out_60 & valid_out_61 & valid_out_62 & valid_out_63 & valid_out_64 & valid_out_65 & valid_out_66 & valid_out_67 & valid_out_68 & valid_out_69 & valid_out_70 & valid_out_71 & valid_out_72 & valid_out_73 & valid_out_74 & valid_out_75 & valid_out_76 & valid_out_77 & valid_out_78 & valid_out_79 & valid_out_80 & valid_out_81 & valid_out_82 & valid_out_83 & valid_out_84 & valid_out_85 & valid_out_86 & valid_out_87 & valid_out_88 & valid_out_89 & valid_out_90 & valid_out_91 & valid_out_92 & valid_out_93 & valid_out_94 & valid_out_95 & valid_out_96 & valid_out_97 & valid_out_98 & valid_out_99 & valid_out_100 & valid_out_101 & valid_out_102 & valid_out_103 & valid_out_104 & valid_out_105 & valid_out_106 & valid_out_107 & valid_out_108 & valid_out_109 & valid_out_110 & valid_out_111 & valid_out_112 & valid_out_113 & valid_out_114 & valid_out_115 & valid_out_116 & valid_out_117 & valid_out_118 & valid_out_119 & valid_out_120 & valid_out_121 & valid_out_122 & valid_out_123 & valid_out_124 & valid_out_125 & valid_out_126 & valid_out_127 & valid_out_128 & valid_out_129 & valid_out_130 & valid_out_131 & valid_out_132 & valid_out_133 & valid_out_134 & valid_out_135 & valid_out_136 & valid_out_137 & valid_out_138 & valid_out_139 & valid_out_140 & valid_out_141 & valid_out_142 & valid_out_143 & valid_out_144 & valid_out_145 & valid_out_146 & valid_out_147 & valid_out_148 & valid_out_149 & valid_out_150 & valid_out_151 & valid_out_152 & valid_out_153 & valid_out_154 & valid_out_155 & valid_out_156 & valid_out_157 & valid_out_158 & valid_out_159 & valid_out_160 & valid_out_161 & valid_out_162 & valid_out_163 & valid_out_164 & valid_out_165 & valid_out_166 & valid_out_167 & valid_out_168 & valid_out_169 & valid_out_170 & valid_out_171 & valid_out_172 & valid_out_173 & valid_out_174 & valid_out_175 & valid_out_176 & valid_out_177 & valid_out_178 & valid_out_179 & valid_out_180 & valid_out_181 & valid_out_182 & valid_out_183 & valid_out_184 & valid_out_185 & valid_out_186 & valid_out_187 & valid_out_188 & valid_out_189 & valid_out_190 & valid_out_191 & valid_out_192 & valid_out_193 & valid_out_194 & valid_out_195 & valid_out_196 & valid_out_197 & valid_out_198 & valid_out_199 & valid_out_200 & valid_out_201 & valid_out_202 & valid_out_203 & valid_out_204 & valid_out_205 & valid_out_206 & valid_out_207 & valid_out_208 & valid_out_209 & valid_out_210 & valid_out_211 & valid_out_212 & valid_out_213 & valid_out_214 & valid_out_215 & valid_out_216 & valid_out_217 & valid_out_218 & valid_out_219 & valid_out_220 & valid_out_221 & valid_out_222 & valid_out_223 & valid_out_224 & valid_out_225 & valid_out_226 & valid_out_227 & valid_out_228 & valid_out_229 & valid_out_230 & valid_out_231 & valid_out_232 & valid_out_233 & valid_out_234 & valid_out_235 & valid_out_236 & valid_out_237 & valid_out_238 & valid_out_239 & valid_out_240 & valid_out_241 & valid_out_242 & valid_out_243 & valid_out_244 & valid_out_245 & valid_out_246 & valid_out_247 & valid_out_248 & valid_out_249 & valid_out_250 & valid_out_251 & valid_out_252 & valid_out_253 & valid_out_254 & valid_out_255;
endmodule