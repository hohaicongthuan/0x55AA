module layer_6_featuremap_33(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bad65),
	.w1(32'hbbfe4f0b),
	.w2(32'hbb9200ea),
	.w3(32'hbb932681),
	.w4(32'h3ba239b2),
	.w5(32'h3bae76e1),
	.w6(32'hbac7ea82),
	.w7(32'h3bd1d947),
	.w8(32'h3bdc7bc4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb437d73),
	.w1(32'hbabfc3f7),
	.w2(32'h3ad5cb11),
	.w3(32'hba5e6764),
	.w4(32'hbb64b213),
	.w5(32'hbb5e1907),
	.w6(32'h3c82ec6e),
	.w7(32'h3c3a1372),
	.w8(32'h3c5edc39),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7230c),
	.w1(32'hbaa47b15),
	.w2(32'hbbf29647),
	.w3(32'hbc1eb96a),
	.w4(32'hbbbd5da9),
	.w5(32'hbc5f524b),
	.w6(32'hbbb89ae7),
	.w7(32'hbc96f0c6),
	.w8(32'hbcc79547),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe019d6),
	.w1(32'h3ad72b64),
	.w2(32'h3b37bf53),
	.w3(32'hbadc8166),
	.w4(32'hbb22eb39),
	.w5(32'hbb22b657),
	.w6(32'hbab7218d),
	.w7(32'hbb1f8f32),
	.w8(32'hbb3cabc9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad046ed),
	.w1(32'hbb9fdedd),
	.w2(32'hbc3071ae),
	.w3(32'h3cad1038),
	.w4(32'h3d37c541),
	.w5(32'h3cf356a5),
	.w6(32'h3cf96bcd),
	.w7(32'h3d69c4e2),
	.w8(32'h3d4d3135),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc201d),
	.w1(32'hbbf39271),
	.w2(32'hbc0f3b34),
	.w3(32'hbc0877e7),
	.w4(32'hbb89ea2a),
	.w5(32'hbb1904a1),
	.w6(32'hbbac0ee8),
	.w7(32'hba89cb0d),
	.w8(32'h3b07bb04),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb1bc),
	.w1(32'h3b39ee77),
	.w2(32'h3c2e678a),
	.w3(32'hbc151de8),
	.w4(32'hbc0ec978),
	.w5(32'hbbfd4418),
	.w6(32'hbb5006e6),
	.w7(32'hba3bf8af),
	.w8(32'hbb21b76e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ccbe1),
	.w1(32'h3c15e2da),
	.w2(32'hba143e9f),
	.w3(32'h3a775117),
	.w4(32'h3c66f4d7),
	.w5(32'h3d0118e4),
	.w6(32'h3caaebd8),
	.w7(32'h3d07b861),
	.w8(32'h3cc70bc4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4794a2),
	.w1(32'hbbe3e6e5),
	.w2(32'hbcd4848c),
	.w3(32'h3c713139),
	.w4(32'h3ca87290),
	.w5(32'h3c5c8b42),
	.w6(32'hbce62fa7),
	.w7(32'hbd6648a0),
	.w8(32'hbd23916d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc441db4),
	.w1(32'hbc60855b),
	.w2(32'hbc49f6a4),
	.w3(32'hbb4e919a),
	.w4(32'h3b629c90),
	.w5(32'h3b3e092d),
	.w6(32'hbc11f59b),
	.w7(32'hbbbd5383),
	.w8(32'hbbf1614d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f67de),
	.w1(32'h39c15599),
	.w2(32'h3b97e604),
	.w3(32'hbc371508),
	.w4(32'hbbb16f31),
	.w5(32'hbbad61de),
	.w6(32'h3ae48fe8),
	.w7(32'h3a931619),
	.w8(32'hbc45abf6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a992161),
	.w1(32'h3bf3a452),
	.w2(32'h3afaeb0d),
	.w3(32'hbad22fb1),
	.w4(32'h3c26935c),
	.w5(32'h3bace042),
	.w6(32'h3b545761),
	.w7(32'h3ba6162a),
	.w8(32'h3ad45817),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff5786),
	.w1(32'hbbb0f02b),
	.w2(32'h3be0bd71),
	.w3(32'hbbb192ea),
	.w4(32'h3b0a1353),
	.w5(32'hbbf6fc0f),
	.w6(32'hbb99e812),
	.w7(32'h3b8568fd),
	.w8(32'hbbaa5f57),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a1b0),
	.w1(32'hbb8b54f0),
	.w2(32'hbc356689),
	.w3(32'hbbbbcc94),
	.w4(32'hbc12a49e),
	.w5(32'hbbf36bc5),
	.w6(32'hbb11f338),
	.w7(32'h3a953828),
	.w8(32'hbb0a1326),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a34ba),
	.w1(32'hbae9a630),
	.w2(32'h3ab22abb),
	.w3(32'h3c16c184),
	.w4(32'h3c396179),
	.w5(32'h3ba53c7b),
	.w6(32'h3bcea0e7),
	.w7(32'h3c1bd9a1),
	.w8(32'hbaabd430),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00eea9),
	.w1(32'hb98243e9),
	.w2(32'h3b9aeed2),
	.w3(32'hba66ac68),
	.w4(32'hbb12d620),
	.w5(32'hbb39d3bb),
	.w6(32'h3b5a40ee),
	.w7(32'h3bd55c79),
	.w8(32'h3c00a8e9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d47f1),
	.w1(32'h3b3d77b2),
	.w2(32'h3c81c0d5),
	.w3(32'h3c8a2680),
	.w4(32'h3b771547),
	.w5(32'hbb3b1351),
	.w6(32'h3c4f7d77),
	.w7(32'h3be52aeb),
	.w8(32'h3c53ea11),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c872c36),
	.w1(32'hbc0772b6),
	.w2(32'hbba96671),
	.w3(32'h3a28570b),
	.w4(32'h3bdad5eb),
	.w5(32'h3bf1c3a9),
	.w6(32'hbb11ae4f),
	.w7(32'hb8e5bf7b),
	.w8(32'h39eaa3e8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a18ce),
	.w1(32'h3a0c36ed),
	.w2(32'hba1c8833),
	.w3(32'hb9aacd21),
	.w4(32'hbb13c837),
	.w5(32'hbb07c664),
	.w6(32'h39c600cf),
	.w7(32'hb9f1e051),
	.w8(32'hba65b7a0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b051ab),
	.w1(32'h3bbbd860),
	.w2(32'hbbd566bd),
	.w3(32'h3a983fb2),
	.w4(32'h3c0d6171),
	.w5(32'hbc2dfca8),
	.w6(32'hbb89815f),
	.w7(32'hbc08aff5),
	.w8(32'hbc5bae7e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e48cd),
	.w1(32'h3889a4d6),
	.w2(32'h3a773ed3),
	.w3(32'h3a5957e6),
	.w4(32'hba2969c7),
	.w5(32'hb9631a9e),
	.w6(32'h3a3e18ab),
	.w7(32'h39da168a),
	.w8(32'hbacc59a7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f901f),
	.w1(32'h3b311333),
	.w2(32'h3b52e535),
	.w3(32'h3add982a),
	.w4(32'h396bfe99),
	.w5(32'h3aff7774),
	.w6(32'h3b1bff86),
	.w7(32'hb9107fc9),
	.w8(32'h3b31b7d0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3c249),
	.w1(32'hbc640e14),
	.w2(32'hbc0675d1),
	.w3(32'hbc9fb50b),
	.w4(32'h3c1841be),
	.w5(32'h3c5a7a15),
	.w6(32'hbc52cd22),
	.w7(32'hbad2086f),
	.w8(32'h3b8bbd33),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8445),
	.w1(32'h3a893ba1),
	.w2(32'h3c2a9861),
	.w3(32'hbc297ef0),
	.w4(32'hbc6e20f6),
	.w5(32'hbc2b2f30),
	.w6(32'hbcf7473b),
	.w7(32'hbd5a9633),
	.w8(32'hbd415482),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a737b),
	.w1(32'h3ad1b09b),
	.w2(32'h3bbb863a),
	.w3(32'hbaba1c32),
	.w4(32'h3ab53d15),
	.w5(32'h3a344761),
	.w6(32'h3c61950e),
	.w7(32'h3c6a839e),
	.w8(32'h3caae421),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38284f14),
	.w1(32'hbbc4f676),
	.w2(32'hbc337c76),
	.w3(32'hbbc93447),
	.w4(32'hbb77b142),
	.w5(32'hbbb33d13),
	.w6(32'hbc3f7360),
	.w7(32'hbc4b212e),
	.w8(32'hbc7cda2f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0959d9),
	.w1(32'hb9d006be),
	.w2(32'hb9a5b8b3),
	.w3(32'hbb9123e4),
	.w4(32'hbbd2dcf0),
	.w5(32'h3b1316d6),
	.w6(32'h3c716f6a),
	.w7(32'h3ca9ce08),
	.w8(32'h3c96a3a1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c8c18),
	.w1(32'h3bc84531),
	.w2(32'h3c1239f2),
	.w3(32'h3a2cf9f1),
	.w4(32'hba931b20),
	.w5(32'hbaf06bde),
	.w6(32'h3b37f632),
	.w7(32'h3b411902),
	.w8(32'h3a643c7e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84bd8c),
	.w1(32'h3b537397),
	.w2(32'hbac07573),
	.w3(32'h3b085669),
	.w4(32'hbb34a57f),
	.w5(32'hbb2178b7),
	.w6(32'h3b3564ce),
	.w7(32'hbaf85078),
	.w8(32'hbabbe599),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be3d9a),
	.w1(32'hbc202278),
	.w2(32'h3afb8e0d),
	.w3(32'hbbe544d0),
	.w4(32'hbc2f6d7b),
	.w5(32'hbbe387b4),
	.w6(32'hbc8a103e),
	.w7(32'hbcae9f78),
	.w8(32'hbc8784cb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33221f),
	.w1(32'h3cce9839),
	.w2(32'h3d3cc9de),
	.w3(32'hbd58bca8),
	.w4(32'hbd992c9b),
	.w5(32'hbd804a08),
	.w6(32'h3c6a1585),
	.w7(32'h3c3f629b),
	.w8(32'h3c7d6f04),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f333a),
	.w1(32'hbb9fa9c5),
	.w2(32'hbbb0274a),
	.w3(32'h3c756b8e),
	.w4(32'h3bdaabab),
	.w5(32'hbabc4783),
	.w6(32'h3c83f789),
	.w7(32'h3c8dddeb),
	.w8(32'h3c49cafd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97daf55),
	.w1(32'hbc575647),
	.w2(32'h3bc22595),
	.w3(32'hbb17183b),
	.w4(32'hbb8858e1),
	.w5(32'hbc16b8cb),
	.w6(32'hbbf1254a),
	.w7(32'hbc3b5837),
	.w8(32'hbc18195d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90eeb52),
	.w1(32'hbc529c02),
	.w2(32'hbc023d9d),
	.w3(32'hba9f486c),
	.w4(32'hb8f40a5a),
	.w5(32'hbbf1379f),
	.w6(32'h38096efa),
	.w7(32'hbba1ce66),
	.w8(32'hbc8c3fc7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ac4ca),
	.w1(32'hbc4c3950),
	.w2(32'hbc6be340),
	.w3(32'hbad511ae),
	.w4(32'h39c84217),
	.w5(32'h3b9602e4),
	.w6(32'hbbc4d26f),
	.w7(32'hbbd7883d),
	.w8(32'hbab3e490),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfac302),
	.w1(32'hbabdcf59),
	.w2(32'hbb87ee70),
	.w3(32'hbb9387b4),
	.w4(32'h3aa3d811),
	.w5(32'h3c020378),
	.w6(32'hbb9775a5),
	.w7(32'hbba560d6),
	.w8(32'h3bd05ec5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4de2d),
	.w1(32'h3a5e3593),
	.w2(32'h3b066013),
	.w3(32'hbad4aaa8),
	.w4(32'h3b8163fd),
	.w5(32'hbac5dc4d),
	.w6(32'h3b0f2586),
	.w7(32'h3c323eb9),
	.w8(32'h3b905bea),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba177e1c),
	.w1(32'h3a0dfa7b),
	.w2(32'hb84ec0ee),
	.w3(32'h3a8b2f65),
	.w4(32'hb99b22c6),
	.w5(32'h3969054f),
	.w6(32'hba14375d),
	.w7(32'hbb214744),
	.w8(32'hba9258d7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4c214),
	.w1(32'h39f98ec3),
	.w2(32'h39eccec5),
	.w3(32'hbc83d219),
	.w4(32'hbce1a1d5),
	.w5(32'hbc7542ba),
	.w6(32'hbb8de8d9),
	.w7(32'hbc547044),
	.w8(32'hbc669884),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b15c03),
	.w1(32'hbb84fb61),
	.w2(32'hbb54ab08),
	.w3(32'h3c8676f9),
	.w4(32'h3c572649),
	.w5(32'h3b2d9403),
	.w6(32'h3b12a5e1),
	.w7(32'h3b5f1bb6),
	.w8(32'h3bbea7ee),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a1aca),
	.w1(32'h3c31b06b),
	.w2(32'hbb8dac75),
	.w3(32'h3abda8d2),
	.w4(32'hbc31298f),
	.w5(32'hbc5a236e),
	.w6(32'hbbc86e58),
	.w7(32'hbcc69d1c),
	.w8(32'hbd219241),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc867037),
	.w1(32'h3a83af60),
	.w2(32'h3b614541),
	.w3(32'hbaf333b6),
	.w4(32'hba897813),
	.w5(32'hba5e10f8),
	.w6(32'hba84968a),
	.w7(32'hb9375177),
	.w8(32'h39563e87),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3ad4),
	.w1(32'h3b3008aa),
	.w2(32'h3ac7756d),
	.w3(32'h3b85dd8b),
	.w4(32'h3c7171c9),
	.w5(32'h3c8815a9),
	.w6(32'h3a83593c),
	.w7(32'h3b82568c),
	.w8(32'h3bc7640f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b166c9d),
	.w1(32'h3bd5751a),
	.w2(32'h3afead9f),
	.w3(32'h3bde6302),
	.w4(32'h3bee7d29),
	.w5(32'hbb3d973a),
	.w6(32'h3cabe119),
	.w7(32'h3cd83a19),
	.w8(32'h3c63a09c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06d79a),
	.w1(32'hba598e9b),
	.w2(32'hba5a15fc),
	.w3(32'h3b71d863),
	.w4(32'h3b8e05bd),
	.w5(32'h3bacc761),
	.w6(32'hbaa49208),
	.w7(32'hbb13c513),
	.w8(32'hbb108f53),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a388a8),
	.w1(32'hbc019314),
	.w2(32'hbcc213b1),
	.w3(32'hbbb91024),
	.w4(32'h397553a9),
	.w5(32'hbbd26de0),
	.w6(32'hbca45fc7),
	.w7(32'hbc3b8b3d),
	.w8(32'hbc595326),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47a0cd),
	.w1(32'h3a3924e3),
	.w2(32'h3c6750b4),
	.w3(32'hbaf11aac),
	.w4(32'hbb15b2ea),
	.w5(32'hbc44cbf8),
	.w6(32'hbb333bc5),
	.w7(32'hbc42334d),
	.w8(32'hbc70334c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c361e98),
	.w1(32'hbb8beeb2),
	.w2(32'hbbec4165),
	.w3(32'h3b067327),
	.w4(32'h3b213d5f),
	.w5(32'h3b466c32),
	.w6(32'hbbc8da71),
	.w7(32'hbc90dad2),
	.w8(32'hbc44fc3c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbca362),
	.w1(32'h3b626e9f),
	.w2(32'h3b15a181),
	.w3(32'hbaea134e),
	.w4(32'hbb7f11ea),
	.w5(32'hbb32f7ad),
	.w6(32'hbb1a08e9),
	.w7(32'hbb7a704a),
	.w8(32'hbb86f89b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b541c0c),
	.w1(32'h3c25d52f),
	.w2(32'h3c542d9a),
	.w3(32'hbcfa35bc),
	.w4(32'hbd02ad11),
	.w5(32'hbcfa51df),
	.w6(32'h3c86ec5f),
	.w7(32'h3d157dfc),
	.w8(32'h3d2a1bbb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8485e8),
	.w1(32'h3b838004),
	.w2(32'h3c421088),
	.w3(32'hb9a9f697),
	.w4(32'h3a783c62),
	.w5(32'hbafc3e65),
	.w6(32'h3a5c4bfc),
	.w7(32'h3a900627),
	.w8(32'hbb992ef2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd38d2),
	.w1(32'hbb848a20),
	.w2(32'h397c01dd),
	.w3(32'hbc2196ea),
	.w4(32'hbbe9f34a),
	.w5(32'h3b4da86b),
	.w6(32'hbc39de06),
	.w7(32'hbbb9277b),
	.w8(32'hba75c7c7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b255f8),
	.w1(32'h3bdad5bc),
	.w2(32'h3c23431c),
	.w3(32'hbb52bd99),
	.w4(32'hbc0f3059),
	.w5(32'hbb9ead45),
	.w6(32'hba714667),
	.w7(32'hbb939213),
	.w8(32'hba9f5e54),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bfcd1),
	.w1(32'h3bcea416),
	.w2(32'h3c70a141),
	.w3(32'hbc243908),
	.w4(32'hbc087b37),
	.w5(32'hbbe2779e),
	.w6(32'hbb93179c),
	.w7(32'hbb13369a),
	.w8(32'h3a12d5ad),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c854fd5),
	.w1(32'h3929676b),
	.w2(32'h3ba45e21),
	.w3(32'hbb0a3f86),
	.w4(32'hbb0f3656),
	.w5(32'hbb580deb),
	.w6(32'hbbe10fb2),
	.w7(32'hbc57c112),
	.w8(32'hbc7d02a1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf41ea),
	.w1(32'hbc7cb4b1),
	.w2(32'hbc900b63),
	.w3(32'h3c652f73),
	.w4(32'h3c8b2eaa),
	.w5(32'h3cb36de8),
	.w6(32'hb95c72b3),
	.w7(32'h3ad92e5e),
	.w8(32'h3c4fd666),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c1d45),
	.w1(32'h3b728d7f),
	.w2(32'h3b815910),
	.w3(32'h3bfa9067),
	.w4(32'h3bde67a1),
	.w5(32'h3bbbb2b0),
	.w6(32'h3bc39c15),
	.w7(32'h3b6f8279),
	.w8(32'h3b762b0b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78ac71),
	.w1(32'hbac223ce),
	.w2(32'hbc850f7b),
	.w3(32'hbba0b6b3),
	.w4(32'h3995f274),
	.w5(32'h3cbc91e7),
	.w6(32'hbbe3c5d6),
	.w7(32'hbd191d87),
	.w8(32'hbcb8b1a9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc758dc),
	.w1(32'h3a55afda),
	.w2(32'h394b8af3),
	.w3(32'hbb8807d4),
	.w4(32'hbbc40ada),
	.w5(32'hbba34d7d),
	.w6(32'hba8f3dfb),
	.w7(32'hba843827),
	.w8(32'hba528055),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e043f5),
	.w1(32'h3a13097b),
	.w2(32'hb9ea6481),
	.w3(32'h3b612d0d),
	.w4(32'h3c311330),
	.w5(32'h3c13a86b),
	.w6(32'hbc284902),
	.w7(32'hbc978a49),
	.w8(32'hbca0a673),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc120367),
	.w1(32'hbb61f1e0),
	.w2(32'h3b242036),
	.w3(32'hbc02c92d),
	.w4(32'hbc0d4a3f),
	.w5(32'hbc319355),
	.w6(32'hbb9a88f8),
	.w7(32'hbb127c38),
	.w8(32'hbc2c2901),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba875fab),
	.w1(32'hb985cf92),
	.w2(32'h3c740d08),
	.w3(32'h3b857fe1),
	.w4(32'h3c4889d4),
	.w5(32'h3b7d2547),
	.w6(32'h3b6acad9),
	.w7(32'hbbbf9d95),
	.w8(32'hbbe860f3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e301),
	.w1(32'hbc9532b6),
	.w2(32'hbcb2f8a5),
	.w3(32'h3b2aa215),
	.w4(32'hbc3e869b),
	.w5(32'hbcd2f623),
	.w6(32'h3c961017),
	.w7(32'h3d428850),
	.w8(32'h3ceb2c43),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19fae1),
	.w1(32'h399af1e4),
	.w2(32'hbb66b67d),
	.w3(32'h3b1c7f44),
	.w4(32'hbc2594c5),
	.w5(32'hbc90a5a8),
	.w6(32'h3b367ea9),
	.w7(32'hb9d0e92e),
	.w8(32'hbb21ac9d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule