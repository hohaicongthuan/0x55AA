module layer_10_featuremap_78(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32e5d9),
	.w1(32'hbb90b01a),
	.w2(32'hba14334a),
	.w3(32'hbc9bacce),
	.w4(32'hbc3779e1),
	.w5(32'hbbcfee3b),
	.w6(32'hbc7504cb),
	.w7(32'h3ae10262),
	.w8(32'hbc399e9f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d094f),
	.w1(32'hbc276fd2),
	.w2(32'hbc4bf80b),
	.w3(32'hbc80d92e),
	.w4(32'hbbb36f6a),
	.w5(32'hbc102dd2),
	.w6(32'hbb627cc0),
	.w7(32'h3b59c33b),
	.w8(32'hbc06091d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e3021),
	.w1(32'h3baf5818),
	.w2(32'h3bd23959),
	.w3(32'h3b6cb23e),
	.w4(32'hbab970ec),
	.w5(32'h3bc1b30d),
	.w6(32'hbbb0c3b5),
	.w7(32'hb9cb92a4),
	.w8(32'hbbc99d8a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49c2d2),
	.w1(32'h3c050360),
	.w2(32'h39213903),
	.w3(32'h3b953c45),
	.w4(32'h3bfe1a49),
	.w5(32'hbb775355),
	.w6(32'h3b04db6e),
	.w7(32'h3aa3a4e7),
	.w8(32'hbb4b65c8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a4fe7),
	.w1(32'h3b708804),
	.w2(32'h3ba5c52c),
	.w3(32'h3b62bfb6),
	.w4(32'h3bbfb469),
	.w5(32'h38ef1cfd),
	.w6(32'h3bfd474b),
	.w7(32'h3c6dccae),
	.w8(32'hbba8f897),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05138a),
	.w1(32'hbc033efb),
	.w2(32'hb9a4a564),
	.w3(32'hbc4c3092),
	.w4(32'hbc036307),
	.w5(32'hb9fae9d3),
	.w6(32'hbc1489f1),
	.w7(32'hbbd9a011),
	.w8(32'hba18c181),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb218fc6),
	.w1(32'hbb3a87af),
	.w2(32'hbb9c2ca1),
	.w3(32'hbaf1d576),
	.w4(32'hbaebd298),
	.w5(32'h3ae10199),
	.w6(32'hba65e468),
	.w7(32'h3aa763c4),
	.w8(32'hbb6b00d6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b127162),
	.w1(32'h3b8562a3),
	.w2(32'h3bbb3d3a),
	.w3(32'h3b84e92b),
	.w4(32'h3bd7f240),
	.w5(32'hbb621bb3),
	.w6(32'h3adfc704),
	.w7(32'h3bface0b),
	.w8(32'hbaa505c4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07881e),
	.w1(32'h3a34b10f),
	.w2(32'hbc8b5fae),
	.w3(32'hbc03d7b9),
	.w4(32'hb99019e0),
	.w5(32'hbb81e2ed),
	.w6(32'hbb92067e),
	.w7(32'h3bdcbdb9),
	.w8(32'hb9f37976),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e73ac),
	.w1(32'h3a869874),
	.w2(32'h3a681cec),
	.w3(32'h3b8e1632),
	.w4(32'hbb020295),
	.w5(32'h39067ac3),
	.w6(32'hbb5faead),
	.w7(32'hbc3af706),
	.w8(32'h3a1d0c8b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b608d),
	.w1(32'h3a6ec438),
	.w2(32'h3bda62e4),
	.w3(32'h3b2685b8),
	.w4(32'h3b937cc3),
	.w5(32'h3bcfef4c),
	.w6(32'h3b72b669),
	.w7(32'h3b65d5f1),
	.w8(32'h3bee2b88),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1bb10),
	.w1(32'hbb5c3ae2),
	.w2(32'h3b0ddf52),
	.w3(32'h3bc0b8a1),
	.w4(32'hba95cf1c),
	.w5(32'hb9a1a93d),
	.w6(32'h3a8fff27),
	.w7(32'h3c0a393b),
	.w8(32'h3adc5795),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb838ea58),
	.w1(32'h3b13d596),
	.w2(32'h3b86431d),
	.w3(32'h3b194253),
	.w4(32'h3a64ec1b),
	.w5(32'h39f7e2fe),
	.w6(32'h3aeeab5b),
	.w7(32'h3981130a),
	.w8(32'hba34853a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a884854),
	.w1(32'hbb1f3f75),
	.w2(32'hbb2ecea0),
	.w3(32'hbb783ada),
	.w4(32'hba924d48),
	.w5(32'hbc5ef5cb),
	.w6(32'hbb5ac159),
	.w7(32'hbade836a),
	.w8(32'hbb6e4219),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc325b9e),
	.w1(32'hbbc188a3),
	.w2(32'h3b23edf3),
	.w3(32'hbc32b63e),
	.w4(32'h3b9757aa),
	.w5(32'hbabf1e6e),
	.w6(32'h3ae9f825),
	.w7(32'h3c2d4aa0),
	.w8(32'h3a9a97ed),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ffa5d),
	.w1(32'h3b31cd5b),
	.w2(32'h3aa2fc02),
	.w3(32'hbb70434f),
	.w4(32'hba6875b4),
	.w5(32'hb9bef030),
	.w6(32'hbb5b4a22),
	.w7(32'h3b7ce5a9),
	.w8(32'h3800d62b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2198b2),
	.w1(32'h3aa08e11),
	.w2(32'hb8f3c229),
	.w3(32'h3a0039ea),
	.w4(32'h3b5afb72),
	.w5(32'h3b001a95),
	.w6(32'h3af08efd),
	.w7(32'h3afc7d27),
	.w8(32'h3b364706),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd1b3f),
	.w1(32'h3ba9d54a),
	.w2(32'hbb95ad96),
	.w3(32'h3bcb7985),
	.w4(32'h3bba1749),
	.w5(32'hbb07c45b),
	.w6(32'h3b335d4d),
	.w7(32'h3bd4c7ec),
	.w8(32'h3a12b94e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ef3c6),
	.w1(32'h3abadf48),
	.w2(32'hbb8007a5),
	.w3(32'h3ae5157c),
	.w4(32'hbb81b590),
	.w5(32'hbc944620),
	.w6(32'h3b3aba41),
	.w7(32'hba42a3e2),
	.w8(32'hbc851c2b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc91dbb),
	.w1(32'hbca2e4ba),
	.w2(32'h3b9a6928),
	.w3(32'hbd105a1e),
	.w4(32'hbcb4b23f),
	.w5(32'h3bbb7fbd),
	.w6(32'hbcb8b40d),
	.w7(32'hbc89f880),
	.w8(32'hb9cdbd5d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb71ccb),
	.w1(32'h3b8cce49),
	.w2(32'h3b357519),
	.w3(32'h3a1630b2),
	.w4(32'h3b64489c),
	.w5(32'h3ae9190f),
	.w6(32'hba8eafad),
	.w7(32'h3ac317c1),
	.w8(32'hbb27b79f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b565b93),
	.w1(32'h3c3ec2bf),
	.w2(32'h3b5d5d03),
	.w3(32'h3b80868a),
	.w4(32'h3c45a9a1),
	.w5(32'hbbf52e41),
	.w6(32'h3937019c),
	.w7(32'h3c06a8d6),
	.w8(32'hbbb5ff60),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5153b3),
	.w1(32'hbbfb8e6d),
	.w2(32'h3ac2e3e0),
	.w3(32'hbc1b55cc),
	.w4(32'hbc2278f2),
	.w5(32'h3a970855),
	.w6(32'hbc290bfa),
	.w7(32'hb88cc8b9),
	.w8(32'h3a3167c0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936c53c),
	.w1(32'hba189042),
	.w2(32'h3a29425d),
	.w3(32'h3b1e703f),
	.w4(32'h3ad191f6),
	.w5(32'hbb2a2fd0),
	.w6(32'hba95044e),
	.w7(32'h39d7e89b),
	.w8(32'hbb938adb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b583f01),
	.w1(32'h3a2bd6e5),
	.w2(32'hbc66c569),
	.w3(32'h39891bbb),
	.w4(32'hbbacdfd3),
	.w5(32'hbcca1948),
	.w6(32'h3afe6e52),
	.w7(32'h3b557f86),
	.w8(32'hbc57a6bf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb883fc),
	.w1(32'hbc390258),
	.w2(32'h3b4e3e75),
	.w3(32'hbcd80682),
	.w4(32'hbc7b70cd),
	.w5(32'hb9368e25),
	.w6(32'hbca50f5c),
	.w7(32'h3ad9a5f9),
	.w8(32'hbb7f67c2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40fe2c),
	.w1(32'hbb92fdcd),
	.w2(32'hbf50ba79),
	.w3(32'hbc0abeb2),
	.w4(32'h3b5cdc98),
	.w5(32'h3e361744),
	.w6(32'hba6f066f),
	.w7(32'h3c290cf8),
	.w8(32'hbe9d2d74),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9159fc),
	.w1(32'hbe8bc15a),
	.w2(32'h3e9187ac),
	.w3(32'hbf32cea6),
	.w4(32'h3eda3a13),
	.w5(32'hbe1c4503),
	.w6(32'hbf808355),
	.w7(32'hbde3d60b),
	.w8(32'h3f60cf1c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbefd627a),
	.w1(32'h3f23b3b8),
	.w2(32'hbfa63c47),
	.w3(32'hbe150aba),
	.w4(32'hbf4da74b),
	.w5(32'h3e766a88),
	.w6(32'hbedcdf8c),
	.w7(32'hbda165be),
	.w8(32'hbeedbc47),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe3d4f28),
	.w1(32'hbf8b1f00),
	.w2(32'hbf4ec090),
	.w3(32'hbf851260),
	.w4(32'h3e523d9e),
	.w5(32'hbe98b1e9),
	.w6(32'hbf8a76d0),
	.w7(32'hbea6e3e1),
	.w8(32'hbee59a71),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf81d812),
	.w1(32'hbf0ca50e),
	.w2(32'h3ecdb5d0),
	.w3(32'hbf99205d),
	.w4(32'hbf494c10),
	.w5(32'hbf032d33),
	.w6(32'hbf157e0a),
	.w7(32'hbf8e8931),
	.w8(32'h3caa2653),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3e27d),
	.w1(32'hbf93d002),
	.w2(32'h3fec909e),
	.w3(32'h3df88f76),
	.w4(32'hbf49d577),
	.w5(32'h3e56268a),
	.w6(32'hbeb070fa),
	.w7(32'hbf0c645c),
	.w8(32'hbccd31d4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf4cc706),
	.w1(32'h3e6d3726),
	.w2(32'h3cb0edf2),
	.w3(32'hbf935387),
	.w4(32'h3d54aa47),
	.w5(32'hbe97ece1),
	.w6(32'hbed9ee17),
	.w7(32'hbe705c44),
	.w8(32'hbf16573a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf9d6198),
	.w1(32'hbe577ead),
	.w2(32'h3d8697ee),
	.w3(32'hbf40999d),
	.w4(32'h3e0bc92f),
	.w5(32'hbf9e8d1e),
	.w6(32'hbe403bf3),
	.w7(32'hbf3db7b2),
	.w8(32'h3f9348ca),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe724534),
	.w1(32'hbf933cdf),
	.w2(32'h3de34846),
	.w3(32'hbe92e162),
	.w4(32'hbda94c05),
	.w5(32'h3cb624c0),
	.w6(32'hbf8ff874),
	.w7(32'h3edb9c51),
	.w8(32'h3de2398a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf25ca2f),
	.w1(32'h3f47f896),
	.w2(32'hbf6d72f2),
	.w3(32'hbebcae04),
	.w4(32'hbf654890),
	.w5(32'hbf8a743b),
	.w6(32'hbf59340f),
	.w7(32'hbf5453ac),
	.w8(32'hbf440ab3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec969c1),
	.w1(32'hbf1b0575),
	.w2(32'hbf01e3ea),
	.w3(32'hbef4aa6c),
	.w4(32'hbe9d3e69),
	.w5(32'hbf58415e),
	.w6(32'hbfa4f934),
	.w7(32'hbf14c80b),
	.w8(32'hbf1f8e52),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3eb80994),
	.w1(32'hbf3b6718),
	.w2(32'hbf0add51),
	.w3(32'h3c7da216),
	.w4(32'hbe1a8247),
	.w5(32'hbf79e1c4),
	.w6(32'hbf7b5b39),
	.w7(32'hbf9986e9),
	.w8(32'h3c777157),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf6a4e9c),
	.w1(32'h3abac90e),
	.w2(32'hbf61a566),
	.w3(32'hbf785072),
	.w4(32'h3f19606c),
	.w5(32'hbf690f98),
	.w6(32'h3f972293),
	.w7(32'hbe6fd75e),
	.w8(32'h3f19b7d2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe76eb24),
	.w1(32'h3d750ade),
	.w2(32'h3f62ff07),
	.w3(32'h3d32aad2),
	.w4(32'hbf32bda9),
	.w5(32'h3e95848e),
	.w6(32'hbe99cf8a),
	.w7(32'hbee230e8),
	.w8(32'h3ece90ec),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe400621),
	.w1(32'hbea6fd6a),
	.w2(32'h3e33de3d),
	.w3(32'hbf28c863),
	.w4(32'h3e42cc2a),
	.w5(32'hbf6c139c),
	.w6(32'hbeff17c8),
	.w7(32'hbf0cdd7b),
	.w8(32'h3f35f3f8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e979562),
	.w1(32'h3f28065d),
	.w2(32'h3ecb5e90),
	.w3(32'h3f8df5b3),
	.w4(32'h3f9c0827),
	.w5(32'h3f121319),
	.w6(32'h3eff145d),
	.w7(32'h3f5bec07),
	.w8(32'h3ea0cfb7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ebe954a),
	.w1(32'h3f2a9515),
	.w2(32'h3fb0410c),
	.w3(32'h3ee5fcfb),
	.w4(32'h3edfbe8b),
	.w5(32'h3eb30998),
	.w6(32'h3f3e2ea9),
	.w7(32'h3f151f13),
	.w8(32'h3f9090b9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f0dc336),
	.w1(32'h3f53e705),
	.w2(32'h3ea18891),
	.w3(32'h3eff0d00),
	.w4(32'h3fa8268d),
	.w5(32'h3f0c8a03),
	.w6(32'h3eb027be),
	.w7(32'h3f765e3f),
	.w8(32'h3f4f18a1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ecc4184),
	.w1(32'h3f847bb5),
	.w2(32'h3f4afd26),
	.w3(32'h3f170448),
	.w4(32'h3ef83412),
	.w5(32'h3f8762bb),
	.w6(32'h3f61c890),
	.w7(32'h3ef86200),
	.w8(32'h3f041b87),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3efe558b),
	.w1(32'h3e98105c),
	.w2(32'h3f37e99a),
	.w3(32'h3f0d1d94),
	.w4(32'h3f020599),
	.w5(32'h3f031a5a),
	.w6(32'h3ee8a0df),
	.w7(32'h3f81f0a3),
	.w8(32'h3f0371e8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f0de608),
	.w1(32'h3f7523bf),
	.w2(32'h3f069cbf),
	.w3(32'h3ef3c291),
	.w4(32'h3ee8d9f0),
	.w5(32'h3f9176c2),
	.w6(32'h3fb396a2),
	.w7(32'h3ea16f7b),
	.w8(32'h3f1a66a4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3744b5),
	.w1(32'h3f544dc4),
	.w2(32'h3e9ce704),
	.w3(32'h3f1e812e),
	.w4(32'h3f5a6054),
	.w5(32'h3f4a2bcb),
	.w6(32'h3f90994e),
	.w7(32'h3f10b179),
	.w8(32'h3eaf2ec7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f94607e),
	.w1(32'h3f35d66d),
	.w2(32'h3ec8b89f),
	.w3(32'h3ebb8fbd),
	.w4(32'h3f7f1b34),
	.w5(32'h3f17a94d),
	.w6(32'h3ec9908b),
	.w7(32'h3f7b3e42),
	.w8(32'h3ee3738f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ea139c8),
	.w1(32'h3f17de25),
	.w2(32'h3f5c919a),
	.w3(32'h3e8c2ef0),
	.w4(32'h3fa9f085),
	.w5(32'h3f4c040e),
	.w6(32'h3f1b5c96),
	.w7(32'h3eb0093b),
	.w8(32'h3f42e466),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f776895),
	.w1(32'h3f23707b),
	.w2(32'h3f18c027),
	.w3(32'h3f3e32a8),
	.w4(32'h3f938a12),
	.w5(32'h3eef56cb),
	.w6(32'h3f023d9a),
	.w7(32'h3f2ad404),
	.w8(32'h3f198c24),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2a5ed4),
	.w1(32'h3ef16f7c),
	.w2(32'h3f23d18e),
	.w3(32'h3f06a7e9),
	.w4(32'h3f61497c),
	.w5(32'h3f8487e6),
	.w6(32'h3edea897),
	.w7(32'h3f21ef2d),
	.w8(32'h3f41ff51),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f6e23b7),
	.w1(32'h3fc02d86),
	.w2(32'h3e80ffa2),
	.w3(32'h3f0668b2),
	.w4(32'h3f06a9a7),
	.w5(32'h3eba7d29),
	.w6(32'h3f9dda71),
	.w7(32'h3eb67de4),
	.w8(32'h3f3dfbf4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f38ac4e),
	.w1(32'h3eb9c344),
	.w2(32'h3f348b2f),
	.w3(32'h3e91d4a7),
	.w4(32'h3f836ada),
	.w5(32'h3f2eadfc),
	.w6(32'h3f29f324),
	.w7(32'h3eb6af1c),
	.w8(32'h3ec75c2a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e818892),
	.w1(32'h3f44b318),
	.w2(32'h3ea30df5),
	.w3(32'h3e86a177),
	.w4(32'h3f2d9a23),
	.w5(32'h3f9c580b),
	.w6(32'h3f32ca1b),
	.w7(32'h3f08b2bf),
	.w8(32'h3f2baf13),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f404d6c),
	.w1(32'hbe6e9100),
	.w2(32'h3d808f83),
	.w3(32'h3d9424d1),
	.w4(32'h3df813b4),
	.w5(32'hbe42f4bb),
	.w6(32'h3d933896),
	.w7(32'h3e1d3309),
	.w8(32'h3dd675ac),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db70d6f),
	.w1(32'h3e161915),
	.w2(32'hbc2ab0cb),
	.w3(32'hbd8e9bae),
	.w4(32'h3e5dd56f),
	.w5(32'hbe4d9a27),
	.w6(32'h3d67608c),
	.w7(32'hbd60edb1),
	.w8(32'hbe0790dd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9836b0),
	.w1(32'h3dffc901),
	.w2(32'h3e13263b),
	.w3(32'h3d9e292f),
	.w4(32'h3d83bfdb),
	.w5(32'hbcc04b1f),
	.w6(32'h3d2043e9),
	.w7(32'h3d86a78f),
	.w8(32'hbc778dbc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d97da67),
	.w1(32'hbc98eca9),
	.w2(32'hbc84b8b2),
	.w3(32'h3d2da8b8),
	.w4(32'h3e85407d),
	.w5(32'h3ce1b380),
	.w6(32'h3bfb844b),
	.w7(32'h3d3dd0ed),
	.w8(32'h3e1ab322),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84a21d),
	.w1(32'h3db3ab2d),
	.w2(32'h3d303e87),
	.w3(32'h3e4e9d5b),
	.w4(32'h3dc4300a),
	.w5(32'h3d2b6068),
	.w6(32'h3d4224f5),
	.w7(32'h3c554644),
	.w8(32'h3e730b67),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce9c483),
	.w1(32'hbdd0697d),
	.w2(32'h3d9945b4),
	.w3(32'h3da40270),
	.w4(32'hbe19db30),
	.w5(32'hbe16c8f5),
	.w6(32'hbe680f4d),
	.w7(32'h3d86075c),
	.w8(32'hbe7dcdcc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe0a5ecd),
	.w1(32'h3d76d535),
	.w2(32'hbdde1684),
	.w3(32'h3e143291),
	.w4(32'h3e01a4a6),
	.w5(32'h3dd17e96),
	.w6(32'hbd2787c5),
	.w7(32'hbe215498),
	.w8(32'h3c3892d3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ddce52d),
	.w1(32'h3dd27489),
	.w2(32'h3e181547),
	.w3(32'hbda41f9a),
	.w4(32'h3d1e1e59),
	.w5(32'h3d1a5cfe),
	.w6(32'h3e3f7ef9),
	.w7(32'hbdd42d60),
	.w8(32'h3cf6fc76),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec6d492),
	.w1(32'h3c6a2da4),
	.w2(32'h3d15ef54),
	.w3(32'h3e285395),
	.w4(32'h3cee4218),
	.w5(32'hbdc4630a),
	.w6(32'hbaa4ccb4),
	.w7(32'h3d3615a0),
	.w8(32'h3e148549),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb55bbe),
	.w1(32'h3d5a5e84),
	.w2(32'hbaa53708),
	.w3(32'h3ceb1e1a),
	.w4(32'h3db278cf),
	.w5(32'h3d02cf63),
	.w6(32'hbc047fca),
	.w7(32'hbcf84ae4),
	.w8(32'hbde220fa),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96ce1d),
	.w1(32'h3cd563fc),
	.w2(32'h3cab367d),
	.w3(32'h3dd75295),
	.w4(32'hbd3b83ac),
	.w5(32'h3dc09f2d),
	.w6(32'h3afc8fa9),
	.w7(32'h3d70e813),
	.w8(32'hbd8fedd5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c410a72),
	.w1(32'h3c87d0d1),
	.w2(32'hbe218407),
	.w3(32'h3e1150de),
	.w4(32'h3db04dd5),
	.w5(32'h3b0ad861),
	.w6(32'h3e02e6d8),
	.w7(32'hbe8e9651),
	.w8(32'hbd5df740),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0fe3d5),
	.w1(32'hbdb26585),
	.w2(32'h3b1dbd3f),
	.w3(32'h3dddfb50),
	.w4(32'hbe57b32d),
	.w5(32'h3d397a93),
	.w6(32'h3d242014),
	.w7(32'hbb73c9ef),
	.w8(32'h3d22661d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe08a54b),
	.w1(32'h3a82bafd),
	.w2(32'h39e3b700),
	.w3(32'hbddd1e77),
	.w4(32'hbdf8c8c5),
	.w5(32'h3d84b601),
	.w6(32'hbcacd800),
	.w7(32'hbbbb04ff),
	.w8(32'hbc9f28a6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe7a9551),
	.w1(32'h3c6cc102),
	.w2(32'h3ce1002c),
	.w3(32'h3da05ba9),
	.w4(32'h3c9fee7a),
	.w5(32'h3c2476af),
	.w6(32'h3d0771bb),
	.w7(32'h3cf61ef1),
	.w8(32'h3cae418a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c875660),
	.w1(32'h3d01c483),
	.w2(32'h3bf2d6af),
	.w3(32'h3d1513a7),
	.w4(32'h3bf7e2b7),
	.w5(32'h3cc85e89),
	.w6(32'h3d15b068),
	.w7(32'h3d9d572e),
	.w8(32'h3bef7bd4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dbaae3c),
	.w1(32'h3c0184b0),
	.w2(32'h3bb80275),
	.w3(32'h3cfa40b9),
	.w4(32'h3d8d0803),
	.w5(32'h3c9ab84a),
	.w6(32'h3c01b57e),
	.w7(32'h3c03f44c),
	.w8(32'h3d16ebe7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b8b44),
	.w1(32'h3c1c9dcc),
	.w2(32'h3c88eb8e),
	.w3(32'h3ced32dc),
	.w4(32'h3bd45bba),
	.w5(32'h3bbe594d),
	.w6(32'h3bd67e0d),
	.w7(32'h3c287805),
	.w8(32'h3bdb0bda),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f6cb),
	.w1(32'h3d8476e9),
	.w2(32'h3ce506c5),
	.w3(32'h3c3538d8),
	.w4(32'h3bd80c49),
	.w5(32'h3ca28f45),
	.w6(32'h3c706bed),
	.w7(32'h3d0e10bf),
	.w8(32'h3c59a0ce),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1084a),
	.w1(32'h3def3340),
	.w2(32'h3d0878c4),
	.w3(32'h3bc43c35),
	.w4(32'h3d62a9a8),
	.w5(32'h3c494038),
	.w6(32'h3c0fcb1b),
	.w7(32'h3cdbecc4),
	.w8(32'h3bfcacbe),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf53dd9),
	.w1(32'h3d079d5d),
	.w2(32'h3c0d79f5),
	.w3(32'h3d47eadf),
	.w4(32'h3c8ae4e5),
	.w5(32'h3c772a03),
	.w6(32'h3d25474e),
	.w7(32'h3bd1a918),
	.w8(32'h3cf09a0d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd37072),
	.w1(32'h3c8239c1),
	.w2(32'h3c0dd2a1),
	.w3(32'h3cbb95b0),
	.w4(32'h3ca37058),
	.w5(32'h3c908579),
	.w6(32'h3ca78bfb),
	.w7(32'h3d6f41c2),
	.w8(32'h3b9cc834),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13f234),
	.w1(32'h3d12d196),
	.w2(32'h3c3dec92),
	.w3(32'h3c16f53f),
	.w4(32'h3c563fa3),
	.w5(32'h3c823379),
	.w6(32'h3da13743),
	.w7(32'h3c87feb4),
	.w8(32'h3d0f8c44),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d39c807),
	.w1(32'h3c8b58db),
	.w2(32'h3ba13029),
	.w3(32'h3c7c7552),
	.w4(32'h3bf52fc5),
	.w5(32'h3c8b882f),
	.w6(32'h3c1226c3),
	.w7(32'h3bdb6dee),
	.w8(32'h3c0e7344),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be475f8),
	.w1(32'h3c03ad13),
	.w2(32'h3d2ba56f),
	.w3(32'h3ca9c864),
	.w4(32'h3c5c818c),
	.w5(32'h3cc37817),
	.w6(32'h3bce1716),
	.w7(32'h3c0414bc),
	.w8(32'h3c03b386),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1eef5a),
	.w1(32'h3c3aa66f),
	.w2(32'h3cf1d738),
	.w3(32'h3c8e5493),
	.w4(32'h3cc34169),
	.w5(32'h3ce659da),
	.w6(32'h3bd8b334),
	.w7(32'h3cbf8f6d),
	.w8(32'h3dd710aa),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56af12),
	.w1(32'h3c09ca01),
	.w2(32'h3d2fa8f0),
	.w3(32'h3ccd04d0),
	.w4(32'h3c5e1061),
	.w5(32'h3c6d74a5),
	.w6(32'h3bb8faf9),
	.w7(32'h3cf2776d),
	.w8(32'h3d1d4d1c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6199fb),
	.w1(32'h3d6e2e04),
	.w2(32'h3c9c4222),
	.w3(32'h3c857af2),
	.w4(32'h3caa09c5),
	.w5(32'h3c59f0c3),
	.w6(32'h3c98bad9),
	.w7(32'h3cc6d9a6),
	.w8(32'h3c766d83),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2eb1f3),
	.w1(32'h3d584a61),
	.w2(32'h3b12d663),
	.w3(32'h3ceaf09c),
	.w4(32'h3c6f01fd),
	.w5(32'hb9bb4568),
	.w6(32'h3d27604b),
	.w7(32'hbafd322c),
	.w8(32'h3bb0d7ce),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91b978),
	.w1(32'hbb4fb48c),
	.w2(32'h3c258732),
	.w3(32'h3b852cd0),
	.w4(32'h3bf27904),
	.w5(32'hba8d3f4b),
	.w6(32'hbae926e5),
	.w7(32'hb90b855e),
	.w8(32'h39ea44e6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab497ec),
	.w1(32'hbb0bbf8b),
	.w2(32'h3acaf72f),
	.w3(32'h39c67241),
	.w4(32'hba014c46),
	.w5(32'h3ae3da5c),
	.w6(32'hbb49c2ca),
	.w7(32'h3b70b8e3),
	.w8(32'hbb2e311d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979cc53),
	.w1(32'hbbe146bc),
	.w2(32'h3b7e4d73),
	.w3(32'hbb375446),
	.w4(32'h3b960913),
	.w5(32'hbb342ee7),
	.w6(32'h3b5c36c0),
	.w7(32'h3996e7f1),
	.w8(32'h39780cb7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38443c8f),
	.w1(32'h3a115920),
	.w2(32'h3a4691cb),
	.w3(32'h3b180d50),
	.w4(32'h392aebab),
	.w5(32'h3c663768),
	.w6(32'h3b8d2aee),
	.w7(32'hbb8e8d92),
	.w8(32'hbabfa89e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa7ea7),
	.w1(32'hbb01b056),
	.w2(32'h3c937c01),
	.w3(32'h3b1d6525),
	.w4(32'hbae0a4d6),
	.w5(32'h3b146c25),
	.w6(32'h3b8343e7),
	.w7(32'h3ab340d1),
	.w8(32'h3b70f7f8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc64fd),
	.w1(32'h3b0b8fee),
	.w2(32'h3a9bf7e2),
	.w3(32'h3a42589f),
	.w4(32'h3b822ae3),
	.w5(32'hbb47d64b),
	.w6(32'hbb53fbd5),
	.w7(32'h3a784e63),
	.w8(32'hbb9cae6d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb96899),
	.w1(32'h3b83fc92),
	.w2(32'h37f7abf5),
	.w3(32'h37c04393),
	.w4(32'h39682d24),
	.w5(32'h3a1de41d),
	.w6(32'hbc0ea64c),
	.w7(32'hbb2c6d99),
	.w8(32'hba785d0e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a45ba),
	.w1(32'h3ae15059),
	.w2(32'hbb87bd97),
	.w3(32'h393f5403),
	.w4(32'hbb90a015),
	.w5(32'h3c9eb56c),
	.w6(32'h3af3e4ef),
	.w7(32'hbb5d562a),
	.w8(32'hbadfc8d6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01805c),
	.w1(32'h39bdd145),
	.w2(32'h3a9aa9cf),
	.w3(32'h3bad4f43),
	.w4(32'hbba55953),
	.w5(32'hbb3601d0),
	.w6(32'h3cbe3af9),
	.w7(32'hbb368644),
	.w8(32'h3b8c1ddc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5295fa),
	.w1(32'hbb835c6a),
	.w2(32'h3bbf73f6),
	.w3(32'h3a8fcedb),
	.w4(32'hbb1ff062),
	.w5(32'hbb836979),
	.w6(32'hbb47ce60),
	.w7(32'h3b053905),
	.w8(32'h3b8afd50),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0de52f),
	.w1(32'hba2b48ed),
	.w2(32'h38bd5853),
	.w3(32'h38da47d6),
	.w4(32'hba819c39),
	.w5(32'hbaa046a5),
	.w6(32'h383cb58d),
	.w7(32'h3c7730ff),
	.w8(32'hbb96a3ff),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf631b),
	.w1(32'h3b1588e5),
	.w2(32'hbb2cfbf6),
	.w3(32'h39a59211),
	.w4(32'hbab040e0),
	.w5(32'h3c763cc7),
	.w6(32'h3c079745),
	.w7(32'h3b911c04),
	.w8(32'h39d8ef52),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2d57),
	.w1(32'h38aece50),
	.w2(32'h3a644d3f),
	.w3(32'hbc66ea31),
	.w4(32'hbb1554e3),
	.w5(32'hba091998),
	.w6(32'hbb4cd081),
	.w7(32'hbaa75d51),
	.w8(32'h36dbe1f7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ea2ac),
	.w1(32'h3b32c00e),
	.w2(32'hba6adc06),
	.w3(32'hb92a8a31),
	.w4(32'hba9c32c2),
	.w5(32'h388930e9),
	.w6(32'h3b6ff6cb),
	.w7(32'hbbcee76e),
	.w8(32'h3b6a0d27),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba76f6b),
	.w1(32'h3cc8dac3),
	.w2(32'hbb87756e),
	.w3(32'h3758076c),
	.w4(32'hbb1e52ad),
	.w5(32'hbb57bdcc),
	.w6(32'hb8c937e6),
	.w7(32'hb915d6b5),
	.w8(32'h3c3db3c5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc198108),
	.w1(32'hb9cda91a),
	.w2(32'hba225380),
	.w3(32'h3adc7e27),
	.w4(32'h3ae65ace),
	.w5(32'h3b444e35),
	.w6(32'hbb65b6ff),
	.w7(32'hba8a8fdf),
	.w8(32'hbbb7cbeb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5688a6),
	.w1(32'hbaf066d7),
	.w2(32'h3b437439),
	.w3(32'hba394031),
	.w4(32'h3a64602c),
	.w5(32'hb8b97d86),
	.w6(32'hbb6b0b2e),
	.w7(32'hb9b86cc2),
	.w8(32'hba6a93a3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0266f6),
	.w1(32'h3bc6d1ac),
	.w2(32'h3c857cc1),
	.w3(32'h3aff2655),
	.w4(32'h39a56f96),
	.w5(32'h36c27de1),
	.w6(32'h3cee1da4),
	.w7(32'h3b163d5f),
	.w8(32'h3b24487b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb082ba1),
	.w1(32'hbb4a924d),
	.w2(32'hbc8e3b0a),
	.w3(32'hbb83db01),
	.w4(32'hbb8c7f81),
	.w5(32'h3bb65ac3),
	.w6(32'hbae1dcfa),
	.w7(32'h3b95c4af),
	.w8(32'hbc5ea9af),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba525cad),
	.w1(32'h3c2cf257),
	.w2(32'hbb968ea7),
	.w3(32'hb98add2a),
	.w4(32'h3b6f5024),
	.w5(32'h3aa1e17f),
	.w6(32'h3b890bf7),
	.w7(32'hbbbcb1ab),
	.w8(32'h3b8e3e24),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895823),
	.w1(32'hbb9f8c7c),
	.w2(32'hbb3ce098),
	.w3(32'h3963ae96),
	.w4(32'hba823a3f),
	.w5(32'h3c49b3ee),
	.w6(32'h3ba7a566),
	.w7(32'hbb488d6d),
	.w8(32'h394b6e8d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30e6e3),
	.w1(32'h3a0de8b4),
	.w2(32'hbaf0e403),
	.w3(32'hbb9c4dcb),
	.w4(32'h3b1b1fd3),
	.w5(32'h3b18b14d),
	.w6(32'hba39bdef),
	.w7(32'hbae33c33),
	.w8(32'h3a7dd5c7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c364aed),
	.w1(32'h3bfe96ca),
	.w2(32'h39bcd384),
	.w3(32'h3bdc6da6),
	.w4(32'hba1361c3),
	.w5(32'hb9e03d64),
	.w6(32'hb9eda84e),
	.w7(32'hb9409210),
	.w8(32'hb9120ff8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09264c),
	.w1(32'hbb76785c),
	.w2(32'h3a1507da),
	.w3(32'hb9d460fc),
	.w4(32'h3a8c694b),
	.w5(32'hbac8fa9f),
	.w6(32'hb960dd89),
	.w7(32'hba5b2ce0),
	.w8(32'h3ace57d6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c32a6),
	.w1(32'h3b04e11e),
	.w2(32'h3bae9a48),
	.w3(32'hbc854e9c),
	.w4(32'h3b95f936),
	.w5(32'hba191079),
	.w6(32'h3b2a6b2d),
	.w7(32'h3b68e2d7),
	.w8(32'hb98c4ecd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb313bda),
	.w1(32'h3b0d04f6),
	.w2(32'hbb4c5947),
	.w3(32'hbaf24ce0),
	.w4(32'h3b41d10d),
	.w5(32'h3b594b49),
	.w6(32'h3b9e904d),
	.w7(32'hbac45ffa),
	.w8(32'hbbaae202),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b778769),
	.w1(32'h3bbacd63),
	.w2(32'h3982db42),
	.w3(32'h3b7a0586),
	.w4(32'h3b94d1a9),
	.w5(32'h3bf2871d),
	.w6(32'h3bccc434),
	.w7(32'h3a9147b5),
	.w8(32'hba70e7b0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf71c23),
	.w1(32'h3b627e59),
	.w2(32'h3ad10113),
	.w3(32'h39fcbfc4),
	.w4(32'h3a62ab65),
	.w5(32'h39a86837),
	.w6(32'h3b3045cc),
	.w7(32'h3ae5d5f9),
	.w8(32'h39e1d1b1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbf35a),
	.w1(32'hbabefc87),
	.w2(32'hbbe28514),
	.w3(32'h3b91c93f),
	.w4(32'hba014d4a),
	.w5(32'hba942251),
	.w6(32'hba90ad9e),
	.w7(32'h3ace4dae),
	.w8(32'hbc8e8419),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b270074),
	.w1(32'h39fd1519),
	.w2(32'h3b0c3d12),
	.w3(32'h3c82850e),
	.w4(32'hbbbc39e2),
	.w5(32'h3a94986e),
	.w6(32'hbaacb535),
	.w7(32'hba3bacd4),
	.w8(32'hba81cec5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc334f09),
	.w1(32'h3b897b9a),
	.w2(32'h3b514bf2),
	.w3(32'h3a54f4f9),
	.w4(32'hbb56698f),
	.w5(32'hba8828f4),
	.w6(32'h39d6acb7),
	.w7(32'hbb93904d),
	.w8(32'h3b831096),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fe884),
	.w1(32'h3adf7fd0),
	.w2(32'hb604cbc6),
	.w3(32'hba530378),
	.w4(32'h3b3d8887),
	.w5(32'h3ad48ac6),
	.w6(32'h3a4f891a),
	.w7(32'h39c137c0),
	.w8(32'hba9d95ee),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9abb88),
	.w1(32'h3abe4433),
	.w2(32'h3a9e725a),
	.w3(32'h3a1ac872),
	.w4(32'h3c06c6b9),
	.w5(32'h3968afdb),
	.w6(32'h3aff63de),
	.w7(32'hbb37c614),
	.w8(32'h3bafb89a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a8ec),
	.w1(32'h3b0cf816),
	.w2(32'hbb6ad756),
	.w3(32'h3b88eddf),
	.w4(32'h3aab6968),
	.w5(32'h3b33c431),
	.w6(32'h3b13a3f0),
	.w7(32'h3b565c36),
	.w8(32'hbb42c0f5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba22788),
	.w1(32'hbb5442fa),
	.w2(32'hbbc2ed84),
	.w3(32'h3abe9200),
	.w4(32'h3b1413dc),
	.w5(32'hbb43441a),
	.w6(32'hbae06ed6),
	.w7(32'hba156d21),
	.w8(32'h3b214d83),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fa3c5),
	.w1(32'hbab2f481),
	.w2(32'h3b2e5e48),
	.w3(32'hbb76d312),
	.w4(32'h3a10d2d7),
	.w5(32'hba53a192),
	.w6(32'h3b8a4d13),
	.w7(32'hb9f02383),
	.w8(32'h39fcc190),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9c570),
	.w1(32'hbb735b75),
	.w2(32'hb9a070eb),
	.w3(32'h3ac67ffe),
	.w4(32'h3b0035ff),
	.w5(32'hbb7a6aae),
	.w6(32'hbb369355),
	.w7(32'h3d23702a),
	.w8(32'h3a606035),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1401d5),
	.w1(32'h3930eb93),
	.w2(32'h3b92edcd),
	.w3(32'hbb2d1be6),
	.w4(32'hbbccd6dc),
	.w5(32'hbbafc3c4),
	.w6(32'hbbc1bbfc),
	.w7(32'hb95a528b),
	.w8(32'hb9addc31),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b7ba1),
	.w1(32'h398c349f),
	.w2(32'hb61ff58a),
	.w3(32'h3cc9a70c),
	.w4(32'hbbd8b7c6),
	.w5(32'hba9f2867),
	.w6(32'h3a5cce14),
	.w7(32'hbb4894a8),
	.w8(32'hbb8518c0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6e747),
	.w1(32'hbc9edfbc),
	.w2(32'hba8537b1),
	.w3(32'h3897de4e),
	.w4(32'h3a2fdccb),
	.w5(32'h3b6fb5f4),
	.w6(32'hbb9c6f99),
	.w7(32'h39895b24),
	.w8(32'hba419fe3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad64395),
	.w1(32'h3a2233e8),
	.w2(32'h3a467261),
	.w3(32'hbb113d94),
	.w4(32'h3a1e2d78),
	.w5(32'hbc00f917),
	.w6(32'hbb8776dc),
	.w7(32'hbc5d3c39),
	.w8(32'hbbaf99a3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39997214),
	.w1(32'hb2eb2f75),
	.w2(32'hbaff8dfd),
	.w3(32'h3aab075a),
	.w4(32'h3b93251a),
	.w5(32'hba600e0c),
	.w6(32'hba09e61d),
	.w7(32'h39220a4e),
	.w8(32'hbaa34fd5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3806e46f),
	.w1(32'h3b80cac3),
	.w2(32'h3aacc569),
	.w3(32'h3a263f8b),
	.w4(32'h3b946fe7),
	.w5(32'h3d02bc6d),
	.w6(32'h39ec2094),
	.w7(32'h3b07bb20),
	.w8(32'hba838c81),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ae461),
	.w1(32'h3bba5df9),
	.w2(32'hbaadae57),
	.w3(32'h3a978e27),
	.w4(32'h3a9f0e8f),
	.w5(32'h3a4e776e),
	.w6(32'hbbcc3e2c),
	.w7(32'h3a53ddaa),
	.w8(32'hbb16fc0b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932ded),
	.w1(32'h3aa2b6a1),
	.w2(32'h3bc21ef4),
	.w3(32'hba98f606),
	.w4(32'h3acdd976),
	.w5(32'h3a15e076),
	.w6(32'h3b19fad8),
	.w7(32'h3b9fc572),
	.w8(32'h3d1b3ef7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18066d),
	.w1(32'h3a8527dc),
	.w2(32'h3c8d97bb),
	.w3(32'hbac2afaa),
	.w4(32'hba1fef56),
	.w5(32'h38cda854),
	.w6(32'h39bf510d),
	.w7(32'h3b0e3270),
	.w8(32'hbb308c86),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b735582),
	.w1(32'h3897e526),
	.w2(32'h3abce50e),
	.w3(32'h3cd2a11d),
	.w4(32'hba6b6b66),
	.w5(32'hba440974),
	.w6(32'hb80ef336),
	.w7(32'hbc959429),
	.w8(32'h39bbb37a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eaa669),
	.w1(32'hbc11ed74),
	.w2(32'h39d2937f),
	.w3(32'hbc48b5e7),
	.w4(32'hbb7fe505),
	.w5(32'h3b4c3a40),
	.w6(32'h3a542394),
	.w7(32'h3a1442b9),
	.w8(32'hba34ea9f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab415ed),
	.w1(32'hbaa8d1e4),
	.w2(32'h3b62b07f),
	.w3(32'h3a34f6aa),
	.w4(32'h3b06aea3),
	.w5(32'hbbbf0d96),
	.w6(32'hba2b27fb),
	.w7(32'h3c030c7a),
	.w8(32'hbadef645),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb6708),
	.w1(32'h3a55caf5),
	.w2(32'hb99cf915),
	.w3(32'h3b129617),
	.w4(32'hbbafdefa),
	.w5(32'h3960f09c),
	.w6(32'h3b2ed702),
	.w7(32'hb9d7772f),
	.w8(32'h3abd8350),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9eb3ac),
	.w1(32'h3b6d311a),
	.w2(32'hb9744652),
	.w3(32'hbb03f376),
	.w4(32'h3b85bfc6),
	.w5(32'hbc1646e5),
	.w6(32'hbb3e3e4b),
	.w7(32'hba07838b),
	.w8(32'h39b1a274),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae10bde),
	.w1(32'hb970d4b8),
	.w2(32'h38b29af6),
	.w3(32'h3b8cb5cf),
	.w4(32'h3b15f8a4),
	.w5(32'hba3ebbb8),
	.w6(32'hbac3bcc5),
	.w7(32'hba126e50),
	.w8(32'h3a8eb529),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08c59c),
	.w1(32'h3a01c18d),
	.w2(32'hbabe5778),
	.w3(32'hb64f31f6),
	.w4(32'hbc3450d6),
	.w5(32'hbb3a6e3f),
	.w6(32'hbb01600a),
	.w7(32'hbb57788c),
	.w8(32'h39e37769),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad17909),
	.w1(32'hba069237),
	.w2(32'hba4278df),
	.w3(32'hbac0000b),
	.w4(32'hbafbe2f3),
	.w5(32'h3aeec9ad),
	.w6(32'hb93e7a0b),
	.w7(32'h3b4b4f12),
	.w8(32'hbaa909a1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3429e),
	.w1(32'h3b714ad3),
	.w2(32'h3949294b),
	.w3(32'h3ab95017),
	.w4(32'h3a0325b0),
	.w5(32'hbb22a173),
	.w6(32'h3b263e9d),
	.w7(32'h3b2499bf),
	.w8(32'h3b1c8288),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba98add),
	.w1(32'hbb484144),
	.w2(32'h3afdeda2),
	.w3(32'hbb84226c),
	.w4(32'h3a9a79bd),
	.w5(32'hbaf9d0ba),
	.w6(32'hbb898acb),
	.w7(32'h399ced64),
	.w8(32'h3b48346e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15682a),
	.w1(32'hb8983f25),
	.w2(32'hbc3f67db),
	.w3(32'h3ac1caf1),
	.w4(32'hbc61a72f),
	.w5(32'h3c1fc911),
	.w6(32'h3b94b3c7),
	.w7(32'hba02f4d7),
	.w8(32'h3b124591),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae34154),
	.w1(32'hbcc78ca2),
	.w2(32'hbab729bf),
	.w3(32'hbbbbd187),
	.w4(32'h3c1482da),
	.w5(32'hb99b0ae9),
	.w6(32'hbc069ce6),
	.w7(32'h3c1f0284),
	.w8(32'hbbc64a89),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4f271),
	.w1(32'h3907fd53),
	.w2(32'h3c3e732a),
	.w3(32'h3bbe291e),
	.w4(32'hbc66d946),
	.w5(32'hbb78bd20),
	.w6(32'hbb4f17a9),
	.w7(32'h3c31c30e),
	.w8(32'h3b01fd26),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fee9b),
	.w1(32'h3b7d169c),
	.w2(32'h3b546bcb),
	.w3(32'h3b0d6b7d),
	.w4(32'hba2c7d68),
	.w5(32'h3b274bef),
	.w6(32'hbccb3164),
	.w7(32'hbc8a1458),
	.w8(32'h3a006bd1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05e32b),
	.w1(32'hbbab69ec),
	.w2(32'hbc2a5aa6),
	.w3(32'hbc039a55),
	.w4(32'h3d45e119),
	.w5(32'hbaaf28a3),
	.w6(32'h3bf3d8ef),
	.w7(32'h3b4e11d2),
	.w8(32'hba5d40cd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97656),
	.w1(32'hbb60e525),
	.w2(32'hbcafe3fa),
	.w3(32'h3b443528),
	.w4(32'h3ad7afb2),
	.w5(32'h3b92c21a),
	.w6(32'hbbb9fddc),
	.w7(32'hbbcec0ed),
	.w8(32'hbad253d8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f88a1),
	.w1(32'h3b27eea8),
	.w2(32'hbb6f0e6c),
	.w3(32'hbbe962e9),
	.w4(32'h3aea9f1e),
	.w5(32'h3aeb162c),
	.w6(32'h37cae89e),
	.w7(32'hbc37cea2),
	.w8(32'hbb07b4b1),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba466171),
	.w1(32'h3b9a23e0),
	.w2(32'hbb6e0830),
	.w3(32'h3d47d17b),
	.w4(32'h3b3769bb),
	.w5(32'h3a711a88),
	.w6(32'hbbfb1323),
	.w7(32'hba41ea7c),
	.w8(32'h3b772a2d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fb81a),
	.w1(32'h3c35676f),
	.w2(32'hbd5f0e34),
	.w3(32'h3af8c598),
	.w4(32'h3ba8fced),
	.w5(32'h398fd181),
	.w6(32'hbad4adac),
	.w7(32'hbab7b1fe),
	.w8(32'h3a62b439),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c13e7),
	.w1(32'hbb9d7edc),
	.w2(32'hbae71748),
	.w3(32'hbc6b021c),
	.w4(32'hbb9284c1),
	.w5(32'h3c0ae409),
	.w6(32'hbc911450),
	.w7(32'h3ba3fd27),
	.w8(32'hbba2428e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab16e99),
	.w1(32'hbadf601d),
	.w2(32'hba1fe488),
	.w3(32'hbb02d64e),
	.w4(32'hb9b567f1),
	.w5(32'hbbc2a6ff),
	.w6(32'h3ba09af4),
	.w7(32'hbc26655b),
	.w8(32'hbbc6e002),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9549e1),
	.w1(32'hbc666b8a),
	.w2(32'hbbf69987),
	.w3(32'hb8ca7f38),
	.w4(32'hbbcc5434),
	.w5(32'hbc0980c7),
	.w6(32'hbd928115),
	.w7(32'hb886723d),
	.w8(32'hb91c2ef5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf73011),
	.w1(32'hbb9f59c0),
	.w2(32'hbc8b0bc6),
	.w3(32'h3ba657ff),
	.w4(32'h3a58052e),
	.w5(32'h3a163869),
	.w6(32'h3b31c7d5),
	.w7(32'h3a2574ed),
	.w8(32'h3b3d0c60),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c113a6c),
	.w1(32'h3aaeab12),
	.w2(32'hbd2abd23),
	.w3(32'h3bb8e2e2),
	.w4(32'hbc10df8f),
	.w5(32'hb67b55d4),
	.w6(32'h3b822912),
	.w7(32'h3b8d4b9d),
	.w8(32'hbd3df413),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39236f28),
	.w1(32'hbbfb3e84),
	.w2(32'hba82aed7),
	.w3(32'hb947571d),
	.w4(32'h3b4cd335),
	.w5(32'hbb6f10f2),
	.w6(32'hbbf2642a),
	.w7(32'hbb8ef754),
	.w8(32'hbbee4f86),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c342660),
	.w1(32'hbc1b6298),
	.w2(32'h3c9ebfa9),
	.w3(32'hbb6fa36e),
	.w4(32'h3c514a5f),
	.w5(32'hbb6f56ba),
	.w6(32'hbb3f3c10),
	.w7(32'hbc79a77c),
	.w8(32'h3bc2522d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab046a9),
	.w1(32'h3b2ad586),
	.w2(32'hbb23fe0e),
	.w3(32'hba93d8f9),
	.w4(32'hba064cde),
	.w5(32'h3a7498e3),
	.w6(32'hbc1a3f21),
	.w7(32'hbb0e5dc9),
	.w8(32'hbc8d5678),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d1526),
	.w1(32'h3c08d0f8),
	.w2(32'h3be0fd31),
	.w3(32'h3bd7dd91),
	.w4(32'h3b5cc777),
	.w5(32'hbbd64065),
	.w6(32'h3babbeda),
	.w7(32'h3bfa13d5),
	.w8(32'h39b44fb4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cacea),
	.w1(32'h3887157b),
	.w2(32'hb672b489),
	.w3(32'hbc91bfcd),
	.w4(32'hbb8fcdb1),
	.w5(32'h39618261),
	.w6(32'hbb289586),
	.w7(32'hbc08531c),
	.w8(32'h3c377dad),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6506b1),
	.w1(32'hbb7a554c),
	.w2(32'hbb86c5af),
	.w3(32'h3ad9bfac),
	.w4(32'hbbe66f43),
	.w5(32'h3cc2dc24),
	.w6(32'hbb60d2c1),
	.w7(32'h3c9bd939),
	.w8(32'hbbc59a6c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d7a72),
	.w1(32'h39bb9ce1),
	.w2(32'h3aa47468),
	.w3(32'h3bf0bbb7),
	.w4(32'hb8ab7a2d),
	.w5(32'hbb1e5ba9),
	.w6(32'hbb98fe00),
	.w7(32'h3c13a8f8),
	.w8(32'hbaa19a3a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc4415),
	.w1(32'h3abbce58),
	.w2(32'hbd4ade47),
	.w3(32'hbb28fcde),
	.w4(32'hbb5569ba),
	.w5(32'h3bf324fb),
	.w6(32'h3c60507e),
	.w7(32'hbc87a6de),
	.w8(32'hbc4f1aef),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba6790),
	.w1(32'h3abfa98f),
	.w2(32'hbaacf749),
	.w3(32'h3c003db2),
	.w4(32'h3c6c3273),
	.w5(32'hbc079a6a),
	.w6(32'h3c19cbda),
	.w7(32'hbb6294c2),
	.w8(32'hbd1d8910),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad21198),
	.w1(32'hbaf126fa),
	.w2(32'h3a35bd6e),
	.w3(32'hba504401),
	.w4(32'h3a3dd757),
	.w5(32'h38a401f8),
	.w6(32'hbd190ed7),
	.w7(32'hbb85c354),
	.w8(32'hbb9f4067),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d95b7),
	.w1(32'hbb869220),
	.w2(32'h3ad96abf),
	.w3(32'h3b9e5d6c),
	.w4(32'h37b806e7),
	.w5(32'hb8cafc62),
	.w6(32'h3c09caed),
	.w7(32'h391634f8),
	.w8(32'hbd477f5d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6c7cb),
	.w1(32'h3a88a4e5),
	.w2(32'h3aa65c6d),
	.w3(32'h3b7920c0),
	.w4(32'h3a5b9fcc),
	.w5(32'hbca517a7),
	.w6(32'hbc2ab579),
	.w7(32'hbc2c92ed),
	.w8(32'hbc1b933c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b556c4c),
	.w1(32'hba8a9c42),
	.w2(32'hbb1e6e9c),
	.w3(32'h3bfba198),
	.w4(32'hbb3f8e70),
	.w5(32'h3b293ca1),
	.w6(32'h3b9ff615),
	.w7(32'h3bf032f0),
	.w8(32'hbba3e5bb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb945e8),
	.w1(32'hbb931e70),
	.w2(32'hbc5b554a),
	.w3(32'h3c24a527),
	.w4(32'hbb9c775f),
	.w5(32'hbb6b60fb),
	.w6(32'hbc64ca69),
	.w7(32'h3a66c463),
	.w8(32'h3c44e975),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b92a3),
	.w1(32'hba997eb0),
	.w2(32'hbb9f689d),
	.w3(32'hbba89b5e),
	.w4(32'h38b2ca5e),
	.w5(32'hba229cee),
	.w6(32'hba51be4f),
	.w7(32'h3b9e9a59),
	.w8(32'h3a9a6c5f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b389f57),
	.w1(32'h3b419a45),
	.w2(32'hbb6f53a6),
	.w3(32'h3aaed2e2),
	.w4(32'h3b081f1c),
	.w5(32'h3bb03ee0),
	.w6(32'hbb253f09),
	.w7(32'hbb3a0f48),
	.w8(32'hbb8669b6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92c36a),
	.w1(32'hbac43749),
	.w2(32'h3ac8c479),
	.w3(32'hbae269e0),
	.w4(32'hbb683788),
	.w5(32'hba8d6bfe),
	.w6(32'hbb975755),
	.w7(32'h3b9f6100),
	.w8(32'h3ce57e8e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4be7bf),
	.w1(32'h3b34feaf),
	.w2(32'h3d143c32),
	.w3(32'h3ba35faf),
	.w4(32'h3a95524e),
	.w5(32'h3b96181c),
	.w6(32'h3b0cb8c0),
	.w7(32'h3a40a89e),
	.w8(32'hb9ce8578),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16e835),
	.w1(32'hba95fd9e),
	.w2(32'h3b6562c9),
	.w3(32'h392fa4ca),
	.w4(32'h3a2a1a0f),
	.w5(32'h3ada071f),
	.w6(32'hbb032870),
	.w7(32'h3abe9112),
	.w8(32'hbb7b831c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff0e13),
	.w1(32'h3aae356a),
	.w2(32'h3b91555f),
	.w3(32'h3b924f4b),
	.w4(32'hbb318f08),
	.w5(32'hbac7dca5),
	.w6(32'hbb647534),
	.w7(32'h3b00e96c),
	.w8(32'hb999ea6f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4efb4e),
	.w1(32'h39e05e6c),
	.w2(32'hba72940e),
	.w3(32'h3b86d43f),
	.w4(32'h3a76e97b),
	.w5(32'hbb4c2a43),
	.w6(32'h3ac177b9),
	.w7(32'hb9ef41e0),
	.w8(32'hb994582b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370ab4bd),
	.w1(32'h3b3400a4),
	.w2(32'h3b226837),
	.w3(32'hbb100e6a),
	.w4(32'hb840bd1c),
	.w5(32'hba34e6a2),
	.w6(32'hbb849679),
	.w7(32'h3baa766e),
	.w8(32'h3bd19117),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98d74e),
	.w1(32'h3adc8f7f),
	.w2(32'hb924e0b9),
	.w3(32'h3b23784b),
	.w4(32'h3b188b3c),
	.w5(32'hbb0e22e0),
	.w6(32'h3a95db16),
	.w7(32'h3b014f85),
	.w8(32'hbad774d8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc21327),
	.w1(32'hbbd5c425),
	.w2(32'h3aa1feb5),
	.w3(32'hbc39c770),
	.w4(32'h3b92c227),
	.w5(32'hbb5484e2),
	.w6(32'hbb5aae83),
	.w7(32'hb9fb3e93),
	.w8(32'h397a7fd9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20121f),
	.w1(32'h3c03eab1),
	.w2(32'h3c2d6e63),
	.w3(32'hb94d7c48),
	.w4(32'h3a84dd52),
	.w5(32'h3b331edb),
	.w6(32'hbbb7dd6e),
	.w7(32'h3b4b8a54),
	.w8(32'hbb8b0ca4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b0e30),
	.w1(32'h3c100b07),
	.w2(32'hbb7a0e48),
	.w3(32'h3bb1ff56),
	.w4(32'h392ed316),
	.w5(32'h3b976b8d),
	.w6(32'hbac00738),
	.w7(32'hb4f8bdd6),
	.w8(32'hbbb31ef1),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e4a006),
	.w1(32'h3be23645),
	.w2(32'h3b61e4c5),
	.w3(32'h3b30dd82),
	.w4(32'h39c395c9),
	.w5(32'h3b8737d4),
	.w6(32'h3c1d68b2),
	.w7(32'h3b67600c),
	.w8(32'h3b08bfd3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec99c0),
	.w1(32'hbab40429),
	.w2(32'h3cd6e5cd),
	.w3(32'hbc4a3f66),
	.w4(32'h3cc99713),
	.w5(32'h3a25f504),
	.w6(32'h3a37fa5f),
	.w7(32'hbb06e90e),
	.w8(32'hba32adb3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba915987),
	.w1(32'h3b17b803),
	.w2(32'h3accc31e),
	.w3(32'h3a143891),
	.w4(32'h3845c095),
	.w5(32'h3a4ed9cc),
	.w6(32'h354d4a50),
	.w7(32'h3a8c56fd),
	.w8(32'hbb8d2e63),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f51cc),
	.w1(32'hbb2677b2),
	.w2(32'hbc7fe826),
	.w3(32'h3ab99b6a),
	.w4(32'h3937c14a),
	.w5(32'hbb13f238),
	.w6(32'h3ab6776e),
	.w7(32'h3488a2d8),
	.w8(32'hbb5d5c77),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae3891),
	.w1(32'h3a3aa1a0),
	.w2(32'hbb5423af),
	.w3(32'h3a2f54ba),
	.w4(32'h3ab30a2a),
	.w5(32'hbb3b3d08),
	.w6(32'hbcf6c1fb),
	.w7(32'h3aab1e6b),
	.w8(32'h3bbdb90c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fcefc),
	.w1(32'h3ac28122),
	.w2(32'h3ad3a291),
	.w3(32'h3b70c452),
	.w4(32'h3b8cb0ee),
	.w5(32'hbb6acfb9),
	.w6(32'h3c077f33),
	.w7(32'hbac71b60),
	.w8(32'hbb8077b1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c492d),
	.w1(32'h3b39a9df),
	.w2(32'h3b7d7291),
	.w3(32'hba8bd670),
	.w4(32'hb7c650b3),
	.w5(32'h3af25601),
	.w6(32'hbb1569f1),
	.w7(32'hbc983181),
	.w8(32'hb98608be),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40b596),
	.w1(32'h3b3a30b2),
	.w2(32'h3a9ae48c),
	.w3(32'hb7b45dc0),
	.w4(32'h3b654c3c),
	.w5(32'hbb820a76),
	.w6(32'h3b5d0567),
	.w7(32'hbbad66ee),
	.w8(32'h3bc304d0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d044530),
	.w1(32'h3c962c2f),
	.w2(32'h3aa10748),
	.w3(32'h3b55c91c),
	.w4(32'h39eb4d7b),
	.w5(32'hba5bb6b5),
	.w6(32'hbae15034),
	.w7(32'hbb532abd),
	.w8(32'h3ab76770),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0d9da),
	.w1(32'hbaccb284),
	.w2(32'h3cf41e12),
	.w3(32'hbac2cd28),
	.w4(32'hbc03e646),
	.w5(32'h3b08ce23),
	.w6(32'h3a574a48),
	.w7(32'hbb7e4c82),
	.w8(32'h3ad7ca9b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc79f6),
	.w1(32'h3a40242d),
	.w2(32'h3a0d36dc),
	.w3(32'h389bef59),
	.w4(32'h3b2bb9d2),
	.w5(32'h3ac52ef6),
	.w6(32'h3b17c8fc),
	.w7(32'hbba3e1fe),
	.w8(32'hbbe190e5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a4175),
	.w1(32'hbc1112b2),
	.w2(32'h3b0144c7),
	.w3(32'h3af8117c),
	.w4(32'h3a0365c0),
	.w5(32'h38a43c4d),
	.w6(32'hba229550),
	.w7(32'h37a58d69),
	.w8(32'h3a8fa901),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38633f),
	.w1(32'h3a928e81),
	.w2(32'hb96d2897),
	.w3(32'h3b338afb),
	.w4(32'hbab50f44),
	.w5(32'h3b13287a),
	.w6(32'h38fa4db2),
	.w7(32'hbb06ad8b),
	.w8(32'hba0e6561),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7949b78),
	.w1(32'hbc15ccab),
	.w2(32'hbb0990f9),
	.w3(32'hbb340255),
	.w4(32'hbb2511e9),
	.w5(32'h3b07ca97),
	.w6(32'h3accfe1a),
	.w7(32'h3a42313b),
	.w8(32'hbb589e98),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ab72a8),
	.w1(32'h3a827bb0),
	.w2(32'h38930b7e),
	.w3(32'h3ade861a),
	.w4(32'h3982fe5b),
	.w5(32'h3a00da2f),
	.w6(32'hbb891c5c),
	.w7(32'hbaf550b2),
	.w8(32'h3b8855d1),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d73c1),
	.w1(32'h3b7603d2),
	.w2(32'h3c019c83),
	.w3(32'h3ac582d2),
	.w4(32'h3a15b31f),
	.w5(32'h3aa1ea0e),
	.w6(32'hb982f1e4),
	.w7(32'hbb733346),
	.w8(32'hbc41b1fa),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b277e80),
	.w1(32'h3b1c2885),
	.w2(32'h3b59d66f),
	.w3(32'hbbb811c4),
	.w4(32'h39018a4c),
	.w5(32'h39ad6f3a),
	.w6(32'h3afba4f8),
	.w7(32'hbb17946d),
	.w8(32'h3b4735e4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a7824),
	.w1(32'h3b8ced98),
	.w2(32'hbbaf1700),
	.w3(32'hbae0f911),
	.w4(32'h3a0d0606),
	.w5(32'h3b3711c9),
	.w6(32'h3a5f2e52),
	.w7(32'h3c185f40),
	.w8(32'h3990cf55),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a315c),
	.w1(32'h3ac5970b),
	.w2(32'h3bb3f86b),
	.w3(32'hba0b2eec),
	.w4(32'hbbb96cca),
	.w5(32'h38febff9),
	.w6(32'h3cc8b964),
	.w7(32'hba4f331b),
	.w8(32'hbb81a935),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050aff),
	.w1(32'h3c00f033),
	.w2(32'h3bc94bac),
	.w3(32'hbb02b88a),
	.w4(32'h3a81c274),
	.w5(32'h3a3748d8),
	.w6(32'h39c94f83),
	.w7(32'hbb14ff21),
	.w8(32'h39e991aa),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12dba6),
	.w1(32'h3b1b037a),
	.w2(32'h3b45b94a),
	.w3(32'h3d07ac23),
	.w4(32'hb8511d75),
	.w5(32'hba8bed8e),
	.w6(32'h3b785508),
	.w7(32'h3aabc5ca),
	.w8(32'hba9a3ac8),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9d598),
	.w1(32'hbab7984f),
	.w2(32'h3b7e85f6),
	.w3(32'hbb7e0416),
	.w4(32'h3b290ccc),
	.w5(32'hbc0b77f1),
	.w6(32'hbb4596c8),
	.w7(32'h3cbb5bd5),
	.w8(32'hba55dd9c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac32fc2),
	.w1(32'h3b18b981),
	.w2(32'h3b628ba5),
	.w3(32'h3b3d0fa4),
	.w4(32'hbbe9c007),
	.w5(32'hbb4cec81),
	.w6(32'h3c2556aa),
	.w7(32'h3bf14543),
	.w8(32'h3b225ba0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf961c4),
	.w1(32'hba7c99c8),
	.w2(32'h39580d92),
	.w3(32'hba43e01c),
	.w4(32'hbb8c3044),
	.w5(32'hba0a1ede),
	.w6(32'hbbbe0915),
	.w7(32'hb9e47b6f),
	.w8(32'hb9467f39),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eeee0),
	.w1(32'h3acdb1e0),
	.w2(32'h3a524121),
	.w3(32'hbadc6472),
	.w4(32'hb7d3ae78),
	.w5(32'hba15ffe1),
	.w6(32'hbbb6b1b9),
	.w7(32'h398f183b),
	.w8(32'hbb849d3d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf4512),
	.w1(32'hbac7cff5),
	.w2(32'h3acdb5cb),
	.w3(32'h3a7db5c7),
	.w4(32'h3ac42cf0),
	.w5(32'h3ab60396),
	.w6(32'hbba819e0),
	.w7(32'h3b4adb94),
	.w8(32'hbb34765b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f4b9),
	.w1(32'h3ae7eaaf),
	.w2(32'hbb1a684d),
	.w3(32'h3b18aa6a),
	.w4(32'h3b6c8d55),
	.w5(32'h3b460409),
	.w6(32'h39f4587b),
	.w7(32'h3a1fbbb8),
	.w8(32'h3aa0a95b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fc6ef),
	.w1(32'h3abf7024),
	.w2(32'hbb99f2ca),
	.w3(32'h3c1cfd57),
	.w4(32'hbbfa2d3a),
	.w5(32'h3b9bdda6),
	.w6(32'h3b1f2e7e),
	.w7(32'h3b0ef3d6),
	.w8(32'h3905153b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aada4d),
	.w1(32'hbbb28c56),
	.w2(32'h3bb03a29),
	.w3(32'hba63f65b),
	.w4(32'h383fc2c3),
	.w5(32'h3a908b98),
	.w6(32'h3b8e318b),
	.w7(32'hbb028011),
	.w8(32'h3ab78684),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54a368),
	.w1(32'h3a10788d),
	.w2(32'hbb0ac3e0),
	.w3(32'hbb5c57a8),
	.w4(32'hb9fed8bb),
	.w5(32'hbb83948a),
	.w6(32'h3bc70d95),
	.w7(32'h3ac4df6c),
	.w8(32'h3b0af5e8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac51bed),
	.w1(32'h3b5ff085),
	.w2(32'h35b3d881),
	.w3(32'h3bfa6bc7),
	.w4(32'hbb31dbf4),
	.w5(32'h3b2c8422),
	.w6(32'h3ad4a405),
	.w7(32'h3c537010),
	.w8(32'hb8a862d0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb019f73),
	.w1(32'hbb5c993f),
	.w2(32'h3b854e36),
	.w3(32'h3c284fc7),
	.w4(32'hbaec0e00),
	.w5(32'hbb5d563d),
	.w6(32'h398bd765),
	.w7(32'h3b9be44f),
	.w8(32'hbbb730db),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf675e2),
	.w1(32'hba6aff3c),
	.w2(32'hbbae5de3),
	.w3(32'hbc50f84e),
	.w4(32'hbb8e7623),
	.w5(32'hb8b2e333),
	.w6(32'h3b83643e),
	.w7(32'h3c86399a),
	.w8(32'h3b045c06),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb5f01),
	.w1(32'hbb551f7d),
	.w2(32'h3be3dab0),
	.w3(32'h3c225df3),
	.w4(32'h3b52df82),
	.w5(32'h3b87d611),
	.w6(32'hbb460204),
	.w7(32'h3b596e9e),
	.w8(32'hbadc8a96),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60bd9f),
	.w1(32'h398b790e),
	.w2(32'hba898325),
	.w3(32'hbad36e61),
	.w4(32'h3b1bbc41),
	.w5(32'hbb20bf6c),
	.w6(32'hbbe70081),
	.w7(32'h39cda1ff),
	.w8(32'h3b5069a8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc199b9e),
	.w1(32'hbbb3da11),
	.w2(32'h3abd0ce1),
	.w3(32'hbb1e2cb2),
	.w4(32'hbb477b10),
	.w5(32'h3905fe32),
	.w6(32'h39109546),
	.w7(32'hb73467a5),
	.w8(32'h3bbceb1e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba874261),
	.w1(32'h3a9e78a7),
	.w2(32'hbadd8e1d),
	.w3(32'hbb899aca),
	.w4(32'h3c6103ed),
	.w5(32'h3cac1229),
	.w6(32'h3ac004d2),
	.w7(32'h3a80c4a9),
	.w8(32'hb94af57a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c69f),
	.w1(32'h3b11f630),
	.w2(32'h3bceac54),
	.w3(32'hbbb01b7b),
	.w4(32'h3b84dceb),
	.w5(32'hbb06b0cf),
	.w6(32'h3b421db8),
	.w7(32'hbb543f24),
	.w8(32'h3c448120),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf751f),
	.w1(32'hba8ecda5),
	.w2(32'hbb7bc703),
	.w3(32'h39c950f3),
	.w4(32'hb72478c3),
	.w5(32'hb919a91b),
	.w6(32'hb7badd7b),
	.w7(32'h3a9f0c34),
	.w8(32'hba7fbb58),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98606cf),
	.w1(32'hbc16a372),
	.w2(32'h3ae1ee75),
	.w3(32'h3b8a2389),
	.w4(32'h3b8816b6),
	.w5(32'hbb53d940),
	.w6(32'h372184a2),
	.w7(32'hbb2b3022),
	.w8(32'h3acccc3c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad095e5),
	.w1(32'hba4574b4),
	.w2(32'h3847e542),
	.w3(32'h3bb8ecca),
	.w4(32'h3b14a674),
	.w5(32'h3b77975f),
	.w6(32'h3ad5723b),
	.w7(32'h3a83a96a),
	.w8(32'h391101f9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21fa79),
	.w1(32'h39c09730),
	.w2(32'hbad5d281),
	.w3(32'h3aaaa563),
	.w4(32'hb8bf91f5),
	.w5(32'h3b913589),
	.w6(32'hb9f4af2b),
	.w7(32'h3b0ed780),
	.w8(32'h3c083571),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24edd5),
	.w1(32'hbb5d40a7),
	.w2(32'h3bb151ee),
	.w3(32'h399d56b6),
	.w4(32'hbb57da89),
	.w5(32'h39a8dfab),
	.w6(32'hbb9eae48),
	.w7(32'h3b90c281),
	.w8(32'h3a07cc25),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdef78),
	.w1(32'h3a6e51e0),
	.w2(32'h3bcc74ac),
	.w3(32'h3a8054ee),
	.w4(32'h3ade30cf),
	.w5(32'hb8b88f82),
	.w6(32'hbadc6fde),
	.w7(32'h3c29b65d),
	.w8(32'hb98992c8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7feaba),
	.w1(32'hba8d4a0e),
	.w2(32'hba47c2dc),
	.w3(32'h3b656d22),
	.w4(32'hbb26d274),
	.w5(32'hba9a0cab),
	.w6(32'h3afe1759),
	.w7(32'h3b651524),
	.w8(32'hbb68ef3d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3241ea),
	.w1(32'h3a141d26),
	.w2(32'hbb3067aa),
	.w3(32'h3b04c288),
	.w4(32'hba4a8176),
	.w5(32'hbac2e58a),
	.w6(32'h3b5296b7),
	.w7(32'h3ae9bf3c),
	.w8(32'h3b14f6d0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8329f34),
	.w1(32'h3a8c72cc),
	.w2(32'hbc232c74),
	.w3(32'hbc4f6165),
	.w4(32'hb92d1047),
	.w5(32'hba529684),
	.w6(32'hbb75bb24),
	.w7(32'h3b933edb),
	.w8(32'h3c1d0285),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7130c),
	.w1(32'hb9262c32),
	.w2(32'hbac782cd),
	.w3(32'hbbabff4c),
	.w4(32'hbb09c206),
	.w5(32'hbc3ee1a0),
	.w6(32'h3a412f0d),
	.w7(32'h3bdff363),
	.w8(32'hbb103be6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe57592),
	.w1(32'hbb09e484),
	.w2(32'hbc972940),
	.w3(32'h3bb3e7f7),
	.w4(32'h3c4ece16),
	.w5(32'hba08651d),
	.w6(32'h3ad0806d),
	.w7(32'h3c7efe7e),
	.w8(32'h3ab8fe7f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ba4ac),
	.w1(32'h3c4416aa),
	.w2(32'hbaab5ea0),
	.w3(32'hbc10e1ac),
	.w4(32'hbc501f46),
	.w5(32'hbd4a9952),
	.w6(32'hbab21e1f),
	.w7(32'hba6f093f),
	.w8(32'hbbcd258e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d442c9a),
	.w1(32'h3c0f6466),
	.w2(32'h3b686913),
	.w3(32'hbb39b02a),
	.w4(32'hbc04ac43),
	.w5(32'hbbe32480),
	.w6(32'h3c42307d),
	.w7(32'h3c4395fc),
	.w8(32'hbbd0fd4f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb756c55),
	.w1(32'h3b9b4002),
	.w2(32'hbb8b9ec3),
	.w3(32'hbc847dfc),
	.w4(32'hbbae0a6b),
	.w5(32'h3bee0521),
	.w6(32'hbad9e67c),
	.w7(32'h3b39e8de),
	.w8(32'h3bfb2fb8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c532a0f),
	.w1(32'hb993fee5),
	.w2(32'hbb0abcae),
	.w3(32'h3abd50fb),
	.w4(32'hbc749253),
	.w5(32'h3c284f94),
	.w6(32'h3a253dae),
	.w7(32'hbc05d220),
	.w8(32'h3b78d0a9),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7622ec),
	.w1(32'h3bb05be4),
	.w2(32'hbbd017fe),
	.w3(32'h3ac9a878),
	.w4(32'hbbdf0cad),
	.w5(32'hba9ee4f8),
	.w6(32'hbab58362),
	.w7(32'hb7a262b2),
	.w8(32'hbaf7b4df),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1b15),
	.w1(32'h3cc820cb),
	.w2(32'hba57ca08),
	.w3(32'h3b81ea89),
	.w4(32'hbc2b33be),
	.w5(32'hbc55cde9),
	.w6(32'h3b405688),
	.w7(32'h3baeb45e),
	.w8(32'hbbd197a5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf34f05),
	.w1(32'h3a9e15d4),
	.w2(32'hbb40d7ff),
	.w3(32'hbaeca773),
	.w4(32'hbc29778e),
	.w5(32'hbb27bb46),
	.w6(32'hbb2ccabe),
	.w7(32'hba9399d2),
	.w8(32'hb9932d24),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d0c44),
	.w1(32'h3ad3e815),
	.w2(32'h3b9b54e2),
	.w3(32'hbbf509b3),
	.w4(32'hb5593653),
	.w5(32'hbc105a33),
	.w6(32'hbb00b3c6),
	.w7(32'h3d14d8ac),
	.w8(32'hb8c58573),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b0708),
	.w1(32'hbb875d86),
	.w2(32'hbbeb17a1),
	.w3(32'hbc767c25),
	.w4(32'hbc2c865e),
	.w5(32'h3c32fa0e),
	.w6(32'h3bd33111),
	.w7(32'hbba9a346),
	.w8(32'hbb637a0c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5fbfc),
	.w1(32'hba350a32),
	.w2(32'hba9efcc7),
	.w3(32'h3af48093),
	.w4(32'h3a7f06f1),
	.w5(32'h3b29aa59),
	.w6(32'h3826305f),
	.w7(32'hbc0fe24b),
	.w8(32'hbac51235),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8da27),
	.w1(32'h380410df),
	.w2(32'hbb4ff70e),
	.w3(32'hb894ec28),
	.w4(32'hbad6bf4c),
	.w5(32'h3c411198),
	.w6(32'h3d0474fd),
	.w7(32'hbba7c89a),
	.w8(32'h3b4ca0d7),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b072b05),
	.w1(32'hbc4b8074),
	.w2(32'h3bce888b),
	.w3(32'h3bec0d71),
	.w4(32'hbb872823),
	.w5(32'h3bafec5d),
	.w6(32'h3ae93df3),
	.w7(32'h3c7cf5c3),
	.w8(32'h3cc0c09f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceb4106),
	.w1(32'hba147852),
	.w2(32'hbbec3d50),
	.w3(32'h3b62a5a9),
	.w4(32'h3b21ef17),
	.w5(32'hbb8b1f00),
	.w6(32'h3b0e7846),
	.w7(32'h3b653377),
	.w8(32'h3aa5c0d9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aed6ed),
	.w1(32'h3aa9cbfa),
	.w2(32'h3c14fcec),
	.w3(32'hbad86e90),
	.w4(32'h3b4ad8b7),
	.w5(32'hbc120dfa),
	.w6(32'h3bd43fa7),
	.w7(32'h3b67c86a),
	.w8(32'h3a08bc6e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ec7ab),
	.w1(32'h3a473f9f),
	.w2(32'hbab066fc),
	.w3(32'hbb212a2a),
	.w4(32'h3a8cfe07),
	.w5(32'hbafa7728),
	.w6(32'hbb76d0e4),
	.w7(32'hbb6bece3),
	.w8(32'h3c055723),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h340f17a3),
	.w1(32'hbbfb831e),
	.w2(32'h3ad759c6),
	.w3(32'hbbc26b34),
	.w4(32'h3b92af71),
	.w5(32'h3bc10ef5),
	.w6(32'hbbf58807),
	.w7(32'h39f73ddf),
	.w8(32'hbb39eb9a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe30faa),
	.w1(32'h3ad15644),
	.w2(32'hbc393e51),
	.w3(32'h3c821676),
	.w4(32'hbafbeb27),
	.w5(32'h3af421e3),
	.w6(32'h3a1727c6),
	.w7(32'h3a1f533f),
	.w8(32'hbc40a1bf),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be702b5),
	.w1(32'h3c3d34d8),
	.w2(32'hbbfcb6dd),
	.w3(32'h3b46d9cb),
	.w4(32'h3bd28d37),
	.w5(32'h3bb3031c),
	.w6(32'hbb3b1429),
	.w7(32'hbbdecdac),
	.w8(32'hba596459),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a0eec),
	.w1(32'h3c5165ba),
	.w2(32'h3a867345),
	.w3(32'h3bd0b51c),
	.w4(32'hbc1e32af),
	.w5(32'h3c04e5b7),
	.w6(32'hbac1a773),
	.w7(32'h3c86cc18),
	.w8(32'hbb8f94cc),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cffac),
	.w1(32'hb918de7b),
	.w2(32'h3ad2a687),
	.w3(32'h3b126eee),
	.w4(32'h3c5c652f),
	.w5(32'hbb474b0e),
	.w6(32'hbb98ba2b),
	.w7(32'hbc35ebf1),
	.w8(32'h3c2ebcd2),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52d7a5),
	.w1(32'hbb57cd59),
	.w2(32'hbba26f02),
	.w3(32'hb8e5a0d6),
	.w4(32'hbbcaf134),
	.w5(32'hbae093ff),
	.w6(32'hbba78b86),
	.w7(32'hba2249a8),
	.w8(32'hb984667a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89ac30),
	.w1(32'h3c90b297),
	.w2(32'hbbb83e7a),
	.w3(32'hbb90d5e1),
	.w4(32'hbbadd2ed),
	.w5(32'hbc0f90b1),
	.w6(32'hbc03d50c),
	.w7(32'hbbee1236),
	.w8(32'h3c159c04),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e43c7),
	.w1(32'h3c464bb8),
	.w2(32'hbb5394cd),
	.w3(32'h3a78efe8),
	.w4(32'hbb86bc5c),
	.w5(32'hbbdca60b),
	.w6(32'h3b9c2807),
	.w7(32'hba98e929),
	.w8(32'hbb95fd3d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef06e4),
	.w1(32'h39c29fb2),
	.w2(32'hbb9cd80b),
	.w3(32'h3c53e21a),
	.w4(32'hbc3093e4),
	.w5(32'hbb770f89),
	.w6(32'h3c03b8be),
	.w7(32'hbbaf5718),
	.w8(32'hbaf00594),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6712e3),
	.w1(32'hbaa0b169),
	.w2(32'h3b8c4548),
	.w3(32'h3ae82ff4),
	.w4(32'hbbbe7cf9),
	.w5(32'h3b0ee1fe),
	.w6(32'hba481ce4),
	.w7(32'hbbe1ce75),
	.w8(32'hbad0aede),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7a0fe),
	.w1(32'h3a306b56),
	.w2(32'hbb6bfcc4),
	.w3(32'hbb7fee50),
	.w4(32'h3b0f79ca),
	.w5(32'h3a610288),
	.w6(32'hbb223655),
	.w7(32'hba867254),
	.w8(32'hb96b4468),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf36465),
	.w1(32'hbc21bde3),
	.w2(32'hbb1c198a),
	.w3(32'hbcb803e4),
	.w4(32'hba89b2d7),
	.w5(32'hbb23e011),
	.w6(32'hbc0f2b76),
	.w7(32'hba221941),
	.w8(32'hb9acf2eb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule