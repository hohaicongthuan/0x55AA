module layer_10_featuremap_377(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc382725),
	.w1(32'h3b495637),
	.w2(32'h3cb1a990),
	.w3(32'hbad8aea4),
	.w4(32'hbada6d93),
	.w5(32'h3bea4038),
	.w6(32'h3c1741c7),
	.w7(32'h3b788b49),
	.w8(32'hbbcbfdda),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3a5f5),
	.w1(32'h3bbd8d56),
	.w2(32'hbb0b8850),
	.w3(32'hbb85d2ce),
	.w4(32'hbbe0cd3c),
	.w5(32'hb82b082e),
	.w6(32'h3b995b96),
	.w7(32'h3b871117),
	.w8(32'h3b0bfbfd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86002d),
	.w1(32'hbaa63c35),
	.w2(32'hbc39d6c1),
	.w3(32'hbc73d9af),
	.w4(32'hbb900594),
	.w5(32'hbc1e1777),
	.w6(32'hbc1fdc4c),
	.w7(32'hbb38d25b),
	.w8(32'hbc09a3b3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cd16e),
	.w1(32'hbcc569d5),
	.w2(32'h3c49dabb),
	.w3(32'hbaa26f9d),
	.w4(32'h3bd301e9),
	.w5(32'h3c787d92),
	.w6(32'hbc25a50c),
	.w7(32'h3bf3ac9d),
	.w8(32'h3c3b6939),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01794e),
	.w1(32'h391f2edd),
	.w2(32'hbc069024),
	.w3(32'hba2148ee),
	.w4(32'h3ba51587),
	.w5(32'h3a6d597a),
	.w6(32'hbbed1b42),
	.w7(32'hb98b3b22),
	.w8(32'hbc50b2e7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16038e),
	.w1(32'hbbece795),
	.w2(32'hbbb39841),
	.w3(32'hbbf9a2e8),
	.w4(32'h3b61acfb),
	.w5(32'h3c4cdbf4),
	.w6(32'hbb5d1784),
	.w7(32'hbc50c471),
	.w8(32'h3c50c279),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e7b22),
	.w1(32'hbbc064b1),
	.w2(32'h3bf9b960),
	.w3(32'hbc8af23f),
	.w4(32'hbc44399e),
	.w5(32'hbb46a865),
	.w6(32'hbb64452b),
	.w7(32'hbc80244e),
	.w8(32'hbbdaabe8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398806ee),
	.w1(32'hbc5b7041),
	.w2(32'h3b9dcb6c),
	.w3(32'hbaa7e5c4),
	.w4(32'h3b995a75),
	.w5(32'h3960ed3d),
	.w6(32'h3c3c8b2e),
	.w7(32'h3a2cbbe4),
	.w8(32'hbba484c9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b0a43),
	.w1(32'hbaf95d08),
	.w2(32'h3c8411c6),
	.w3(32'hbba056dc),
	.w4(32'hbbe9109b),
	.w5(32'hbc5d05eb),
	.w6(32'h3c2f7378),
	.w7(32'h3bbccdc3),
	.w8(32'hbb402e49),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc120c3),
	.w1(32'h3b081b2a),
	.w2(32'hbb13903b),
	.w3(32'h3c14454b),
	.w4(32'hbc4300cd),
	.w5(32'hbab4c9e9),
	.w6(32'hbc15d6ae),
	.w7(32'hbba217d2),
	.w8(32'hba7d03e2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61a0e2),
	.w1(32'h3c9a5c1a),
	.w2(32'hbbcd4c28),
	.w3(32'hbbbe2d0e),
	.w4(32'h3a064f74),
	.w5(32'h3b8e44b8),
	.w6(32'h3c3ab086),
	.w7(32'hbb367105),
	.w8(32'hbb1d5a2b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03d9dc),
	.w1(32'hba514eca),
	.w2(32'hbb603774),
	.w3(32'h39d30003),
	.w4(32'hbaa9c9ee),
	.w5(32'h3b3418bd),
	.w6(32'hbbb713aa),
	.w7(32'h39d926ac),
	.w8(32'hbb55736c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa8190),
	.w1(32'h3c4ae564),
	.w2(32'h3b05072a),
	.w3(32'h3ba61565),
	.w4(32'h3c327485),
	.w5(32'h3cbfedcb),
	.w6(32'hbc4b229e),
	.w7(32'h3bb10b30),
	.w8(32'hbc08f028),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fbe04),
	.w1(32'h3b923c93),
	.w2(32'hbd0d204d),
	.w3(32'hbb8c6d78),
	.w4(32'h3bb9d656),
	.w5(32'h371f8a70),
	.w6(32'hbb6465f4),
	.w7(32'hbb2499e0),
	.w8(32'h3c272946),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe71376),
	.w1(32'h39867478),
	.w2(32'hbb731715),
	.w3(32'h3ab7fff4),
	.w4(32'hbb357bd8),
	.w5(32'h3c28e9d1),
	.w6(32'hbc6d361d),
	.w7(32'hbb7bf760),
	.w8(32'h3a923e78),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caef660),
	.w1(32'h3b842320),
	.w2(32'hbae4bbbd),
	.w3(32'hb99f84a2),
	.w4(32'h3b2ae8af),
	.w5(32'h3c16fabc),
	.w6(32'h3b8763bc),
	.w7(32'hbbd9fd1f),
	.w8(32'hbb8df6af),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97efa0),
	.w1(32'h3c1c0110),
	.w2(32'hbc34b543),
	.w3(32'h3b425b96),
	.w4(32'h39b2dfb2),
	.w5(32'hbb1ee2f0),
	.w6(32'hbbef01d9),
	.w7(32'h3c6fbc5f),
	.w8(32'hbb69ea10),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c431543),
	.w1(32'h3bdabfc9),
	.w2(32'hbc30b160),
	.w3(32'hbc6842af),
	.w4(32'hbbe6f7ab),
	.w5(32'h3bd660b1),
	.w6(32'h3bcded4a),
	.w7(32'hba9d31d6),
	.w8(32'h3be3fe8f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11fa9c),
	.w1(32'hbb6a3559),
	.w2(32'h3c3c8d5c),
	.w3(32'hbc1165a6),
	.w4(32'h3beba16d),
	.w5(32'hbc3f9eec),
	.w6(32'hbc4bdc0e),
	.w7(32'h3c5aba6f),
	.w8(32'hbc2075c1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38472b),
	.w1(32'hbbbbaa42),
	.w2(32'h3c08ee20),
	.w3(32'hbc285fe7),
	.w4(32'hbb168d27),
	.w5(32'h3bafa47d),
	.w6(32'hbc807714),
	.w7(32'hbaba4a7f),
	.w8(32'h3baf1115),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b7e3),
	.w1(32'h3bb252d7),
	.w2(32'h3c915447),
	.w3(32'h3c065248),
	.w4(32'hbbe2eeef),
	.w5(32'hbbb6d5bd),
	.w6(32'hbb97c9fe),
	.w7(32'h3b19f821),
	.w8(32'hbb9a6440),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcecde4),
	.w1(32'hbbbdbb23),
	.w2(32'h3b9fe049),
	.w3(32'hbb38652d),
	.w4(32'h3b2cda3b),
	.w5(32'hbca8e90c),
	.w6(32'h3b3e95ff),
	.w7(32'h3a924273),
	.w8(32'hbad5003f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb3fc3),
	.w1(32'h3a059840),
	.w2(32'h3c75a214),
	.w3(32'h3ac6a2fb),
	.w4(32'h3a951ccc),
	.w5(32'hbc1ececb),
	.w6(32'hba385659),
	.w7(32'hbc776102),
	.w8(32'hbb70f46d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e7684),
	.w1(32'h3ac9be09),
	.w2(32'h3c1377f9),
	.w3(32'hb9978889),
	.w4(32'hba6e2e5d),
	.w5(32'hbb59dcab),
	.w6(32'hbc50fa4b),
	.w7(32'hbbabdac5),
	.w8(32'h3c1a747d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c1ab9),
	.w1(32'h3a2dbebe),
	.w2(32'h3c6ef6a8),
	.w3(32'hbc60457f),
	.w4(32'h39324d13),
	.w5(32'h3ceb53bd),
	.w6(32'hbbd76c59),
	.w7(32'hbb943fbd),
	.w8(32'h3b40b45f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817550),
	.w1(32'h3b44a0aa),
	.w2(32'hbadd554d),
	.w3(32'h3c3cdd20),
	.w4(32'h3c351c77),
	.w5(32'h3b83a76c),
	.w6(32'h3a3a8080),
	.w7(32'h3c5efc56),
	.w8(32'hbb0c0830),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15fb21),
	.w1(32'hbc21bb10),
	.w2(32'hbb34ef5a),
	.w3(32'h3cbb7c9c),
	.w4(32'hbba491b2),
	.w5(32'hba89702e),
	.w6(32'h3c8b0bf9),
	.w7(32'hbbe153ed),
	.w8(32'h3b5af97b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08081),
	.w1(32'h3c94b175),
	.w2(32'h3c9a5883),
	.w3(32'h3c8edcda),
	.w4(32'hbc9c45a8),
	.w5(32'h3bc2ff76),
	.w6(32'h3c189e24),
	.w7(32'hbb81e7cf),
	.w8(32'hbaa88e7e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adeaf1),
	.w1(32'hba8d19d9),
	.w2(32'h3cc79526),
	.w3(32'h3c9a68b4),
	.w4(32'h3b9334d2),
	.w5(32'hbb38e217),
	.w6(32'hbbe71007),
	.w7(32'hbb1d9149),
	.w8(32'hbbdb33a8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c0fdd),
	.w1(32'h3c7dd049),
	.w2(32'h3c1c069c),
	.w3(32'hbbf3f9d1),
	.w4(32'hbc12366c),
	.w5(32'hbb1b7b51),
	.w6(32'h3d042c88),
	.w7(32'h3b8e76c8),
	.w8(32'hbb0856b7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c9b72),
	.w1(32'h3b105538),
	.w2(32'h3ba7bfea),
	.w3(32'hbcaf730d),
	.w4(32'h3bf03a5a),
	.w5(32'h3b9d70c5),
	.w6(32'hbb124f17),
	.w7(32'h3bd4ddd7),
	.w8(32'h3bd7dc14),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ead45),
	.w1(32'hbb0e00c1),
	.w2(32'h3c23c90b),
	.w3(32'hbbb7429f),
	.w4(32'h3bddcd76),
	.w5(32'h3cf68b4e),
	.w6(32'hb9f513e0),
	.w7(32'h3aa2ae89),
	.w8(32'hbaa9d705),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17faa6),
	.w1(32'hbbfe7ece),
	.w2(32'h3bccef75),
	.w3(32'hbc366edf),
	.w4(32'h3c145eb1),
	.w5(32'h3b1b6e53),
	.w6(32'hbc0e0410),
	.w7(32'h3c7f0a7c),
	.w8(32'h3c197b87),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d9675),
	.w1(32'h3c8a3a57),
	.w2(32'h3b440943),
	.w3(32'hbc24839a),
	.w4(32'hbc53ec04),
	.w5(32'h3cb974d8),
	.w6(32'h3ba0a642),
	.w7(32'hbab5e3c0),
	.w8(32'hbbeeea52),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba782ca),
	.w1(32'hbb9dc2ff),
	.w2(32'h3b4a514d),
	.w3(32'hbb4d46fc),
	.w4(32'h3bb942c8),
	.w5(32'h3c92cc68),
	.w6(32'h39b6176d),
	.w7(32'h3c9feff5),
	.w8(32'h3d153275),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc288c17),
	.w1(32'h39dd3876),
	.w2(32'hbc97b9a4),
	.w3(32'h3c6afa45),
	.w4(32'hbb949155),
	.w5(32'h3ca6d7c4),
	.w6(32'h3b3f8707),
	.w7(32'hbba00179),
	.w8(32'h3c99e61b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf43c),
	.w1(32'h3bb8268c),
	.w2(32'hbc04e806),
	.w3(32'h3a64c18c),
	.w4(32'h3c7555f7),
	.w5(32'h3b4e249a),
	.w6(32'h3b480f8a),
	.w7(32'h3cae1087),
	.w8(32'h3c638423),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d75815),
	.w1(32'h3b8a3f65),
	.w2(32'h3d115cb6),
	.w3(32'h3c8b6359),
	.w4(32'h3c8e7f88),
	.w5(32'hbbbb006c),
	.w6(32'hbad0e36e),
	.w7(32'h3c40bb94),
	.w8(32'hbb38392e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9402477),
	.w1(32'h3cfed36e),
	.w2(32'h3a198e0c),
	.w3(32'h3b0c380b),
	.w4(32'h3c1d490e),
	.w5(32'h3cb30067),
	.w6(32'hbb98d5de),
	.w7(32'h3c5f07f3),
	.w8(32'hbc119c53),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bce93),
	.w1(32'h3b6980e5),
	.w2(32'h3b081019),
	.w3(32'hbb8ee0f6),
	.w4(32'h3b842b78),
	.w5(32'h3c19cbcb),
	.w6(32'hbc363f89),
	.w7(32'hb95eb525),
	.w8(32'hbbe6f879),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17d807),
	.w1(32'h3cfc39c3),
	.w2(32'h39da22a5),
	.w3(32'hbbc2ca8a),
	.w4(32'h3be052ed),
	.w5(32'hbba8f15f),
	.w6(32'hba8313b4),
	.w7(32'h3aa0b1ae),
	.w8(32'h3b98ed9b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e675e),
	.w1(32'hbbba6afc),
	.w2(32'h3b3fd0fe),
	.w3(32'hba8ca6b2),
	.w4(32'h3bba5834),
	.w5(32'h3b046194),
	.w6(32'hbb0bab18),
	.w7(32'hbba084ff),
	.w8(32'h3c2b6e91),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecfe09),
	.w1(32'h3b3a3483),
	.w2(32'hbc338e3b),
	.w3(32'h3c88b6dd),
	.w4(32'h3bd79f76),
	.w5(32'h3b81eeb2),
	.w6(32'h3cad6459),
	.w7(32'hbbc5c318),
	.w8(32'h3c3e521d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3b666),
	.w1(32'hbb398bf9),
	.w2(32'hbb018969),
	.w3(32'h3ab4f9af),
	.w4(32'h3b82ed1e),
	.w5(32'hbb0f0993),
	.w6(32'h3a93537c),
	.w7(32'hbabe3387),
	.w8(32'hbb885109),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b65bc),
	.w1(32'h3c53a946),
	.w2(32'h3c58cc2f),
	.w3(32'h3b920a07),
	.w4(32'h3cabc4b4),
	.w5(32'h3c417668),
	.w6(32'h3be71abd),
	.w7(32'h3c99b92d),
	.w8(32'h398e4880),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb7b9a),
	.w1(32'h3b9840aa),
	.w2(32'h3c19a13a),
	.w3(32'hb9bd294c),
	.w4(32'hbb97aa78),
	.w5(32'h3cfb947f),
	.w6(32'h3c1e5a1d),
	.w7(32'hbc63ea49),
	.w8(32'h3cb1d5cb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b8129),
	.w1(32'h3aa6cad4),
	.w2(32'hbb1b8305),
	.w3(32'h3c621848),
	.w4(32'h3c09cb3a),
	.w5(32'hbaad582b),
	.w6(32'hbadf5ed5),
	.w7(32'h3b9ba869),
	.w8(32'hbac018cb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ecb8a),
	.w1(32'h3bab7834),
	.w2(32'h3ae874f1),
	.w3(32'h3c478b5e),
	.w4(32'hbb9bd227),
	.w5(32'h3982d9ff),
	.w6(32'hbb301f2c),
	.w7(32'h3b922ee9),
	.w8(32'h3cf8acaa),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6831ab),
	.w1(32'hb8b80756),
	.w2(32'h3c040fb9),
	.w3(32'hbbf633f6),
	.w4(32'hbba491ea),
	.w5(32'h3b1d4930),
	.w6(32'h3b775265),
	.w7(32'hbb150ff9),
	.w8(32'hbc519fe2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19f472),
	.w1(32'h3aef6085),
	.w2(32'h3d07ec39),
	.w3(32'h3c89bf99),
	.w4(32'h3bd5abff),
	.w5(32'hbb6b3231),
	.w6(32'hbc6a6d3a),
	.w7(32'h3b33c9ee),
	.w8(32'h3bdfb9b7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b561d4d),
	.w1(32'h3bac0b83),
	.w2(32'hba3011aa),
	.w3(32'hbc3118d4),
	.w4(32'h3bf1bec2),
	.w5(32'h3a435e63),
	.w6(32'h3cea1f80),
	.w7(32'h3b48517e),
	.w8(32'hbba2c462),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb0c8b),
	.w1(32'h3bcec78d),
	.w2(32'hbb7cf827),
	.w3(32'h3becc03c),
	.w4(32'h3cf6c624),
	.w5(32'h3b7a3e0d),
	.w6(32'hbc6fc354),
	.w7(32'hbb77a17c),
	.w8(32'hb87ade2a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf0d41),
	.w1(32'hb99efbf8),
	.w2(32'hbbdad9c9),
	.w3(32'hbbd89a8e),
	.w4(32'hbbe664d8),
	.w5(32'h3c03974e),
	.w6(32'hbbfe1bc5),
	.w7(32'hbb27e838),
	.w8(32'h3c632e62),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c374cc6),
	.w1(32'h3d2a7395),
	.w2(32'hbc672450),
	.w3(32'h3b861191),
	.w4(32'h3c04a565),
	.w5(32'hbb0fa223),
	.w6(32'h3bd22e45),
	.w7(32'h3be0d1ec),
	.w8(32'h3b099db1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fa65d),
	.w1(32'hb867b3df),
	.w2(32'h3c79e676),
	.w3(32'h3bb6edf9),
	.w4(32'hbc00e749),
	.w5(32'hbc8f5889),
	.w6(32'h3c3ed581),
	.w7(32'hba14ca17),
	.w8(32'h3c11fc0d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce2e5d),
	.w1(32'h3c2fc921),
	.w2(32'h3c471feb),
	.w3(32'h3c68834f),
	.w4(32'hbb3cfc28),
	.w5(32'hbc2a9787),
	.w6(32'hba406608),
	.w7(32'hbc223e37),
	.w8(32'h3b2155c7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc325f0),
	.w1(32'h3bae6727),
	.w2(32'h3b64b9bb),
	.w3(32'hbcdb3066),
	.w4(32'hbc3e9e27),
	.w5(32'hbc29371a),
	.w6(32'h3b94bee3),
	.w7(32'h3c3ab040),
	.w8(32'hb813c9d7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1043d),
	.w1(32'hbc33707f),
	.w2(32'hbace15ab),
	.w3(32'h3ad1c51b),
	.w4(32'hbc833c01),
	.w5(32'h3a55b539),
	.w6(32'hbc81a780),
	.w7(32'h3ca04e84),
	.w8(32'h3bccf120),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b20ab),
	.w1(32'hbbaf26b9),
	.w2(32'hbbb5c23d),
	.w3(32'hbbd76af9),
	.w4(32'hbc71321e),
	.w5(32'hbbd913f6),
	.w6(32'h3c8b726c),
	.w7(32'h3b880c2a),
	.w8(32'hbad91138),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4b1a4),
	.w1(32'hbbb8a249),
	.w2(32'hbc0d92ca),
	.w3(32'h3c14ba7f),
	.w4(32'h3c32b381),
	.w5(32'hbc58f394),
	.w6(32'hbc4e1ca6),
	.w7(32'h3cf3cc25),
	.w8(32'h3c8bb8e3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf84505),
	.w1(32'hbc352877),
	.w2(32'hbc9b07c7),
	.w3(32'hbc653755),
	.w4(32'h3afcfbde),
	.w5(32'hbc155b6c),
	.w6(32'h3c5bc0f2),
	.w7(32'hbb337cc3),
	.w8(32'h3ce47e09),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b015c15),
	.w1(32'h3c1093fc),
	.w2(32'h3afa5b9a),
	.w3(32'h3cf2271b),
	.w4(32'hbb0b2bf2),
	.w5(32'h3c29d509),
	.w6(32'h3b9f7260),
	.w7(32'hbc5cd06a),
	.w8(32'hba88d3a2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d4c24),
	.w1(32'h3b313f6d),
	.w2(32'h3c7ca200),
	.w3(32'hb904365d),
	.w4(32'h3c1bf62d),
	.w5(32'h3c6ed5bb),
	.w6(32'hbcf08a9d),
	.w7(32'hbbe33b73),
	.w8(32'hbc0f3fd6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71b61d),
	.w1(32'h3c987345),
	.w2(32'hbbf128dc),
	.w3(32'hbad49b7c),
	.w4(32'hbc364f0f),
	.w5(32'h3ba50937),
	.w6(32'h3c63bf2a),
	.w7(32'h3ba950af),
	.w8(32'hbc08046d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc3f23),
	.w1(32'h3bb84ce7),
	.w2(32'hbbb4f391),
	.w3(32'hbc021133),
	.w4(32'hb9e8fd20),
	.w5(32'hbbf1bd09),
	.w6(32'hbb4c8b49),
	.w7(32'hbbcca315),
	.w8(32'hbaf4c0b2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e458f),
	.w1(32'hbc59dd01),
	.w2(32'h3aa4827a),
	.w3(32'h3a6948e5),
	.w4(32'hbb3c8c12),
	.w5(32'hbc010fa5),
	.w6(32'hbbc318af),
	.w7(32'hbbbb92a1),
	.w8(32'h3c8c06ef),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cf6d9),
	.w1(32'h3b9015c2),
	.w2(32'h3a8c8463),
	.w3(32'h3a8727b9),
	.w4(32'h3a082fbe),
	.w5(32'h3b511407),
	.w6(32'h37d0d8c1),
	.w7(32'hbc3ff4f7),
	.w8(32'h3ba84e30),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e5917),
	.w1(32'h3b8c48d2),
	.w2(32'h3ac74a08),
	.w3(32'hbbed029b),
	.w4(32'h3ac8a4c2),
	.w5(32'h3c353dbb),
	.w6(32'hba25c00e),
	.w7(32'hbbc9d782),
	.w8(32'h3ba17564),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffaa13),
	.w1(32'hbc4c3a2a),
	.w2(32'h3b0c84b3),
	.w3(32'hbb2b9baf),
	.w4(32'hb9fe05fa),
	.w5(32'hbccca06c),
	.w6(32'hba844901),
	.w7(32'hbc299333),
	.w8(32'hbbee6c0a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b593862),
	.w1(32'h3ba6c046),
	.w2(32'hbc7f5991),
	.w3(32'hbb595942),
	.w4(32'h3afd5073),
	.w5(32'hbc091621),
	.w6(32'h3c47485e),
	.w7(32'h3b40aa28),
	.w8(32'h3b812e72),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc201192),
	.w1(32'hbbf25488),
	.w2(32'hbc721d4c),
	.w3(32'h3c25870a),
	.w4(32'hbb327fdd),
	.w5(32'h3c0233fa),
	.w6(32'hbc341324),
	.w7(32'h3cd12b91),
	.w8(32'hbc26acc3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba24d0b),
	.w1(32'hbc0308a9),
	.w2(32'h3cbdc1f0),
	.w3(32'h3c8c2f18),
	.w4(32'h3c24dcb2),
	.w5(32'h3b0450ea),
	.w6(32'h3c4d0cd4),
	.w7(32'h3aa61eca),
	.w8(32'hbbd94800),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9dba3),
	.w1(32'hb9c005ce),
	.w2(32'h39ecab15),
	.w3(32'h3ba700d5),
	.w4(32'hbb937d7e),
	.w5(32'hbb07c6ed),
	.w6(32'h3b9a800c),
	.w7(32'hbc048e30),
	.w8(32'hbbd7b672),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8548e1),
	.w1(32'h3929eeb2),
	.w2(32'hbb3cf3e4),
	.w3(32'h3c238577),
	.w4(32'hb969bace),
	.w5(32'h3b185b9e),
	.w6(32'h3c15fd57),
	.w7(32'h3b607ed7),
	.w8(32'h3b84fa0a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfa0e73),
	.w1(32'hba4b26db),
	.w2(32'hbb1c0b5c),
	.w3(32'hbc1e3d58),
	.w4(32'hb8fd1583),
	.w5(32'hbb2b04f2),
	.w6(32'h3bed440f),
	.w7(32'hbaa422e3),
	.w8(32'h3c15ec1f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a083e),
	.w1(32'hbbd04526),
	.w2(32'hbb71bbab),
	.w3(32'h3b29479e),
	.w4(32'h3c72c881),
	.w5(32'hbc0147ab),
	.w6(32'h3b61e940),
	.w7(32'h3c0d859d),
	.w8(32'hbc095524),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e3d7d),
	.w1(32'hbbea4f46),
	.w2(32'h3a48a2c6),
	.w3(32'h3c092cbf),
	.w4(32'h3b8726a5),
	.w5(32'h3b17f848),
	.w6(32'hba6bc6d7),
	.w7(32'hbb357e04),
	.w8(32'hb824d9e4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd40c9b),
	.w1(32'h3cbe072c),
	.w2(32'h3bdfec1d),
	.w3(32'h3b91e97c),
	.w4(32'h3c232c4f),
	.w5(32'h3c48acbd),
	.w6(32'hbb8da792),
	.w7(32'hbb5ac3d4),
	.w8(32'hba5f60b8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50e6f8),
	.w1(32'h3bec355f),
	.w2(32'hbc364b11),
	.w3(32'hbc840d3e),
	.w4(32'h3ab4dfb2),
	.w5(32'hbc34ec45),
	.w6(32'hbc3d2b23),
	.w7(32'hbbbc2155),
	.w8(32'hbbd779f5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0fd7d),
	.w1(32'h3bfcd1a6),
	.w2(32'hbc710472),
	.w3(32'h3af471f3),
	.w4(32'hbc9370b0),
	.w5(32'h3b6758a7),
	.w6(32'hb8337f01),
	.w7(32'hbc271e2f),
	.w8(32'h3c3c691e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7aeba0),
	.w1(32'h3a8b1d1a),
	.w2(32'hbc1c6130),
	.w3(32'h3b04a1ea),
	.w4(32'h3c86d487),
	.w5(32'hbc62436d),
	.w6(32'h3bf53cd1),
	.w7(32'hbb7c96b1),
	.w8(32'hbb0547ee),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd506f2),
	.w1(32'h3c04b58e),
	.w2(32'hbb5d8473),
	.w3(32'hbb221f53),
	.w4(32'hbbd20397),
	.w5(32'hbc30a657),
	.w6(32'hbc6667bf),
	.w7(32'hba227340),
	.w8(32'h3bf17dcf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7fb5d),
	.w1(32'hba2cf30f),
	.w2(32'h3a82926b),
	.w3(32'hba9d9ec1),
	.w4(32'hbb01a044),
	.w5(32'h3bcf5cf1),
	.w6(32'hbc50294a),
	.w7(32'hb92ba96d),
	.w8(32'hbc560a23),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2e3a2),
	.w1(32'hbb8dfa66),
	.w2(32'hba367edf),
	.w3(32'hba043a05),
	.w4(32'hbc3f94da),
	.w5(32'h3baebefb),
	.w6(32'h3acaa6e6),
	.w7(32'h3bc8e083),
	.w8(32'h3bbd6e3b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9bdce),
	.w1(32'hbaccbfb7),
	.w2(32'hbc2ac7e3),
	.w3(32'h3c7d7ab8),
	.w4(32'hbc5aab49),
	.w5(32'h3b1a4f81),
	.w6(32'h3c0a315f),
	.w7(32'hbad14f83),
	.w8(32'h3bc6a3b1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3da3b2),
	.w1(32'h3cb3e66e),
	.w2(32'hbc0adf3b),
	.w3(32'hbc44bbc2),
	.w4(32'hba3f1838),
	.w5(32'hbc3e3124),
	.w6(32'hbbb8cad8),
	.w7(32'h3b220204),
	.w8(32'hba2b27e2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb9238),
	.w1(32'hbc947716),
	.w2(32'hbc26cafc),
	.w3(32'h3d14b88b),
	.w4(32'hbbb1838f),
	.w5(32'h3c58c449),
	.w6(32'h3b8a708b),
	.w7(32'h3bff01a8),
	.w8(32'hbcf98127),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850263),
	.w1(32'hba34faf8),
	.w2(32'h3b5702db),
	.w3(32'hbb252e66),
	.w4(32'h3bd375d1),
	.w5(32'h3c133839),
	.w6(32'hbc42df7f),
	.w7(32'hbc244beb),
	.w8(32'h3cde8131),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c804b78),
	.w1(32'h3c77e7c0),
	.w2(32'h3c4c56c7),
	.w3(32'h3a0c7460),
	.w4(32'hbc92fce1),
	.w5(32'hbb64c9e6),
	.w6(32'hb9a6b3df),
	.w7(32'hbc68e546),
	.w8(32'hbc355171),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25ed44),
	.w1(32'h3ac1e74b),
	.w2(32'hba283032),
	.w3(32'h3c316e0d),
	.w4(32'hbb656c50),
	.w5(32'h3c9ed0ef),
	.w6(32'h3b942f1b),
	.w7(32'h3a0dd929),
	.w8(32'hbb800e14),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d1959),
	.w1(32'hbc4e99a6),
	.w2(32'hbab59ed0),
	.w3(32'h3ba7438b),
	.w4(32'h3bb5a090),
	.w5(32'h3b49ccf4),
	.w6(32'hbc77bea9),
	.w7(32'hbc2162b4),
	.w8(32'h3b96ce40),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89741b),
	.w1(32'hbad0a988),
	.w2(32'hbae8bc56),
	.w3(32'h3cd9ba1c),
	.w4(32'h3c6ad898),
	.w5(32'hba23de7a),
	.w6(32'hbc09d1bf),
	.w7(32'h3ba1b4e5),
	.w8(32'hbbe7cbea),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b808d6c),
	.w1(32'h3c33846d),
	.w2(32'h3c048ba2),
	.w3(32'h3c3bc3fc),
	.w4(32'h3bc1da56),
	.w5(32'hbbd60297),
	.w6(32'h3c0fd5f6),
	.w7(32'hbbff7646),
	.w8(32'hbbacdc55),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03fabc),
	.w1(32'hbb6226ef),
	.w2(32'h3b01a217),
	.w3(32'hbbbdbef6),
	.w4(32'h3b6a52cb),
	.w5(32'h3b0afe92),
	.w6(32'hbc6cf1f0),
	.w7(32'hbc3c693a),
	.w8(32'hbc13c7f4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc618037),
	.w1(32'hbbed85fd),
	.w2(32'h3a92a87e),
	.w3(32'hbb04908f),
	.w4(32'h3bcaccaf),
	.w5(32'hbc162b61),
	.w6(32'hb967572c),
	.w7(32'h3b386852),
	.w8(32'hbc9ff947),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc446458),
	.w1(32'hbbacdc51),
	.w2(32'hbab3f668),
	.w3(32'hbbd3cea1),
	.w4(32'h3c6e44e8),
	.w5(32'hbb687045),
	.w6(32'h3c48fe07),
	.w7(32'hbc6b8e92),
	.w8(32'h3b9693f7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4710df),
	.w1(32'h3a4c3f1b),
	.w2(32'h3c455d5c),
	.w3(32'h3c0e6cf9),
	.w4(32'hbb127878),
	.w5(32'hbc9889d6),
	.w6(32'hbbb369de),
	.w7(32'h3abe7cfd),
	.w8(32'hb9fbf7b7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf61760),
	.w1(32'hbccfee76),
	.w2(32'h3bbc6cb4),
	.w3(32'hbb86c76a),
	.w4(32'hbc0523e2),
	.w5(32'h39b56d6e),
	.w6(32'hbc508da2),
	.w7(32'hbb3b0003),
	.w8(32'h3b24d15c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c771c),
	.w1(32'hbcf86700),
	.w2(32'hbc60ded2),
	.w3(32'h3c1124a5),
	.w4(32'hbc7b5ec6),
	.w5(32'h3bd6281f),
	.w6(32'h3b26b73b),
	.w7(32'hbab50a65),
	.w8(32'hbc957c41),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90d38b),
	.w1(32'h3c5babc6),
	.w2(32'h3bf0d9cd),
	.w3(32'h3a504c65),
	.w4(32'hbb131083),
	.w5(32'h3cee76de),
	.w6(32'h3c60e891),
	.w7(32'hbc1d53c8),
	.w8(32'hbbfd656b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb932a),
	.w1(32'h3c86de15),
	.w2(32'h3c2376fb),
	.w3(32'h3b8cfa78),
	.w4(32'hbb5d0943),
	.w5(32'hbb49c7a9),
	.w6(32'h3b64fee6),
	.w7(32'hbb353d25),
	.w8(32'h3c07195a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdae8b2),
	.w1(32'h3be59641),
	.w2(32'h3b2544c0),
	.w3(32'h3b0ac4bb),
	.w4(32'hba80d757),
	.w5(32'h3a273a23),
	.w6(32'hbc0aa754),
	.w7(32'h3c6acf35),
	.w8(32'hbb5c0a94),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fafcc),
	.w1(32'h3b0f11aa),
	.w2(32'hbcabd959),
	.w3(32'hbc83d387),
	.w4(32'hbb3ff788),
	.w5(32'h3c6c94b6),
	.w6(32'hbbf38508),
	.w7(32'h3bc4c2a7),
	.w8(32'hbb9f50bd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393118ae),
	.w1(32'h3d1082cf),
	.w2(32'h3cab60e5),
	.w3(32'h3b9374c9),
	.w4(32'hbb7d0771),
	.w5(32'h3a2db28c),
	.w6(32'h3ad74131),
	.w7(32'h3ba0bd5b),
	.w8(32'hbb218b72),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42cb59),
	.w1(32'h3c31a21e),
	.w2(32'h3c1f4579),
	.w3(32'h3c482342),
	.w4(32'hbc9a7268),
	.w5(32'hbc629758),
	.w6(32'h3c4fcec6),
	.w7(32'h3caafc9e),
	.w8(32'hbc12e36a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29000c),
	.w1(32'h3c0ae106),
	.w2(32'hbc198085),
	.w3(32'h3c1143a2),
	.w4(32'h3bfd3025),
	.w5(32'h3b645481),
	.w6(32'h3a5bef35),
	.w7(32'hb983d402),
	.w8(32'hbc5dca80),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb5c8d),
	.w1(32'hbc6790f4),
	.w2(32'hbbd116b2),
	.w3(32'hbc63b886),
	.w4(32'h3c0258b5),
	.w5(32'hbb1df1c3),
	.w6(32'h3d12f51e),
	.w7(32'h3b283893),
	.w8(32'h3b308090),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6d5b2),
	.w1(32'h3bbe5449),
	.w2(32'hb9c7eb9b),
	.w3(32'hbb99808c),
	.w4(32'hbac4655f),
	.w5(32'h3bb08854),
	.w6(32'h3c39c4bd),
	.w7(32'hba86d4a1),
	.w8(32'h3af0fdfc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b3e2e),
	.w1(32'h3a60a810),
	.w2(32'h3cb807d0),
	.w3(32'hbcabd09f),
	.w4(32'hbad1244a),
	.w5(32'h3c8990d0),
	.w6(32'hbc47498d),
	.w7(32'hbc1b8acc),
	.w8(32'h3c0cd653),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a327b),
	.w1(32'hbadb5fc9),
	.w2(32'hbcc4d893),
	.w3(32'h3b7a7f3b),
	.w4(32'h3c259b2c),
	.w5(32'h3c3f5de7),
	.w6(32'hba89e155),
	.w7(32'hbc3157f6),
	.w8(32'hbc5f3d86),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb753a0e),
	.w1(32'h3c2bd328),
	.w2(32'hbc1f1f02),
	.w3(32'h3c7456d5),
	.w4(32'h3a0e7484),
	.w5(32'hba9c2b78),
	.w6(32'hbba86fe1),
	.w7(32'hbc566aa1),
	.w8(32'h38f48bd8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0b5391),
	.w1(32'h3c6970e0),
	.w2(32'h3c5265a1),
	.w3(32'h3bbcf2ce),
	.w4(32'h3c240ee8),
	.w5(32'hba8b3b7a),
	.w6(32'h3bb95a31),
	.w7(32'h3bf57058),
	.w8(32'h3bec0d4a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe6d6e),
	.w1(32'hbb2da113),
	.w2(32'h3bc9de06),
	.w3(32'h3b4812c1),
	.w4(32'h3bb7a689),
	.w5(32'hbc1a15d3),
	.w6(32'hbb22a7b7),
	.w7(32'h3b516137),
	.w8(32'h3b849c24),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e3b92),
	.w1(32'hbaffd7e8),
	.w2(32'hbb258922),
	.w3(32'hbc5506ab),
	.w4(32'h3bd62a8b),
	.w5(32'h3c265020),
	.w6(32'hbb5aa86d),
	.w7(32'h3bd4b670),
	.w8(32'hbb914cea),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b4eaa),
	.w1(32'hbac3c13d),
	.w2(32'h3c0973eb),
	.w3(32'h3a5a24e6),
	.w4(32'hbbe3574d),
	.w5(32'h3ba06634),
	.w6(32'hbc26fd8c),
	.w7(32'h3c70fa67),
	.w8(32'hbb173ec1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1203f),
	.w1(32'h39807678),
	.w2(32'h3b3cbefd),
	.w3(32'hbc27dd80),
	.w4(32'hbbbfc62c),
	.w5(32'hbb53fc1f),
	.w6(32'hbc0307e4),
	.w7(32'h3b2955ba),
	.w8(32'hbb047679),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc05b66),
	.w1(32'hba04a557),
	.w2(32'h3b2e4563),
	.w3(32'hbb7cac26),
	.w4(32'h3b83436d),
	.w5(32'h3bf2f3e3),
	.w6(32'h3c8b45fc),
	.w7(32'hbb37cd89),
	.w8(32'h3c42d3f4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7db02d),
	.w1(32'hbac42aff),
	.w2(32'hbbc7ddb0),
	.w3(32'hbba689c7),
	.w4(32'hb99841da),
	.w5(32'hbc2d23fe),
	.w6(32'hbc932d20),
	.w7(32'hbaa16ede),
	.w8(32'hbbeee484),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a025b59),
	.w1(32'hbb0dcf09),
	.w2(32'h3cc8c6ae),
	.w3(32'hbb9c8216),
	.w4(32'h3b697670),
	.w5(32'hbb6c28bc),
	.w6(32'h3bd4f4c7),
	.w7(32'h3a2ccf94),
	.w8(32'hb8ed2662),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba5b5e),
	.w1(32'h3a4a7f33),
	.w2(32'h3ba8ce5b),
	.w3(32'h3c18c114),
	.w4(32'hbab834a3),
	.w5(32'h3a8faaf9),
	.w6(32'hba35a486),
	.w7(32'h3bd8f2d4),
	.w8(32'h3b367d86),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e5065),
	.w1(32'h3b70c7da),
	.w2(32'h3bda717c),
	.w3(32'h3ca5f74c),
	.w4(32'h3b825586),
	.w5(32'hbc3c9192),
	.w6(32'hbd3118aa),
	.w7(32'h3a3c22ef),
	.w8(32'h39d119f4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba47ac),
	.w1(32'h3b1fd83c),
	.w2(32'h3bda8e98),
	.w3(32'hbbdbad5e),
	.w4(32'h3c201497),
	.w5(32'h3b275643),
	.w6(32'h391ca016),
	.w7(32'hbb4b902c),
	.w8(32'h39169ebd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e1301),
	.w1(32'hbbbf2a73),
	.w2(32'h3aa227c5),
	.w3(32'h3a07bc57),
	.w4(32'hbc7abafb),
	.w5(32'hbc877281),
	.w6(32'hbc4d9ad4),
	.w7(32'hbbc9382e),
	.w8(32'h3bb13dce),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f0fa4),
	.w1(32'hbc411370),
	.w2(32'hbb32ba3a),
	.w3(32'hbbbb2b4e),
	.w4(32'hbc4aba91),
	.w5(32'hbb9293ed),
	.w6(32'hbb951df7),
	.w7(32'hbc0de65d),
	.w8(32'h3b18fff3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa36c0),
	.w1(32'hbb2f3477),
	.w2(32'h3bcf6bbb),
	.w3(32'h3bc0d01c),
	.w4(32'hba935dfc),
	.w5(32'hbac9e749),
	.w6(32'hbbb92320),
	.w7(32'hbba46871),
	.w8(32'hba509d61),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93a276),
	.w1(32'hba4df5dc),
	.w2(32'h3ac46ff5),
	.w3(32'hbbc285e8),
	.w4(32'h3c1f9880),
	.w5(32'hbc1d22dc),
	.w6(32'hbce0b6aa),
	.w7(32'h3b11cfb1),
	.w8(32'hbab49f82),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91421f),
	.w1(32'h3b005994),
	.w2(32'hbb6c13e1),
	.w3(32'h3bacdcca),
	.w4(32'hbc111930),
	.w5(32'hbc003574),
	.w6(32'hbb8b32e7),
	.w7(32'hbc262b08),
	.w8(32'h3c03ba26),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60a1f2),
	.w1(32'hba326876),
	.w2(32'hbc11b3f5),
	.w3(32'h3ba6df84),
	.w4(32'hb936305a),
	.w5(32'h3c166556),
	.w6(32'h3ba3faa1),
	.w7(32'hbc765193),
	.w8(32'h3973e634),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73ff6e),
	.w1(32'h3b468407),
	.w2(32'h3b20bee4),
	.w3(32'hbb8a6a02),
	.w4(32'h3b61c189),
	.w5(32'h3c128631),
	.w6(32'h3b0c33a5),
	.w7(32'h3ad5efbb),
	.w8(32'hbbd8a846),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ef34b),
	.w1(32'hbc153c2b),
	.w2(32'h3d1e21fd),
	.w3(32'h3aba7b11),
	.w4(32'hbbd0c8d7),
	.w5(32'h3bf2c4fc),
	.w6(32'hbb7e3c4c),
	.w7(32'hbbe89415),
	.w8(32'h3affb32d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29368a),
	.w1(32'hbb94cc04),
	.w2(32'h3b6e7cbc),
	.w3(32'hbbcd44c9),
	.w4(32'h3b1ff3c5),
	.w5(32'h3b5e0f84),
	.w6(32'h39075559),
	.w7(32'hbc3ad828),
	.w8(32'hbbd890ce),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58b141),
	.w1(32'h3ced06c3),
	.w2(32'h3ad1bb95),
	.w3(32'hbcd2beeb),
	.w4(32'h3bb2c253),
	.w5(32'h3b15503d),
	.w6(32'h3c915573),
	.w7(32'hbb8d603c),
	.w8(32'hbb9ef47e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f9f5e),
	.w1(32'hbbe68e82),
	.w2(32'hbab85d25),
	.w3(32'h39cc5ecc),
	.w4(32'hbb87a361),
	.w5(32'hbbc90e73),
	.w6(32'hbc4ce3db),
	.w7(32'h3b9b8c4d),
	.w8(32'hbad786c6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b195ce9),
	.w1(32'hbbf0a843),
	.w2(32'h3b434ca2),
	.w3(32'h3b8e788c),
	.w4(32'hbc42ab29),
	.w5(32'hbba8dad2),
	.w6(32'hbc8c9ab3),
	.w7(32'hbba81aae),
	.w8(32'hbae9a76a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c042274),
	.w1(32'h3b3c89d5),
	.w2(32'h392f45c7),
	.w3(32'hbbd55fe5),
	.w4(32'hbcb5fab3),
	.w5(32'hbc24f437),
	.w6(32'h3b197a5b),
	.w7(32'hbbeea6bc),
	.w8(32'hbbb2d122),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05423b),
	.w1(32'h3b2a0977),
	.w2(32'h3b9db78f),
	.w3(32'hbb03d742),
	.w4(32'hba1d7fd3),
	.w5(32'h3b864c3c),
	.w6(32'hba469bac),
	.w7(32'h3b050c95),
	.w8(32'hbb350d2a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b32cc4),
	.w1(32'hbbb022df),
	.w2(32'h3bb71296),
	.w3(32'hb92ff756),
	.w4(32'h3d52d8bf),
	.w5(32'hbb797823),
	.w6(32'h3b5d6b70),
	.w7(32'h3a61f829),
	.w8(32'h3bc248e2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb979043),
	.w1(32'hbc3918dc),
	.w2(32'h39d79c9a),
	.w3(32'hbbdd1720),
	.w4(32'hbc986aa5),
	.w5(32'hbb1d8c64),
	.w6(32'hbc5a073d),
	.w7(32'hbb7cf537),
	.w8(32'h3b91a816),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b103da5),
	.w1(32'h3bad93be),
	.w2(32'h3b2f1f60),
	.w3(32'h3bc5944d),
	.w4(32'h3b35ed59),
	.w5(32'h3abb60c3),
	.w6(32'h3be20844),
	.w7(32'h3a7cc29a),
	.w8(32'hbb2131ed),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44f37e),
	.w1(32'h3a93033e),
	.w2(32'hbba092de),
	.w3(32'hbc4a05f0),
	.w4(32'h3c3767bc),
	.w5(32'hbc4e34b0),
	.w6(32'hbc3afb22),
	.w7(32'hbb81765a),
	.w8(32'h3b8a3971),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba990b5),
	.w1(32'h3bc76c48),
	.w2(32'hb9d7895e),
	.w3(32'h3b42cd72),
	.w4(32'hbb8e23b5),
	.w5(32'hba9a0b29),
	.w6(32'h3b5ed23d),
	.w7(32'hbb6f79d9),
	.w8(32'hba6d48ce),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7414),
	.w1(32'h3cb0b54b),
	.w2(32'h3b46c1ce),
	.w3(32'hbc623041),
	.w4(32'hbd42559d),
	.w5(32'h3b9045b4),
	.w6(32'h3ae17122),
	.w7(32'hbd91152d),
	.w8(32'h3b6bdbb4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc212d06),
	.w1(32'hbbb832bc),
	.w2(32'hbb4fdb96),
	.w3(32'hbb415364),
	.w4(32'h3c0c203f),
	.w5(32'h3bd6868c),
	.w6(32'hbc570620),
	.w7(32'hba3fdcd9),
	.w8(32'h3b534bf6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba790b28),
	.w1(32'hbb8c49ea),
	.w2(32'hbb4c3166),
	.w3(32'hbc14e4c6),
	.w4(32'hbbedd12b),
	.w5(32'h3beffce0),
	.w6(32'hbcc7a95f),
	.w7(32'hbb0499c5),
	.w8(32'h3b97ca1f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c046792),
	.w1(32'h3b4ff0a4),
	.w2(32'h3c6b7f2c),
	.w3(32'hbb34c264),
	.w4(32'h3bc8d8da),
	.w5(32'hb98cec02),
	.w6(32'hbad68cb9),
	.w7(32'hbb4956de),
	.w8(32'h3b44956e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e7a0b),
	.w1(32'h3c45db30),
	.w2(32'hbc832f84),
	.w3(32'h3ad71ea2),
	.w4(32'hbbd17e07),
	.w5(32'h3beb8509),
	.w6(32'h38875367),
	.w7(32'h3d088af5),
	.w8(32'h3c0067b8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9af1e2),
	.w1(32'hbc22e038),
	.w2(32'h3a630063),
	.w3(32'h3b013018),
	.w4(32'hba6b7c45),
	.w5(32'hbc461250),
	.w6(32'h3c307578),
	.w7(32'hbc40c220),
	.w8(32'h3b42a524),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb119356),
	.w1(32'hbb572640),
	.w2(32'h3bc0c47b),
	.w3(32'hbd5c3fd3),
	.w4(32'h3ce8fcbb),
	.w5(32'h3b8e73fc),
	.w6(32'h3b8e1b5e),
	.w7(32'hbcdabd14),
	.w8(32'hb9a56a5b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b978c),
	.w1(32'hbc072a1f),
	.w2(32'h3d489afe),
	.w3(32'hbc775641),
	.w4(32'hbb609f7d),
	.w5(32'h3c14b97b),
	.w6(32'h3bea69a0),
	.w7(32'hbad18d30),
	.w8(32'hbc164ead),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd66528),
	.w1(32'hbbd1cb69),
	.w2(32'h3bf3f917),
	.w3(32'hbc17540a),
	.w4(32'h3b3418b1),
	.w5(32'hbc57ed35),
	.w6(32'h3c320348),
	.w7(32'h3b993136),
	.w8(32'h3c4fe3c8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82657a),
	.w1(32'h3bddcc22),
	.w2(32'h3c0b1ed7),
	.w3(32'hbbd0b2d6),
	.w4(32'hbbb9d1ac),
	.w5(32'hbba9a198),
	.w6(32'hbce049d1),
	.w7(32'h3b46eece),
	.w8(32'hbd4ac152),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc91597),
	.w1(32'hbc3715b6),
	.w2(32'h3a34af2b),
	.w3(32'hbb48a01c),
	.w4(32'h3bb2075a),
	.w5(32'hbc144741),
	.w6(32'hbca08913),
	.w7(32'h3bda01f1),
	.w8(32'hbb156cb3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb75466),
	.w1(32'h3c316712),
	.w2(32'hbc37aab7),
	.w3(32'h3b421ed4),
	.w4(32'h3b2f5b0a),
	.w5(32'h3ad9300b),
	.w6(32'hbc66f839),
	.w7(32'hbbc38af8),
	.w8(32'hbb4ea476),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdfb7d),
	.w1(32'hbc10e83d),
	.w2(32'h3b8b03fe),
	.w3(32'hbbae5a4d),
	.w4(32'h39a27a02),
	.w5(32'hb90aea90),
	.w6(32'h3b89527e),
	.w7(32'hbad4d0c0),
	.w8(32'hbbe5c4af),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a33b9f),
	.w1(32'hbc33c8ab),
	.w2(32'h35b3019a),
	.w3(32'h3b4c21a5),
	.w4(32'h3c0e3ab8),
	.w5(32'h3bacf120),
	.w6(32'h3b8b9f5f),
	.w7(32'hbb07edbd),
	.w8(32'h3c161b37),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2498de),
	.w1(32'h3c1ade91),
	.w2(32'h3c6812f2),
	.w3(32'h3b897b17),
	.w4(32'hbca3ae89),
	.w5(32'hbbf798a9),
	.w6(32'h3cad34d0),
	.w7(32'hbbf04ece),
	.w8(32'h3c1d7d34),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97aab8c),
	.w1(32'h3b1f1095),
	.w2(32'hba34f5d1),
	.w3(32'hbb1b1192),
	.w4(32'hbc85d337),
	.w5(32'hbac47298),
	.w6(32'hbb4159d1),
	.w7(32'hbc0a946c),
	.w8(32'h3baba249),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74ead7),
	.w1(32'h3ca6ec38),
	.w2(32'hbbd0d26c),
	.w3(32'h3bb24f1c),
	.w4(32'h3be4593b),
	.w5(32'h3a15d2a8),
	.w6(32'h3af16964),
	.w7(32'h3b94ec14),
	.w8(32'hbad5d1bc),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd35dd5),
	.w1(32'hbc5166cd),
	.w2(32'h39f1a550),
	.w3(32'h3ce1d83f),
	.w4(32'hbbf693ad),
	.w5(32'hb990ba02),
	.w6(32'h38a9d54b),
	.w7(32'hbc84e8c0),
	.w8(32'h3b97d555),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c351025),
	.w1(32'hbc1b2eae),
	.w2(32'h3c69858c),
	.w3(32'h3a267b1f),
	.w4(32'h3c317253),
	.w5(32'hbd561fa1),
	.w6(32'hbbb82332),
	.w7(32'hbc29f153),
	.w8(32'h3ac35a8b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6203f3),
	.w1(32'hbb2c368c),
	.w2(32'h3950fe4f),
	.w3(32'h3b66cfbf),
	.w4(32'hbc64491f),
	.w5(32'h3be4e7dc),
	.w6(32'h3c31502e),
	.w7(32'h3bb55dda),
	.w8(32'h39d87e26),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb0eef),
	.w1(32'hbc2f39bb),
	.w2(32'h3cd0d58f),
	.w3(32'h3aeccf38),
	.w4(32'h3b199d0e),
	.w5(32'hbb6edf26),
	.w6(32'hbc096ae2),
	.w7(32'h3b67e6da),
	.w8(32'h3bab20e0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd20338),
	.w1(32'h3c2f9751),
	.w2(32'h3bbc48a4),
	.w3(32'hbb495e51),
	.w4(32'h3bd16446),
	.w5(32'h3c0c4801),
	.w6(32'hba968074),
	.w7(32'hbc3224f8),
	.w8(32'h3c5184ca),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810c2f),
	.w1(32'hbbed9196),
	.w2(32'hbb8c16fb),
	.w3(32'hbc287bc5),
	.w4(32'h3c11acd3),
	.w5(32'h3a28faad),
	.w6(32'hbceb0b96),
	.w7(32'h3a25d9ff),
	.w8(32'h3b9b351c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5f4d3),
	.w1(32'hbc4fa729),
	.w2(32'hbaf98516),
	.w3(32'h3933c983),
	.w4(32'hbb5263eb),
	.w5(32'hbc201449),
	.w6(32'h3bb48bb6),
	.w7(32'hb896d874),
	.w8(32'hbc9424f2),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc683f5),
	.w1(32'h3b93c191),
	.w2(32'h3c47b5c0),
	.w3(32'hbb79f972),
	.w4(32'h3bfac453),
	.w5(32'hba2786f9),
	.w6(32'hbc90faca),
	.w7(32'h3ba9be24),
	.w8(32'h3a18b16c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcc2bd),
	.w1(32'h3b29e57b),
	.w2(32'hbc83c318),
	.w3(32'hbba57efb),
	.w4(32'h3c1dd488),
	.w5(32'hbbaefafa),
	.w6(32'h3c28ce31),
	.w7(32'h3c6ba275),
	.w8(32'hbc0a22e8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb348b61),
	.w1(32'h3b0eff87),
	.w2(32'h3c851ade),
	.w3(32'hbbfd005d),
	.w4(32'hbc77fbd4),
	.w5(32'hbc2e44fd),
	.w6(32'h3c2078bc),
	.w7(32'h3be669a4),
	.w8(32'hbb937586),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb157993),
	.w1(32'hbbac4064),
	.w2(32'h3b65287a),
	.w3(32'h3b05ef89),
	.w4(32'h3c4bd4a6),
	.w5(32'hbbd29577),
	.w6(32'h3c99f6e6),
	.w7(32'hbbed0c49),
	.w8(32'h3bf68304),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c63ec1),
	.w1(32'hbbe44a61),
	.w2(32'h3b98a0d9),
	.w3(32'hbbd30f3d),
	.w4(32'h3b9d9c98),
	.w5(32'h3b7b0a54),
	.w6(32'hbaaf15f4),
	.w7(32'hbc5473e7),
	.w8(32'h3cb7f884),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51ae29),
	.w1(32'h3b7b084c),
	.w2(32'hb9ea073d),
	.w3(32'hbad559cc),
	.w4(32'h3aee8d93),
	.w5(32'hbc25befb),
	.w6(32'h3b01d5eb),
	.w7(32'hbba54376),
	.w8(32'hbc51205d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd3d71),
	.w1(32'hbc2d2b51),
	.w2(32'hbb3eae6a),
	.w3(32'h3b5c1da9),
	.w4(32'h3cd92951),
	.w5(32'hbbe750bb),
	.w6(32'h3bef4f9a),
	.w7(32'hba8c573b),
	.w8(32'h3bb8a523),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc822762),
	.w1(32'hba78eba4),
	.w2(32'h3b1d0133),
	.w3(32'hbc0073c9),
	.w4(32'hbab87662),
	.w5(32'h3c9a0976),
	.w6(32'hbb906ed5),
	.w7(32'hbbe7b8c4),
	.w8(32'hbb77d56a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6379b9),
	.w1(32'hbc8a2796),
	.w2(32'hbc21a70a),
	.w3(32'hba43a522),
	.w4(32'h3a690a47),
	.w5(32'hbba35e09),
	.w6(32'h3b765a4d),
	.w7(32'hba9249cb),
	.w8(32'h3b87cab3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8abec4),
	.w1(32'hbbf9f09f),
	.w2(32'hbae0c07f),
	.w3(32'h399629a1),
	.w4(32'hbbc0ac7e),
	.w5(32'hbbe06418),
	.w6(32'h3bb9e477),
	.w7(32'hbb34c4de),
	.w8(32'hbc79e20b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcda5e6),
	.w1(32'hb9c0692e),
	.w2(32'h3b893ab1),
	.w3(32'h3bcf0f49),
	.w4(32'h3af17527),
	.w5(32'h3b11413c),
	.w6(32'h3bd7d881),
	.w7(32'h3c60e0ef),
	.w8(32'hbad4de36),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18508d),
	.w1(32'h3badf636),
	.w2(32'h3bae214b),
	.w3(32'hbb39a2ff),
	.w4(32'h3c3c2bcb),
	.w5(32'hbcd5eeb0),
	.w6(32'hbac5fd1a),
	.w7(32'hbac25474),
	.w8(32'hbb61e2ba),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfff40e),
	.w1(32'h3b31de22),
	.w2(32'hba32edbc),
	.w3(32'h3a592a6a),
	.w4(32'hbc4dec7a),
	.w5(32'h3ad20b0f),
	.w6(32'h3b9f177b),
	.w7(32'h3c0bbcc4),
	.w8(32'hbc9b154c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6b0db),
	.w1(32'hbbcea903),
	.w2(32'h3bd49bd0),
	.w3(32'h3c9755f9),
	.w4(32'hba58d2c7),
	.w5(32'h3c2153ab),
	.w6(32'hbc6e0b73),
	.w7(32'h3c52bf96),
	.w8(32'hbc0486b5),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd64fd),
	.w1(32'h3c3210d8),
	.w2(32'hbb58c535),
	.w3(32'h3c1eaa2e),
	.w4(32'h3c0823da),
	.w5(32'h3ba30e5e),
	.w6(32'hbbf65005),
	.w7(32'h3a08c428),
	.w8(32'hbadded58),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33ec83),
	.w1(32'hbbdf9a18),
	.w2(32'hbbac886d),
	.w3(32'hbb73eff3),
	.w4(32'hbb980abb),
	.w5(32'h3c824e34),
	.w6(32'h3bd6ffc0),
	.w7(32'hbabd501b),
	.w8(32'hbc484c00),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b4525),
	.w1(32'h3b9b3b26),
	.w2(32'hbb8dbc83),
	.w3(32'h3c178cbb),
	.w4(32'hbc04b839),
	.w5(32'h3ba95fce),
	.w6(32'hbc0b2992),
	.w7(32'h3c01578d),
	.w8(32'h3b80c0c0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b7761),
	.w1(32'hbc337c08),
	.w2(32'hbbbb27e4),
	.w3(32'h3b6eb21a),
	.w4(32'h39ae5063),
	.w5(32'h3b0b6e2d),
	.w6(32'h3851f46b),
	.w7(32'hbb68accf),
	.w8(32'h3c878696),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301e97),
	.w1(32'hbbacc174),
	.w2(32'h3b974e78),
	.w3(32'h3bc2ae86),
	.w4(32'hbd0b6b7d),
	.w5(32'hbc21fc46),
	.w6(32'hbbfd7987),
	.w7(32'hba0579d3),
	.w8(32'hbc9288a4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51fde8),
	.w1(32'h3cb18891),
	.w2(32'hb985153a),
	.w3(32'h3ac656cb),
	.w4(32'hb89c5cf4),
	.w5(32'hbc80706f),
	.w6(32'hbacaa43a),
	.w7(32'h3a0d4c6a),
	.w8(32'hbce3f35c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b193b0c),
	.w1(32'h3b83f0c3),
	.w2(32'hba26d19c),
	.w3(32'hbb4ecefa),
	.w4(32'h3c4e88b0),
	.w5(32'h3bb22c7e),
	.w6(32'h3c268dcc),
	.w7(32'h3aad93d0),
	.w8(32'hbc1210ef),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0214b),
	.w1(32'hbbf1c282),
	.w2(32'hbba97c67),
	.w3(32'hbba438ec),
	.w4(32'hbc3a0f4c),
	.w5(32'h3bab6a38),
	.w6(32'hb9a7684d),
	.w7(32'h3bab2fe1),
	.w8(32'hb93e2f1e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ad9c1),
	.w1(32'h3bfce070),
	.w2(32'hbba460f4),
	.w3(32'h39c63d2b),
	.w4(32'hbb54a5cb),
	.w5(32'h3c340f5f),
	.w6(32'h3b373270),
	.w7(32'h3b948c21),
	.w8(32'hba10f9df),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba02809),
	.w1(32'hbb3c9993),
	.w2(32'h3bfa5373),
	.w3(32'h3afde1b0),
	.w4(32'h3b980440),
	.w5(32'h3c27dd99),
	.w6(32'h3bd318ba),
	.w7(32'hbb123463),
	.w8(32'hba9b0c3f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ea806),
	.w1(32'hbc4578ae),
	.w2(32'hbb9314c9),
	.w3(32'hbc51a8c2),
	.w4(32'hbbb6ebed),
	.w5(32'h3bf98baa),
	.w6(32'hbc27f4bf),
	.w7(32'hbb5cff1b),
	.w8(32'hbbe32547),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f50f5),
	.w1(32'h3b95f7fd),
	.w2(32'hba911308),
	.w3(32'hbab34f9d),
	.w4(32'hbbaece07),
	.w5(32'hbc4b1c62),
	.w6(32'hbc05f757),
	.w7(32'hbc094398),
	.w8(32'hba79c3fc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3192cc),
	.w1(32'hbc4c6227),
	.w2(32'h3be246f6),
	.w3(32'hbc1bf0c7),
	.w4(32'hbb6b09b8),
	.w5(32'h3bb8e3c8),
	.w6(32'h3bb51f47),
	.w7(32'hbc049251),
	.w8(32'h3a612f4e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc222254),
	.w1(32'h3af09f12),
	.w2(32'h3aef4900),
	.w3(32'h3b8931d5),
	.w4(32'hbb427205),
	.w5(32'h3b4c791a),
	.w6(32'h3b66edbe),
	.w7(32'hbbbefe27),
	.w8(32'h3b22e592),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9596a85),
	.w1(32'hbc2a41dc),
	.w2(32'hb9a11fa2),
	.w3(32'hbaea4550),
	.w4(32'h3bdede8c),
	.w5(32'hbb89e074),
	.w6(32'hbb4da783),
	.w7(32'hbbc8f877),
	.w8(32'hbb002b15),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ce51),
	.w1(32'h3c206c60),
	.w2(32'hbc1de27a),
	.w3(32'hbba7ede5),
	.w4(32'hbb9850bc),
	.w5(32'hbb6374db),
	.w6(32'hbc1519c0),
	.w7(32'h3b18592c),
	.w8(32'h3c35238d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8b1b3),
	.w1(32'h3b7bfa88),
	.w2(32'hbc04e5d7),
	.w3(32'h3cc7acef),
	.w4(32'hbbb1f0de),
	.w5(32'h3b1ffbe4),
	.w6(32'h3bc1e3fa),
	.w7(32'h3b423abe),
	.w8(32'h3acfd289),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967312),
	.w1(32'h3bc5f647),
	.w2(32'hbc02ab71),
	.w3(32'h3c1097ed),
	.w4(32'h3b70a1b8),
	.w5(32'h3bf6c471),
	.w6(32'hbb8326fb),
	.w7(32'h3c110fa7),
	.w8(32'h3c03edef),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13f23a),
	.w1(32'hbc3c6a07),
	.w2(32'hbbf3d431),
	.w3(32'h3aa8eb54),
	.w4(32'hbbb31422),
	.w5(32'hbc2820eb),
	.w6(32'hba47326f),
	.w7(32'h3b0aef69),
	.w8(32'hbb607c3a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc146492),
	.w1(32'hbc0f3b33),
	.w2(32'hbbda68c7),
	.w3(32'h3be445c9),
	.w4(32'h3c118d6c),
	.w5(32'hba1d71a6),
	.w6(32'hbc960dc1),
	.w7(32'h3b660517),
	.w8(32'hbaf46025),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a5417),
	.w1(32'h3a5549e6),
	.w2(32'h3be27e6a),
	.w3(32'h3b21e627),
	.w4(32'hbb04b39f),
	.w5(32'hbb065ba9),
	.w6(32'hbbd3047d),
	.w7(32'hbc57f625),
	.w8(32'h3cf9ce1b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beabfb9),
	.w1(32'hbb0037a2),
	.w2(32'hbbe53383),
	.w3(32'hbc82aecd),
	.w4(32'hba4b9327),
	.w5(32'hbc83b952),
	.w6(32'hbbc5ec8d),
	.w7(32'hbb2c90cb),
	.w8(32'h3ba202f7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becf823),
	.w1(32'hbb5555a8),
	.w2(32'hbc39f46c),
	.w3(32'h3ad15387),
	.w4(32'hbb730b23),
	.w5(32'hba7c954e),
	.w6(32'h3c186652),
	.w7(32'hbc2c5859),
	.w8(32'h3b9de1c8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2764),
	.w1(32'hbc00ae1f),
	.w2(32'h3a9d3675),
	.w3(32'hbc0a6162),
	.w4(32'hbb8ff930),
	.w5(32'hbb8859fc),
	.w6(32'hbb861af3),
	.w7(32'hbb93759c),
	.w8(32'h3a3498a5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e71f2),
	.w1(32'h3af2ccef),
	.w2(32'hbc56e685),
	.w3(32'hbb36d0dc),
	.w4(32'hbc081da9),
	.w5(32'h36f0641b),
	.w6(32'hbce9f229),
	.w7(32'h3c47435f),
	.w8(32'h3b210343),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd093d6a),
	.w1(32'h3c82dd84),
	.w2(32'hbc1d38c5),
	.w3(32'h39b1ed3d),
	.w4(32'hbb29e0a7),
	.w5(32'h3b4c450e),
	.w6(32'h3b7a80da),
	.w7(32'hbbc9dd81),
	.w8(32'h3c058f0c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe4d77),
	.w1(32'hbc282935),
	.w2(32'h3b8671fd),
	.w3(32'hbc7b7096),
	.w4(32'hb99b1d7c),
	.w5(32'hbad25722),
	.w6(32'h3c1dd5f7),
	.w7(32'h3c8c246d),
	.w8(32'h3bb4aa2b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea5dfe),
	.w1(32'hbcea10d2),
	.w2(32'h3c22fd85),
	.w3(32'hbbadf920),
	.w4(32'h3b97c9eb),
	.w5(32'hba1ae9fc),
	.w6(32'hbadef259),
	.w7(32'hbc110e35),
	.w8(32'hba3ccca0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d9760),
	.w1(32'hbbecde68),
	.w2(32'h3b7899b7),
	.w3(32'hbbd857bb),
	.w4(32'hbc793593),
	.w5(32'hbc19f1de),
	.w6(32'h3c1ad158),
	.w7(32'hbc87be00),
	.w8(32'hbc4c2a55),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96fb0c),
	.w1(32'h3aff8a61),
	.w2(32'hbc187a55),
	.w3(32'hbbde7840),
	.w4(32'hbbbf72af),
	.w5(32'hbc1d4e75),
	.w6(32'h3bceb6e1),
	.w7(32'h3b94f161),
	.w8(32'h3b72304f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11cb3c),
	.w1(32'hba8b6374),
	.w2(32'hbc10619d),
	.w3(32'hbc4dae11),
	.w4(32'hbb97fed2),
	.w5(32'hbbb93376),
	.w6(32'h3ba0de43),
	.w7(32'hbb9dcf97),
	.w8(32'hbb8d2eda),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa00d96),
	.w1(32'h3a40ea33),
	.w2(32'hb9bbe29b),
	.w3(32'hbc1e6f2a),
	.w4(32'hbc0c2e13),
	.w5(32'hbc35d9d8),
	.w6(32'h3af4e396),
	.w7(32'h3c414baf),
	.w8(32'h3b0145fa),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2188cf),
	.w1(32'h3c712368),
	.w2(32'hbc3337db),
	.w3(32'h3b3fdc87),
	.w4(32'h3bcc2722),
	.w5(32'hbc09cff6),
	.w6(32'h3c8eebcb),
	.w7(32'hbbf1c9b7),
	.w8(32'h3b4b4328),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc819735),
	.w1(32'hbc52b62e),
	.w2(32'h3aee742e),
	.w3(32'hbc1ac374),
	.w4(32'h3c326184),
	.w5(32'hbaf89dbe),
	.w6(32'h3ac17054),
	.w7(32'h3c7c57d5),
	.w8(32'hbc555924),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cbd1b),
	.w1(32'hbcd13b34),
	.w2(32'h3b7d5d89),
	.w3(32'h3c902072),
	.w4(32'hbae2e4f4),
	.w5(32'h3be527aa),
	.w6(32'hbc463625),
	.w7(32'h3c4110af),
	.w8(32'hbc3c3fb4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f3221),
	.w1(32'hbb800986),
	.w2(32'h3a3a095f),
	.w3(32'h3bc0ff1b),
	.w4(32'hbb80d544),
	.w5(32'hbc79c4f4),
	.w6(32'h3c275f0a),
	.w7(32'h3b245eb4),
	.w8(32'hbbec0f8a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7b7c7),
	.w1(32'hbb05b12b),
	.w2(32'hbbc23384),
	.w3(32'hbc180dca),
	.w4(32'hbb2b931e),
	.w5(32'hbb5e11b3),
	.w6(32'h3b04691e),
	.w7(32'h3a345d4a),
	.w8(32'hbb7357d0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf5608),
	.w1(32'hba9fe20e),
	.w2(32'hbc7f40f6),
	.w3(32'h3bc58d1c),
	.w4(32'hbb9b484c),
	.w5(32'hbcb6fa35),
	.w6(32'hbb59842f),
	.w7(32'hbd07bb23),
	.w8(32'h389cc581),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab62589),
	.w1(32'hbac00cd9),
	.w2(32'h3be9712e),
	.w3(32'h3b790d0f),
	.w4(32'hbc7f069b),
	.w5(32'h3b0747e0),
	.w6(32'hbbd2f9cc),
	.w7(32'hbc7e3c68),
	.w8(32'h3c116eae),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920342),
	.w1(32'hbb1a0037),
	.w2(32'hbc01ac47),
	.w3(32'hbaf053c6),
	.w4(32'hbba9f062),
	.w5(32'h3b9f144b),
	.w6(32'h3aba78f0),
	.w7(32'hbae8e677),
	.w8(32'h3b98d4b9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e14ea9),
	.w1(32'hbc622419),
	.w2(32'h3b6ae40a),
	.w3(32'h3c20c5a9),
	.w4(32'h392745b7),
	.w5(32'hbbbdf503),
	.w6(32'hbc11c13b),
	.w7(32'hbb4c70fd),
	.w8(32'h3b810447),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add288a),
	.w1(32'hbce0d495),
	.w2(32'h3ac115bb),
	.w3(32'hbc93bdb9),
	.w4(32'h3bff8f19),
	.w5(32'hbb5f3508),
	.w6(32'h3ad37bc4),
	.w7(32'h3baa4113),
	.w8(32'hbbcef458),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f7ed1),
	.w1(32'h3bf11f34),
	.w2(32'hbc13368b),
	.w3(32'hbc348c56),
	.w4(32'hb9a3dab0),
	.w5(32'hbc952991),
	.w6(32'hbb7236c5),
	.w7(32'hbb0f2979),
	.w8(32'h3cc1714a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c166788),
	.w1(32'hbaacbbb5),
	.w2(32'h3bbc2cd4),
	.w3(32'hbba531cf),
	.w4(32'h3b64b666),
	.w5(32'hba7d9ece),
	.w6(32'hbc04ce33),
	.w7(32'hbc4cea97),
	.w8(32'hbc5ae7c3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63750b),
	.w1(32'hbb6b30cb),
	.w2(32'h3a8a8281),
	.w3(32'hbc857e7c),
	.w4(32'h3ad863f1),
	.w5(32'h3b6ef885),
	.w6(32'hbb87f2b2),
	.w7(32'h3c832aff),
	.w8(32'hbb848d53),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeed356),
	.w1(32'h3a6d3844),
	.w2(32'h3bbefa4e),
	.w3(32'h3c7bae8a),
	.w4(32'hbc9ceec8),
	.w5(32'h36bd148d),
	.w6(32'h3b45faea),
	.w7(32'hbccf94c1),
	.w8(32'hbba3ba51),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1854aa),
	.w1(32'h3bb91489),
	.w2(32'hbbc33c8e),
	.w3(32'hbcac2eb7),
	.w4(32'hbb468e34),
	.w5(32'hbb747bc8),
	.w6(32'h3b17aae2),
	.w7(32'hbbdc25dc),
	.w8(32'h3b1584b3),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06aa4b),
	.w1(32'hbb176e3f),
	.w2(32'h3bc7a358),
	.w3(32'hbc092e5b),
	.w4(32'hbc9f00e5),
	.w5(32'hbcdf8adb),
	.w6(32'hbbc4d4c4),
	.w7(32'h3b7d04ef),
	.w8(32'h3c18d706),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b733961),
	.w1(32'hbaf50d43),
	.w2(32'hbb154eeb),
	.w3(32'h3bc98816),
	.w4(32'hbb0672d4),
	.w5(32'hbc2e5882),
	.w6(32'hbc582589),
	.w7(32'hbad0adda),
	.w8(32'hb6a31e6d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52f8bc),
	.w1(32'h3c2b9b2f),
	.w2(32'hba8db5c2),
	.w3(32'hbbfb41c2),
	.w4(32'h3bb0ec9f),
	.w5(32'hbc00c747),
	.w6(32'h3989b80a),
	.w7(32'h3c01164f),
	.w8(32'hbc00c27c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e44d7),
	.w1(32'h3bd0962a),
	.w2(32'hbbf61003),
	.w3(32'hbc20da67),
	.w4(32'hb9fabd0a),
	.w5(32'hbc1a30e5),
	.w6(32'h3b231893),
	.w7(32'hbbaf3f2a),
	.w8(32'hb9d7068e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aebf7),
	.w1(32'h3bdef8b2),
	.w2(32'hbb72ba7a),
	.w3(32'hbb4ac2df),
	.w4(32'h3ba9f116),
	.w5(32'hbc078859),
	.w6(32'hbbec5537),
	.w7(32'hbc7e17e2),
	.w8(32'hbb32e261),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc963ed1),
	.w1(32'h3c2c812e),
	.w2(32'hbc0f7727),
	.w3(32'h3b17b1e2),
	.w4(32'hbadc74cf),
	.w5(32'hba7b2825),
	.w6(32'h3ae38e34),
	.w7(32'hba531862),
	.w8(32'hbca18d32),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab515d3),
	.w1(32'h39f241b5),
	.w2(32'h3bf9c805),
	.w3(32'hb9caf55c),
	.w4(32'h3d1e2d87),
	.w5(32'hbb29e5fa),
	.w6(32'h3bd5296f),
	.w7(32'h3bd5539a),
	.w8(32'hbc81a21d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47aea),
	.w1(32'h3c3cd242),
	.w2(32'hbab37b12),
	.w3(32'hba859059),
	.w4(32'h3c5f5462),
	.w5(32'h3bf3272d),
	.w6(32'hbb18a1a6),
	.w7(32'hbc47041b),
	.w8(32'hbaefa774),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee86c5),
	.w1(32'h3b9b82f9),
	.w2(32'hbbe1af06),
	.w3(32'h3aeb56c5),
	.w4(32'hba4279ad),
	.w5(32'h3bcdf5fd),
	.w6(32'h3bf64667),
	.w7(32'h3c622325),
	.w8(32'h3b38a655),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3effb8),
	.w1(32'h3b80c353),
	.w2(32'h3c10f5ec),
	.w3(32'h3c2a764c),
	.w4(32'hbbf21c5b),
	.w5(32'hbc1ecebb),
	.w6(32'hbb14b9c0),
	.w7(32'h3c59e27a),
	.w8(32'h3c53968a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000b6c),
	.w1(32'h3ba6e6fe),
	.w2(32'h3c261645),
	.w3(32'hb9b74b1f),
	.w4(32'h3b8acdd6),
	.w5(32'hbcaa1026),
	.w6(32'h3b18d637),
	.w7(32'h3a21724f),
	.w8(32'h398b622c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fb59e),
	.w1(32'h3b9171d5),
	.w2(32'h3b3c5350),
	.w3(32'hbb97cc32),
	.w4(32'hbca97c5b),
	.w5(32'hbbf2ed7b),
	.w6(32'h3be1b56a),
	.w7(32'hbc3fa987),
	.w8(32'hbce6a6ea),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc874869),
	.w1(32'h3c23a258),
	.w2(32'hbba974ce),
	.w3(32'h3b97c0f9),
	.w4(32'hbb95adcf),
	.w5(32'h3c0bb929),
	.w6(32'h3b2bc42d),
	.w7(32'h3a110cc4),
	.w8(32'h39e5c435),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35ea6d),
	.w1(32'h3aae7dfc),
	.w2(32'hbb4ea5bd),
	.w3(32'h39b4494f),
	.w4(32'h3b544526),
	.w5(32'h3c957f88),
	.w6(32'h3c351acb),
	.w7(32'hbbc39c51),
	.w8(32'hbb2074e3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57adf4),
	.w1(32'h3b8c828e),
	.w2(32'h3b39d90f),
	.w3(32'h3af73be2),
	.w4(32'h3c57552e),
	.w5(32'h3b7d004e),
	.w6(32'h3c3431cf),
	.w7(32'h3a20b124),
	.w8(32'hbbe4fc4c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf81b32),
	.w1(32'hbd28b18b),
	.w2(32'h3aead060),
	.w3(32'h3c1ebaa3),
	.w4(32'hbb7cf175),
	.w5(32'hb9e36d99),
	.w6(32'hbb08bb11),
	.w7(32'hbc121143),
	.w8(32'h3c1a1c39),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab982d0),
	.w1(32'h3b199be9),
	.w2(32'h39925e34),
	.w3(32'hbb990b1a),
	.w4(32'h39d03793),
	.w5(32'hbbc144ce),
	.w6(32'hb9f8164b),
	.w7(32'hbbf59448),
	.w8(32'hbaa6a936),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4b98a),
	.w1(32'h3b98ddf2),
	.w2(32'h3c3a1f46),
	.w3(32'hbbc3a945),
	.w4(32'hbc94ff74),
	.w5(32'h3a75e7af),
	.w6(32'h3c5567d7),
	.w7(32'h3c419fac),
	.w8(32'h3c30c9ea),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cd673),
	.w1(32'hbb1459a4),
	.w2(32'h3c30eedb),
	.w3(32'h3b951e20),
	.w4(32'hba25ab97),
	.w5(32'hbb8c91a8),
	.w6(32'hbad04cfa),
	.w7(32'h3bcb27f6),
	.w8(32'hbc5342b4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc095ed),
	.w1(32'hbb9f7934),
	.w2(32'h3c070705),
	.w3(32'h3d41f58d),
	.w4(32'h3c89fa28),
	.w5(32'hbcaf522a),
	.w6(32'hbbbed47d),
	.w7(32'h3ae54cce),
	.w8(32'h3b1ffce8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f7c440),
	.w1(32'h3c36a2a8),
	.w2(32'hbba9a779),
	.w3(32'hbc47a783),
	.w4(32'h3b90d705),
	.w5(32'h3be970e0),
	.w6(32'hbc048795),
	.w7(32'h3c83acfa),
	.w8(32'hbbc974b0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6f9e70),
	.w1(32'hbb9e1191),
	.w2(32'hba701ece),
	.w3(32'h3be45683),
	.w4(32'hbc0dcdee),
	.w5(32'h39321f5c),
	.w6(32'hbc1dfc85),
	.w7(32'hbc139ecf),
	.w8(32'hbb3c2e72),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f8dd7),
	.w1(32'h3baf48fd),
	.w2(32'hba6889fd),
	.w3(32'h3b6d57ab),
	.w4(32'hbba85ad0),
	.w5(32'hbbf47caa),
	.w6(32'hbd095450),
	.w7(32'hbc12a17f),
	.w8(32'hbb510c7d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d560d),
	.w1(32'h3b980df0),
	.w2(32'h3a3184ae),
	.w3(32'h3a8ca855),
	.w4(32'h3a9af3eb),
	.w5(32'hba9ea06c),
	.w6(32'hba14ddb9),
	.w7(32'h3af7db8a),
	.w8(32'hb8cb23fa),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35b2b0),
	.w1(32'h3d06c49d),
	.w2(32'h3c958c0c),
	.w3(32'h3bc5d919),
	.w4(32'hbc4d16f2),
	.w5(32'h3bdabc8b),
	.w6(32'h3c9a7edf),
	.w7(32'hbc2fff88),
	.w8(32'hbbc4076c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b87e42),
	.w1(32'h3be0e6cb),
	.w2(32'hbbadc357),
	.w3(32'hbb4e264e),
	.w4(32'h3b931ad1),
	.w5(32'h39f28587),
	.w6(32'hb7a97e34),
	.w7(32'h3c4dcb94),
	.w8(32'hbb213469),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2a2c1),
	.w1(32'hbbe02e05),
	.w2(32'hbbb5d104),
	.w3(32'hbb329483),
	.w4(32'hbd27924f),
	.w5(32'h3a535712),
	.w6(32'h3ad45e1d),
	.w7(32'hbc4e0678),
	.w8(32'hbb151168),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15b6d6),
	.w1(32'hbae648e1),
	.w2(32'h3b7c0c8f),
	.w3(32'hbbc4c259),
	.w4(32'h3c41c13d),
	.w5(32'h3bb17750),
	.w6(32'hbb59fa6e),
	.w7(32'h3bd8e288),
	.w8(32'h3a978d7f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9913031),
	.w1(32'hbc34f0f8),
	.w2(32'h3be192ea),
	.w3(32'hbb870d97),
	.w4(32'hbbf8ee5a),
	.w5(32'hbbc6cac0),
	.w6(32'hb9c53e25),
	.w7(32'hbc16e16a),
	.w8(32'h3c4d3acb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88fcc9),
	.w1(32'h3c131f3c),
	.w2(32'h3be61dc3),
	.w3(32'h3cd4a281),
	.w4(32'h3a44f209),
	.w5(32'hbbba0a06),
	.w6(32'hbaf803a6),
	.w7(32'hbba3172a),
	.w8(32'h3bbdecd9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule