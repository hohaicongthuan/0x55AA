module layer_10_featuremap_446(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc6dbb),
	.w1(32'h3b4e0a44),
	.w2(32'h3b3cab49),
	.w3(32'h3a99b753),
	.w4(32'h3986dbc5),
	.w5(32'h3a603fd1),
	.w6(32'hbb60c73b),
	.w7(32'h3a8fbc7b),
	.w8(32'hbb4dace0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36c99d),
	.w1(32'hbaa4bf1c),
	.w2(32'hba47b77e),
	.w3(32'h3b881320),
	.w4(32'hbb7e499c),
	.w5(32'hbaa3d851),
	.w6(32'hb9d698e8),
	.w7(32'hba9b9c98),
	.w8(32'hbb296404),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9ca8e),
	.w1(32'hba1bd1a2),
	.w2(32'hbba282ab),
	.w3(32'hbb37a6d7),
	.w4(32'hba9bfd8a),
	.w5(32'hbb883138),
	.w6(32'hbada713a),
	.w7(32'hbb622bfb),
	.w8(32'hbb95842c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6f86f),
	.w1(32'hbb859d8c),
	.w2(32'hb9d172ae),
	.w3(32'hbb72acb3),
	.w4(32'h3bc1df9d),
	.w5(32'h3c9ab101),
	.w6(32'hb7c62d81),
	.w7(32'h3bb66322),
	.w8(32'hbb750c50),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac47867),
	.w1(32'h3afd2909),
	.w2(32'hba2dab1f),
	.w3(32'h3b5608a4),
	.w4(32'h3a97a090),
	.w5(32'hbace5751),
	.w6(32'hbb583971),
	.w7(32'h38dbe550),
	.w8(32'hbb82023a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8f727),
	.w1(32'h3aeae1d5),
	.w2(32'h3af2f311),
	.w3(32'hba55d07f),
	.w4(32'h3acbd422),
	.w5(32'h3ae60d65),
	.w6(32'hbaa426e7),
	.w7(32'h3a096f5f),
	.w8(32'h3ba4f584),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33d29c),
	.w1(32'h3c1dc93a),
	.w2(32'h3b72a9c9),
	.w3(32'h3c162a44),
	.w4(32'h3bc0fb47),
	.w5(32'hbb9c0383),
	.w6(32'h3bec70a9),
	.w7(32'hbb242b51),
	.w8(32'hbbea47b6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985130f),
	.w1(32'hba153276),
	.w2(32'hbc0da094),
	.w3(32'hbb29c456),
	.w4(32'hbbbe38b1),
	.w5(32'hba54ff6e),
	.w6(32'hbb1ab648),
	.w7(32'hbbfabb8e),
	.w8(32'hbaa32a9b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec043a),
	.w1(32'h3b984cfb),
	.w2(32'h3aee47f1),
	.w3(32'hbb8fd195),
	.w4(32'h3a83acd7),
	.w5(32'hbb0ea477),
	.w6(32'h3b0a15e6),
	.w7(32'hb8cbdec3),
	.w8(32'h3a06d1e1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46fb7f),
	.w1(32'hb8fa7e25),
	.w2(32'hb98f320c),
	.w3(32'hbadf0c53),
	.w4(32'h3bda050e),
	.w5(32'h3bf182bd),
	.w6(32'h3b695110),
	.w7(32'h3b2acd38),
	.w8(32'hb995d482),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8e294),
	.w1(32'h39324e49),
	.w2(32'h3b6b72c1),
	.w3(32'h3c01dcd6),
	.w4(32'h3b2df072),
	.w5(32'h3b7da901),
	.w6(32'h3be95d3a),
	.w7(32'h3abf2d78),
	.w8(32'h3a117551),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e3087),
	.w1(32'h3c06c3b3),
	.w2(32'hbb1eb267),
	.w3(32'h3c32fb66),
	.w4(32'h3b524231),
	.w5(32'hbbf43475),
	.w6(32'h3bdd9719),
	.w7(32'hba0517dd),
	.w8(32'hbb7e136a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f5d54),
	.w1(32'hbba4e6c3),
	.w2(32'hbc056cc8),
	.w3(32'h3ac27513),
	.w4(32'hbb98f086),
	.w5(32'hbb63d87a),
	.w6(32'h3c0f2af4),
	.w7(32'hbb516bd2),
	.w8(32'hbbdb5197),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dcaa0),
	.w1(32'hb88c8f6e),
	.w2(32'h3b0d1be2),
	.w3(32'hbb066fb6),
	.w4(32'hba9bf289),
	.w5(32'h3b539f27),
	.w6(32'hbb2c80b7),
	.w7(32'h3b17ab8e),
	.w8(32'h3bf45288),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adede67),
	.w1(32'hb9fbc65b),
	.w2(32'h3a423699),
	.w3(32'h3ba15b0e),
	.w4(32'h3b9f1420),
	.w5(32'hbab566ea),
	.w6(32'h3bdf8e4d),
	.w7(32'h3be80881),
	.w8(32'h3bc1aea0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad45113),
	.w1(32'hbb88e218),
	.w2(32'hbb7f2f15),
	.w3(32'h3a00e96c),
	.w4(32'hbba85cf6),
	.w5(32'hbbee0433),
	.w6(32'h3a9a6f8f),
	.w7(32'hbb7acd68),
	.w8(32'h3952ad11),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc5905),
	.w1(32'h3ba0bf88),
	.w2(32'h3b7b9d7a),
	.w3(32'hbb0e41a3),
	.w4(32'hb8be3302),
	.w5(32'h3a5b68a2),
	.w6(32'h38873ec8),
	.w7(32'h3b689a9e),
	.w8(32'h3b8f6f4a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dc99a),
	.w1(32'hbb364ad3),
	.w2(32'hbc052b1d),
	.w3(32'hba63ffba),
	.w4(32'hbc17c881),
	.w5(32'hbc255118),
	.w6(32'h3b1b099e),
	.w7(32'hbc3cb3c3),
	.w8(32'hbc019b5d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae82a2),
	.w1(32'hbbdb67ff),
	.w2(32'hbc08a79a),
	.w3(32'hbb2c1560),
	.w4(32'hbbcf7ca0),
	.w5(32'hbc456e2b),
	.w6(32'hbaeafa39),
	.w7(32'hbb9c05ce),
	.w8(32'hbbcf095a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7368),
	.w1(32'h3a9144e3),
	.w2(32'h3bd12683),
	.w3(32'hbb86e2ca),
	.w4(32'hbab7e5c2),
	.w5(32'h3902ae22),
	.w6(32'hba2176f5),
	.w7(32'h3b0ad3d4),
	.w8(32'hbb05d6e0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0bd8b),
	.w1(32'hbbcc78de),
	.w2(32'hbba141b6),
	.w3(32'h3b8cee07),
	.w4(32'hbb890b0e),
	.w5(32'hbb00d0ee),
	.w6(32'hba570c8d),
	.w7(32'h39d36f8a),
	.w8(32'h3b634e68),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4a53),
	.w1(32'hbba9b3d8),
	.w2(32'h387ead23),
	.w3(32'hb9e1be99),
	.w4(32'h3ad9b98f),
	.w5(32'hb9ef06ff),
	.w6(32'h3b1cc7f6),
	.w7(32'hbaf9e09b),
	.w8(32'h38040bc9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c2e06),
	.w1(32'hbbd54c49),
	.w2(32'hbc91ea1c),
	.w3(32'h3ba4a2ee),
	.w4(32'hbb87f290),
	.w5(32'hbc5217d1),
	.w6(32'hba46fa4b),
	.w7(32'hbc5c2bd6),
	.w8(32'hbc7203c0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ad01b),
	.w1(32'hbb4d3f3c),
	.w2(32'hbb914f4f),
	.w3(32'hbaf9ce7d),
	.w4(32'hbaf24e6a),
	.w5(32'hbaef509b),
	.w6(32'hbb3f2638),
	.w7(32'h3a48552f),
	.w8(32'hbb71f5fb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdccb0),
	.w1(32'h3a8ff24d),
	.w2(32'h3bea94fc),
	.w3(32'h3a43698e),
	.w4(32'h3ba500f1),
	.w5(32'hbb1d0787),
	.w6(32'h38c88d10),
	.w7(32'h3b1ba24e),
	.w8(32'h3b43dc49),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6551c0),
	.w1(32'h3a7d0ee9),
	.w2(32'h39a56a78),
	.w3(32'hbbb64b05),
	.w4(32'h3b4429b0),
	.w5(32'h3b9f52e2),
	.w6(32'hbaf9c2f4),
	.w7(32'h3b6d9743),
	.w8(32'h3ae5e4e9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2a5e9),
	.w1(32'h3c1e211e),
	.w2(32'h3b961a06),
	.w3(32'hb8e4e862),
	.w4(32'h3b1f763f),
	.w5(32'hb898a431),
	.w6(32'h3bd7a111),
	.w7(32'h3afa90d5),
	.w8(32'h3c1ca9b5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9b22f),
	.w1(32'h3b162fc3),
	.w2(32'h3ab34b85),
	.w3(32'h3b40568b),
	.w4(32'h3bae6f41),
	.w5(32'hbb5294db),
	.w6(32'h3c4cadef),
	.w7(32'hba248782),
	.w8(32'hb9ad34b5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9559aa),
	.w1(32'h3c1505d2),
	.w2(32'h3c2c0c8d),
	.w3(32'h3acf52df),
	.w4(32'h3bc29d25),
	.w5(32'h3a86e551),
	.w6(32'h3b80fda3),
	.w7(32'h39544cb8),
	.w8(32'h3be3268b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ab374),
	.w1(32'h3bb90aad),
	.w2(32'h3b4f9925),
	.w3(32'h3a060464),
	.w4(32'h3ae5ec0c),
	.w5(32'h3b8a7fca),
	.w6(32'h3b9ec357),
	.w7(32'h3ab620d1),
	.w8(32'h3bc61e4d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8521f25),
	.w1(32'h3b10494b),
	.w2(32'h3a9a49f1),
	.w3(32'h3b177dfd),
	.w4(32'hbb7b1a60),
	.w5(32'hbb13e565),
	.w6(32'hba6a15a8),
	.w7(32'hbb3c83d9),
	.w8(32'hbb556e67),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bd76f),
	.w1(32'h3b00de55),
	.w2(32'h3963cbcd),
	.w3(32'h3a720c1f),
	.w4(32'hbb4e5400),
	.w5(32'hbbcd8fbc),
	.w6(32'h3a662652),
	.w7(32'hbb592251),
	.w8(32'hbb123431),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba523c89),
	.w1(32'h3ad3108d),
	.w2(32'hbac56c0d),
	.w3(32'hbb9c3427),
	.w4(32'hbb957b4a),
	.w5(32'hbc0e45da),
	.w6(32'hbb18c8c4),
	.w7(32'hbb092f0e),
	.w8(32'hbb40cd9a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d9392),
	.w1(32'h39339b38),
	.w2(32'h3b10766f),
	.w3(32'hbbd6ecd0),
	.w4(32'hbab14cc9),
	.w5(32'hbbc87cc8),
	.w6(32'h3899c1b2),
	.w7(32'hba02b211),
	.w8(32'h39e0a9bd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97fb72),
	.w1(32'hbc0281dc),
	.w2(32'hbbca68fe),
	.w3(32'hbb88f69d),
	.w4(32'hbb82a78e),
	.w5(32'hbb0d55f9),
	.w6(32'hb9e4f67d),
	.w7(32'h3a8ccc87),
	.w8(32'h3b5d2445),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eae90),
	.w1(32'h3b4e1e9f),
	.w2(32'h3b45aee3),
	.w3(32'h3b6056ed),
	.w4(32'h3acb4116),
	.w5(32'h3ba1d938),
	.w6(32'h3b09a906),
	.w7(32'h3ae3ce48),
	.w8(32'hba4293b1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb08e6d),
	.w1(32'h3c27fff6),
	.w2(32'hbb9f271b),
	.w3(32'h3c25e354),
	.w4(32'h3c5fdf76),
	.w5(32'h3bfef0a4),
	.w6(32'h3bf6ddbd),
	.w7(32'h3c79a138),
	.w8(32'hba71a489),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad20685),
	.w1(32'h3b849dc5),
	.w2(32'h3bd8af4f),
	.w3(32'h3b0a33d8),
	.w4(32'h3b634c19),
	.w5(32'h3b3c2515),
	.w6(32'hb9b7316f),
	.w7(32'h3b23adde),
	.w8(32'hb971802b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6653f),
	.w1(32'hbba3dd9b),
	.w2(32'h3b369db2),
	.w3(32'hbb4eb5b9),
	.w4(32'hbb0ada2e),
	.w5(32'hbbf6b87d),
	.w6(32'h3b4ab77e),
	.w7(32'hbb0b4214),
	.w8(32'hba8614ed),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4722a4),
	.w1(32'hba68a72b),
	.w2(32'h3adaf8d1),
	.w3(32'hbb0ef824),
	.w4(32'h3a8d18bb),
	.w5(32'h3b04b96b),
	.w6(32'hbb298d05),
	.w7(32'hba3ad44f),
	.w8(32'hbb20bdd4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb900c22),
	.w1(32'h3b9e8d2c),
	.w2(32'h3b08b240),
	.w3(32'hbb1d4df8),
	.w4(32'hb9af2078),
	.w5(32'h3a5b6f2d),
	.w6(32'h3b232465),
	.w7(32'h3b89dc66),
	.w8(32'h3aa30834),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a0965),
	.w1(32'hbac10ced),
	.w2(32'hbb6ce726),
	.w3(32'hbb295859),
	.w4(32'hbae763e0),
	.w5(32'hbb87ca59),
	.w6(32'h3a6eced0),
	.w7(32'h3a956410),
	.w8(32'h3ac58781),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81b3ce),
	.w1(32'h3a47e45f),
	.w2(32'h3b13d389),
	.w3(32'hbb442c32),
	.w4(32'h3aeac897),
	.w5(32'h3c10cef8),
	.w6(32'hbb9490c9),
	.w7(32'hbb355150),
	.w8(32'hbb44b165),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54b83f),
	.w1(32'hbc578109),
	.w2(32'hbb15e85e),
	.w3(32'hbb86e1a0),
	.w4(32'hbbcc4544),
	.w5(32'hbaa0b13f),
	.w6(32'hbbd43e62),
	.w7(32'h3b8ba53b),
	.w8(32'h3acfc890),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af93c9a),
	.w1(32'h3b970735),
	.w2(32'h3a883ff5),
	.w3(32'hbb8688da),
	.w4(32'h3a3e47f1),
	.w5(32'hbb582cfa),
	.w6(32'hb9f68394),
	.w7(32'h3ae5ed53),
	.w8(32'hb9a0fca8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6d82f),
	.w1(32'hbacf22d8),
	.w2(32'hba88ec52),
	.w3(32'h39a4f45c),
	.w4(32'hbb51e0d5),
	.w5(32'hbb5f357c),
	.w6(32'h3c0cd426),
	.w7(32'hba6ca302),
	.w8(32'h3b9d1d06),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24f2d6),
	.w1(32'hbc10c2d1),
	.w2(32'hbbc3f42a),
	.w3(32'hbb21f412),
	.w4(32'hbab2af5b),
	.w5(32'h3be99d98),
	.w6(32'hbb2c8e49),
	.w7(32'hbac52807),
	.w8(32'hbb84c1ac),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace8d77),
	.w1(32'hbbedcf1d),
	.w2(32'hbc629a3e),
	.w3(32'hbaf14d52),
	.w4(32'hbbe47d96),
	.w5(32'hbc5ef687),
	.w6(32'hbbb4cac9),
	.w7(32'hbc0e69e1),
	.w8(32'hbc2aef56),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39897e0a),
	.w1(32'h3b8ed2ca),
	.w2(32'h3bc4c670),
	.w3(32'hb93138ad),
	.w4(32'h3b74cb84),
	.w5(32'h3b7a64ea),
	.w6(32'h3a09c0e6),
	.w7(32'h3b2fafda),
	.w8(32'h3ba55b3a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b226ded),
	.w1(32'h3a2e5526),
	.w2(32'h3b2bfff5),
	.w3(32'h3a912777),
	.w4(32'h389132a2),
	.w5(32'hba421d4a),
	.w6(32'h3a30d6f9),
	.w7(32'h3af22c22),
	.w8(32'hba22aa7d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5578d4),
	.w1(32'hb94fdeca),
	.w2(32'hba6a8b42),
	.w3(32'hbb289fdc),
	.w4(32'hb95f0367),
	.w5(32'hbbaf0295),
	.w6(32'hbac82b63),
	.w7(32'hba29e8b2),
	.w8(32'hbb62fd6d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fadc5),
	.w1(32'hbb872d01),
	.w2(32'hbb7ea797),
	.w3(32'hbbbb0b1e),
	.w4(32'h3a3281a1),
	.w5(32'hbb08ac8e),
	.w6(32'hba8359b5),
	.w7(32'hba4552ce),
	.w8(32'h3ae6c061),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e8308),
	.w1(32'hb9c08364),
	.w2(32'hbae4f577),
	.w3(32'h3b020d64),
	.w4(32'hbbaad577),
	.w5(32'hbb9f6d6b),
	.w6(32'h3b762a8a),
	.w7(32'hbba815d3),
	.w8(32'hbabbafe1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc97f3e),
	.w1(32'hbc2627b3),
	.w2(32'hbc9740e7),
	.w3(32'hbbf77c16),
	.w4(32'hbc477673),
	.w5(32'hbc46caa2),
	.w6(32'hbb069876),
	.w7(32'hbc334593),
	.w8(32'hbc0713ac),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fe035),
	.w1(32'hba9370a1),
	.w2(32'hbb6571fd),
	.w3(32'hbc0eab93),
	.w4(32'hba62815e),
	.w5(32'hba5cc37a),
	.w6(32'hbad33345),
	.w7(32'h3b137c27),
	.w8(32'h39d5479b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4175),
	.w1(32'h3a75f19d),
	.w2(32'hba08f98d),
	.w3(32'hbb097ec7),
	.w4(32'hbb90f4a2),
	.w5(32'hbbcb3223),
	.w6(32'hb9fd4213),
	.w7(32'hbbf0f2bc),
	.w8(32'hbbce2c90),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb900e02),
	.w1(32'hb96df3e7),
	.w2(32'hbb5f1557),
	.w3(32'hbb96e750),
	.w4(32'hb7a2b734),
	.w5(32'hba5794ba),
	.w6(32'hba97b6d1),
	.w7(32'h3a4ef9e3),
	.w8(32'h3a74c25e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68887),
	.w1(32'hbaffbd81),
	.w2(32'h3a59ca99),
	.w3(32'h3a6ef14b),
	.w4(32'hbb38ddaa),
	.w5(32'h38834136),
	.w6(32'h3ab03576),
	.w7(32'hbb12a402),
	.w8(32'h3b1483c2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db3e4b),
	.w1(32'h3bba9bff),
	.w2(32'hba209b9c),
	.w3(32'h3a53f08b),
	.w4(32'h3b607183),
	.w5(32'hbb28ca0d),
	.w6(32'hbb66f05f),
	.w7(32'h3b041627),
	.w8(32'hbb3f7b03),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c7f346),
	.w1(32'hbb19088e),
	.w2(32'h39f89a79),
	.w3(32'h398b88ad),
	.w4(32'hbb1d87f7),
	.w5(32'hbbb9fa53),
	.w6(32'hba0130cb),
	.w7(32'h3b86fe4c),
	.w8(32'h3b014458),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d8e83),
	.w1(32'hbb2418a5),
	.w2(32'hbb7062fe),
	.w3(32'hbbbabf26),
	.w4(32'hbc0f1c8b),
	.w5(32'hbc2aa40f),
	.w6(32'hb9e8de59),
	.w7(32'hbaeaa2fb),
	.w8(32'hbb5aa2c3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba669b64),
	.w1(32'h3aa9280c),
	.w2(32'h3ba3af60),
	.w3(32'hbc063c6e),
	.w4(32'h3af27ce3),
	.w5(32'hbb0e43e0),
	.w6(32'hbb9f49a2),
	.w7(32'hb985283f),
	.w8(32'h3a878f1b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9723a),
	.w1(32'hbada4461),
	.w2(32'hb91ed694),
	.w3(32'h3bf08bb5),
	.w4(32'h3b170594),
	.w5(32'h3a2b68d5),
	.w6(32'h3b9cb8eb),
	.w7(32'h3a39d566),
	.w8(32'hbbe977c5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0438d),
	.w1(32'h3afc08f9),
	.w2(32'hb99d6655),
	.w3(32'hbc01365b),
	.w4(32'hbb186672),
	.w5(32'hbb20903a),
	.w6(32'hbbce550b),
	.w7(32'hbb1df8a7),
	.w8(32'hbb854072),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43a537),
	.w1(32'h3aebfce6),
	.w2(32'h3adef144),
	.w3(32'h3a940d2b),
	.w4(32'h3aeaf6bd),
	.w5(32'h3ba5553c),
	.w6(32'h3a3daa7f),
	.w7(32'h3b3ce276),
	.w8(32'h3b324ef7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b565c2f),
	.w1(32'h3ac58607),
	.w2(32'h3b2fae64),
	.w3(32'h3b8873fc),
	.w4(32'hbb928942),
	.w5(32'hbb770385),
	.w6(32'h3ba3af0a),
	.w7(32'hbabb5555),
	.w8(32'h3b0ae697),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5341),
	.w1(32'hbb193e7b),
	.w2(32'hbbe8c3b9),
	.w3(32'h3b0cd447),
	.w4(32'h39dc00eb),
	.w5(32'h3aec0cc7),
	.w6(32'h3b6e2a17),
	.w7(32'hb97fd32b),
	.w8(32'h3b430bae),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa208fd),
	.w1(32'h3b1f88de),
	.w2(32'h3abb77d5),
	.w3(32'h3ba2b293),
	.w4(32'h3b548e40),
	.w5(32'hb8aab0ea),
	.w6(32'h3bdf8e61),
	.w7(32'h3b877193),
	.w8(32'h3a91277d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87967d),
	.w1(32'hbbcab49d),
	.w2(32'h39e17a9e),
	.w3(32'h394699e1),
	.w4(32'h3b5f958d),
	.w5(32'hbb3df2ef),
	.w6(32'hbb4230fa),
	.w7(32'h3926cd52),
	.w8(32'hba884a3e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a308cf8),
	.w1(32'h3c0c1a9d),
	.w2(32'hba897b08),
	.w3(32'h3b3bb2ec),
	.w4(32'h3c0bd801),
	.w5(32'hbbe78270),
	.w6(32'h3b4903f6),
	.w7(32'h3c7b8e4a),
	.w8(32'hbbf1fb5d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59c43f),
	.w1(32'h3c01776a),
	.w2(32'h3c90dc83),
	.w3(32'hbc4846a2),
	.w4(32'h3c91e253),
	.w5(32'h3c6cb76a),
	.w6(32'hbbe8ff11),
	.w7(32'h3c7451b6),
	.w8(32'h3cf4793e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c882328),
	.w1(32'h3c6b307c),
	.w2(32'hba233ed5),
	.w3(32'h3d0212c4),
	.w4(32'hbbb02d4b),
	.w5(32'h3ba559fe),
	.w6(32'h3c299fd1),
	.w7(32'h3b30ae91),
	.w8(32'h3a4b26ad),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac696d),
	.w1(32'h3b9b1834),
	.w2(32'h3c0c6f2d),
	.w3(32'hbbfce3b6),
	.w4(32'h3b2bbf25),
	.w5(32'h3bd1db51),
	.w6(32'h3ba22eac),
	.w7(32'h3b42ee09),
	.w8(32'h3affd09b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082a95),
	.w1(32'hbc200692),
	.w2(32'h3a7353a2),
	.w3(32'hbc8a5497),
	.w4(32'hb944a55f),
	.w5(32'h3ba50e45),
	.w6(32'hbc3b9853),
	.w7(32'hbb6c97d4),
	.w8(32'hbb4f3f35),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8fc6),
	.w1(32'h39d1261a),
	.w2(32'h3814dfd8),
	.w3(32'h3bab2e80),
	.w4(32'h3be878cd),
	.w5(32'h3c9e9930),
	.w6(32'h3a062a40),
	.w7(32'h3a33434e),
	.w8(32'hbbf2fc0a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d4eec),
	.w1(32'h3a11b1a2),
	.w2(32'hbba08b70),
	.w3(32'h3c333bce),
	.w4(32'h3b08a800),
	.w5(32'hbabed2be),
	.w6(32'hbbb0e80f),
	.w7(32'hbb2a686b),
	.w8(32'hbc2d3dda),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ae43a),
	.w1(32'h3bcb2774),
	.w2(32'hbbd8fc1c),
	.w3(32'hbb6d858e),
	.w4(32'h3a324435),
	.w5(32'hbc79b3ab),
	.w6(32'hbb3845ae),
	.w7(32'h3bb56b95),
	.w8(32'hbc412d90),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b4d00),
	.w1(32'hbbc40836),
	.w2(32'h3ad6443e),
	.w3(32'hbb45958a),
	.w4(32'hba84e583),
	.w5(32'hbbaf3f53),
	.w6(32'h3b0e72d7),
	.w7(32'h3b838df7),
	.w8(32'h3bbcc416),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc206ec3),
	.w1(32'hbc5ba1e4),
	.w2(32'hbbc0a391),
	.w3(32'hbc32dcbd),
	.w4(32'hbb869430),
	.w5(32'h3aefa73f),
	.w6(32'hbbf36313),
	.w7(32'hbb940394),
	.w8(32'hbb863ce0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947fd2),
	.w1(32'hbaae825a),
	.w2(32'hbb2bd531),
	.w3(32'hba59b1ae),
	.w4(32'hbbf71e0e),
	.w5(32'hbc0d4a9c),
	.w6(32'hbb585358),
	.w7(32'hbc031317),
	.w8(32'hbc5f188b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc282fe6),
	.w1(32'hbc30faa1),
	.w2(32'hbc3b9389),
	.w3(32'hbc5c52e3),
	.w4(32'hbb8d419b),
	.w5(32'hbc42b2a8),
	.w6(32'hbc6292b2),
	.w7(32'hbb5a3deb),
	.w8(32'hbace5e2e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f542e2),
	.w1(32'hb935ec09),
	.w2(32'h3b3e9e20),
	.w3(32'h3b6316db),
	.w4(32'h3b552de2),
	.w5(32'hbae76cd5),
	.w6(32'h3cb128bd),
	.w7(32'h3b323111),
	.w8(32'h3c016dfd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67b59c),
	.w1(32'hbbdf0b81),
	.w2(32'hbb321b6e),
	.w3(32'h3c64db47),
	.w4(32'hbc0f06c7),
	.w5(32'h3b22b7de),
	.w6(32'h3c45ca48),
	.w7(32'hba2edabb),
	.w8(32'h3b2a4e81),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5332fb),
	.w1(32'h3bbd6a03),
	.w2(32'hba9682a6),
	.w3(32'h3b5df72a),
	.w4(32'h3b66776c),
	.w5(32'h3b537527),
	.w6(32'h3b681f1b),
	.w7(32'h3c0464ff),
	.w8(32'h3c02a480),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae99714),
	.w1(32'h3a93e403),
	.w2(32'h3c1bd043),
	.w3(32'h3c26058a),
	.w4(32'hbb11ab0d),
	.w5(32'hb963e567),
	.w6(32'hbc056180),
	.w7(32'hb9876b78),
	.w8(32'h3c168525),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1b9c7),
	.w1(32'h3c08612f),
	.w2(32'h3b4523ed),
	.w3(32'h3bb65665),
	.w4(32'h3b409054),
	.w5(32'h3d02cdea),
	.w6(32'h3bec7602),
	.w7(32'h3b84b9d5),
	.w8(32'h3c39a2e8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39befe88),
	.w1(32'h3bb59297),
	.w2(32'h3b92b58d),
	.w3(32'hbb386300),
	.w4(32'h3b7c27ec),
	.w5(32'hbb75e24e),
	.w6(32'hbbbdac3b),
	.w7(32'h3a9a0d65),
	.w8(32'hbc7cb304),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab52e29),
	.w1(32'hbbd5fbb6),
	.w2(32'hbaf8eb3d),
	.w3(32'h3b92f818),
	.w4(32'hbbbfb350),
	.w5(32'hbb66f8e0),
	.w6(32'hbbf9eb7f),
	.w7(32'hb9e39952),
	.w8(32'hbc2ae9bc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e611c),
	.w1(32'hbb6f2896),
	.w2(32'hbbc3a9f3),
	.w3(32'h3a9cccc7),
	.w4(32'h3b6296bc),
	.w5(32'hba75b686),
	.w6(32'hbc2ccef9),
	.w7(32'h3c05bdd9),
	.w8(32'h3c494e37),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba667d38),
	.w1(32'hbb91cc45),
	.w2(32'hbc6a06e6),
	.w3(32'h3c99143b),
	.w4(32'hbc01217f),
	.w5(32'hbc773c7d),
	.w6(32'hba707d45),
	.w7(32'hbc1ad913),
	.w8(32'hbc2e708f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f9e8),
	.w1(32'hbc0b6439),
	.w2(32'h3b508e66),
	.w3(32'hbb3d5c32),
	.w4(32'hb9a5a3ec),
	.w5(32'h3c0b5fb7),
	.w6(32'hbbc8f6f7),
	.w7(32'h3954c99b),
	.w8(32'h3c8683f5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c431e),
	.w1(32'h3b1aac2f),
	.w2(32'hbc4bf892),
	.w3(32'h3d149dfc),
	.w4(32'h3c8718eb),
	.w5(32'h3b6194c5),
	.w6(32'h3cbc8ac6),
	.w7(32'hbc28cf96),
	.w8(32'hbc81e2de),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90d09),
	.w1(32'hba1b7a52),
	.w2(32'hbb72a8fb),
	.w3(32'h3c9dbacf),
	.w4(32'hbb818c09),
	.w5(32'hbbad76f3),
	.w6(32'hbadf865f),
	.w7(32'hbc0c2ac9),
	.w8(32'hbaafde77),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1122bb),
	.w1(32'hbc1dcf10),
	.w2(32'hbc75ecdf),
	.w3(32'hbb4d781b),
	.w4(32'hb91413a1),
	.w5(32'hbbe349db),
	.w6(32'h3a99d026),
	.w7(32'hbbee4784),
	.w8(32'hbba0667c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde2fba),
	.w1(32'h3bcd5e07),
	.w2(32'hbbebc6a1),
	.w3(32'h3b29537d),
	.w4(32'h3c7850eb),
	.w5(32'h3c646e26),
	.w6(32'h3bdb0405),
	.w7(32'h3bdfc19f),
	.w8(32'h3c4ebd71),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104ad2),
	.w1(32'h3994325e),
	.w2(32'hbba1bd67),
	.w3(32'h3ca89572),
	.w4(32'h3b227ae8),
	.w5(32'h3bade1ad),
	.w6(32'h3bda61f1),
	.w7(32'h3aa6b2a4),
	.w8(32'hbb2bf353),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64ccf3),
	.w1(32'h3b56b06a),
	.w2(32'h3a23c796),
	.w3(32'hba17cd25),
	.w4(32'h3b5201a4),
	.w5(32'h3be8f39b),
	.w6(32'hb9c94c80),
	.w7(32'h3b3999d2),
	.w8(32'h3c0ea229),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390597),
	.w1(32'h398adee4),
	.w2(32'hbb8846b4),
	.w3(32'hbbb21585),
	.w4(32'hba92428a),
	.w5(32'hbad5b9be),
	.w6(32'hbc8a2a5f),
	.w7(32'h3afb09ba),
	.w8(32'hbbd088bd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387d28f1),
	.w1(32'h3c1523ff),
	.w2(32'hbbff1c80),
	.w3(32'hbaa22ef3),
	.w4(32'h3bcaa087),
	.w5(32'h3ac0eb7b),
	.w6(32'h38d650a4),
	.w7(32'h3b23b3e9),
	.w8(32'hbbe37865),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17570b),
	.w1(32'h3972fa90),
	.w2(32'hbb98abe9),
	.w3(32'h3bdf9a52),
	.w4(32'hb98b35fa),
	.w5(32'hbc0e221f),
	.w6(32'h3b00ec96),
	.w7(32'hbb9e7426),
	.w8(32'hbc8d9af0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf7cc1),
	.w1(32'hbb39c96b),
	.w2(32'h3ad181e4),
	.w3(32'hbc4258ec),
	.w4(32'h3c0f66f7),
	.w5(32'h3c84740e),
	.w6(32'hbc9270bf),
	.w7(32'h3b5e9e1d),
	.w8(32'h3c5b1512),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9a477),
	.w1(32'hbbab818c),
	.w2(32'hbb8a86ce),
	.w3(32'h3c80ac87),
	.w4(32'hbb8aad42),
	.w5(32'hbb57d197),
	.w6(32'h3c1e5a43),
	.w7(32'hbb88afcb),
	.w8(32'h3a8eaf95),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba14c98),
	.w1(32'h3b807b05),
	.w2(32'hbbeb4690),
	.w3(32'hbbc1dc4d),
	.w4(32'h3b925db8),
	.w5(32'h3b98b72f),
	.w6(32'hbbde9abd),
	.w7(32'h3bc2b126),
	.w8(32'hbc093bf9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8ff3a),
	.w1(32'hb851e993),
	.w2(32'h3c0d55b9),
	.w3(32'hbb20f3ea),
	.w4(32'hb994b8aa),
	.w5(32'h3bbf4dee),
	.w6(32'hbc303a68),
	.w7(32'hbb32d4f5),
	.w8(32'h3c29e646),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93e549),
	.w1(32'hbc835567),
	.w2(32'hbc980a1f),
	.w3(32'hbbc96bdc),
	.w4(32'hbb60d1e5),
	.w5(32'hbc38f054),
	.w6(32'hbab37266),
	.w7(32'h3b174291),
	.w8(32'h3b558f4b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35359c),
	.w1(32'hb9cf3c8a),
	.w2(32'hbb9969bc),
	.w3(32'h3c4ae473),
	.w4(32'h3b93874b),
	.w5(32'h391eca34),
	.w6(32'h3c29503d),
	.w7(32'h3c51a19d),
	.w8(32'h3b2fdcee),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb58e2b),
	.w1(32'hbb0cf244),
	.w2(32'hba573136),
	.w3(32'h3abf2759),
	.w4(32'h3a93d094),
	.w5(32'h3a12ae34),
	.w6(32'h3b17eaa7),
	.w7(32'h3b805842),
	.w8(32'h3c160bbe),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad743e2),
	.w1(32'hbc170d18),
	.w2(32'hbad4adf1),
	.w3(32'h3ad77bf5),
	.w4(32'hb94e39c1),
	.w5(32'hbb7fde97),
	.w6(32'hbb18b68a),
	.w7(32'h3a4a15cc),
	.w8(32'h3af8266d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa951d),
	.w1(32'hbbcd9783),
	.w2(32'hbb404d69),
	.w3(32'hbc649210),
	.w4(32'hbba768fb),
	.w5(32'hbbb450f0),
	.w6(32'hbc05fe52),
	.w7(32'hbb71f15f),
	.w8(32'hbc06ea8f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba31bc6),
	.w1(32'hbc51b734),
	.w2(32'hbc392a70),
	.w3(32'hbb063141),
	.w4(32'hbb412a1e),
	.w5(32'hbc4ccd42),
	.w6(32'h3abf26d8),
	.w7(32'hbb19a5cd),
	.w8(32'hbb71a73f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42d7cf),
	.w1(32'h3c53a395),
	.w2(32'hbbeb0381),
	.w3(32'hbb957dbf),
	.w4(32'h3b10bc45),
	.w5(32'h39951da1),
	.w6(32'hbc42fc5a),
	.w7(32'hbb0adc19),
	.w8(32'h3c1a22fb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbca8ca),
	.w1(32'h3bea55bb),
	.w2(32'hb9ab5f99),
	.w3(32'hb903322a),
	.w4(32'h3bdc1fee),
	.w5(32'hbc2d8e4a),
	.w6(32'h3bc4da36),
	.w7(32'h393c1288),
	.w8(32'hbbcff80f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca03d5),
	.w1(32'h3b09b347),
	.w2(32'hb9bc9219),
	.w3(32'hbc96b2b0),
	.w4(32'h3b90270d),
	.w5(32'hb9560a86),
	.w6(32'hbc3dea88),
	.w7(32'h3c31fdf1),
	.w8(32'h3b01aad1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b209e7d),
	.w1(32'hbb00f94e),
	.w2(32'hbc0c6f28),
	.w3(32'h3b19896b),
	.w4(32'h3c189cd5),
	.w5(32'hbb83cb41),
	.w6(32'hbb0b85ba),
	.w7(32'hbc043732),
	.w8(32'hbba970e9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb953f52),
	.w1(32'hbb475398),
	.w2(32'hbc0a9bad),
	.w3(32'hbb77497e),
	.w4(32'hbb9559a8),
	.w5(32'hbb978139),
	.w6(32'hbb3fe8d3),
	.w7(32'hbb29f4a6),
	.w8(32'hbc37db61),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed08c),
	.w1(32'h3c3c8e30),
	.w2(32'h3ca0c333),
	.w3(32'hba4fc5ea),
	.w4(32'h3c6c277c),
	.w5(32'h3c86f029),
	.w6(32'h3ab171f4),
	.w7(32'h3c9e9676),
	.w8(32'h3c6d5b03),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4b94f),
	.w1(32'hb9179fb9),
	.w2(32'hba925611),
	.w3(32'h3c3df2e5),
	.w4(32'h3b401f93),
	.w5(32'h3be04aba),
	.w6(32'h3be38e74),
	.w7(32'h3b565ff6),
	.w8(32'h39a9d9bb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20990f),
	.w1(32'h3ac96455),
	.w2(32'h3a18136f),
	.w3(32'h3c0002d2),
	.w4(32'h3b665ec1),
	.w5(32'hbb6ae3d7),
	.w6(32'h3be5c000),
	.w7(32'h3b3e1d2f),
	.w8(32'hbb90bbc2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b195d9c),
	.w1(32'hbb448e1b),
	.w2(32'hbbad93fd),
	.w3(32'hba0bee11),
	.w4(32'hbc47a9f7),
	.w5(32'hbbbf0bfa),
	.w6(32'h3c044fc1),
	.w7(32'hbbf9d9b6),
	.w8(32'hbbe38618),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f3f4b),
	.w1(32'hbb859e6e),
	.w2(32'hbbb7988b),
	.w3(32'hbc2e186a),
	.w4(32'hb996cd17),
	.w5(32'h3bce8a21),
	.w6(32'hbc0534b8),
	.w7(32'h3b14bc5e),
	.w8(32'hbba04601),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6e4de),
	.w1(32'hbb7cd72e),
	.w2(32'h3b30e1ae),
	.w3(32'hbbf35c91),
	.w4(32'hbb31bb48),
	.w5(32'hbc03907a),
	.w6(32'hbc09d991),
	.w7(32'hba9b3f5f),
	.w8(32'hbbbe79da),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29b7f6),
	.w1(32'hbb928f27),
	.w2(32'hbbb22f18),
	.w3(32'h3c4d9371),
	.w4(32'hbaad44c3),
	.w5(32'hbc3849b5),
	.w6(32'h3bce8be9),
	.w7(32'hbc0041d2),
	.w8(32'hbc12d586),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08ef94),
	.w1(32'h3bee1cc5),
	.w2(32'h3c40b210),
	.w3(32'hbc3b6cb5),
	.w4(32'h3c11f876),
	.w5(32'h3c7d1f6e),
	.w6(32'hbc98749d),
	.w7(32'h3c51995f),
	.w8(32'h3cb9f923),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84c383),
	.w1(32'hbc02e0c6),
	.w2(32'hbb0960eb),
	.w3(32'h3cad8781),
	.w4(32'h3a22e839),
	.w5(32'h3bf7967b),
	.w6(32'hb918905a),
	.w7(32'hb9d4ee1e),
	.w8(32'h3bf91ff7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3834b6bc),
	.w1(32'h3c6520d6),
	.w2(32'h3c174757),
	.w3(32'h3a36c0c2),
	.w4(32'h3bfe0fd5),
	.w5(32'hba447bc4),
	.w6(32'hbb6b46fa),
	.w7(32'h3bf43dc2),
	.w8(32'h3b30ee1c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09098e),
	.w1(32'hbbd9a8a7),
	.w2(32'h3adf41f0),
	.w3(32'hbc2d9cc9),
	.w4(32'hbb092c66),
	.w5(32'h3c39d5ee),
	.w6(32'h3baa4991),
	.w7(32'hb9f082c5),
	.w8(32'h3b1a6387),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b069b10),
	.w1(32'hbacd7e2e),
	.w2(32'hbb91cbb0),
	.w3(32'h39be0fc0),
	.w4(32'hbb604731),
	.w5(32'hbb815d5c),
	.w6(32'hbbcd09f2),
	.w7(32'hbc79ad0b),
	.w8(32'hbc69cca9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba47d51),
	.w1(32'h3c750a56),
	.w2(32'h3c412c41),
	.w3(32'h3b243837),
	.w4(32'h3c1679c9),
	.w5(32'h3c092544),
	.w6(32'hbc39baa8),
	.w7(32'h3c79d07b),
	.w8(32'h3c89d76c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62966b),
	.w1(32'h3a9d694c),
	.w2(32'hbbe56a7c),
	.w3(32'h3c6e7b24),
	.w4(32'h3b66d547),
	.w5(32'h3a9f061a),
	.w6(32'h3b5db4dc),
	.w7(32'h3a696d03),
	.w8(32'hbb6b04b0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07bf33),
	.w1(32'hbb1279c7),
	.w2(32'hbbb86f7d),
	.w3(32'h3be79c62),
	.w4(32'hbbbdae6d),
	.w5(32'h3adf0af7),
	.w6(32'h3c526e20),
	.w7(32'hba165a4b),
	.w8(32'hbb02c44d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9080b),
	.w1(32'h3a1fe1ca),
	.w2(32'hbbee4447),
	.w3(32'hbb7ab979),
	.w4(32'h3b1ebc3f),
	.w5(32'hbc5930bb),
	.w6(32'hbbf314f7),
	.w7(32'h3b855348),
	.w8(32'hbbf6177f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c9de9),
	.w1(32'h3bfb12e8),
	.w2(32'hbb11deba),
	.w3(32'hbc54f292),
	.w4(32'h3a7967fa),
	.w5(32'hbbb230e2),
	.w6(32'hbb9b9198),
	.w7(32'h3a9d39f6),
	.w8(32'hbb10ef0e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a839956),
	.w1(32'hbb87f875),
	.w2(32'hbb12a7b9),
	.w3(32'hbb2cd4a9),
	.w4(32'hb9f50d61),
	.w5(32'h3a4c9e54),
	.w6(32'hba960f69),
	.w7(32'hbbb9163f),
	.w8(32'hbab31356),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5792ee),
	.w1(32'hbb5ae765),
	.w2(32'hbc4ddc30),
	.w3(32'hbc001005),
	.w4(32'hbba9d8db),
	.w5(32'hbc34f141),
	.w6(32'hbb59e32f),
	.w7(32'hbbfbe653),
	.w8(32'hbc1a6ae5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bf480),
	.w1(32'hbb8999c8),
	.w2(32'hbc55e934),
	.w3(32'hbbfce407),
	.w4(32'hbc241235),
	.w5(32'hbc4a1ba9),
	.w6(32'h3b2d3b68),
	.w7(32'hbc175391),
	.w8(32'hbc34a2bf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8018b),
	.w1(32'h3bb2741b),
	.w2(32'hbabcee24),
	.w3(32'hbc473639),
	.w4(32'h3c3041b7),
	.w5(32'hbc132182),
	.w6(32'hbad7e019),
	.w7(32'h3a97f54b),
	.w8(32'h3af9f031),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39027dc6),
	.w1(32'hbb5b1b17),
	.w2(32'h3b6a514d),
	.w3(32'h3b9538a3),
	.w4(32'h3bd0d549),
	.w5(32'h3c2f7c59),
	.w6(32'h3c04bdb4),
	.w7(32'hbb62b1e9),
	.w8(32'h3b2ee70c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af06f9a),
	.w1(32'h3b419ba1),
	.w2(32'hbbc6cfa0),
	.w3(32'h3b09eecc),
	.w4(32'h3b7923da),
	.w5(32'hbc2a244d),
	.w6(32'h3a2e4b2e),
	.w7(32'hbc0a467e),
	.w8(32'hbb6ca396),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9a8d4),
	.w1(32'h3ba9eaf8),
	.w2(32'h3ba373f3),
	.w3(32'hbabc046a),
	.w4(32'h3bc7b54d),
	.w5(32'h3b797236),
	.w6(32'h3a51c3c3),
	.w7(32'hb9f91e18),
	.w8(32'hbb00471e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af2c25),
	.w1(32'hba8c6197),
	.w2(32'hbb06e1c2),
	.w3(32'hb8526741),
	.w4(32'hbabb6bfd),
	.w5(32'hbc3c3cb3),
	.w6(32'hbb9c311a),
	.w7(32'h3b2c6bde),
	.w8(32'hbbe2a94d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27a761),
	.w1(32'hbb70fff0),
	.w2(32'h3c2226fa),
	.w3(32'hbb856074),
	.w4(32'hb9721a51),
	.w5(32'h3bdababc),
	.w6(32'hbba2add0),
	.w7(32'h3bffc78e),
	.w8(32'h3cc6f50f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c219164),
	.w1(32'hbbc90cd0),
	.w2(32'hba09ccfe),
	.w3(32'h3c3b8b87),
	.w4(32'hbb7a2e5c),
	.w5(32'hbc116f95),
	.w6(32'h3b98b69d),
	.w7(32'h3b1a2797),
	.w8(32'hbb758d07),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3f672),
	.w1(32'h3bdbc042),
	.w2(32'h3c26ad25),
	.w3(32'hb804cc71),
	.w4(32'h3bf8dbcd),
	.w5(32'h3b486283),
	.w6(32'hb9d57d04),
	.w7(32'h3c287e5b),
	.w8(32'h3c4cbedd),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3e184),
	.w1(32'h3bf79ae7),
	.w2(32'h3c000769),
	.w3(32'hbb2399e3),
	.w4(32'h3c026406),
	.w5(32'hbbb3e78d),
	.w6(32'h38a8452c),
	.w7(32'h3c3dcbbc),
	.w8(32'h3badd9c7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b299e),
	.w1(32'hbbeea2d2),
	.w2(32'h3b5a09c7),
	.w3(32'h3a574cb4),
	.w4(32'hbc0f8fd4),
	.w5(32'hbb8c5a6f),
	.w6(32'hbbe9c5f2),
	.w7(32'hbb93ca8c),
	.w8(32'hbc03581b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804e32),
	.w1(32'hbaba24d3),
	.w2(32'hbbb4ff59),
	.w3(32'hbc19903e),
	.w4(32'h3b3d99e7),
	.w5(32'hba509b20),
	.w6(32'hbb8bcfda),
	.w7(32'h3b464087),
	.w8(32'hbbf482a5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1bb95),
	.w1(32'h3ba0ad80),
	.w2(32'h3bed7ef3),
	.w3(32'hbbc97b5b),
	.w4(32'h3c6bb5e4),
	.w5(32'h3b4950e7),
	.w6(32'hbb110b5b),
	.w7(32'h3c25ebbf),
	.w8(32'h3c674c4e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b297117),
	.w1(32'h3b3b69ac),
	.w2(32'hbb6803f0),
	.w3(32'h3b5ebc64),
	.w4(32'h3bc8beeb),
	.w5(32'hbbead598),
	.w6(32'hbafbc680),
	.w7(32'hbb56dc06),
	.w8(32'hbbbc05a9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1234bb),
	.w1(32'hbb86aa21),
	.w2(32'hbbe3483e),
	.w3(32'h3b5dcca7),
	.w4(32'hbbc27e82),
	.w5(32'hbbc9b212),
	.w6(32'h3b82e000),
	.w7(32'hbc2aca4f),
	.w8(32'hba930863),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c8e10),
	.w1(32'hba99605a),
	.w2(32'h3c035ef1),
	.w3(32'h3a85d46f),
	.w4(32'hbb8e92f7),
	.w5(32'h3a4a09a9),
	.w6(32'h39e8f2db),
	.w7(32'hbbf0b0d1),
	.w8(32'h3ad53974),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a686a96),
	.w1(32'hbb97c247),
	.w2(32'h3c3dc278),
	.w3(32'h3ace6220),
	.w4(32'hbb82cbbb),
	.w5(32'hbc4ba9fb),
	.w6(32'h3c02592f),
	.w7(32'hbc15c595),
	.w8(32'hbc904b31),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ed3f7),
	.w1(32'hba92b6e2),
	.w2(32'hbc9a34e9),
	.w3(32'hbc36c487),
	.w4(32'hb9e3e30a),
	.w5(32'hbc375b37),
	.w6(32'h3b7fae1e),
	.w7(32'hbc129e09),
	.w8(32'hbca91cf0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc289e50),
	.w1(32'hbbde0fdd),
	.w2(32'hbc159140),
	.w3(32'hbc7e300a),
	.w4(32'h3a9abbad),
	.w5(32'hbbd2372a),
	.w6(32'hbc777aaf),
	.w7(32'hbb1329a9),
	.w8(32'hbb7fad6f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d4269),
	.w1(32'hbbb776ad),
	.w2(32'hbbaf876a),
	.w3(32'hbaa3cf56),
	.w4(32'hba85e612),
	.w5(32'h3c0216ca),
	.w6(32'h39a17dfc),
	.w7(32'hbc02f6d1),
	.w8(32'hbb3f4820),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1190c6),
	.w1(32'h3ac94951),
	.w2(32'h3b644840),
	.w3(32'h3b44af3f),
	.w4(32'h3c5e576d),
	.w5(32'h3c51c232),
	.w6(32'h3bce3c2f),
	.w7(32'h3c4bf7a6),
	.w8(32'h3bcb29e3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0818e),
	.w1(32'hbbc0a8a3),
	.w2(32'hba6894ec),
	.w3(32'h3b421e34),
	.w4(32'hbb78014a),
	.w5(32'h3ae5c058),
	.w6(32'hbbf85e47),
	.w7(32'h3ac72205),
	.w8(32'h3bfb1ae0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5a4ba),
	.w1(32'h3c672ea3),
	.w2(32'hbc4313af),
	.w3(32'hbafc2c87),
	.w4(32'hbc1ca6a7),
	.w5(32'hbc27fccd),
	.w6(32'hba3389bf),
	.w7(32'hbb93148a),
	.w8(32'hbc1701f3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de2827),
	.w1(32'hbbe4d5bc),
	.w2(32'h3a37def4),
	.w3(32'h3a94c8c8),
	.w4(32'h38e3a306),
	.w5(32'hbac03d45),
	.w6(32'h3b5f62d1),
	.w7(32'h3ad85708),
	.w8(32'h3a97cba2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eb2d2),
	.w1(32'hbb10bfa5),
	.w2(32'hbbd60f50),
	.w3(32'hbc0f5432),
	.w4(32'hbb7a3b03),
	.w5(32'hbc4b7fd4),
	.w6(32'hbb1eaeb8),
	.w7(32'hbb6bc7b4),
	.w8(32'hbc7c4499),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc152088),
	.w1(32'hbb1b0977),
	.w2(32'hbb09ec91),
	.w3(32'hbc63e0b1),
	.w4(32'hbbccb27e),
	.w5(32'h3a665671),
	.w6(32'hbb934924),
	.w7(32'hbafa4636),
	.w8(32'hb9bd83d2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d4b45),
	.w1(32'h3b8ffbdc),
	.w2(32'hbb8bcf96),
	.w3(32'h3aa04b61),
	.w4(32'h3bf07dce),
	.w5(32'hbb16fa22),
	.w6(32'h3b2f97a4),
	.w7(32'h3c131bbb),
	.w8(32'h3b71b3ab),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2456ae),
	.w1(32'hbb44843b),
	.w2(32'hbb856eb8),
	.w3(32'h3c4d4f0a),
	.w4(32'h3bbb89d2),
	.w5(32'h3b24426b),
	.w6(32'h3c525a7d),
	.w7(32'h3bab3468),
	.w8(32'h39d91f34),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95130b),
	.w1(32'h3aec004d),
	.w2(32'h3aa27d89),
	.w3(32'h3ac45074),
	.w4(32'h3ac66109),
	.w5(32'hbc10981d),
	.w6(32'h3bace05f),
	.w7(32'hb9b018d6),
	.w8(32'hba115a1d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4768fa),
	.w1(32'hb9110003),
	.w2(32'h3a49aee6),
	.w3(32'hbb5d7ce5),
	.w4(32'h398d66ce),
	.w5(32'hbba9d39f),
	.w6(32'hbb4cda4d),
	.w7(32'hbb4338fd),
	.w8(32'hbc6bd4eb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae005d1),
	.w1(32'h3ac523d1),
	.w2(32'hbb88c4b4),
	.w3(32'hbba6969f),
	.w4(32'h3b2a798f),
	.w5(32'h39dbf10d),
	.w6(32'hbb237247),
	.w7(32'hba21fe1a),
	.w8(32'hbbe1d5e6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c890e),
	.w1(32'hbc1cf3aa),
	.w2(32'hbb9dd0a9),
	.w3(32'hbbe0b84a),
	.w4(32'hbbe45986),
	.w5(32'hbb49d9b8),
	.w6(32'hbc3e033f),
	.w7(32'hbb831ee5),
	.w8(32'hbaeef0f2),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb080a),
	.w1(32'hb930d492),
	.w2(32'hbc0fc8a1),
	.w3(32'h3bbda8f6),
	.w4(32'hbc0dd0f6),
	.w5(32'hbc02b14d),
	.w6(32'h3b947485),
	.w7(32'hbc164bad),
	.w8(32'hbc1dcfd4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb082fcc),
	.w1(32'hba233a2d),
	.w2(32'h3a9486ad),
	.w3(32'hbaa343fd),
	.w4(32'h39fda74b),
	.w5(32'hba2732ca),
	.w6(32'hbb959f8a),
	.w7(32'hbc07589f),
	.w8(32'hbb54a415),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e947d),
	.w1(32'hbb9b518b),
	.w2(32'h3af5f693),
	.w3(32'hbb974dd8),
	.w4(32'hbbe90b3d),
	.w5(32'h3bae4be8),
	.w6(32'hbbed530a),
	.w7(32'hbbfa29ec),
	.w8(32'h3ad4000f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb643701),
	.w1(32'hbbbce12e),
	.w2(32'hbb5d9355),
	.w3(32'h3c1196f4),
	.w4(32'hbabdf49a),
	.w5(32'h3a3f3f64),
	.w6(32'hbacf158f),
	.w7(32'hbb1812df),
	.w8(32'h3b86467d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbddbb3),
	.w1(32'h3b8351ee),
	.w2(32'hbbfaf4aa),
	.w3(32'hbc125102),
	.w4(32'hbbaa0808),
	.w5(32'h3b986337),
	.w6(32'hbc564baa),
	.w7(32'h3aa5a240),
	.w8(32'h3b9f954d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5de4ac),
	.w1(32'h3c1edc31),
	.w2(32'hbc18c1f0),
	.w3(32'hbb88c127),
	.w4(32'h3b854803),
	.w5(32'hbc25031b),
	.w6(32'hbbaee262),
	.w7(32'hbb33e12f),
	.w8(32'hbc17feeb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9293bf7),
	.w1(32'h3b85c5dd),
	.w2(32'h3c7163ab),
	.w3(32'h3c018519),
	.w4(32'h3c87f40f),
	.w5(32'h3caefa5e),
	.w6(32'h3c7682dd),
	.w7(32'h3c03c5b9),
	.w8(32'h3c9f17fe),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a29d8),
	.w1(32'h3c024a0b),
	.w2(32'h3c0d639a),
	.w3(32'h3bbb7f7d),
	.w4(32'h3c016eb1),
	.w5(32'h3a1bdf73),
	.w6(32'h389402ef),
	.w7(32'h3c15b1cb),
	.w8(32'h3be3d6ab),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41d584),
	.w1(32'hbbdae1ab),
	.w2(32'hbbde63c9),
	.w3(32'hbbd4652b),
	.w4(32'hbc7722e1),
	.w5(32'hbc5f223e),
	.w6(32'hbc668b67),
	.w7(32'hbbd04afc),
	.w8(32'hbab0fdcf),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeeeb09),
	.w1(32'h3b7af7cd),
	.w2(32'hbb926edd),
	.w3(32'hbbad7d5b),
	.w4(32'hbc1a13d0),
	.w5(32'hbc1045f9),
	.w6(32'hbc37c1ed),
	.w7(32'hbb1e5b4f),
	.w8(32'hbc0ad921),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b67d),
	.w1(32'hbab6e2d9),
	.w2(32'h3afd3a97),
	.w3(32'hbb723c50),
	.w4(32'h3b12f2ef),
	.w5(32'hbaf668c1),
	.w6(32'hbab145c4),
	.w7(32'hbc0aa8a6),
	.w8(32'hbbf3a80f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a19350),
	.w1(32'hb7a37a81),
	.w2(32'hbb8fed38),
	.w3(32'hb97713a7),
	.w4(32'hbb78dea0),
	.w5(32'hbbc6b586),
	.w6(32'hbb1b6b4b),
	.w7(32'hbbb6dc6f),
	.w8(32'hbc3e318b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bcd57),
	.w1(32'h3b2e99e6),
	.w2(32'h3b8c2716),
	.w3(32'hbbda22da),
	.w4(32'hbb313fcf),
	.w5(32'hb9bbd17e),
	.w6(32'hbbef5465),
	.w7(32'hbaa5ea31),
	.w8(32'hbc22cb7c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e70fc2),
	.w1(32'h3acfded5),
	.w2(32'hbb61135c),
	.w3(32'hbc3d97bc),
	.w4(32'h3b21588f),
	.w5(32'hbc2ff8c5),
	.w6(32'hbbf298d6),
	.w7(32'h3b489d3a),
	.w8(32'hbba4cdc8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb924777),
	.w1(32'hbc5b250c),
	.w2(32'hbc0bf88f),
	.w3(32'hb82d3fe7),
	.w4(32'hbbb52911),
	.w5(32'hbc10ef82),
	.w6(32'hbbb6b6bc),
	.w7(32'hbc2dd160),
	.w8(32'hbc0fd1fc),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0f77),
	.w1(32'hbb139ce9),
	.w2(32'hbbadc470),
	.w3(32'hbb10635f),
	.w4(32'h3bd2435d),
	.w5(32'hbb2b5f91),
	.w6(32'hbb478c7e),
	.w7(32'h3bb98586),
	.w8(32'h3c40fdc6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e8b83),
	.w1(32'hbb0f88b9),
	.w2(32'hbafea0dd),
	.w3(32'h3bef5c00),
	.w4(32'hbb913a33),
	.w5(32'hbba75a37),
	.w6(32'h3c3608be),
	.w7(32'hbbe0ee59),
	.w8(32'hbb166954),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb9742),
	.w1(32'h3aa32f57),
	.w2(32'h3b359983),
	.w3(32'h3b0fe6d0),
	.w4(32'h3a9bb95c),
	.w5(32'hbaef4b8e),
	.w6(32'hba4c23d4),
	.w7(32'h3b8a9a3a),
	.w8(32'h3b515f14),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacfee5),
	.w1(32'h392e6337),
	.w2(32'hba01ec61),
	.w3(32'hbb88c815),
	.w4(32'h3c6a6199),
	.w5(32'hbc2b2ef0),
	.w6(32'h3a9375c9),
	.w7(32'h3bb6dd08),
	.w8(32'hbbbbda17),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7861e),
	.w1(32'h3a24afdb),
	.w2(32'hbbbbf802),
	.w3(32'hbae1e0b2),
	.w4(32'hbac2ad08),
	.w5(32'h3aad50b7),
	.w6(32'hbbc747b0),
	.w7(32'hbc18b48b),
	.w8(32'h3a23d5d7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd06d),
	.w1(32'hbb534cc2),
	.w2(32'h3b129930),
	.w3(32'hbb83be52),
	.w4(32'hbb5f9baf),
	.w5(32'h3bc722ea),
	.w6(32'hbbf4f467),
	.w7(32'hba83afaa),
	.w8(32'h3b4af27d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47db2b),
	.w1(32'hbc0e9495),
	.w2(32'hbc49c07d),
	.w3(32'hbc5f9a16),
	.w4(32'hbc8cdc3c),
	.w5(32'hbcb5e906),
	.w6(32'hb9e99004),
	.w7(32'hbbc8f7a9),
	.w8(32'hbb949bb0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f231f),
	.w1(32'h3c10a17f),
	.w2(32'hb7f0e3ca),
	.w3(32'hbc85ab66),
	.w4(32'h3b1ec2da),
	.w5(32'hbc48dfec),
	.w6(32'hbbba0227),
	.w7(32'hbbf0bef5),
	.w8(32'hb9b8fce3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b34a8c),
	.w1(32'hbb829c19),
	.w2(32'hbbb28684),
	.w3(32'hbc0dfe63),
	.w4(32'h3b67aba7),
	.w5(32'hbb04b2e4),
	.w6(32'h3be35d8a),
	.w7(32'h3a1135b3),
	.w8(32'h3a85fccc),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b241678),
	.w1(32'h3b0c2ffc),
	.w2(32'hbb2db5e4),
	.w3(32'h3c042e38),
	.w4(32'h3b98df7b),
	.w5(32'h3acb08d1),
	.w6(32'h3bdea69b),
	.w7(32'hbab6dd03),
	.w8(32'hbc37fce3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47b7a6),
	.w1(32'h3b94f60e),
	.w2(32'h3c07e0fa),
	.w3(32'hbc05ab1e),
	.w4(32'h3c62d2ef),
	.w5(32'hb9ec35df),
	.w6(32'hbbfb3817),
	.w7(32'h3c528c32),
	.w8(32'h3c74471d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4b007),
	.w1(32'hbb83ba6b),
	.w2(32'hbacdda7b),
	.w3(32'h3a277675),
	.w4(32'h3b54ecea),
	.w5(32'hbb90b72a),
	.w6(32'hbae2aa17),
	.w7(32'h3b4d96ae),
	.w8(32'h3b91cc38),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b0b14),
	.w1(32'hbb5742dc),
	.w2(32'hbb9c24e1),
	.w3(32'h3c877d21),
	.w4(32'hbabaacea),
	.w5(32'h3ba3cbb3),
	.w6(32'h3cc7325c),
	.w7(32'hbbc68376),
	.w8(32'hbbcfee22),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813a3f),
	.w1(32'hbbbd082d),
	.w2(32'hbc28a63f),
	.w3(32'hb9c175e6),
	.w4(32'h3a99efdb),
	.w5(32'h3b64698c),
	.w6(32'hbc57e7c5),
	.w7(32'h3a862aa1),
	.w8(32'h39943dfc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbd014),
	.w1(32'hbbab488c),
	.w2(32'hbc31fcb9),
	.w3(32'hbb1d4531),
	.w4(32'h39676687),
	.w5(32'hbc324a00),
	.w6(32'h3ba85bf3),
	.w7(32'h3be4b440),
	.w8(32'hbbdd73c1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74e7fd),
	.w1(32'hbb644536),
	.w2(32'hbc90a797),
	.w3(32'hbc2073bd),
	.w4(32'hbc972c1e),
	.w5(32'hbc483663),
	.w6(32'hbc2b9c20),
	.w7(32'hbc17d1eb),
	.w8(32'hbc8bf899),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad11945),
	.w1(32'hbb23f143),
	.w2(32'hbbb7b2d1),
	.w3(32'h3af4e0b7),
	.w4(32'h39f9ff11),
	.w5(32'hbc65ae8a),
	.w6(32'h3b995322),
	.w7(32'h3bb025eb),
	.w8(32'hbaf6915b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba491a80),
	.w1(32'h3b1916ac),
	.w2(32'hbba79cbf),
	.w3(32'h3b0c792a),
	.w4(32'h39ef517d),
	.w5(32'hbb89d02f),
	.w6(32'h3a80cefb),
	.w7(32'h3b010a84),
	.w8(32'h3aee2cd2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f71b6),
	.w1(32'h3b466cd9),
	.w2(32'h3b32411d),
	.w3(32'h3a5ce1a1),
	.w4(32'h3b955780),
	.w5(32'hbbf1ec1e),
	.w6(32'hba7be893),
	.w7(32'hbc02acf6),
	.w8(32'h3ba8dd04),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25104f),
	.w1(32'h3a7b217c),
	.w2(32'hbb720770),
	.w3(32'hb980642a),
	.w4(32'hbad1b9d1),
	.w5(32'h39792e84),
	.w6(32'h3b0ad226),
	.w7(32'hbb5d19a6),
	.w8(32'h3ba09e45),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3baf3c),
	.w1(32'hbb556177),
	.w2(32'hb9ceba84),
	.w3(32'h3b60742b),
	.w4(32'hba948712),
	.w5(32'h3c68d5e6),
	.w6(32'h3c0204c1),
	.w7(32'h3b48d7a9),
	.w8(32'h3b9af4a8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a5ebc),
	.w1(32'hbac3f116),
	.w2(32'hbb489709),
	.w3(32'h3a792047),
	.w4(32'hbb0e540e),
	.w5(32'hbc5854c8),
	.w6(32'hbb3a81b8),
	.w7(32'h3b84a9ac),
	.w8(32'hbb4a8263),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bcf3e),
	.w1(32'h3ab21eb5),
	.w2(32'hbab6e48c),
	.w3(32'hbb985b4d),
	.w4(32'h3ba01990),
	.w5(32'h3bb8b345),
	.w6(32'hbb6e2a2e),
	.w7(32'h3ba9ec88),
	.w8(32'h3c1bf721),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39612534),
	.w1(32'h3b84109a),
	.w2(32'h3a99b9a8),
	.w3(32'h3ab0fe01),
	.w4(32'h38779e3c),
	.w5(32'h3c2f1616),
	.w6(32'h3b051ee2),
	.w7(32'hbb89bb22),
	.w8(32'hbc0178ce),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966800),
	.w1(32'hb8cb139b),
	.w2(32'hbb85bb65),
	.w3(32'h3b48e2b8),
	.w4(32'hba2b262f),
	.w5(32'h3bdb4fd3),
	.w6(32'hba48d91d),
	.w7(32'hbaf031f6),
	.w8(32'hbc290c58),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9efde),
	.w1(32'hbb8593a2),
	.w2(32'hbbc6d35a),
	.w3(32'hbbc7db43),
	.w4(32'hbb4925a9),
	.w5(32'hbb3ed33a),
	.w6(32'hb8841d01),
	.w7(32'hbaa3cc56),
	.w8(32'h39c948a2),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad0205),
	.w1(32'hbb2a3278),
	.w2(32'hb8c06fcb),
	.w3(32'hbb942014),
	.w4(32'hbc14cce8),
	.w5(32'hbbf72b78),
	.w6(32'hbb0e0751),
	.w7(32'h3a9c7b15),
	.w8(32'hbc013731),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1cd5f),
	.w1(32'hba90bf1c),
	.w2(32'h3ba26f7b),
	.w3(32'hbbca5d6c),
	.w4(32'hbb07f861),
	.w5(32'h3b946cae),
	.w6(32'h3aad5313),
	.w7(32'hbae8e16d),
	.w8(32'h3b90254c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12ce03),
	.w1(32'h3ba03c30),
	.w2(32'h3abe8ba9),
	.w3(32'h3962b2cd),
	.w4(32'h3b57c0f3),
	.w5(32'h3a1d3682),
	.w6(32'h3ace1af4),
	.w7(32'h3a339308),
	.w8(32'h3b2ed600),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a17b7),
	.w1(32'hbaad87ae),
	.w2(32'hbb37776a),
	.w3(32'hb9059ef0),
	.w4(32'hbbca7e7c),
	.w5(32'hbc8b72a0),
	.w6(32'h3ae1c840),
	.w7(32'h3ae6606b),
	.w8(32'h3b8191b0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc710),
	.w1(32'h3c3930a2),
	.w2(32'h3bbbbdc1),
	.w3(32'h39ccc1ac),
	.w4(32'h3bdac578),
	.w5(32'h3b1fb6e8),
	.w6(32'h3c2fa92a),
	.w7(32'hbb7f4f70),
	.w8(32'hbb4d8d16),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb754946),
	.w1(32'hba98fbe4),
	.w2(32'hba0acb57),
	.w3(32'h3b2e5fef),
	.w4(32'hbb127bdf),
	.w5(32'h3a9f839b),
	.w6(32'h3beac8a8),
	.w7(32'hbbb022c6),
	.w8(32'hba562c2e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a345fe),
	.w1(32'hbb4ed7f7),
	.w2(32'h3bd3eb57),
	.w3(32'h3b163bae),
	.w4(32'h3bd8b9c9),
	.w5(32'h3b299262),
	.w6(32'h3b869ae9),
	.w7(32'h3c29298d),
	.w8(32'hba861fd5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b989110),
	.w1(32'h3854581a),
	.w2(32'hbb81aef5),
	.w3(32'hbad297fa),
	.w4(32'hbba3775b),
	.w5(32'hbbf90e79),
	.w6(32'h3c1e0f21),
	.w7(32'hbb8dd559),
	.w8(32'hbc7b4bda),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac818cb),
	.w1(32'hbb6487e3),
	.w2(32'hbb561486),
	.w3(32'hbc52ab84),
	.w4(32'hbc68bc38),
	.w5(32'hbbc4d91b),
	.w6(32'hbc33ab74),
	.w7(32'h3a86ad9c),
	.w8(32'hbc04f8d7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc169684),
	.w1(32'h3b078764),
	.w2(32'hbaafea96),
	.w3(32'hbc42aa83),
	.w4(32'hbb59ac9b),
	.w5(32'h3bc1992f),
	.w6(32'hbb92f26d),
	.w7(32'hbc162c52),
	.w8(32'hbbe2cf97),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee1fa3),
	.w1(32'h3c6d3fb6),
	.w2(32'hbb1060ab),
	.w3(32'hba9a390d),
	.w4(32'h3bdeb5eb),
	.w5(32'hbb8330ad),
	.w6(32'hba439ee8),
	.w7(32'h3ba0eeba),
	.w8(32'hbbc3e1d7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2a674),
	.w1(32'h39b2d4ba),
	.w2(32'hbb15d066),
	.w3(32'h3a217944),
	.w4(32'hbb584b8a),
	.w5(32'hbc0688cf),
	.w6(32'h3bb86209),
	.w7(32'hbc2c2ece),
	.w8(32'hbc4f0d35),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac8b5e),
	.w1(32'hba96169c),
	.w2(32'h3a8b86f3),
	.w3(32'h3aecc98e),
	.w4(32'h3bce32a2),
	.w5(32'h3c003253),
	.w6(32'h3b00d77d),
	.w7(32'h3bdae0bd),
	.w8(32'hbc4ce5b8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924130e),
	.w1(32'hbb2485ab),
	.w2(32'h3b7d28f5),
	.w3(32'hba9e87e5),
	.w4(32'hbc1e20a4),
	.w5(32'hbc8d1f8b),
	.w6(32'h3ba2609b),
	.w7(32'hbb75a02c),
	.w8(32'h3be04578),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ed78a),
	.w1(32'hbb1903c3),
	.w2(32'h3baae5c5),
	.w3(32'hbb82913f),
	.w4(32'h38690afd),
	.w5(32'h3c52c9f9),
	.w6(32'h3b456a4b),
	.w7(32'h3b24b9cf),
	.w8(32'h3bd2f21e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a636da7),
	.w1(32'h3a590433),
	.w2(32'h3a7e3881),
	.w3(32'h3829009c),
	.w4(32'hbc4529e0),
	.w5(32'hbbc2e7e2),
	.w6(32'h3b18aa70),
	.w7(32'h3ab1c3a9),
	.w8(32'hbc2cfb78),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfdde),
	.w1(32'hbb31e99e),
	.w2(32'hbc2c1477),
	.w3(32'hbbc7a9da),
	.w4(32'hbb92c573),
	.w5(32'hbbfdda0e),
	.w6(32'hbae13240),
	.w7(32'hbbca2b3d),
	.w8(32'hbc81ae4b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0d2b),
	.w1(32'hbadc7896),
	.w2(32'hbbe61a59),
	.w3(32'hbc32f2ea),
	.w4(32'hbc27a34e),
	.w5(32'hbb103c83),
	.w6(32'hbc551597),
	.w7(32'hb6a67c60),
	.w8(32'h3af2aefb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70e942),
	.w1(32'h3b643229),
	.w2(32'h3acacae2),
	.w3(32'hbbc80917),
	.w4(32'hbabcd6ba),
	.w5(32'h3afc866d),
	.w6(32'hbb89c29b),
	.w7(32'hbb024632),
	.w8(32'h3bd70f7c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beea015),
	.w1(32'hbbe6a3eb),
	.w2(32'hbc379d2d),
	.w3(32'h3b46c36b),
	.w4(32'h3a88ae55),
	.w5(32'hbb81a991),
	.w6(32'h3c001b19),
	.w7(32'hb9b95e2b),
	.w8(32'h3a885d2b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b3e79),
	.w1(32'hbb916248),
	.w2(32'hbae8e049),
	.w3(32'hbb37d518),
	.w4(32'hbbe0b754),
	.w5(32'hbc7fce59),
	.w6(32'h3b91c954),
	.w7(32'h3b14fcec),
	.w8(32'h3b9c0c4c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9193f3),
	.w1(32'hbac28f37),
	.w2(32'hbb6bd4f4),
	.w3(32'hbb0d3e9c),
	.w4(32'hbc1d0ebe),
	.w5(32'hbb993bc4),
	.w6(32'hbbb8556e),
	.w7(32'hbb4e38d2),
	.w8(32'hbc00884c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ed700),
	.w1(32'hbbce8b53),
	.w2(32'hbb720d65),
	.w3(32'hbc433fa1),
	.w4(32'h3a19e274),
	.w5(32'hbbd8f150),
	.w6(32'hbbf2ebd3),
	.w7(32'hbc0f5a4a),
	.w8(32'h3a5bda11),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b3ec5),
	.w1(32'h3aa5f219),
	.w2(32'hbc2b2a83),
	.w3(32'hbb93e6ff),
	.w4(32'h3b0fe51d),
	.w5(32'hbb3988d6),
	.w6(32'h3a6f147d),
	.w7(32'h3afec04b),
	.w8(32'hbc575100),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec0bb6),
	.w1(32'hbb88d78c),
	.w2(32'hbb2c3915),
	.w3(32'hbbd83b9a),
	.w4(32'hbb282da6),
	.w5(32'hbaa4ce41),
	.w6(32'hbb4e409d),
	.w7(32'hbbb070b8),
	.w8(32'hbbb1762f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba297a3),
	.w1(32'hbc0bad99),
	.w2(32'hbc2e4e51),
	.w3(32'h398a6692),
	.w4(32'hbc3929e1),
	.w5(32'hbca2c15f),
	.w6(32'h3b26076d),
	.w7(32'hbc35051f),
	.w8(32'hbc0c1079),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc558d9e),
	.w1(32'hbbedf8d3),
	.w2(32'hbb865dd7),
	.w3(32'hbbcab428),
	.w4(32'hbb9d11df),
	.w5(32'hbb9e819a),
	.w6(32'hbc27f4d1),
	.w7(32'hbb9b85dc),
	.w8(32'hbbe25dc3),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4d085),
	.w1(32'h3bb6bbc7),
	.w2(32'hbc043037),
	.w3(32'hbab3ec43),
	.w4(32'h3b9da265),
	.w5(32'hbadb8e95),
	.w6(32'hbb2fffdf),
	.w7(32'h3bbe4d4f),
	.w8(32'h3ba3ba61),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01dd0c),
	.w1(32'h3abd08cf),
	.w2(32'hb8899df3),
	.w3(32'hba69beef),
	.w4(32'h3b953fad),
	.w5(32'hbc11d999),
	.w6(32'h3c12b784),
	.w7(32'hbb63ad7f),
	.w8(32'h3ba8241f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3504c0),
	.w1(32'hbbcb7a99),
	.w2(32'hbb396bdb),
	.w3(32'h3b04e7a8),
	.w4(32'hba01a2a2),
	.w5(32'hbc9ab85d),
	.w6(32'hbba9d6f3),
	.w7(32'h3b75c8ef),
	.w8(32'h3c9b9e29),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a268a90),
	.w1(32'hbbbe77c9),
	.w2(32'hbc0f45b2),
	.w3(32'h3acd435e),
	.w4(32'hbbc9f9cd),
	.w5(32'hbc4f04fe),
	.w6(32'h3b6d9ece),
	.w7(32'hbc165162),
	.w8(32'hbbc0dcc1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadff45),
	.w1(32'h3b50d23c),
	.w2(32'h3b1b9581),
	.w3(32'hbc507a20),
	.w4(32'h3ba2ef42),
	.w5(32'h3b3f80f0),
	.w6(32'hbc6b17fe),
	.w7(32'h39fea23f),
	.w8(32'hbaa5f33c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d9bcf),
	.w1(32'hbb1dff94),
	.w2(32'hbbb3b87b),
	.w3(32'h3bb7b01d),
	.w4(32'hbb41afcd),
	.w5(32'hbab772af),
	.w6(32'h3b155ef3),
	.w7(32'hbc1e4ce2),
	.w8(32'hbc046ec9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3409),
	.w1(32'hbc1e9496),
	.w2(32'hbbe1621f),
	.w3(32'hbbba6ac7),
	.w4(32'hbb4b8389),
	.w5(32'h3b9ee2b7),
	.w6(32'hbbcbb3b3),
	.w7(32'h3bab0ddf),
	.w8(32'hbb884dfe),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae102cd),
	.w1(32'h3932615b),
	.w2(32'h3b061709),
	.w3(32'hbb877b46),
	.w4(32'hbbe42102),
	.w5(32'hba08cdf9),
	.w6(32'hbba1c34f),
	.w7(32'hbc0942d8),
	.w8(32'h3af1eab4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2d76a),
	.w1(32'h3b1905a6),
	.w2(32'h3c3ac6ad),
	.w3(32'hbb34f23d),
	.w4(32'h39ed11f7),
	.w5(32'h3c4f2f7a),
	.w6(32'h38923d1c),
	.w7(32'h3c51e52c),
	.w8(32'h3c4062ee),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c001317),
	.w1(32'hbb3259ee),
	.w2(32'h3b024b02),
	.w3(32'h3c37d32a),
	.w4(32'hbbaa1617),
	.w5(32'h3a53c92e),
	.w6(32'h3c00e816),
	.w7(32'hbbaea031),
	.w8(32'hbb5f9be5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9942c3c),
	.w1(32'hb97bca7b),
	.w2(32'h3a203f4f),
	.w3(32'h3b9fe47e),
	.w4(32'h3b33be1c),
	.w5(32'h3c13fcc4),
	.w6(32'h3a6ef56c),
	.w7(32'hbb11cae6),
	.w8(32'hbb7cfdb3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd00a5),
	.w1(32'hbb8ccda0),
	.w2(32'h3aa56142),
	.w3(32'h3b7bfc04),
	.w4(32'hba561048),
	.w5(32'h3b6eaf02),
	.w6(32'h3b49f742),
	.w7(32'hbb72dd17),
	.w8(32'h3c0b94c1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c0ebae),
	.w1(32'h3b9dee53),
	.w2(32'h3c1514da),
	.w3(32'h3b62e0d1),
	.w4(32'h3aa2c753),
	.w5(32'h3c87f394),
	.w6(32'hb7ed2c1a),
	.w7(32'h3b24ec99),
	.w8(32'h3c13efd1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdd5b8),
	.w1(32'hbb67a84f),
	.w2(32'hbbe558c9),
	.w3(32'h3b639246),
	.w4(32'hbb904be7),
	.w5(32'hbc3f33c9),
	.w6(32'h3b805634),
	.w7(32'hbbc416f5),
	.w8(32'hbbcff2b0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc170ca4),
	.w1(32'h3b686df2),
	.w2(32'hb9e97bae),
	.w3(32'hbc039edf),
	.w4(32'hbb18f57a),
	.w5(32'h3aea5d8e),
	.w6(32'hbbf9d3fe),
	.w7(32'hbbca49e9),
	.w8(32'hbbd557a8),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1cd2),
	.w1(32'hbc2da48d),
	.w2(32'hba70acb2),
	.w3(32'hbc01ad80),
	.w4(32'h3adebfef),
	.w5(32'hbc04ee7c),
	.w6(32'hbb64dbc7),
	.w7(32'h3c2902b1),
	.w8(32'hb9cd476a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bb04b),
	.w1(32'hbb1c773e),
	.w2(32'hbbd143df),
	.w3(32'hbb8f81c5),
	.w4(32'hbc0bafa4),
	.w5(32'hbb469bad),
	.w6(32'h3bc50f45),
	.w7(32'hbaf72201),
	.w8(32'hbbdf447f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08d1c),
	.w1(32'hbc3a66ee),
	.w2(32'hbba909ea),
	.w3(32'hbb424fa3),
	.w4(32'hbb8b454b),
	.w5(32'h3a8dd7a1),
	.w6(32'hbac18228),
	.w7(32'h3b85f844),
	.w8(32'h3b37b8b3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73b0c5),
	.w1(32'h3a22f2f4),
	.w2(32'h3affd1b8),
	.w3(32'hbbba15a2),
	.w4(32'h3b8afcb6),
	.w5(32'hbbb175df),
	.w6(32'hbbd62292),
	.w7(32'hbc2f0426),
	.w8(32'h3b5b5712),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf35840),
	.w1(32'hbbdd0dbe),
	.w2(32'hbbb9f61b),
	.w3(32'hb9abc27f),
	.w4(32'hbb2a7167),
	.w5(32'hbc505477),
	.w6(32'hbc2fa916),
	.w7(32'hbc50684f),
	.w8(32'hbc0f747d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8257d5),
	.w1(32'h3bcd06c3),
	.w2(32'hb9931386),
	.w3(32'hbb134aac),
	.w4(32'h3b6b2410),
	.w5(32'h3ba9a2c1),
	.w6(32'hbc0a56e4),
	.w7(32'h3b9428c1),
	.w8(32'hbb4c3948),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9687656),
	.w1(32'hbaf3a275),
	.w2(32'h3a81f7cd),
	.w3(32'hbb0ef1ab),
	.w4(32'hbb033c93),
	.w5(32'hbbfd7c52),
	.w6(32'hbbdd79ba),
	.w7(32'hbb946e87),
	.w8(32'hbbaac7c2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule