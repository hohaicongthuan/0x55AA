module layer_8_featuremap_136(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc53d9a),
	.w1(32'hbbece4e0),
	.w2(32'hbb084bc3),
	.w3(32'hbb256f7e),
	.w4(32'hbc98a478),
	.w5(32'hba59d471),
	.w6(32'hba8b4a3e),
	.w7(32'hbcaac91b),
	.w8(32'h3cc98e0d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17c06f),
	.w1(32'hbb00cca3),
	.w2(32'hbbf1efca),
	.w3(32'h3ca1af08),
	.w4(32'h3ca237fa),
	.w5(32'h3b68410a),
	.w6(32'h3ce082cf),
	.w7(32'h3c10af37),
	.w8(32'h3c2529e7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53832d),
	.w1(32'h3ba3398d),
	.w2(32'h3cee308a),
	.w3(32'h3c20b960),
	.w4(32'h3c294d90),
	.w5(32'h3cb43d24),
	.w6(32'h3c35ad2b),
	.w7(32'h3baf8859),
	.w8(32'h3d1888a7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f9de6),
	.w1(32'hbcc862b7),
	.w2(32'hbc2b7ee1),
	.w3(32'hbb653067),
	.w4(32'h3aded88b),
	.w5(32'h3c8016b6),
	.w6(32'hbc788f9d),
	.w7(32'hbb304792),
	.w8(32'h3c09cca5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc081121),
	.w1(32'h3a2a67c8),
	.w2(32'hbc65b6ee),
	.w3(32'hbb155c44),
	.w4(32'h3a87ccb8),
	.w5(32'h3c445963),
	.w6(32'hbbb89a32),
	.w7(32'hbb970269),
	.w8(32'hbc8bd906),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc375641),
	.w1(32'hbb991a29),
	.w2(32'hbc084cbb),
	.w3(32'hbbd233a3),
	.w4(32'h3bf23c47),
	.w5(32'hbb955e7b),
	.w6(32'hbba8e426),
	.w7(32'h3ce41a57),
	.w8(32'hbc5fc7e2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ae4bd),
	.w1(32'h3b5722b3),
	.w2(32'hbc240d6f),
	.w3(32'hbc9f4302),
	.w4(32'hbb13ee30),
	.w5(32'h3bd2bc32),
	.w6(32'hbbc5782d),
	.w7(32'h3c8bb47d),
	.w8(32'hb8d407d3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba45609),
	.w1(32'hbb8d39a6),
	.w2(32'h3bc39bb2),
	.w3(32'hbb420445),
	.w4(32'h3ce84939),
	.w5(32'h3c86a63b),
	.w6(32'h3ca937f0),
	.w7(32'h3d436efd),
	.w8(32'hbca077ca),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72caf0),
	.w1(32'hb98d6e6f),
	.w2(32'hbc114495),
	.w3(32'hbc63fdf3),
	.w4(32'h39017adc),
	.w5(32'h3c5953d6),
	.w6(32'h3b7d46ff),
	.w7(32'hbbb4d48d),
	.w8(32'h3bb535f2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbae0d),
	.w1(32'hbc36d168),
	.w2(32'hbab5fcf9),
	.w3(32'h3c20ca7d),
	.w4(32'h3cf2de28),
	.w5(32'h3b76169c),
	.w6(32'hbaab6677),
	.w7(32'h3c727b04),
	.w8(32'hbc8b0de0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e3c77),
	.w1(32'hbab7e734),
	.w2(32'hbbfa6887),
	.w3(32'hbc84ad99),
	.w4(32'h3b4ed683),
	.w5(32'h3cd100ed),
	.w6(32'hbc8f8c70),
	.w7(32'hbc4d91a1),
	.w8(32'h3ba8ab84),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89fd14),
	.w1(32'hbc9f152d),
	.w2(32'hbba62d27),
	.w3(32'hbc1d4d6c),
	.w4(32'h3cb5cc0a),
	.w5(32'h3c667357),
	.w6(32'hbcb394ee),
	.w7(32'h3d49594d),
	.w8(32'hbb836906),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a626b),
	.w1(32'h3b94f05b),
	.w2(32'h3bcda575),
	.w3(32'h3c16d3d6),
	.w4(32'h3a4e03c7),
	.w5(32'h3c556083),
	.w6(32'h3cd24435),
	.w7(32'hbaafde61),
	.w8(32'hbb06a66b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad340d4),
	.w1(32'h3a49cdb4),
	.w2(32'hbae80217),
	.w3(32'h3bee91bf),
	.w4(32'h397dc5b6),
	.w5(32'hb9947915),
	.w6(32'h3bc156f3),
	.w7(32'hba2a9e69),
	.w8(32'h3b405a19),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991922f),
	.w1(32'h3be09451),
	.w2(32'h3b82943a),
	.w3(32'h3b827ab2),
	.w4(32'h3aa7b970),
	.w5(32'h3b376ce6),
	.w6(32'h3bb85507),
	.w7(32'h3b243baa),
	.w8(32'h3b72571a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ce76),
	.w1(32'h3c20b81a),
	.w2(32'h3b42656c),
	.w3(32'h3adf0fd9),
	.w4(32'h3c1f8afe),
	.w5(32'h3c0eb870),
	.w6(32'h3c091405),
	.w7(32'hbbb66431),
	.w8(32'hbaba2322),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5f59c),
	.w1(32'h3b1541fc),
	.w2(32'h3c1da629),
	.w3(32'hba2dda49),
	.w4(32'h3b493944),
	.w5(32'h3c2a32eb),
	.w6(32'hbb2a420f),
	.w7(32'hbbd5854d),
	.w8(32'hbc89a678),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc242fb3),
	.w1(32'hbbab3517),
	.w2(32'h3b74836c),
	.w3(32'hbbc13de4),
	.w4(32'hbc428776),
	.w5(32'hbc80815c),
	.w6(32'hbb468ce9),
	.w7(32'h3c296af7),
	.w8(32'hba16ffac),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5adef),
	.w1(32'hbc80ffe5),
	.w2(32'hbc2caa86),
	.w3(32'hbc861138),
	.w4(32'hbc298c3c),
	.w5(32'hbc620e97),
	.w6(32'h3c11ee08),
	.w7(32'hbc7765f0),
	.w8(32'hbce4a3c5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f9a94),
	.w1(32'h39cd380c),
	.w2(32'hbc8209c1),
	.w3(32'h3b401557),
	.w4(32'h3bf94b46),
	.w5(32'hbc75e28b),
	.w6(32'hbc488200),
	.w7(32'h3bc5071d),
	.w8(32'hbb5d6c0f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc378c08),
	.w1(32'h3bb74cdd),
	.w2(32'h3cb8f109),
	.w3(32'hbc60cf93),
	.w4(32'hba1fa9ca),
	.w5(32'h3c36db91),
	.w6(32'hbb55cf5f),
	.w7(32'hbccc0893),
	.w8(32'hbd3aa7af),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7af54c),
	.w1(32'h3c562455),
	.w2(32'h3b743f3d),
	.w3(32'h3c9546e2),
	.w4(32'h3ae231bc),
	.w5(32'h3c74507d),
	.w6(32'hbc4bfbb8),
	.w7(32'hbbed9770),
	.w8(32'h3c8e4ccb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48a27f),
	.w1(32'hbc1d0238),
	.w2(32'h3cc02f81),
	.w3(32'h3bdd1378),
	.w4(32'h3c630985),
	.w5(32'h3c765a6b),
	.w6(32'h3c6031e0),
	.w7(32'h3cc03cef),
	.w8(32'h3cc6c5ce),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8227c2),
	.w1(32'h3bcc29bb),
	.w2(32'h3b461956),
	.w3(32'hb7f8db1d),
	.w4(32'h3bf2256c),
	.w5(32'h3b3442c8),
	.w6(32'h3c18ebc3),
	.w7(32'h3b951e60),
	.w8(32'h3c35a7de),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be04d56),
	.w1(32'h3c0723d3),
	.w2(32'h3bab35c1),
	.w3(32'h3a4bfc81),
	.w4(32'h3b5790e4),
	.w5(32'hbac092a7),
	.w6(32'h3bd2d623),
	.w7(32'h3b8f3ec2),
	.w8(32'hbb78740d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc8eef),
	.w1(32'hb85bd421),
	.w2(32'hbb04f7b1),
	.w3(32'hbbf97b41),
	.w4(32'h3bfc9878),
	.w5(32'h3cb2f4db),
	.w6(32'hbbbd4cce),
	.w7(32'hbbfd2ee5),
	.w8(32'h3cb0b754),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5de3f),
	.w1(32'hbb927058),
	.w2(32'hbaf744f4),
	.w3(32'hbb0f8545),
	.w4(32'hbc4154f0),
	.w5(32'hbcb162bc),
	.w6(32'hbbb3d5cb),
	.w7(32'h3bc00abc),
	.w8(32'hba9fecab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7d0641),
	.w1(32'h3c96d2df),
	.w2(32'hbd608514),
	.w3(32'h3aed729a),
	.w4(32'h3c944b25),
	.w5(32'hbc509ebb),
	.w6(32'hbd31c592),
	.w7(32'h3bc9636e),
	.w8(32'h3d8631e0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39870e45),
	.w1(32'h3b50ff31),
	.w2(32'hbc89feb4),
	.w3(32'hbd193931),
	.w4(32'hbb01b888),
	.w5(32'hbc4362c0),
	.w6(32'h3c6918f4),
	.w7(32'hbb829902),
	.w8(32'h3c17898d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9183d),
	.w1(32'h3c668d0f),
	.w2(32'h3c618d0c),
	.w3(32'hbc82a6de),
	.w4(32'hbc746af7),
	.w5(32'hbcc191e5),
	.w6(32'hbbf06cf7),
	.w7(32'h3caed23d),
	.w8(32'hbc628d25),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cedf87e),
	.w1(32'h3abdd7e4),
	.w2(32'h3c02c8cd),
	.w3(32'h3c7895d7),
	.w4(32'h3bd2efee),
	.w5(32'h3c110eed),
	.w6(32'hbd287a8e),
	.w7(32'h3bafe34b),
	.w8(32'h3c1ca6da),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9249fa),
	.w1(32'h3c834a1d),
	.w2(32'h3c7991fd),
	.w3(32'h3c1c4653),
	.w4(32'h3bd66326),
	.w5(32'h3ca949c1),
	.w6(32'h3c4c18e4),
	.w7(32'hbbc753de),
	.w8(32'hbd1f6258),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd3a2d),
	.w1(32'hbba9b4e7),
	.w2(32'h3cf11b36),
	.w3(32'h3ca306ab),
	.w4(32'hbc2da13a),
	.w5(32'h3c589108),
	.w6(32'h3b183c05),
	.w7(32'hbcddd54a),
	.w8(32'hbd31d24d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb72a80),
	.w1(32'hbc57b5a5),
	.w2(32'h3ca2a8f5),
	.w3(32'h3d1bdbd3),
	.w4(32'hbbc805bf),
	.w5(32'h3c89370c),
	.w6(32'h3ae9f401),
	.w7(32'hba97d679),
	.w8(32'hbcdd46e1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7186e8),
	.w1(32'hb9f8f635),
	.w2(32'h3c101a9f),
	.w3(32'h3cc9d10c),
	.w4(32'h3abeb5c9),
	.w5(32'h3b81146f),
	.w6(32'hbb912839),
	.w7(32'hbc090ab6),
	.w8(32'hbbc05f3e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8366a0),
	.w1(32'h3c40d7b0),
	.w2(32'h3b9e5a53),
	.w3(32'hba8ebb11),
	.w4(32'hbd17b0ff),
	.w5(32'hbccb7435),
	.w6(32'h3b353eb0),
	.w7(32'h3c96bcfe),
	.w8(32'h3b54f9fa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e18f6),
	.w1(32'hbc0d022e),
	.w2(32'h3b0c9f5a),
	.w3(32'hbb95a81f),
	.w4(32'hbc8fb760),
	.w5(32'h3b945163),
	.w6(32'h3cfeab78),
	.w7(32'hbbcc5e58),
	.w8(32'h3cfed4c0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c95304),
	.w1(32'h3b2f8bdd),
	.w2(32'h3b9502a6),
	.w3(32'h3acf7593),
	.w4(32'h3c93ca0b),
	.w5(32'h3c695fcd),
	.w6(32'h3cb68adf),
	.w7(32'h3c127792),
	.w8(32'h3c99f8cc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d462f),
	.w1(32'hbc3519d3),
	.w2(32'h3c937b2c),
	.w3(32'h3c217cc0),
	.w4(32'hb99e7059),
	.w5(32'h3cb17947),
	.w6(32'h3b27baf3),
	.w7(32'h3b8ca00c),
	.w8(32'hbcd399f4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8006ce),
	.w1(32'hbbf56634),
	.w2(32'h3b17c76f),
	.w3(32'hbb6e6f7e),
	.w4(32'h3c39eb9c),
	.w5(32'h3c5f686f),
	.w6(32'h3c07bed5),
	.w7(32'h3c14bfef),
	.w8(32'h3ca58ca0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb770ffe),
	.w1(32'hbc49a48f),
	.w2(32'hbc4121d5),
	.w3(32'h3afea212),
	.w4(32'h3c9f84ce),
	.w5(32'h3c35ad28),
	.w6(32'h3b3fa8b6),
	.w7(32'h3beee404),
	.w8(32'hba080c32),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c268a40),
	.w1(32'h3c9704cb),
	.w2(32'hbc02cc0e),
	.w3(32'hba397dd2),
	.w4(32'hbae2ab02),
	.w5(32'hbcafe2b9),
	.w6(32'hbbcb14e7),
	.w7(32'h3ca24b45),
	.w8(32'h3d2ae438),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c273674),
	.w1(32'h3b852067),
	.w2(32'h3c0df140),
	.w3(32'hbcb61d7b),
	.w4(32'hbc328b59),
	.w5(32'h3b7a142f),
	.w6(32'hba0dae06),
	.w7(32'hbc27bfb2),
	.w8(32'hbce071cc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a95a3),
	.w1(32'hbc2d1cd4),
	.w2(32'h3940ccaa),
	.w3(32'h3c02b05b),
	.w4(32'h39e4c203),
	.w5(32'h3c1059fc),
	.w6(32'h395e49a7),
	.w7(32'hbbbf9c43),
	.w8(32'hbb2badc5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf5caa),
	.w1(32'hbbfc58c0),
	.w2(32'hbc978c97),
	.w3(32'hbb357213),
	.w4(32'h3c1bbcce),
	.w5(32'h3c4cfe42),
	.w6(32'h3b2e7780),
	.w7(32'hbc19aa57),
	.w8(32'hbbd102ec),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ccfb7),
	.w1(32'hbae863a8),
	.w2(32'hbb433a83),
	.w3(32'hbc571ab4),
	.w4(32'hbb6795ed),
	.w5(32'hbc71d63d),
	.w6(32'hbbd1a8b9),
	.w7(32'h3c6f946e),
	.w8(32'h3d04fbd0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4839b4),
	.w1(32'hbbcff89f),
	.w2(32'hbbcc784b),
	.w3(32'hbc33e489),
	.w4(32'h3c429df9),
	.w5(32'h3c4071c8),
	.w6(32'h3d07b085),
	.w7(32'hbbe17f4b),
	.w8(32'h3d1af58f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a1f57),
	.w1(32'h3c252183),
	.w2(32'hbb0db8c2),
	.w3(32'hbcbb89c8),
	.w4(32'h3a2ca57e),
	.w5(32'hbbadb2ee),
	.w6(32'h3c7bf3b9),
	.w7(32'hbb9aabbf),
	.w8(32'hbc326a13),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7d2cc),
	.w1(32'h3b9922d0),
	.w2(32'hbb930227),
	.w3(32'h3b70a8af),
	.w4(32'h3a7ffaf4),
	.w5(32'h3b0e4d6b),
	.w6(32'h3bd15df8),
	.w7(32'h3b371215),
	.w8(32'hba1e2200),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc815bfb),
	.w1(32'hbcaf75dc),
	.w2(32'hbcdf5062),
	.w3(32'h3bca08ac),
	.w4(32'hbcb1265c),
	.w5(32'hbb1a5444),
	.w6(32'hbc29ae6a),
	.w7(32'hbc89dc35),
	.w8(32'hbbfc3fa0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbf9ae),
	.w1(32'hbd00d368),
	.w2(32'hbce17cdd),
	.w3(32'hbbc838e5),
	.w4(32'h3c9c7f8c),
	.w5(32'hbcaa9d1b),
	.w6(32'h3a492e89),
	.w7(32'h3d0c1c70),
	.w8(32'h3d881417),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfca22),
	.w1(32'hbbedae2d),
	.w2(32'hbcdf2246),
	.w3(32'hbd53b019),
	.w4(32'h3bb7d377),
	.w5(32'h3bf70550),
	.w6(32'hba645417),
	.w7(32'hbd0aa20c),
	.w8(32'hbccf7479),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21d7b4),
	.w1(32'h3acf2357),
	.w2(32'hbba308d7),
	.w3(32'h3c561bde),
	.w4(32'h3c0fdfd7),
	.w5(32'hbbeba754),
	.w6(32'hbc86c85e),
	.w7(32'h3c19b02e),
	.w8(32'hbb58589a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a06cd),
	.w1(32'hba8762e4),
	.w2(32'hbafbfdea),
	.w3(32'hba4d7dd8),
	.w4(32'h3a161404),
	.w5(32'h3c2b384b),
	.w6(32'hbb0a7599),
	.w7(32'hbb7a2367),
	.w8(32'h3ae9c628),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af33a9),
	.w1(32'h3b304775),
	.w2(32'hbc363802),
	.w3(32'h39c1f2ed),
	.w4(32'h3ba8e3a2),
	.w5(32'h3ca43d7f),
	.w6(32'h3bd03dd9),
	.w7(32'hbbb64075),
	.w8(32'h3cfcbe79),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ea3ad),
	.w1(32'hbc04b80f),
	.w2(32'hbc076aaf),
	.w3(32'hbc11bd92),
	.w4(32'h3c40f02f),
	.w5(32'h3c16437a),
	.w6(32'hbc068d8a),
	.w7(32'hbb0565f6),
	.w8(32'h3ca458aa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d9bd5),
	.w1(32'hb9b33cd6),
	.w2(32'h3a2c536d),
	.w3(32'hbc684f79),
	.w4(32'hbbb2c2ac),
	.w5(32'hbb161b85),
	.w6(32'h3bfc6eb1),
	.w7(32'hbbe4eec3),
	.w8(32'h3a6f33a0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88a7c2),
	.w1(32'h3bbd6ad0),
	.w2(32'hbcbae9df),
	.w3(32'h3acf2fc8),
	.w4(32'hbb77c05e),
	.w5(32'hbd378f10),
	.w6(32'h3bad4af9),
	.w7(32'h3cf79fb6),
	.w8(32'h3ca9cd90),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce97cb0),
	.w1(32'h3baa0eec),
	.w2(32'h3a9cde29),
	.w3(32'hbd3a730b),
	.w4(32'h3aa9c431),
	.w5(32'h3bf320e3),
	.w6(32'hbc7c9e16),
	.w7(32'hbafef489),
	.w8(32'h3b0b4f59),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70dd8a),
	.w1(32'hbb576afc),
	.w2(32'hba96d478),
	.w3(32'hba8784f5),
	.w4(32'h3c665b74),
	.w5(32'h3c0fb818),
	.w6(32'h3bfcb319),
	.w7(32'hbc7c4567),
	.w8(32'h3ad6b8c8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bfaeb),
	.w1(32'hbbf56411),
	.w2(32'h3b42e15c),
	.w3(32'hb96a7b8a),
	.w4(32'hbc824d75),
	.w5(32'hbd137b1c),
	.w6(32'h3c0def7d),
	.w7(32'h3ca3f86a),
	.w8(32'h3c1cc54f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce7ab95),
	.w1(32'h3c3c141c),
	.w2(32'hb9d4701c),
	.w3(32'hbc99e1a0),
	.w4(32'hb9bb0b74),
	.w5(32'h3c2a9de2),
	.w6(32'hbcdca28a),
	.w7(32'hbb0a9a81),
	.w8(32'h3b91d203),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72b6fa),
	.w1(32'hbc62c4f1),
	.w2(32'hbc5126b4),
	.w3(32'h3b859f71),
	.w4(32'hbb7c1126),
	.w5(32'h3bd12478),
	.w6(32'h3bbb16ac),
	.w7(32'h39d2f3ce),
	.w8(32'hbcadb28e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104610),
	.w1(32'hbad21973),
	.w2(32'h3b831a1f),
	.w3(32'h3d017526),
	.w4(32'hbb6f491d),
	.w5(32'h3baf475b),
	.w6(32'hbbb6a536),
	.w7(32'hbb0ae330),
	.w8(32'hbcb4d452),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb032f70),
	.w1(32'hbc1ebb6d),
	.w2(32'h3a27f2a3),
	.w3(32'hbb81f0b0),
	.w4(32'hbc939bca),
	.w5(32'h3b784e17),
	.w6(32'hbb657a84),
	.w7(32'hbc3074d7),
	.w8(32'h3c2b6617),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdd2fe),
	.w1(32'hbbd8c806),
	.w2(32'h3c973972),
	.w3(32'hbb2e8219),
	.w4(32'hbb8fd956),
	.w5(32'h3ac6818d),
	.w6(32'hbc0cee8e),
	.w7(32'h3b9f03a5),
	.w8(32'hbbafe2cd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae9c63),
	.w1(32'h3c05956a),
	.w2(32'hbc871e5d),
	.w3(32'h3bd38833),
	.w4(32'h3be55895),
	.w5(32'hbc446ff0),
	.w6(32'hba10e20d),
	.w7(32'h3c59a192),
	.w8(32'h3c1be295),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5702d),
	.w1(32'h3acc93be),
	.w2(32'h3d0946b9),
	.w3(32'hbb57e825),
	.w4(32'hbc404492),
	.w5(32'h3c322097),
	.w6(32'hbca6fbbd),
	.w7(32'hbc92aaa9),
	.w8(32'hbd2241ee),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62b3d1),
	.w1(32'h3b624fa8),
	.w2(32'h3baa845d),
	.w3(32'h3cd96560),
	.w4(32'hbbf98aca),
	.w5(32'hbc554bb8),
	.w6(32'hba8d8bbb),
	.w7(32'hbbf03b50),
	.w8(32'h3b53c7c4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6b323),
	.w1(32'hba9fe794),
	.w2(32'h3c4062c0),
	.w3(32'hbce03701),
	.w4(32'hbcb3296c),
	.w5(32'hbc9bb5a3),
	.w6(32'hbb717be7),
	.w7(32'h3c5adb00),
	.w8(32'hbcbb88fc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0eb42),
	.w1(32'h3b82811f),
	.w2(32'h3cd7fc0c),
	.w3(32'h3c92b10e),
	.w4(32'hbb58280f),
	.w5(32'hbc6ce744),
	.w6(32'hbc83c795),
	.w7(32'h3c2776a6),
	.w8(32'hbc81dba1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c850dae),
	.w1(32'h3bbe4e1d),
	.w2(32'h3b1413bd),
	.w3(32'h3c4efe05),
	.w4(32'h397f2b67),
	.w5(32'h3c12bb11),
	.w6(32'hbc6f54b7),
	.w7(32'h3bf44b08),
	.w8(32'hbcf71db0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcce323),
	.w1(32'hbb176a28),
	.w2(32'h3aa86b2d),
	.w3(32'hb9691024),
	.w4(32'hbb828226),
	.w5(32'h3c68237f),
	.w6(32'h3b797666),
	.w7(32'hbbde3cd8),
	.w8(32'hbc29243b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d9fe2),
	.w1(32'hbcad7515),
	.w2(32'hbc274a1f),
	.w3(32'h3bd94a15),
	.w4(32'h3cacbf9e),
	.w5(32'h3d3f97e5),
	.w6(32'h3a2bd78b),
	.w7(32'hbc4b5738),
	.w8(32'h3b74bb8b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc362b80),
	.w1(32'hbb0b89bf),
	.w2(32'hbcdaeedb),
	.w3(32'h3c02ae40),
	.w4(32'hbb4c1235),
	.w5(32'hbc852ce4),
	.w6(32'h3c725a89),
	.w7(32'h3c84c900),
	.w8(32'h3d19eec5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8ac92),
	.w1(32'hbb8df8b0),
	.w2(32'h3bb7083c),
	.w3(32'h3cafae72),
	.w4(32'hbb978504),
	.w5(32'h3c2f287a),
	.w6(32'hbc4bf04e),
	.w7(32'hbb0a98e4),
	.w8(32'hbbdffc73),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac764),
	.w1(32'h3b89b804),
	.w2(32'hba4cc67b),
	.w3(32'hbbb12dc8),
	.w4(32'h3b027d63),
	.w5(32'h3b82bf93),
	.w6(32'h3c9e2298),
	.w7(32'h3bc57df4),
	.w8(32'h3b9f1748),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16b7ab),
	.w1(32'hbba4e85a),
	.w2(32'hbb2660cc),
	.w3(32'h3b58223e),
	.w4(32'hbb943d1d),
	.w5(32'hbc1b341e),
	.w6(32'hbb2763b9),
	.w7(32'h3b4174fa),
	.w8(32'hbbb43d83),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf92612),
	.w1(32'hbbaa09d0),
	.w2(32'hbb847ac3),
	.w3(32'hbb8cc9f5),
	.w4(32'hbbe9ad88),
	.w5(32'hbc000128),
	.w6(32'hbbb9aa8b),
	.w7(32'hbb79759a),
	.w8(32'hbb90f605),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ab566),
	.w1(32'hbaa2b043),
	.w2(32'hbc351a09),
	.w3(32'hbb7a2fe9),
	.w4(32'h3c8da2ae),
	.w5(32'h3c873a2b),
	.w6(32'hba10d4ec),
	.w7(32'h3c33fcc8),
	.w8(32'hbac14f0a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83eeba),
	.w1(32'hbbc80b5b),
	.w2(32'h3bda9e4b),
	.w3(32'h3b208d22),
	.w4(32'hbc11c2aa),
	.w5(32'hbc7b95ad),
	.w6(32'hbbbd591d),
	.w7(32'hbb776c4f),
	.w8(32'h3a94e764),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b991fb0),
	.w1(32'h3c152c28),
	.w2(32'h3b1575e6),
	.w3(32'h3ba9fc11),
	.w4(32'h3c6ec5ff),
	.w5(32'h3acdd3ed),
	.w6(32'h3ba2a373),
	.w7(32'hbc1c0fc3),
	.w8(32'hbc8b4997),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab75e7c),
	.w1(32'hbc57450c),
	.w2(32'h3c26f632),
	.w3(32'h3c1ff7d7),
	.w4(32'h3a4d3ca4),
	.w5(32'h3a6e78d4),
	.w6(32'hbc554240),
	.w7(32'h3ab70926),
	.w8(32'hbc5d2cf2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd12f828),
	.w1(32'hbd3a7209),
	.w2(32'hbcaa46d6),
	.w3(32'hbb158427),
	.w4(32'h3bb479d5),
	.w5(32'h3c149712),
	.w6(32'h3b03f9d2),
	.w7(32'h3c8e2c92),
	.w8(32'h3a3599e8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3365a4),
	.w1(32'hbc23c037),
	.w2(32'h3c0eb224),
	.w3(32'hbc668183),
	.w4(32'h3c193d1b),
	.w5(32'h3c6eb8c4),
	.w6(32'hbbcd6aeb),
	.w7(32'h3c5705bc),
	.w8(32'h3ad4e686),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc804017),
	.w1(32'hbc88375d),
	.w2(32'hbc1759f2),
	.w3(32'hba26fbe5),
	.w4(32'h36d913b4),
	.w5(32'hbaf3e4fb),
	.w6(32'hbbc98687),
	.w7(32'h3c2bdb63),
	.w8(32'hbc45e72e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd68f53),
	.w1(32'hbc46b4fc),
	.w2(32'h3b4d94a8),
	.w3(32'hbc05b03a),
	.w4(32'hbc6d1c61),
	.w5(32'hbc550f74),
	.w6(32'hbc23d305),
	.w7(32'hbb6aad8b),
	.w8(32'h3b49301a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0474b5),
	.w1(32'hbb0f78e8),
	.w2(32'h3b47650d),
	.w3(32'hbb74780c),
	.w4(32'h3ca1cbfb),
	.w5(32'h3bb830d0),
	.w6(32'h3c0d24b9),
	.w7(32'h3bcd8e01),
	.w8(32'hb9f7c2e5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21fe8c),
	.w1(32'hbaf7a3d1),
	.w2(32'h397e752a),
	.w3(32'hbb4c29d2),
	.w4(32'hbc6552c1),
	.w5(32'hbc997047),
	.w6(32'hbb2eca5f),
	.w7(32'hbc9b7ab3),
	.w8(32'hbc4b6aee),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ac5de),
	.w1(32'hbbe0f7e9),
	.w2(32'h3c747413),
	.w3(32'hbc475854),
	.w4(32'hbce64b6a),
	.w5(32'hbca7baef),
	.w6(32'hbc217e68),
	.w7(32'hbb068c99),
	.w8(32'h3d12747c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f9a5d),
	.w1(32'h3bd91c2d),
	.w2(32'hbbab5d56),
	.w3(32'h3c5b2cce),
	.w4(32'h3aa31bc2),
	.w5(32'hbc4325a2),
	.w6(32'h3c91074b),
	.w7(32'hbc35672e),
	.w8(32'hbcd06f51),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80a67b),
	.w1(32'hbc301f68),
	.w2(32'hbc6c82e0),
	.w3(32'hbcbf1d1a),
	.w4(32'hbc1cdd15),
	.w5(32'hbc3d58b8),
	.w6(32'hbc74d44b),
	.w7(32'hbc5b75bc),
	.w8(32'hbd087dde),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc368ebb),
	.w1(32'hbaa49c5d),
	.w2(32'hbb135356),
	.w3(32'h3c604a5c),
	.w4(32'hb985501e),
	.w5(32'h3b786107),
	.w6(32'h3b9fbc0f),
	.w7(32'h3bf45831),
	.w8(32'h3c797315),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d1f0b),
	.w1(32'hbc47a1b8),
	.w2(32'hbc049339),
	.w3(32'hbb12432a),
	.w4(32'h3c5cc9ed),
	.w5(32'h3b08e250),
	.w6(32'h3bc2119e),
	.w7(32'h3af9fb94),
	.w8(32'hbc88bc9a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f9974),
	.w1(32'h39f5d6dd),
	.w2(32'h3ba1f2a3),
	.w3(32'h3b95efb0),
	.w4(32'hba84304d),
	.w5(32'hbb0434fe),
	.w6(32'h3a90ecb9),
	.w7(32'hb987ecc7),
	.w8(32'h3a06dd89),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3b1b7),
	.w1(32'h373007cd),
	.w2(32'hbd2bbb2e),
	.w3(32'hbb6b01c8),
	.w4(32'h3d06168f),
	.w5(32'h3d478792),
	.w6(32'h3ae1944e),
	.w7(32'h3d018952),
	.w8(32'h3c656712),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd30bf91),
	.w1(32'hbd22aba2),
	.w2(32'hbbd7ff49),
	.w3(32'h3c465b72),
	.w4(32'h3ce82ca8),
	.w5(32'h3c773043),
	.w6(32'hbc705110),
	.w7(32'h3c3112fd),
	.w8(32'h3cc3eff4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af134),
	.w1(32'hbc159370),
	.w2(32'h3c09ce01),
	.w3(32'hbc940078),
	.w4(32'h3c096d8e),
	.w5(32'hbcae948b),
	.w6(32'hbc281df1),
	.w7(32'hbbe483d2),
	.w8(32'h3bd3c222),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9127ea),
	.w1(32'h3c06a4e5),
	.w2(32'h3bdec99b),
	.w3(32'hbb1d380f),
	.w4(32'hbc27617f),
	.w5(32'hbbbe0f42),
	.w6(32'h3ad0d880),
	.w7(32'h387ab4d3),
	.w8(32'h3be88c94),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fde46),
	.w1(32'h3c8d31fd),
	.w2(32'hbc2e12e2),
	.w3(32'h3b8ffd08),
	.w4(32'h3bd366c0),
	.w5(32'h3c90be85),
	.w6(32'h3c7293b1),
	.w7(32'hbb9e920a),
	.w8(32'h3c8ac9bb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aff1a),
	.w1(32'hbbedac35),
	.w2(32'hbaf2f44b),
	.w3(32'hbb15b104),
	.w4(32'h3c2407be),
	.w5(32'h3c4137ad),
	.w6(32'h3babff5d),
	.w7(32'h3ba282e2),
	.w8(32'h3a281ed1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76c3bc),
	.w1(32'hbccaeb2c),
	.w2(32'h3beb2d9b),
	.w3(32'hbc20a927),
	.w4(32'hbc392008),
	.w5(32'h3b9e3429),
	.w6(32'hbd0018a2),
	.w7(32'hbabb3bb5),
	.w8(32'h3b759e3f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd549b0),
	.w1(32'hbb5d0bec),
	.w2(32'hbc89bd75),
	.w3(32'h3ab28673),
	.w4(32'h3ce3a79d),
	.w5(32'h3c962107),
	.w6(32'hb959f381),
	.w7(32'h3c222d06),
	.w8(32'h3c1f7d8f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5c765),
	.w1(32'hbc86a977),
	.w2(32'hbab1f58b),
	.w3(32'h3c075157),
	.w4(32'h3cae3dfa),
	.w5(32'h3c89a480),
	.w6(32'hbb96b408),
	.w7(32'h3ca78245),
	.w8(32'h3c8c6621),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ec585),
	.w1(32'hbb846434),
	.w2(32'h3aa46008),
	.w3(32'h3a8df541),
	.w4(32'h3cf237e3),
	.w5(32'h3cf6f4f5),
	.w6(32'h3c366f65),
	.w7(32'h3c9b210b),
	.w8(32'h3b1e3f42),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeeb429),
	.w1(32'h3c00fcab),
	.w2(32'hbc57df4c),
	.w3(32'h3c465a5c),
	.w4(32'h3bfb1919),
	.w5(32'h3b9c6cb1),
	.w6(32'hbbcb24c7),
	.w7(32'hbc2222cd),
	.w8(32'hbc08b76c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae88b93),
	.w1(32'h3c00c4c9),
	.w2(32'h3b83a3c3),
	.w3(32'h3b9171e3),
	.w4(32'h3c3a6e38),
	.w5(32'h3bca2bfb),
	.w6(32'h3c87dc11),
	.w7(32'hbbc88acd),
	.w8(32'hbbdf3193),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf61233),
	.w1(32'hba27304c),
	.w2(32'h3bb6d4c4),
	.w3(32'hbb518075),
	.w4(32'h3b5aecda),
	.w5(32'h3b5fb8fa),
	.w6(32'hbb92647c),
	.w7(32'h3bdc70e3),
	.w8(32'h3bb9d032),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab621a2),
	.w1(32'hb9c678e3),
	.w2(32'hbc7c9fa6),
	.w3(32'h3bed1b1e),
	.w4(32'hba5dbb6d),
	.w5(32'hba51c84f),
	.w6(32'h3aa4952b),
	.w7(32'hbc0aa39d),
	.w8(32'hbaa47f9e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe42da5),
	.w1(32'h3b37cafa),
	.w2(32'hbc1dfb50),
	.w3(32'h3c2aa58f),
	.w4(32'h3c2ab5cb),
	.w5(32'h3bf72658),
	.w6(32'h3c318876),
	.w7(32'h3c110c66),
	.w8(32'h3c607d5b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85d657),
	.w1(32'h3a90411d),
	.w2(32'hba11ca22),
	.w3(32'hbb83a5de),
	.w4(32'h3c9377fc),
	.w5(32'h3bfa73dd),
	.w6(32'hbb4db491),
	.w7(32'hbc0e7aab),
	.w8(32'hbbba8bf8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dcdaa),
	.w1(32'hbc08dac3),
	.w2(32'h3c884d8b),
	.w3(32'hbaa278ce),
	.w4(32'h3b1cfaf7),
	.w5(32'hbc0d7641),
	.w6(32'hbb9c523f),
	.w7(32'h3982ff59),
	.w8(32'h39975524),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c174e31),
	.w1(32'h3aff511b),
	.w2(32'hbcb1b5b5),
	.w3(32'hbc3d4e0c),
	.w4(32'h3d5949ac),
	.w5(32'h3ca8317c),
	.w6(32'hbc2b3d7a),
	.w7(32'h3b61a8b4),
	.w8(32'hbc1e61b1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd00b700),
	.w1(32'hbd07ac17),
	.w2(32'hbd1d58ae),
	.w3(32'h3b8ca5c1),
	.w4(32'h3d658552),
	.w5(32'h3d1f4ca0),
	.w6(32'hbc6b4f1c),
	.w7(32'h3c6bbcf7),
	.w8(32'hbc24ed26),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd50232b),
	.w1(32'hbd82fb0f),
	.w2(32'h3cb0cb57),
	.w3(32'hbac864b0),
	.w4(32'hbb38f499),
	.w5(32'hbb1418a4),
	.w6(32'hbd3aa1ff),
	.w7(32'h3c6c2e2b),
	.w8(32'h3bc31c43),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02e57b),
	.w1(32'hbbbf16a8),
	.w2(32'h3c418ae5),
	.w3(32'h3c152473),
	.w4(32'hbcb6984a),
	.w5(32'hbd16ccc7),
	.w6(32'h3c6edf78),
	.w7(32'h3b3ca7e5),
	.w8(32'hbbbc49dc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca73e46),
	.w1(32'h3c9b289c),
	.w2(32'hbbfcc3af),
	.w3(32'hbc97144f),
	.w4(32'hbc6baf7d),
	.w5(32'h3c45b3b3),
	.w6(32'h3bfb8d8a),
	.w7(32'h3c92a105),
	.w8(32'h3cbf9d56),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc629df4),
	.w1(32'hbc4a6324),
	.w2(32'hbb90ea87),
	.w3(32'h3c859825),
	.w4(32'hbb447839),
	.w5(32'hbb20e7b9),
	.w6(32'h3ba14c55),
	.w7(32'h3bd70aab),
	.w8(32'h3b280f3a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb40568),
	.w1(32'hbb52ef4b),
	.w2(32'h3c5cc5d8),
	.w3(32'h3b365fc0),
	.w4(32'h3c0b0052),
	.w5(32'h3b90e005),
	.w6(32'hbb17fa9a),
	.w7(32'h3b5e5000),
	.w8(32'h3c0315de),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd837fb),
	.w1(32'hbc587fc2),
	.w2(32'hbbce76a1),
	.w3(32'hbb3402ff),
	.w4(32'h3c939bd1),
	.w5(32'h3c9264a4),
	.w6(32'hbc2f87ae),
	.w7(32'h3c12956e),
	.w8(32'hbbd109d9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb4bba2),
	.w1(32'hbcab57f8),
	.w2(32'hbb8fb423),
	.w3(32'h3bb22602),
	.w4(32'h3bb00d10),
	.w5(32'h3b00db62),
	.w6(32'hbc624940),
	.w7(32'h3babff70),
	.w8(32'h3b237034),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96a1a5),
	.w1(32'hbcd3099f),
	.w2(32'h3cd6aa56),
	.w3(32'hbc4f3dfb),
	.w4(32'hbd5f9454),
	.w5(32'hbd260e35),
	.w6(32'hbc974b46),
	.w7(32'hbd1bd5b0),
	.w8(32'hbd03ce60),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc007c9),
	.w1(32'h3ccb7bde),
	.w2(32'hba84ed93),
	.w3(32'h3c42dd5c),
	.w4(32'hbb65120d),
	.w5(32'hbb41aa71),
	.w6(32'h3c7399b1),
	.w7(32'hb956fcb6),
	.w8(32'hbac97bc5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5bb1e),
	.w1(32'hb9ef45eb),
	.w2(32'hbb3c8582),
	.w3(32'h3bb53c28),
	.w4(32'hbb411067),
	.w5(32'h3c36bc53),
	.w6(32'h3a8fbf7f),
	.w7(32'h3a0189ad),
	.w8(32'h3a3ce132),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44d3ed),
	.w1(32'h3b82b303),
	.w2(32'hbc99749a),
	.w3(32'h3c48246a),
	.w4(32'hba0b3bbb),
	.w5(32'h3cc90a33),
	.w6(32'h3b938a41),
	.w7(32'h3a9a9456),
	.w8(32'h3afc05b1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34c38e),
	.w1(32'hb9245462),
	.w2(32'hbacb5790),
	.w3(32'h3c4cef51),
	.w4(32'hb9eaf7b1),
	.w5(32'h3a2e3135),
	.w6(32'h3a061069),
	.w7(32'hbc1033c4),
	.w8(32'hbc2c22a2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba92a80),
	.w1(32'hbbfdb50b),
	.w2(32'h3c62e435),
	.w3(32'h3bbad9e2),
	.w4(32'h3c6fcc7f),
	.w5(32'h3c888422),
	.w6(32'hbc0eb565),
	.w7(32'hbaba8c77),
	.w8(32'hbc615d4f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc790a),
	.w1(32'hbc81cb45),
	.w2(32'hbbd13d75),
	.w3(32'h3c258561),
	.w4(32'h3bb1e313),
	.w5(32'h3b5c0d2b),
	.w6(32'hbc56fc84),
	.w7(32'h3ca2be9f),
	.w8(32'h3c82563e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule