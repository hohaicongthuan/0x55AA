module layer_8_featuremap_47(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadafff),
	.w1(32'h3b858a61),
	.w2(32'hbb84e954),
	.w3(32'h3b24265b),
	.w4(32'h3c387430),
	.w5(32'hba37dbe9),
	.w6(32'hba88c110),
	.w7(32'h3ba11efb),
	.w8(32'hba82cefa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb310ee),
	.w1(32'hbbc7502c),
	.w2(32'hbb45fabe),
	.w3(32'hbb1315d9),
	.w4(32'hbba9852f),
	.w5(32'h3aa5411b),
	.w6(32'h3b98448c),
	.w7(32'hba40bfc1),
	.w8(32'h3bce9891),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb802de0),
	.w1(32'hbc193d9c),
	.w2(32'hbc2b4711),
	.w3(32'hbb7c938c),
	.w4(32'hbbc58375),
	.w5(32'hbba23c5c),
	.w6(32'h3b9133e6),
	.w7(32'hbb047551),
	.w8(32'hbbb1a63e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc32d97),
	.w1(32'h3aa3300f),
	.w2(32'h3b994de3),
	.w3(32'h3c6ec242),
	.w4(32'h3bfc627b),
	.w5(32'h3a1ad42a),
	.w6(32'h3c0615c4),
	.w7(32'h3c049652),
	.w8(32'h3b8a2a60),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dbfef),
	.w1(32'h3a7ec6fa),
	.w2(32'h3bbc35ea),
	.w3(32'hba425844),
	.w4(32'h3a47952f),
	.w5(32'h3c03defc),
	.w6(32'h3a1c82ee),
	.w7(32'h3ac7cc3e),
	.w8(32'h3c1232e4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc467190),
	.w1(32'hbc47f68a),
	.w2(32'h3bca5143),
	.w3(32'hbb1bf120),
	.w4(32'hbc242143),
	.w5(32'h3bb6425c),
	.w6(32'hbb09d861),
	.w7(32'hba22e578),
	.w8(32'h3c501de3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29559a),
	.w1(32'hb9c200a2),
	.w2(32'hba05d7d0),
	.w3(32'hbaa0df48),
	.w4(32'hb9ef7b15),
	.w5(32'hb8600565),
	.w6(32'hba077330),
	.w7(32'hba5d301c),
	.w8(32'hba68ab37),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06e3ed),
	.w1(32'h3b3cba7d),
	.w2(32'hbb950c68),
	.w3(32'h3c484e31),
	.w4(32'h3c289b11),
	.w5(32'h3b933e1e),
	.w6(32'h3c61c17b),
	.w7(32'h3c0d49af),
	.w8(32'h3c104b24),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f7c75),
	.w1(32'hbaf6e278),
	.w2(32'h3b5da5ed),
	.w3(32'hbb2fe89d),
	.w4(32'h3aec3832),
	.w5(32'h3ba7f5d0),
	.w6(32'h3bf60b8a),
	.w7(32'h3bf0ff54),
	.w8(32'h3bc44a64),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b330874),
	.w1(32'h3a254919),
	.w2(32'hbc51b8dc),
	.w3(32'h3b6339d3),
	.w4(32'hbb91adb4),
	.w5(32'hbc560e9b),
	.w6(32'h3a726029),
	.w7(32'hbae4d064),
	.w8(32'hbc0096d3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b7e1b),
	.w1(32'h3b528699),
	.w2(32'hbbfd1c4f),
	.w3(32'h3be5ab33),
	.w4(32'h3c74735c),
	.w5(32'hbb2bbe07),
	.w6(32'h3a8e4b78),
	.w7(32'h3bf0c1b1),
	.w8(32'hb9b87979),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53d757),
	.w1(32'h3bb7e24b),
	.w2(32'h3b4ff87f),
	.w3(32'h3bb6282c),
	.w4(32'h3c034c41),
	.w5(32'h3c0d5423),
	.w6(32'hbb587cdc),
	.w7(32'hbbb79f8c),
	.w8(32'h3b6b7131),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f4b5f),
	.w1(32'hbb86b591),
	.w2(32'hbb7dd48f),
	.w3(32'hbb4fca3a),
	.w4(32'hbbd32e79),
	.w5(32'hbbc04e9b),
	.w6(32'h3afb8e8b),
	.w7(32'hba5389ae),
	.w8(32'h3b17a954),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9738ea7),
	.w1(32'hba3cb40f),
	.w2(32'h38eac962),
	.w3(32'hba8f3486),
	.w4(32'hba90d6a5),
	.w5(32'hb9e17220),
	.w6(32'h3996d8f1),
	.w7(32'h3a943cee),
	.w8(32'hb8548210),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38721cd3),
	.w1(32'h3a375df5),
	.w2(32'h3a861f63),
	.w3(32'hb955b510),
	.w4(32'h3a47b27b),
	.w5(32'h3a8f6820),
	.w6(32'h3a87f14c),
	.w7(32'h3adba5b9),
	.w8(32'h39bf2c49),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a9a6b),
	.w1(32'h3abed1d3),
	.w2(32'hb94d8c17),
	.w3(32'h3a2fcd0b),
	.w4(32'h39e48625),
	.w5(32'hba8ae63e),
	.w6(32'hba47f63e),
	.w7(32'hb9f6f708),
	.w8(32'hbb201b6b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e076f),
	.w1(32'hba78c46c),
	.w2(32'hb998e9f9),
	.w3(32'h3b3f50ae),
	.w4(32'h3ae6d33c),
	.w5(32'hbb9814c5),
	.w6(32'h3a3545b5),
	.w7(32'h3c354f42),
	.w8(32'h3bc63521),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55b3fd),
	.w1(32'h3bb8d2be),
	.w2(32'hbac96d12),
	.w3(32'h3c287f8c),
	.w4(32'h3ba9315d),
	.w5(32'h39f33714),
	.w6(32'h3be361bd),
	.w7(32'hba1ca0a9),
	.w8(32'hbaefacb8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d28b39e),
	.w1(32'h3d09e9a4),
	.w2(32'hbcc1275f),
	.w3(32'h3d3ddc7e),
	.w4(32'h3d818e2e),
	.w5(32'hbc45009b),
	.w6(32'hbc223c9f),
	.w7(32'hbb43572c),
	.w8(32'hbd31e80c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba57f09),
	.w1(32'h3b947833),
	.w2(32'h3be73803),
	.w3(32'hbc02c342),
	.w4(32'hbbabed4a),
	.w5(32'h3bbaaf3f),
	.w6(32'hbc3818db),
	.w7(32'hbbb2f55c),
	.w8(32'h3c6c1f31),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee3628),
	.w1(32'h3bf853de),
	.w2(32'h3c7c6c7b),
	.w3(32'hbb07d00c),
	.w4(32'h3beb7f82),
	.w5(32'h3cb1b37a),
	.w6(32'hbc499e18),
	.w7(32'hbb442d41),
	.w8(32'h3c824830),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0e8b1),
	.w1(32'hbcf00e92),
	.w2(32'hbca5418c),
	.w3(32'hbcbf8193),
	.w4(32'hbcde8cc3),
	.w5(32'hbc83b2ca),
	.w6(32'hbc5c75ae),
	.w7(32'hbc914ccd),
	.w8(32'hbbdb9fac),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba628e6),
	.w1(32'h3c8fb516),
	.w2(32'hbc0a9711),
	.w3(32'h3c1538d5),
	.w4(32'h3d1e5f15),
	.w5(32'h3b915f6e),
	.w6(32'h3a7002e9),
	.w7(32'h3cc5cb3c),
	.w8(32'hb8af0720),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05dbf2),
	.w1(32'hbb9fa53b),
	.w2(32'hbad79516),
	.w3(32'hbc29155d),
	.w4(32'hbc238d9e),
	.w5(32'hbb625853),
	.w6(32'hbba10edb),
	.w7(32'hbac8c92c),
	.w8(32'hba5f73a2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e961d),
	.w1(32'h3a9674ce),
	.w2(32'hbac37acf),
	.w3(32'h3b48e12c),
	.w4(32'h3b53a85c),
	.w5(32'h3ad59591),
	.w6(32'hba162a5c),
	.w7(32'hbaf8066b),
	.w8(32'h3bc2c84e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fd65a),
	.w1(32'hbaec5217),
	.w2(32'hbae3c184),
	.w3(32'h3aca75c4),
	.w4(32'h3c1277ce),
	.w5(32'h3c6489dc),
	.w6(32'hbbb62daf),
	.w7(32'h3be7a7d6),
	.w8(32'h3c4c086f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838402),
	.w1(32'h3b0f78f9),
	.w2(32'h3b4778f7),
	.w3(32'h3b4cd4c1),
	.w4(32'h3ac4ed5b),
	.w5(32'h3b18fc62),
	.w6(32'h3a2a533e),
	.w7(32'h389e970b),
	.w8(32'h3ba3035e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e14c83d),
	.w1(32'h3d800b12),
	.w2(32'h3cc733cc),
	.w3(32'h3defdba0),
	.w4(32'h3dd19034),
	.w5(32'h3e10743e),
	.w6(32'h3c214df5),
	.w7(32'h3da72524),
	.w8(32'h3d8ac59b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfd6e),
	.w1(32'hba6751cb),
	.w2(32'hbbe02568),
	.w3(32'h3bef1270),
	.w4(32'h3c181588),
	.w5(32'hb84c1ae4),
	.w6(32'hbc09df83),
	.w7(32'hba2131ea),
	.w8(32'hbb168910),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac76556),
	.w1(32'hbb1ad36b),
	.w2(32'hb9c63c35),
	.w3(32'hb96c22df),
	.w4(32'h3923250f),
	.w5(32'h3ac8cacc),
	.w6(32'h3af1f3e2),
	.w7(32'h3af80b49),
	.w8(32'h3b722447),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff864),
	.w1(32'h3b11a454),
	.w2(32'h3bde63cd),
	.w3(32'h3beff69d),
	.w4(32'h3ba04e85),
	.w5(32'h3b5b1c10),
	.w6(32'h39a4d21d),
	.w7(32'h37608d7f),
	.w8(32'h3bb8f5e1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68db8f),
	.w1(32'h39155674),
	.w2(32'h3c28cb54),
	.w3(32'hbb89af29),
	.w4(32'hbaa8729d),
	.w5(32'h3c4a4d03),
	.w6(32'hbaa222de),
	.w7(32'hbb3f80e8),
	.w8(32'h3bd8a4b7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad11a34),
	.w1(32'hbb4d2e5c),
	.w2(32'hba28c7aa),
	.w3(32'hbacd71d9),
	.w4(32'hbb0b7e9c),
	.w5(32'hbb27b870),
	.w6(32'hbb08eb3d),
	.w7(32'h39a81a5c),
	.w8(32'h3b07e39e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb6c68),
	.w1(32'h3b09028b),
	.w2(32'hb9f6d60d),
	.w3(32'hbabbefb9),
	.w4(32'hbb5be1e8),
	.w5(32'hba68ec58),
	.w6(32'h3b861325),
	.w7(32'hb9d25fe6),
	.w8(32'h3a5f3ec3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ef3f4),
	.w1(32'hb9bd31f6),
	.w2(32'h3b226969),
	.w3(32'hbc070567),
	.w4(32'hbc38d7ab),
	.w5(32'hbc021c38),
	.w6(32'hbbaaa686),
	.w7(32'hbc277b3a),
	.w8(32'hbc18895e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc9ab5),
	.w1(32'h3c99cf0b),
	.w2(32'h3a84629d),
	.w3(32'h3cb1cee1),
	.w4(32'h3ca69195),
	.w5(32'h3bf590af),
	.w6(32'h3c706d3c),
	.w7(32'h3bf2d094),
	.w8(32'hba4c23a3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39419e),
	.w1(32'hb9c0cff1),
	.w2(32'hbb0d4d06),
	.w3(32'hb8e44869),
	.w4(32'hba70bfc0),
	.w5(32'hbadfc16d),
	.w6(32'hba25a52e),
	.w7(32'hbaa79e4b),
	.w8(32'h3aae8c6e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cdd4c),
	.w1(32'hbbcc6d36),
	.w2(32'hbb63043e),
	.w3(32'hbb675522),
	.w4(32'hbb79b05e),
	.w5(32'hba215a09),
	.w6(32'h3af6ae76),
	.w7(32'h3aa5cc80),
	.w8(32'h3bcc5b42),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a418438),
	.w1(32'h3b0a78df),
	.w2(32'h3b210389),
	.w3(32'hb91475db),
	.w4(32'h3b0bc4c5),
	.w5(32'h3b2c5fa8),
	.w6(32'h3afee185),
	.w7(32'h3b6bb454),
	.w8(32'h3a8242ff),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba046205),
	.w1(32'hbabce78a),
	.w2(32'hbb7a334d),
	.w3(32'hbb16b12c),
	.w4(32'hbaa1a51c),
	.w5(32'hbb8b9a5c),
	.w6(32'hbb6d8b45),
	.w7(32'hbb30d3a5),
	.w8(32'hbb3d38e3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ab1c7),
	.w1(32'h3c4fe0ad),
	.w2(32'h3c441128),
	.w3(32'h3d11d49c),
	.w4(32'h3cf94c5e),
	.w5(32'h3ceb6f70),
	.w6(32'h3cb5b49d),
	.w7(32'h3c74ecac),
	.w8(32'h3ccc92dc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c42f1),
	.w1(32'h3bef73de),
	.w2(32'hba0a0e07),
	.w3(32'h3c373be4),
	.w4(32'h3c1b87a2),
	.w5(32'h392fe540),
	.w6(32'h3b8bce19),
	.w7(32'h3b40fd2e),
	.w8(32'hbb541d40),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ace6b),
	.w1(32'hbb899a63),
	.w2(32'h3a95970b),
	.w3(32'hbac25bbe),
	.w4(32'hbb9582fd),
	.w5(32'h393a79b2),
	.w6(32'hbb8f1c9a),
	.w7(32'hbb2341b9),
	.w8(32'hb985fc96),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba840f9),
	.w1(32'h3bbb0782),
	.w2(32'h3b6bfcb7),
	.w3(32'h3c178187),
	.w4(32'h3c574c28),
	.w5(32'h3c16764e),
	.w6(32'h3be3cc83),
	.w7(32'h3c1927cd),
	.w8(32'h3bf7a9ea),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d9d29),
	.w1(32'hbb00f1b9),
	.w2(32'hbc558682),
	.w3(32'h3afa6453),
	.w4(32'h3c3a7c35),
	.w5(32'hbbc36f74),
	.w6(32'hbc374a33),
	.w7(32'hbb65b15f),
	.w8(32'hbc802711),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c802262),
	.w1(32'h3c608e60),
	.w2(32'hb7ee4c02),
	.w3(32'h3c5b5ee8),
	.w4(32'h3c6d7e3f),
	.w5(32'hbaac2ee6),
	.w6(32'h3be94d71),
	.w7(32'h3b71e9c4),
	.w8(32'hbbebacb6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947dc85),
	.w1(32'h39e3a9e8),
	.w2(32'hba8a3cf3),
	.w3(32'h3a29caa1),
	.w4(32'h393d119b),
	.w5(32'hba85858e),
	.w6(32'hba177ee7),
	.w7(32'hb96068f1),
	.w8(32'h3a19dd4e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9072bc),
	.w1(32'h3c16e4fb),
	.w2(32'h3a3e98d6),
	.w3(32'hbb805070),
	.w4(32'h3c70fdeb),
	.w5(32'h3b8ffaa3),
	.w6(32'hbc13050f),
	.w7(32'h3bcd1ee3),
	.w8(32'hba321066),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb93569),
	.w1(32'hba6e9129),
	.w2(32'hbb3ac2b2),
	.w3(32'h3babeacb),
	.w4(32'hbb1ce3c5),
	.w5(32'hbae865a5),
	.w6(32'h3a7a9186),
	.w7(32'hbab9c52a),
	.w8(32'hbb24da1e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c6e68),
	.w1(32'hbac86938),
	.w2(32'hbbb249ab),
	.w3(32'h3bbae21f),
	.w4(32'h3c157f01),
	.w5(32'hbb06531d),
	.w6(32'hbba083d4),
	.w7(32'hbae7e002),
	.w8(32'hbb0df618),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcef38c9),
	.w1(32'hbc9fc751),
	.w2(32'h3b9c4f02),
	.w3(32'hbca0b643),
	.w4(32'hbc8013b3),
	.w5(32'h3c1ccbe8),
	.w6(32'hbc684f94),
	.w7(32'hbc883750),
	.w8(32'h3bd7daea),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03a489),
	.w1(32'hbac1f756),
	.w2(32'hbc9129a9),
	.w3(32'h3d100295),
	.w4(32'h3d261bb1),
	.w5(32'hbb403b8b),
	.w6(32'h3a714dd9),
	.w7(32'h3cbd8b1c),
	.w8(32'hbc7fe08d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa86795),
	.w1(32'h3a8b44fb),
	.w2(32'h3b8dca76),
	.w3(32'h3ba456ce),
	.w4(32'h3c18f801),
	.w5(32'h3c212329),
	.w6(32'h3b19c977),
	.w7(32'h3c6cb21b),
	.w8(32'h3c318113),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c439262),
	.w1(32'h3c98dd8f),
	.w2(32'h3bb5f7d1),
	.w3(32'h3c20b27a),
	.w4(32'h3c33e023),
	.w5(32'hbb04e9e2),
	.w6(32'h3b57be25),
	.w7(32'hba4a5175),
	.w8(32'hbc668d73),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3882ee),
	.w1(32'hba1b754e),
	.w2(32'h388c3340),
	.w3(32'hba32b799),
	.w4(32'hb8a8f3d0),
	.w5(32'hb9cc6762),
	.w6(32'hba0a8c9f),
	.w7(32'hba82b51a),
	.w8(32'h3ae811c4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4991d),
	.w1(32'h3d0b2a3f),
	.w2(32'h3c902e0a),
	.w3(32'h3c0538bf),
	.w4(32'h3ced13ce),
	.w5(32'h3c90fd2c),
	.w6(32'h3b0449de),
	.w7(32'h3c1e64b4),
	.w8(32'h3a821658),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf05899),
	.w1(32'hbbda7911),
	.w2(32'hbc17ac1d),
	.w3(32'h3b0d6f63),
	.w4(32'hbbcb522b),
	.w5(32'hbc25fccf),
	.w6(32'hbba28072),
	.w7(32'hbb101afa),
	.w8(32'hbb3dfb95),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78ee36),
	.w1(32'hba4b7724),
	.w2(32'hbc6125d8),
	.w3(32'h3cf20e41),
	.w4(32'h3c980ee4),
	.w5(32'hbb72cad1),
	.w6(32'h3c97b51a),
	.w7(32'h3c27e42b),
	.w8(32'h3b1f79d5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aea59),
	.w1(32'h3b9bd5e7),
	.w2(32'h394c5648),
	.w3(32'h3b64d78d),
	.w4(32'h3c5fd914),
	.w5(32'h3b99c8bc),
	.w6(32'hbadfb725),
	.w7(32'h3c421448),
	.w8(32'hb8d66767),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a674e),
	.w1(32'hbb5888fa),
	.w2(32'h3b0d48af),
	.w3(32'h39d23179),
	.w4(32'h3aa86b0d),
	.w5(32'h3b78e40e),
	.w6(32'h3a7ad292),
	.w7(32'h3bcb2cbe),
	.w8(32'h3bc8bd50),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b9d90),
	.w1(32'h3b3fbe8d),
	.w2(32'h3ae738ac),
	.w3(32'h3b3238e1),
	.w4(32'h3a8a896c),
	.w5(32'h3ad6c9d9),
	.w6(32'h3acbbccc),
	.w7(32'h3b3ea983),
	.w8(32'h3b836328),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3181f8),
	.w1(32'h3b183854),
	.w2(32'h3b0174a3),
	.w3(32'hb8727f1e),
	.w4(32'h3b502851),
	.w5(32'h3a47c8d1),
	.w6(32'h3a23d4e5),
	.w7(32'h3b4d5fe1),
	.w8(32'hbb0c2c9d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2946a0),
	.w1(32'h3c8657ad),
	.w2(32'h3c25c294),
	.w3(32'h3cb0ff0a),
	.w4(32'h3ccbd4cc),
	.w5(32'h3c89480e),
	.w6(32'h3af409ab),
	.w7(32'h3adee880),
	.w8(32'h3bd4730b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34843a),
	.w1(32'hb92d6d86),
	.w2(32'hbb581147),
	.w3(32'h3b2355ce),
	.w4(32'h3b97b582),
	.w5(32'h3a405e9a),
	.w6(32'h3ba34650),
	.w7(32'h3b8170ae),
	.w8(32'h3a2c1960),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71dbc7),
	.w1(32'h3a9229e3),
	.w2(32'h3b3b6cd8),
	.w3(32'hb7896a9e),
	.w4(32'h3b098c16),
	.w5(32'h3b940201),
	.w6(32'hba565e4e),
	.w7(32'h3b2939e6),
	.w8(32'h3bb7d61a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09c12a),
	.w1(32'h3b914948),
	.w2(32'hbb1d3246),
	.w3(32'h3c18fda6),
	.w4(32'h3c168cd5),
	.w5(32'h3b90135f),
	.w6(32'h3be736c4),
	.w7(32'h3bc753c1),
	.w8(32'h3b43d317),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb519387),
	.w1(32'hba84809a),
	.w2(32'h3b9de1af),
	.w3(32'hba94feec),
	.w4(32'h3b51aee4),
	.w5(32'h3bdd9e80),
	.w6(32'h3b2cd33f),
	.w7(32'h3b7bec72),
	.w8(32'h3bcd22df),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcd161),
	.w1(32'h3bd96e72),
	.w2(32'h3be6cd93),
	.w3(32'h3bb193b5),
	.w4(32'h3c07745d),
	.w5(32'h3c095231),
	.w6(32'hbb9dbf87),
	.w7(32'hbbad7642),
	.w8(32'hba8c0af9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac615d7),
	.w1(32'h3b09aac0),
	.w2(32'h3b153ba8),
	.w3(32'h3ab25e2c),
	.w4(32'h3b1f7a39),
	.w5(32'h3acf62f5),
	.w6(32'h3a3e319b),
	.w7(32'h3aabe787),
	.w8(32'h3bbfc92c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31153d),
	.w1(32'h3c89a025),
	.w2(32'h3c051044),
	.w3(32'h3c9c5e8d),
	.w4(32'h3d2fc90c),
	.w5(32'h3cbf0507),
	.w6(32'h3c4e45d6),
	.w7(32'h3d1314ec),
	.w8(32'h3c312b6f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d2b56),
	.w1(32'h3a3f39b1),
	.w2(32'h3a0b45ba),
	.w3(32'h3a9040b0),
	.w4(32'h3a31cc64),
	.w5(32'h3951de57),
	.w6(32'h3a1ce3fc),
	.w7(32'hb9246562),
	.w8(32'hba71584b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc981e),
	.w1(32'h37eadff6),
	.w2(32'h3b2e6927),
	.w3(32'hba93e0dd),
	.w4(32'h3b837395),
	.w5(32'h3c1ae98d),
	.w6(32'h3b99f9e8),
	.w7(32'h3c2b7a7c),
	.w8(32'h3c486d49),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c6630),
	.w1(32'h3b4f9bdb),
	.w2(32'h3b5532ca),
	.w3(32'h3b464f1d),
	.w4(32'h3b77568e),
	.w5(32'h3b2b4174),
	.w6(32'h3b4771aa),
	.w7(32'h3b7c8849),
	.w8(32'h3b8b1030),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d734c),
	.w1(32'h3c369b80),
	.w2(32'h3bdbe8f0),
	.w3(32'h3c76c70e),
	.w4(32'h3c3597dd),
	.w5(32'h3c57ca5b),
	.w6(32'h3c0a81b9),
	.w7(32'h38277f46),
	.w8(32'h3c0d51cf),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4975d),
	.w1(32'h3a391206),
	.w2(32'h3a88ef03),
	.w3(32'h38ba446e),
	.w4(32'h3aba38b4),
	.w5(32'h3a841f39),
	.w6(32'hb9a370c7),
	.w7(32'h37a4e356),
	.w8(32'h391b5056),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac18eb),
	.w1(32'h3a1d8782),
	.w2(32'h3a3f1901),
	.w3(32'h3c0d8029),
	.w4(32'h3be1f74e),
	.w5(32'h3ae77e38),
	.w6(32'h3b31b51a),
	.w7(32'h3c161f20),
	.w8(32'h3bd60193),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eea352),
	.w1(32'h3a32fcbf),
	.w2(32'h3a5fef92),
	.w3(32'hb9b6a262),
	.w4(32'h3a106c09),
	.w5(32'h39bf9f74),
	.w6(32'h38865672),
	.w7(32'h3a0131e0),
	.w8(32'h3be3b1d5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44a9e4),
	.w1(32'h3c0a5dcf),
	.w2(32'hbab59370),
	.w3(32'h3cb96ec2),
	.w4(32'h3cd977e3),
	.w5(32'h3c463475),
	.w6(32'h3c1d67d5),
	.w7(32'h3c61433f),
	.w8(32'h3bd86293),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0cce6),
	.w1(32'h3c9342ff),
	.w2(32'hba37f928),
	.w3(32'h3c4e8c79),
	.w4(32'h3c3834ff),
	.w5(32'hbb25c3d4),
	.w6(32'h3bbe5f57),
	.w7(32'h3b638b40),
	.w8(32'hbbc5ee4b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bb5d8),
	.w1(32'hb8bb037f),
	.w2(32'hba3651ee),
	.w3(32'h3b9118c0),
	.w4(32'h3aa95a14),
	.w5(32'hb83b18b3),
	.w6(32'h3af56c01),
	.w7(32'h3ab58cbc),
	.w8(32'h39ffd084),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11b79c),
	.w1(32'h3a55ec05),
	.w2(32'hb9519319),
	.w3(32'hb8f5987f),
	.w4(32'h3accedfa),
	.w5(32'h3a8d32a9),
	.w6(32'h3af5b086),
	.w7(32'h3a165b33),
	.w8(32'hb8e73529),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb466ae9),
	.w1(32'h3a80dd5a),
	.w2(32'h3b19fb09),
	.w3(32'h39ae8647),
	.w4(32'h3b8b4f43),
	.w5(32'h3b98bf93),
	.w6(32'h3be02e96),
	.w7(32'h3c710c9f),
	.w8(32'h3c48ece3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6512),
	.w1(32'hbbac91b6),
	.w2(32'hbbf173a2),
	.w3(32'h3aafeccf),
	.w4(32'h3c4eb27c),
	.w5(32'h3c0e4388),
	.w6(32'hbbf11297),
	.w7(32'h3b2d822b),
	.w8(32'h3c214a9c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a8f6c),
	.w1(32'h3c28a79c),
	.w2(32'h3d06b25d),
	.w3(32'h3d208bab),
	.w4(32'h3c26008b),
	.w5(32'h3ce6fe43),
	.w6(32'h3c6ac2b0),
	.w7(32'h389883e1),
	.w8(32'h3c76c6a5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a2ddb),
	.w1(32'h3cc48694),
	.w2(32'h3bd9705a),
	.w3(32'h3d05df43),
	.w4(32'h3d3e990e),
	.w5(32'h3cd98d8c),
	.w6(32'h3c2e7d54),
	.w7(32'h3cc8995b),
	.w8(32'h3c8f8d7b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb7763),
	.w1(32'h3b9a8e04),
	.w2(32'h3a7f937a),
	.w3(32'h3c3e5160),
	.w4(32'h3c4dde36),
	.w5(32'h3b64e6c9),
	.w6(32'hb9862996),
	.w7(32'h3c8ce974),
	.w8(32'h3ca5e196),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0363c8),
	.w1(32'hbac62a45),
	.w2(32'hba8d24c3),
	.w3(32'h39e8bc03),
	.w4(32'hbb46a374),
	.w5(32'hbad55011),
	.w6(32'hba21c0ae),
	.w7(32'h3a98d7ae),
	.w8(32'hba4cd1a6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a509905),
	.w1(32'h3a7add3b),
	.w2(32'h37b1249a),
	.w3(32'h3a8b3574),
	.w4(32'h3a4b4395),
	.w5(32'hb954bcd8),
	.w6(32'hba0f9aa1),
	.w7(32'hba314d60),
	.w8(32'hba167df8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba612d33),
	.w1(32'hbb24c4d1),
	.w2(32'hbaef2a1d),
	.w3(32'hbb0f6d04),
	.w4(32'hbb5077bd),
	.w5(32'hbb310b51),
	.w6(32'hbb698fbc),
	.w7(32'hbb27e5c9),
	.w8(32'h3b5b8600),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17c1ab),
	.w1(32'h38b93061),
	.w2(32'h3b64982b),
	.w3(32'h3a49c446),
	.w4(32'h3ae26b8f),
	.w5(32'h3b5bb047),
	.w6(32'h3a903056),
	.w7(32'h3c205d5d),
	.w8(32'h3c4462df),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19031b),
	.w1(32'h3b5be112),
	.w2(32'h3bac6392),
	.w3(32'h3b81a988),
	.w4(32'h3bb199d2),
	.w5(32'h3be87081),
	.w6(32'h39b73a04),
	.w7(32'h3bde67f7),
	.w8(32'h3be21661),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd225f),
	.w1(32'h3a32d72d),
	.w2(32'h3a901fdd),
	.w3(32'h3a78e5d6),
	.w4(32'hba734e10),
	.w5(32'hba9eeac7),
	.w6(32'h39fe6ce4),
	.w7(32'hb952db2b),
	.w8(32'h3b823241),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a053406),
	.w1(32'hbc082a75),
	.w2(32'h3ad0fd8c),
	.w3(32'h3bcfa29c),
	.w4(32'hbb5b938a),
	.w5(32'hbaab0536),
	.w6(32'h3be6d38a),
	.w7(32'h3c08ea25),
	.w8(32'h3ae303a9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb260c8d),
	.w1(32'h3b2202b7),
	.w2(32'h3a95a1ef),
	.w3(32'h3b47c758),
	.w4(32'h3bf189b4),
	.w5(32'h3ba85f9a),
	.w6(32'h393c1ba5),
	.w7(32'h3a7b5a5d),
	.w8(32'h3c0ad9dd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc221851),
	.w1(32'hbc1126f5),
	.w2(32'hbbfa9af4),
	.w3(32'hbc6795c1),
	.w4(32'hbc48cde0),
	.w5(32'hbbdd1dbf),
	.w6(32'hbbb6fdf7),
	.w7(32'hbbdc150d),
	.w8(32'hbc2b69a1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fff6f),
	.w1(32'h3a1413f4),
	.w2(32'hba54f51e),
	.w3(32'hbb9e90cd),
	.w4(32'h3b251cb7),
	.w5(32'hba6bc776),
	.w6(32'hbc097d25),
	.w7(32'hbb70b9a6),
	.w8(32'hbb3cf881),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab21e18),
	.w1(32'h3baecaea),
	.w2(32'h3b275a4b),
	.w3(32'h3c63d306),
	.w4(32'h3c9de958),
	.w5(32'h3c0aeb70),
	.w6(32'h3be66e11),
	.w7(32'h3ca09ae8),
	.w8(32'h3c66df5a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62fa297),
	.w1(32'h39e88bff),
	.w2(32'h3939671d),
	.w3(32'h3aac0470),
	.w4(32'h3983df3b),
	.w5(32'hba365740),
	.w6(32'hb9a5bc74),
	.w7(32'h3a36db74),
	.w8(32'h3bbe5df6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d9098),
	.w1(32'h3a298da7),
	.w2(32'h39f58b95),
	.w3(32'h3b5c7700),
	.w4(32'h3a25db27),
	.w5(32'hb7b36076),
	.w6(32'h3aa18f83),
	.w7(32'h3af54e3d),
	.w8(32'h38d06635),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2e785),
	.w1(32'h39c0943a),
	.w2(32'hb8b8d6d2),
	.w3(32'h3a14a13a),
	.w4(32'h38897d04),
	.w5(32'hba22c231),
	.w6(32'hba03a101),
	.w7(32'hb994edc2),
	.w8(32'h3983688f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad83336),
	.w1(32'h3a983e04),
	.w2(32'h3acc8ba4),
	.w3(32'h3ac3a7c7),
	.w4(32'h3a712dc1),
	.w5(32'h3a9d7504),
	.w6(32'h3a159d74),
	.w7(32'h3aedec6a),
	.w8(32'h3a89d9ca),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5fffc),
	.w1(32'hbb1f090c),
	.w2(32'h39daf76c),
	.w3(32'hbbbdd98c),
	.w4(32'hbb34ba37),
	.w5(32'hb8833228),
	.w6(32'hbb07a941),
	.w7(32'hbb02e188),
	.w8(32'h3b59aebf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf109cf),
	.w1(32'h3c08629e),
	.w2(32'h3bf45e95),
	.w3(32'h3c03626c),
	.w4(32'h3bbed7dd),
	.w5(32'h3b90cc43),
	.w6(32'h3a8a7c4c),
	.w7(32'h3ac13ecb),
	.w8(32'h3aeb41a5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b0726),
	.w1(32'hbbd4e587),
	.w2(32'hbb5ed50d),
	.w3(32'hb8fab8cb),
	.w4(32'hbc05919c),
	.w5(32'hbbec07e0),
	.w6(32'h3bae8a1f),
	.w7(32'h3b0d9752),
	.w8(32'h3ad2d2f6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85244f),
	.w1(32'hbb68ff96),
	.w2(32'hba948c89),
	.w3(32'hbbae112e),
	.w4(32'hbc0b0b34),
	.w5(32'hbb7c3909),
	.w6(32'hbb01d8da),
	.w7(32'hbb4b3311),
	.w8(32'hbb4d7da5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04158a),
	.w1(32'h3c39c50f),
	.w2(32'h3ba9cc27),
	.w3(32'h3c42161a),
	.w4(32'h3cc6a75f),
	.w5(32'h3bf2212c),
	.w6(32'h3be5a984),
	.w7(32'h3ca5073f),
	.w8(32'hba2436ba),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ee2b6),
	.w1(32'hba61d2a1),
	.w2(32'hbbecbe0d),
	.w3(32'hbc8bfe61),
	.w4(32'h3ab21c27),
	.w5(32'h3ac6aa3d),
	.w6(32'hbc0e7580),
	.w7(32'h3b821df0),
	.w8(32'h3c0174b6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8031f1),
	.w1(32'hbbacccd0),
	.w2(32'h3c03a81a),
	.w3(32'hbc2777f8),
	.w4(32'hbc397496),
	.w5(32'hbbe4d943),
	.w6(32'hbba66208),
	.w7(32'hbb3de368),
	.w8(32'hbbabe252),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb5b6),
	.w1(32'hbb096884),
	.w2(32'h3b438bcb),
	.w3(32'hbc0402e6),
	.w4(32'hbba90899),
	.w5(32'hbb25d305),
	.w6(32'h39f51fed),
	.w7(32'hbb59062c),
	.w8(32'hbae4f8d8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc303ac6),
	.w1(32'hba016664),
	.w2(32'hbb0e2cc5),
	.w3(32'hb6e9dd3b),
	.w4(32'h3aad370d),
	.w5(32'hbbab5024),
	.w6(32'h3b92c4ca),
	.w7(32'hbb6596f5),
	.w8(32'h3c505127),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b989e47),
	.w1(32'hbc4c42db),
	.w2(32'h3c924556),
	.w3(32'hbcc2e23b),
	.w4(32'hbcb2c7a6),
	.w5(32'hbaba0d21),
	.w6(32'hbc6cec53),
	.w7(32'hbd20d7bd),
	.w8(32'hbc72ea53),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8843b2),
	.w1(32'h3c2d8e2f),
	.w2(32'h3a7a8941),
	.w3(32'h3c1c1c32),
	.w4(32'h3b14dd76),
	.w5(32'hbbe8b660),
	.w6(32'hbb1f4d6d),
	.w7(32'hbc313b12),
	.w8(32'h3cbbfd37),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0fe41f),
	.w1(32'hbc8753f4),
	.w2(32'hbd317b74),
	.w3(32'h3c1cd820),
	.w4(32'hbcbbe48d),
	.w5(32'hbd055363),
	.w6(32'hbc216900),
	.w7(32'hbcd74f62),
	.w8(32'hbc65ef6e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27e98a),
	.w1(32'h3b92cc3b),
	.w2(32'h3b970f47),
	.w3(32'hbba96c36),
	.w4(32'h3a9a3690),
	.w5(32'hba21f4ae),
	.w6(32'h3a784e92),
	.w7(32'h3a31fc37),
	.w8(32'hbb44b270),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f8e2),
	.w1(32'h3b2f6080),
	.w2(32'h3ba74ff0),
	.w3(32'hb9e54544),
	.w4(32'h3ba2b26f),
	.w5(32'h3b180d5b),
	.w6(32'h3b4f3de3),
	.w7(32'h3ba1179d),
	.w8(32'hbb96c78a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bbdd9),
	.w1(32'h3bd89264),
	.w2(32'h3c6b8cf4),
	.w3(32'hbb25e0a7),
	.w4(32'h3bb30f2b),
	.w5(32'h3b81d945),
	.w6(32'h3bf76b29),
	.w7(32'h3c0f66be),
	.w8(32'hb8fdb94e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba49801),
	.w1(32'hbaa14a34),
	.w2(32'hbc80abfe),
	.w3(32'hbcb0c02b),
	.w4(32'hbcce8b7c),
	.w5(32'hbc71f754),
	.w6(32'hbcb37fb3),
	.w7(32'hbb931c0b),
	.w8(32'h3c0690f9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85e559),
	.w1(32'h3b898820),
	.w2(32'hbc0a9a0d),
	.w3(32'h3c51b573),
	.w4(32'h3c709737),
	.w5(32'h3c007bee),
	.w6(32'h3b81477d),
	.w7(32'hba5593ea),
	.w8(32'hbc9a3da8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc964596),
	.w1(32'hbc0907df),
	.w2(32'hbc2a7d28),
	.w3(32'hbc54e42d),
	.w4(32'hbc5f690e),
	.w5(32'hbc0c69a4),
	.w6(32'hbc7e4275),
	.w7(32'hbc8055a6),
	.w8(32'h3c12ad2a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc004b7a),
	.w1(32'h3bf87a34),
	.w2(32'h3c981c20),
	.w3(32'h3c32e548),
	.w4(32'h3c36530b),
	.w5(32'h3c398223),
	.w6(32'h3ab9f325),
	.w7(32'h3b74ffe7),
	.w8(32'h3b9b12b2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba924c63),
	.w1(32'hbbc37dba),
	.w2(32'hbabfd033),
	.w3(32'hbc2a9c5b),
	.w4(32'hbc196df4),
	.w5(32'hbc1c41d2),
	.w6(32'hbc5f8c85),
	.w7(32'h3c20fc72),
	.w8(32'hbc73d7ad),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a9d26),
	.w1(32'h3b3473e0),
	.w2(32'h3c257558),
	.w3(32'h3ca19e70),
	.w4(32'hba71b65d),
	.w5(32'hbc74a3b7),
	.w6(32'hbc1039a8),
	.w7(32'hbba6556c),
	.w8(32'hbb09aa54),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56407f),
	.w1(32'h3ae11e9e),
	.w2(32'h3bdffebf),
	.w3(32'h3b528641),
	.w4(32'hbbcbc0e7),
	.w5(32'hbb8b2a36),
	.w6(32'hbbc5f9bd),
	.w7(32'hbb4dcc9d),
	.w8(32'hbbb1a194),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c9b24),
	.w1(32'hbb09c75b),
	.w2(32'hba27c2e4),
	.w3(32'hbc0e5794),
	.w4(32'hbc0c2182),
	.w5(32'h3b012d6e),
	.w6(32'hbc1adeff),
	.w7(32'hb9cf3fc0),
	.w8(32'hba8a2e93),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c102961),
	.w1(32'hb9d8b907),
	.w2(32'h3b367770),
	.w3(32'hbcdf06cf),
	.w4(32'hbb1e6506),
	.w5(32'hbb22e525),
	.w6(32'hbc9d6757),
	.w7(32'hbc3c7b76),
	.w8(32'hbb85e609),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc92fc),
	.w1(32'h3c181d97),
	.w2(32'h3c8c880a),
	.w3(32'hbc347b77),
	.w4(32'hbae063bf),
	.w5(32'hbb651338),
	.w6(32'h3b93e6e6),
	.w7(32'h3b9c7d3c),
	.w8(32'hbb84dc55),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd99502),
	.w1(32'h3bbd811d),
	.w2(32'h3c539f78),
	.w3(32'hbbe168f7),
	.w4(32'h3af22deb),
	.w5(32'h3c28ef99),
	.w6(32'h3bf828b5),
	.w7(32'h3bcdcf37),
	.w8(32'hbc9fb8a8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b99b5),
	.w1(32'h3bc0fcd4),
	.w2(32'h3baf28ce),
	.w3(32'h3b3824cc),
	.w4(32'h3b45fd06),
	.w5(32'hbc5c19de),
	.w6(32'hbb0bab35),
	.w7(32'h3c8d7cde),
	.w8(32'h3b9734aa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule