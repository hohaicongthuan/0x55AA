module layer_10_featuremap_38(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb9f76),
	.w1(32'hba750006),
	.w2(32'hbb1a5af4),
	.w3(32'h3b5b7af2),
	.w4(32'hbbdb6389),
	.w5(32'h39f47f54),
	.w6(32'hbc23602e),
	.w7(32'hbbe11857),
	.w8(32'h3b2bf003),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac2721),
	.w1(32'h3b8c70f6),
	.w2(32'hbb832c7a),
	.w3(32'h3b2e7f1c),
	.w4(32'h3c65971c),
	.w5(32'h3b1955b7),
	.w6(32'h3aed98cc),
	.w7(32'h3abf3d7e),
	.w8(32'h3ba84404),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc53b4),
	.w1(32'hbaa9f4eb),
	.w2(32'hba76d23c),
	.w3(32'h3c0625fc),
	.w4(32'hba997da2),
	.w5(32'h3bff9a83),
	.w6(32'hb99c12d3),
	.w7(32'hb885e274),
	.w8(32'h39ae84b7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e392),
	.w1(32'hbb372836),
	.w2(32'h3c317122),
	.w3(32'h3b92ce5b),
	.w4(32'h3aa58d0e),
	.w5(32'h3c05a7f7),
	.w6(32'h3afc6621),
	.w7(32'h3bb18b03),
	.w8(32'hbb40a177),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51ac84),
	.w1(32'h3b3ff657),
	.w2(32'h3b65590c),
	.w3(32'h3a41d2a4),
	.w4(32'h3b135d3c),
	.w5(32'h3bd5ce18),
	.w6(32'hbbab69b4),
	.w7(32'hbba2bfa1),
	.w8(32'h3b65a34e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c259a53),
	.w1(32'hbb81e25c),
	.w2(32'hbbe4f97c),
	.w3(32'h3b84b6e1),
	.w4(32'hbba17c02),
	.w5(32'h3a8e72d2),
	.w6(32'h3b3f5d75),
	.w7(32'hbbb6acf8),
	.w8(32'hbc1efce5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb52de5),
	.w1(32'hbba1d555),
	.w2(32'h3a7b154b),
	.w3(32'h3c863dc3),
	.w4(32'hbac48c2a),
	.w5(32'h3b35ba9d),
	.w6(32'h3bf7bf09),
	.w7(32'hbc0f5f6c),
	.w8(32'hbb98c2e3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3802dc),
	.w1(32'h3bd93224),
	.w2(32'hbadee994),
	.w3(32'h3c0b03d5),
	.w4(32'h3c1e861a),
	.w5(32'h3b414dfc),
	.w6(32'hbaf181af),
	.w7(32'hbb82af26),
	.w8(32'h3bac04b4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10bca0),
	.w1(32'h3c114eeb),
	.w2(32'hbb20a51e),
	.w3(32'h3b8348af),
	.w4(32'h3b93e1b7),
	.w5(32'hbaf9adc5),
	.w6(32'h3bd0b6cc),
	.w7(32'h3bbdfea0),
	.w8(32'h3afe6d80),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d453e),
	.w1(32'h3b9527de),
	.w2(32'hbb272864),
	.w3(32'hbad771cf),
	.w4(32'h3bc45821),
	.w5(32'hbc04a0bc),
	.w6(32'h3b75c362),
	.w7(32'h3bfb8e8b),
	.w8(32'hbc1b43b9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63f6d5),
	.w1(32'h3b100ebb),
	.w2(32'h3b1f154a),
	.w3(32'hbc82207e),
	.w4(32'hbbffe4ef),
	.w5(32'hbabf7fd9),
	.w6(32'hbc8594ff),
	.w7(32'hbc1f9dac),
	.w8(32'hba7ee541),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3dc39),
	.w1(32'h3bbab5c6),
	.w2(32'h3cc2a22f),
	.w3(32'h3be0f17b),
	.w4(32'h3b082c4c),
	.w5(32'h3d3259c3),
	.w6(32'h3bf134fe),
	.w7(32'h3b75db47),
	.w8(32'h3d3544a7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2b249d),
	.w1(32'h3d00eb9d),
	.w2(32'hbc70cd47),
	.w3(32'h3d83e162),
	.w4(32'h3d5780e3),
	.w5(32'hbc2e8b7a),
	.w6(32'h3d79f773),
	.w7(32'h3d4991d2),
	.w8(32'hbbbd1a4a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc100a72),
	.w1(32'hbc3ee3ba),
	.w2(32'hbc2cf589),
	.w3(32'hbc53a604),
	.w4(32'hbc30dfbe),
	.w5(32'hba9b15be),
	.w6(32'hbc6f8fd3),
	.w7(32'hbc319400),
	.w8(32'hbb0ecbff),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c1b0e),
	.w1(32'hbbc4be52),
	.w2(32'hbafd642c),
	.w3(32'h3acd2afa),
	.w4(32'hbbbc0632),
	.w5(32'hbaea2be2),
	.w6(32'h3bc4ae81),
	.w7(32'h3b198d65),
	.w8(32'h3b394a3c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f3299),
	.w1(32'h3b2dc445),
	.w2(32'hbacc8638),
	.w3(32'h3a541594),
	.w4(32'h39d362ab),
	.w5(32'hbc4fc955),
	.w6(32'h3a7c2130),
	.w7(32'h39249688),
	.w8(32'hbc3b1fd8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd82df7),
	.w1(32'hba840cc4),
	.w2(32'h392abccc),
	.w3(32'hbd001486),
	.w4(32'hbc9b439c),
	.w5(32'h3b28b20b),
	.w6(32'hbce63937),
	.w7(32'hbc8f9dec),
	.w8(32'h3b1542ad),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c278464),
	.w1(32'hbb0688cb),
	.w2(32'hbbe68fd3),
	.w3(32'h3bfd8bfd),
	.w4(32'h3aeb9629),
	.w5(32'hbba14ebe),
	.w6(32'h3be20f81),
	.w7(32'hba437234),
	.w8(32'hbbb7e4ce),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca2ae9),
	.w1(32'hbc3518aa),
	.w2(32'hbc25b1e4),
	.w3(32'hbc4448a7),
	.w4(32'hbc219ef8),
	.w5(32'hbadb9a83),
	.w6(32'hbc0e93cb),
	.w7(32'hbc37858c),
	.w8(32'h39af3a32),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed8c4),
	.w1(32'hbc4a18f2),
	.w2(32'h3c27be16),
	.w3(32'h3c0719d9),
	.w4(32'hbbead6b7),
	.w5(32'h3c006e03),
	.w6(32'h3b4eed9b),
	.w7(32'h3b93ef1e),
	.w8(32'h3c04c678),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10ba83),
	.w1(32'h3bb4f39a),
	.w2(32'hbafeb163),
	.w3(32'h3bfd4304),
	.w4(32'h3c2b7f91),
	.w5(32'hbabbd121),
	.w6(32'h3c1695be),
	.w7(32'h3bc2e2dc),
	.w8(32'hbab80ba8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0075c),
	.w1(32'h3a4e6c96),
	.w2(32'hbc0047e8),
	.w3(32'h3aa882ff),
	.w4(32'h37e86b1f),
	.w5(32'h3a093078),
	.w6(32'h3b8643e8),
	.w7(32'h3b080f90),
	.w8(32'hbbac72c3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0393),
	.w1(32'hbb62ce9a),
	.w2(32'hbca71495),
	.w3(32'h3c445e57),
	.w4(32'h3b7a6c47),
	.w5(32'hbaf8d58d),
	.w6(32'h3839623d),
	.w7(32'hba8680dd),
	.w8(32'hbc24ca41),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1f25f),
	.w1(32'hbc3f3e71),
	.w2(32'hbc0c0c62),
	.w3(32'h3c6a9699),
	.w4(32'h3b4289c4),
	.w5(32'hbb96e32e),
	.w6(32'h3b751e16),
	.w7(32'hbb8dca6b),
	.w8(32'hbbe388f1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc151597),
	.w1(32'hbc048cf1),
	.w2(32'hbb923481),
	.w3(32'hbc52936c),
	.w4(32'hbc0ab76f),
	.w5(32'h3844fe93),
	.w6(32'hbba596cf),
	.w7(32'hbc21fdb0),
	.w8(32'h3b1faeab),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf66339),
	.w1(32'h3b86aae8),
	.w2(32'hbb4c0933),
	.w3(32'h3a363399),
	.w4(32'h3a1b3e00),
	.w5(32'hbb74baa9),
	.w6(32'hbab5683d),
	.w7(32'hbab92bac),
	.w8(32'h3b54cc4e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd59d8),
	.w1(32'hbb8524d2),
	.w2(32'h399dbcff),
	.w3(32'hbaadec55),
	.w4(32'h3aba268d),
	.w5(32'h3943f096),
	.w6(32'h3b9c3f24),
	.w7(32'h3a89d087),
	.w8(32'h39d92b22),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e309f),
	.w1(32'h39b07f15),
	.w2(32'hba9e6e03),
	.w3(32'h3ad873b7),
	.w4(32'hb9522bd4),
	.w5(32'hbb1edd70),
	.w6(32'h3b969728),
	.w7(32'h3a864ed4),
	.w8(32'hbaeb4b81),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71e874),
	.w1(32'h3adfba7d),
	.w2(32'h391ae806),
	.w3(32'h39da00f1),
	.w4(32'h3ad017ee),
	.w5(32'h3b05153f),
	.w6(32'h3aa1d9dc),
	.w7(32'h3b1eb2dd),
	.w8(32'h3b11d49c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb051398),
	.w1(32'hbaf6de81),
	.w2(32'hba51c308),
	.w3(32'hba97b172),
	.w4(32'hbb376cc1),
	.w5(32'hbac95cad),
	.w6(32'h39ca3d61),
	.w7(32'hbac7dfde),
	.w8(32'hbb1690ee),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa1f14),
	.w1(32'h398d213b),
	.w2(32'h39b15d57),
	.w3(32'hba02a56a),
	.w4(32'hb9932fd7),
	.w5(32'h3acdd27b),
	.w6(32'hb9c34b47),
	.w7(32'h3826946b),
	.w8(32'h3a663942),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba022dee),
	.w1(32'hbb21513c),
	.w2(32'hbaf2feba),
	.w3(32'h3a5bfb46),
	.w4(32'hba1a27a1),
	.w5(32'h3aabb109),
	.w6(32'h3a50c33f),
	.w7(32'hba8d3ab2),
	.w8(32'h385f51d0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11bb01),
	.w1(32'hbb4bbeae),
	.w2(32'hbad66cf6),
	.w3(32'hbb21aab3),
	.w4(32'hbb50adb9),
	.w5(32'hbace2e99),
	.w6(32'hbabf0587),
	.w7(32'hbb531c7a),
	.w8(32'hbb02c7ad),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabda8a1),
	.w1(32'hbab86faa),
	.w2(32'hbacc0ead),
	.w3(32'hbaf07dc7),
	.w4(32'hbafc2614),
	.w5(32'hbaa61fd7),
	.w6(32'hbab873b5),
	.w7(32'hbacc371a),
	.w8(32'hbb2aa446),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25a7c0),
	.w1(32'h3b17bf70),
	.w2(32'hba8dfa2c),
	.w3(32'h3ae46a5e),
	.w4(32'h3b1937be),
	.w5(32'hba8ce5bb),
	.w6(32'h3b3b16d3),
	.w7(32'h3a465117),
	.w8(32'hba9fdcb7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b3a50),
	.w1(32'hbaa75438),
	.w2(32'hba797256),
	.w3(32'hba80cbde),
	.w4(32'hba48b041),
	.w5(32'hb90255aa),
	.w6(32'hbaaabb13),
	.w7(32'hbabe16ab),
	.w8(32'hba7676d3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fda14),
	.w1(32'h3adc1900),
	.w2(32'hbac22a34),
	.w3(32'hbb1c927f),
	.w4(32'h3afedd36),
	.w5(32'h3a9d3451),
	.w6(32'hbb8dba8a),
	.w7(32'hbaac65c8),
	.w8(32'h3b2d7193),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2c07b),
	.w1(32'h3a9ba57d),
	.w2(32'h3b991b3a),
	.w3(32'h3a84007b),
	.w4(32'h3ad3c321),
	.w5(32'h3b4a32ee),
	.w6(32'h3b043a84),
	.w7(32'h3b5a9f14),
	.w8(32'h3b5fad5b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a39d9),
	.w1(32'h38f66b55),
	.w2(32'h3ac4bddc),
	.w3(32'h3b394f96),
	.w4(32'hba90379f),
	.w5(32'h3adf7b6a),
	.w6(32'h3b7143d3),
	.w7(32'h39cd35fb),
	.w8(32'h3b18d21d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3858d2db),
	.w1(32'hba83e13d),
	.w2(32'h3a8c57fe),
	.w3(32'hba810bb2),
	.w4(32'hbb1a644e),
	.w5(32'h3b03a577),
	.w6(32'hb9bbfc2d),
	.w7(32'hbb092625),
	.w8(32'h3a885944),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b806985),
	.w1(32'h3a56337a),
	.w2(32'hb99dded8),
	.w3(32'h3b7e7ab6),
	.w4(32'h3a5bbf15),
	.w5(32'hbaf987d3),
	.w6(32'h3b801986),
	.w7(32'h39f85aee),
	.w8(32'hbacbd69f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dac0a7),
	.w1(32'h39bb7be9),
	.w2(32'h3b58b7fe),
	.w3(32'hb9d8f0d3),
	.w4(32'hbaa318eb),
	.w5(32'h39f499c3),
	.w6(32'hb99f04f5),
	.w7(32'hba66478d),
	.w8(32'h38e57119),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b1fd6),
	.w1(32'hb97e3899),
	.w2(32'hba7cf6f3),
	.w3(32'hba85d611),
	.w4(32'h3926c0d0),
	.w5(32'hba85b88d),
	.w6(32'h39df2d0b),
	.w7(32'h3b0931d5),
	.w8(32'hba7fd5ab),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a3509),
	.w1(32'hba972638),
	.w2(32'hbbcb21ac),
	.w3(32'h3b2b0bb5),
	.w4(32'h393cb4e2),
	.w5(32'hbb8cafcb),
	.w6(32'h3ac9012a),
	.w7(32'hbad5b1c3),
	.w8(32'hbbb393e3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb252688),
	.w1(32'hba91b38e),
	.w2(32'hbb58b7fb),
	.w3(32'hbab97f31),
	.w4(32'hbade6125),
	.w5(32'hbaca62ba),
	.w6(32'hbad8a2b1),
	.w7(32'hbb0f7ed4),
	.w8(32'hbb46a387),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70718b7),
	.w1(32'hb749c05e),
	.w2(32'hbb256397),
	.w3(32'h3936309b),
	.w4(32'h3a91f780),
	.w5(32'hb9d1d76a),
	.w6(32'hba15b72c),
	.w7(32'h3a40bbed),
	.w8(32'hba975384),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7fea1),
	.w1(32'hbb1d575d),
	.w2(32'hbb9f658e),
	.w3(32'hbb293515),
	.w4(32'hba07f45a),
	.w5(32'hbbb955fa),
	.w6(32'hbb2220a4),
	.w7(32'hba5f1433),
	.w8(32'hbbd89fc2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa05cf7),
	.w1(32'hbafc1703),
	.w2(32'hbb9ffaf5),
	.w3(32'h3af2ba67),
	.w4(32'h39e6f1cb),
	.w5(32'hbb4385ac),
	.w6(32'hba12ce5c),
	.w7(32'hbb1bbd80),
	.w8(32'hbb8405f7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398907b9),
	.w1(32'hb888bfdb),
	.w2(32'hbb1e7dc6),
	.w3(32'h3a38f6e8),
	.w4(32'h3a1b6639),
	.w5(32'hbb15c1c8),
	.w6(32'h3a051a53),
	.w7(32'h39cff3f1),
	.w8(32'hbb14e02c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24f301),
	.w1(32'hbb2cc06c),
	.w2(32'hbb0596e2),
	.w3(32'hbaa618ac),
	.w4(32'hbac861d5),
	.w5(32'hbbc0e6e4),
	.w6(32'hbb46bcbb),
	.w7(32'hbb462486),
	.w8(32'hbb928b38),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a58d),
	.w1(32'hba3304f5),
	.w2(32'hbacc7c6f),
	.w3(32'hbb2efeb3),
	.w4(32'hbb6a9560),
	.w5(32'hba2756bf),
	.w6(32'hbb8180c5),
	.w7(32'hbb71c563),
	.w8(32'hba0dfa65),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5a52b),
	.w1(32'hbb36d524),
	.w2(32'hbac15909),
	.w3(32'h3a29a813),
	.w4(32'hba95b46e),
	.w5(32'hbb1e1900),
	.w6(32'h3aa73707),
	.w7(32'h398744d1),
	.w8(32'hbb94b2d5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacff21c),
	.w1(32'hba069211),
	.w2(32'h3a8b10d0),
	.w3(32'hbb2256c6),
	.w4(32'hbaa6d34d),
	.w5(32'hb8fca17a),
	.w6(32'hbb9acfa0),
	.w7(32'hbb66b37c),
	.w8(32'h39958be6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387410ea),
	.w1(32'hbb3d94f2),
	.w2(32'hbbb4e344),
	.w3(32'h3aada286),
	.w4(32'hb914ff0f),
	.w5(32'hbb966342),
	.w6(32'hb9611bf1),
	.w7(32'hba20f365),
	.w8(32'hbb8d84c8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94c754),
	.w1(32'h39ea15d7),
	.w2(32'hbab71de9),
	.w3(32'hba7bff87),
	.w4(32'h3ab62379),
	.w5(32'h39fd56da),
	.w6(32'hbad5ed40),
	.w7(32'h38eba303),
	.w8(32'hb9813dba),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9560ff3),
	.w1(32'h3aa4618b),
	.w2(32'hbb7053bf),
	.w3(32'hb9b93083),
	.w4(32'hb941361b),
	.w5(32'hbb4d6399),
	.w6(32'h3a630146),
	.w7(32'h38c44632),
	.w8(32'hbb05e891),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a5102),
	.w1(32'hbb0700df),
	.w2(32'hbaa7f120),
	.w3(32'hbb6f5210),
	.w4(32'hbb173f39),
	.w5(32'hbafa9859),
	.w6(32'hbb83eea3),
	.w7(32'hbab4c9ce),
	.w8(32'hbaeff489),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac5725),
	.w1(32'h3a611632),
	.w2(32'h39d46154),
	.w3(32'h3a252c6d),
	.w4(32'h39216977),
	.w5(32'h383163f7),
	.w6(32'h3a42e304),
	.w7(32'h398a0831),
	.w8(32'hb9fbdba5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b6e8b),
	.w1(32'h395ced15),
	.w2(32'h3a3a0916),
	.w3(32'hb8df2ee8),
	.w4(32'hb9b4a9d7),
	.w5(32'hb9fc0e33),
	.w6(32'h3a0a2f94),
	.w7(32'hb94eb151),
	.w8(32'hb9337932),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a1551),
	.w1(32'h3976cd9f),
	.w2(32'hba93a54c),
	.w3(32'h381f3204),
	.w4(32'hba5cf152),
	.w5(32'hbae790af),
	.w6(32'h3a88ddd1),
	.w7(32'h393e9fb2),
	.w8(32'hbaf323e6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa472e4),
	.w1(32'hba11fbcd),
	.w2(32'hbb02ab10),
	.w3(32'hb986cc6f),
	.w4(32'hbaec89c1),
	.w5(32'hb67d747d),
	.w6(32'hb832a904),
	.w7(32'hbae50abf),
	.w8(32'hbab4ea3d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae1aca),
	.w1(32'hb984f06a),
	.w2(32'hb86d03db),
	.w3(32'hb983ee14),
	.w4(32'h3adc2e62),
	.w5(32'h3a07f08a),
	.w6(32'h3a39a0f8),
	.w7(32'h3b319c04),
	.w8(32'h3a94f77e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8239ed),
	.w1(32'h3a291e5a),
	.w2(32'h3a853932),
	.w3(32'h3ab1d82b),
	.w4(32'h3a6794da),
	.w5(32'h3a13f0d8),
	.w6(32'h3b319d71),
	.w7(32'h3b4b999e),
	.w8(32'h3ac4d675),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca54a0),
	.w1(32'h3a6166b1),
	.w2(32'hbb2899c7),
	.w3(32'hba35a70b),
	.w4(32'h3a1bea74),
	.w5(32'hbb34fff9),
	.w6(32'h3a057be7),
	.w7(32'h3a47eb7e),
	.w8(32'hbb12f361),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade60b7),
	.w1(32'hba726599),
	.w2(32'hba5ea309),
	.w3(32'hb9cbc145),
	.w4(32'h38a0ff0a),
	.w5(32'hba8bd242),
	.w6(32'hba6229df),
	.w7(32'hb952faaa),
	.w8(32'hba838774),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18a4e2),
	.w1(32'h3a1469b6),
	.w2(32'hbaa1fce6),
	.w3(32'h39541369),
	.w4(32'h39d329c5),
	.w5(32'hbabe9288),
	.w6(32'h38ec71c6),
	.w7(32'h38b33af7),
	.w8(32'hba8fc9d2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b261b12),
	.w1(32'hba6bfad5),
	.w2(32'hbbaf5b0b),
	.w3(32'h3b493d9e),
	.w4(32'hb91b0132),
	.w5(32'hbbbbff02),
	.w6(32'h3b3c23ef),
	.w7(32'h3b0b5d6f),
	.w8(32'hbbb2a76d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94de35c),
	.w1(32'hbb2b2847),
	.w2(32'hbb7e2eb7),
	.w3(32'h38f6727e),
	.w4(32'hba460525),
	.w5(32'hbb5c35db),
	.w6(32'hba8b5ef9),
	.w7(32'hbb878118),
	.w8(32'hbbcf4c84),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384bbe83),
	.w1(32'hbaef2c93),
	.w2(32'h3a9ddf97),
	.w3(32'hb9fb6b36),
	.w4(32'hbb02ccfd),
	.w5(32'h3b29683d),
	.w6(32'hbad3fabe),
	.w7(32'hbb494c11),
	.w8(32'h3ad126ad),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e57df),
	.w1(32'hba296f64),
	.w2(32'hbb030282),
	.w3(32'hba32bed2),
	.w4(32'hba89e7d3),
	.w5(32'hbb25d417),
	.w6(32'h3a6130a0),
	.w7(32'hba131ef5),
	.w8(32'hbb40ea3c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78d90e),
	.w1(32'h3a66491f),
	.w2(32'h39d8bebe),
	.w3(32'h3a290171),
	.w4(32'hb9f56d92),
	.w5(32'h39122b0f),
	.w6(32'h391fad19),
	.w7(32'hb99ff867),
	.w8(32'h39db7499),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a298b28),
	.w1(32'h3a814088),
	.w2(32'h3a6539af),
	.w3(32'h3a023861),
	.w4(32'h3a4781b4),
	.w5(32'h3b183b05),
	.w6(32'h37b0e171),
	.w7(32'h39c878c6),
	.w8(32'h3b32154a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addd3fb),
	.w1(32'hba1e13f0),
	.w2(32'hbb4699d3),
	.w3(32'h3b48e705),
	.w4(32'h39831cbc),
	.w5(32'hbb3c9f65),
	.w6(32'h3b9a1289),
	.w7(32'h39182144),
	.w8(32'hbb59b4a9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a035784),
	.w1(32'h3b865bdc),
	.w2(32'h3a0ce99b),
	.w3(32'h391941bc),
	.w4(32'h3bb20d88),
	.w5(32'h39c7414b),
	.w6(32'hbab64614),
	.w7(32'h3b896407),
	.w8(32'hb95975dc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a5419),
	.w1(32'h3a807c40),
	.w2(32'h3a24142d),
	.w3(32'h3a000848),
	.w4(32'h3aa7bebd),
	.w5(32'h396c58e7),
	.w6(32'h39c8809e),
	.w7(32'h3a7ebde1),
	.w8(32'h38d570a4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20bcd9),
	.w1(32'h384f955b),
	.w2(32'hbb613600),
	.w3(32'h39c9ac43),
	.w4(32'h3a1b69c4),
	.w5(32'hbb5d9f8d),
	.w6(32'h38c572f1),
	.w7(32'h3a42a9f7),
	.w8(32'hbb1b34c6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2757ae),
	.w1(32'hbb28839d),
	.w2(32'hbbcc7f05),
	.w3(32'hbb423974),
	.w4(32'hba152458),
	.w5(32'hbbaa374e),
	.w6(32'hbab50898),
	.w7(32'hbb671f8e),
	.w8(32'hbb42919a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5130e2),
	.w1(32'hbbaa70ef),
	.w2(32'hbb6da4f3),
	.w3(32'hbb88143c),
	.w4(32'hbba3353d),
	.w5(32'hbb9b9b80),
	.w6(32'hbb1568bd),
	.w7(32'hbbc26d00),
	.w8(32'hbba1ccf8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76d634),
	.w1(32'hbadad63e),
	.w2(32'hba0fda0a),
	.w3(32'h39ea102d),
	.w4(32'hbb1993e0),
	.w5(32'hb9b51633),
	.w6(32'h3aa7d4e2),
	.w7(32'hbb1b7889),
	.w8(32'hba33d4bc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d932f),
	.w1(32'h39bd873b),
	.w2(32'hbafff426),
	.w3(32'h3b2fb090),
	.w4(32'h39a9fe55),
	.w5(32'hbb1cbd8a),
	.w6(32'h3b41a2dc),
	.w7(32'h3ab4688a),
	.w8(32'hbaf7fe36),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c15b09),
	.w1(32'hb9900c0b),
	.w2(32'hbaa1343e),
	.w3(32'hba134249),
	.w4(32'hba6eb18d),
	.w5(32'hbafdd1bd),
	.w6(32'hba1a7d4f),
	.w7(32'hba924f8b),
	.w8(32'hbac3e0f8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47af1),
	.w1(32'h390dd41f),
	.w2(32'hba820116),
	.w3(32'h3a367024),
	.w4(32'hb83d502f),
	.w5(32'hb9dce4b1),
	.w6(32'h3a0b9869),
	.w7(32'hb90b459b),
	.w8(32'hba69f686),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc24eb),
	.w1(32'hb95cd96f),
	.w2(32'hbb2a148f),
	.w3(32'h3a5964f5),
	.w4(32'h394da5b5),
	.w5(32'hbb4513e3),
	.w6(32'h3a938e4e),
	.w7(32'h3a78f345),
	.w8(32'hbb1ab8ac),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25d4dd),
	.w1(32'hbad14db4),
	.w2(32'h3b27f53a),
	.w3(32'hba97a403),
	.w4(32'hbb281ba1),
	.w5(32'h3b4d7bc2),
	.w6(32'hba3bc225),
	.w7(32'hbae91640),
	.w8(32'h3b7bb208),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd528f),
	.w1(32'h3ab6a2d3),
	.w2(32'hbaa49789),
	.w3(32'h3ac6ae76),
	.w4(32'h3a7e8a48),
	.w5(32'hba560f05),
	.w6(32'h3b8132f8),
	.w7(32'h3b2e3edc),
	.w8(32'h3a31303d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08241a),
	.w1(32'hb90679a0),
	.w2(32'hb9419cfc),
	.w3(32'h3a129143),
	.w4(32'h3a82ef51),
	.w5(32'hb9979ecd),
	.w6(32'h3a1a8e31),
	.w7(32'h3aea2725),
	.w8(32'h38a20e26),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccb2f0),
	.w1(32'hba4275ae),
	.w2(32'hba86017e),
	.w3(32'hb937a071),
	.w4(32'hb8fd0ab4),
	.w5(32'h39f20235),
	.w6(32'h3a3fccd0),
	.w7(32'h3935fe8e),
	.w8(32'h38bb49e9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42ab15),
	.w1(32'h3a8a0e4f),
	.w2(32'hb78a03b4),
	.w3(32'h3a39f7eb),
	.w4(32'h3a867164),
	.w5(32'hbb213507),
	.w6(32'h3a4f1587),
	.w7(32'h3a8dad43),
	.w8(32'hbb089287),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e500e),
	.w1(32'hb9629c47),
	.w2(32'h3a605368),
	.w3(32'hbb658201),
	.w4(32'hbb6aa66f),
	.w5(32'h3a41493c),
	.w6(32'hbb97fdc7),
	.w7(32'hbb4fc8bd),
	.w8(32'h3a5687d2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8afcdb),
	.w1(32'hba0519dd),
	.w2(32'hba1248c5),
	.w3(32'h3b0e2b37),
	.w4(32'h3b07f411),
	.w5(32'hba2b0e49),
	.w6(32'h3a073fb6),
	.w7(32'h38dbe46a),
	.w8(32'hb9fa5513),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f0ea6),
	.w1(32'h3ab07ace),
	.w2(32'h3b1eafa5),
	.w3(32'h39aa24af),
	.w4(32'h3aab1a46),
	.w5(32'h3b0b752e),
	.w6(32'h3ae457f3),
	.w7(32'h3b12fc25),
	.w8(32'h3b0f1bfb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8dc0a),
	.w1(32'h3a807005),
	.w2(32'hbb15d61a),
	.w3(32'h3a330c39),
	.w4(32'hba9c3e54),
	.w5(32'hbaca6f89),
	.w6(32'h3a311f24),
	.w7(32'hba232d78),
	.w8(32'hbb3da1de),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadf602),
	.w1(32'h3b041ec8),
	.w2(32'h3a7fbf42),
	.w3(32'h3a09cec3),
	.w4(32'h3aaad7af),
	.w5(32'h398e1568),
	.w6(32'hba0fd2ae),
	.w7(32'h3a0d2c77),
	.w8(32'hb96c2df0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ef4cd),
	.w1(32'hbad489ae),
	.w2(32'hbbce229d),
	.w3(32'h3a68e2fa),
	.w4(32'hba520c88),
	.w5(32'hbbd4ca8a),
	.w6(32'h3a117913),
	.w7(32'hb9877fcf),
	.w8(32'hbbd5a742),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba379608),
	.w1(32'hbb0fac1d),
	.w2(32'hbb579c4c),
	.w3(32'hba4012e8),
	.w4(32'hbb7093c3),
	.w5(32'hbb03ada6),
	.w6(32'hbb39225a),
	.w7(32'hbb60f5cf),
	.w8(32'hbac826fe),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e12e8),
	.w1(32'hbb55ccca),
	.w2(32'hb98e7313),
	.w3(32'hb8f0c45f),
	.w4(32'hbb307b2c),
	.w5(32'hba7b7278),
	.w6(32'hb8686747),
	.w7(32'hbb49a7d6),
	.w8(32'hb9411199),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6658ac),
	.w1(32'hb9af5986),
	.w2(32'h3ba6f00a),
	.w3(32'h3a356dfc),
	.w4(32'h3a4d73e7),
	.w5(32'h3ba14afc),
	.w6(32'h39e0c2ca),
	.w7(32'h3ab4fad5),
	.w8(32'h3bbc4b8c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f2d70),
	.w1(32'h3a2c737e),
	.w2(32'hbb977e42),
	.w3(32'h3b082004),
	.w4(32'h3b334645),
	.w5(32'hbb1fb803),
	.w6(32'h3b8e99c4),
	.w7(32'h3abc7e75),
	.w8(32'hbb1cd146),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e7af7),
	.w1(32'h3a16f2d8),
	.w2(32'h3ab3f5ae),
	.w3(32'h3a4a34a0),
	.w4(32'h3a862c01),
	.w5(32'hb98b5df1),
	.w6(32'h3a8d7018),
	.w7(32'h3adcdeee),
	.w8(32'hba5530d2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a45b82),
	.w1(32'h3b806df0),
	.w2(32'h3ab6788d),
	.w3(32'hb9dc1ed3),
	.w4(32'h3b94b439),
	.w5(32'h3c003f70),
	.w6(32'hba91938c),
	.w7(32'h3b126004),
	.w8(32'h3bb73bae),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997b5d),
	.w1(32'h39c8fec9),
	.w2(32'h3a42fa7f),
	.w3(32'hbac50058),
	.w4(32'h3b39994a),
	.w5(32'h3b3ea0b4),
	.w6(32'h3a056076),
	.w7(32'h3b293ae9),
	.w8(32'h3b15a2b3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31d81b),
	.w1(32'hbb0d4740),
	.w2(32'hbae053a3),
	.w3(32'h3a14ab44),
	.w4(32'hba3d4ab9),
	.w5(32'hbb3c7012),
	.w6(32'h3a29ece8),
	.w7(32'hbb41dd2e),
	.w8(32'hbb1c5ba4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac070d0),
	.w1(32'hb96bc9ad),
	.w2(32'hbb0f6b1c),
	.w3(32'hbaec1655),
	.w4(32'h3861cdcf),
	.w5(32'h3a1d2cc0),
	.w6(32'h3a06c6c8),
	.w7(32'h3ad089bc),
	.w8(32'h3a7c718f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f15e90),
	.w1(32'h380f6a72),
	.w2(32'hba939fe6),
	.w3(32'h397b471b),
	.w4(32'h3a3dd239),
	.w5(32'hba165cd9),
	.w6(32'hb9f5e085),
	.w7(32'h3a75fae3),
	.w8(32'hba4f51ef),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a0630),
	.w1(32'hba2c336f),
	.w2(32'hbb963311),
	.w3(32'hbb4a3a0e),
	.w4(32'hbab033df),
	.w5(32'h3a42c55a),
	.w6(32'hbb9486ed),
	.w7(32'hbb0f3770),
	.w8(32'h3b0b12c3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed66ad),
	.w1(32'h398b8cec),
	.w2(32'hbb3ca0ca),
	.w3(32'hba87c1f2),
	.w4(32'hbaafeee0),
	.w5(32'hbafa5f6c),
	.w6(32'h3962a120),
	.w7(32'hb9927539),
	.w8(32'hbaeac983),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5be653),
	.w1(32'hb9a22bf7),
	.w2(32'hb864dbee),
	.w3(32'hba836c3b),
	.w4(32'hb95570c3),
	.w5(32'hba1a20ae),
	.w6(32'hba7611aa),
	.w7(32'hb9cdb0d3),
	.w8(32'hba949a13),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c4836),
	.w1(32'hba89babd),
	.w2(32'hb6e35590),
	.w3(32'hba721310),
	.w4(32'hba9c01e1),
	.w5(32'h3ac0fdd5),
	.w6(32'hbaa0ff91),
	.w7(32'hbab5f495),
	.w8(32'h3aff52e2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a28c2),
	.w1(32'h39253371),
	.w2(32'hbb0f5500),
	.w3(32'hba770f68),
	.w4(32'hba3289b2),
	.w5(32'hbae95d98),
	.w6(32'h3a6743d6),
	.w7(32'hbb10b481),
	.w8(32'hbb378e26),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a293a4a),
	.w1(32'hba96d5df),
	.w2(32'h3b58a768),
	.w3(32'h3ac897db),
	.w4(32'hba6a1fcc),
	.w5(32'h3a33ecaf),
	.w6(32'h3a9356a7),
	.w7(32'hbad5ec28),
	.w8(32'h3aa75a0b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27b404),
	.w1(32'h3b822d0a),
	.w2(32'hb8fe5fb9),
	.w3(32'h3b0e42a9),
	.w4(32'h3af6f8fb),
	.w5(32'hb97ccddd),
	.w6(32'h3b70b07d),
	.w7(32'h3bbf0801),
	.w8(32'h39d6af7d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d7b76),
	.w1(32'h3aa4a8c2),
	.w2(32'h3a180bbe),
	.w3(32'hba50c29e),
	.w4(32'h3b14ac4b),
	.w5(32'hb961f14f),
	.w6(32'h39031d16),
	.w7(32'h3ab4da1b),
	.w8(32'hb92aef98),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b552a17),
	.w1(32'h3b2dcd7a),
	.w2(32'h3a4c778e),
	.w3(32'h3b12d44f),
	.w4(32'h3b33c679),
	.w5(32'h3b0b5547),
	.w6(32'h3b70dafa),
	.w7(32'h3a4c5de9),
	.w8(32'h3a638973),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eac486),
	.w1(32'hbb52f4cd),
	.w2(32'hbb4a7d6f),
	.w3(32'hba95389b),
	.w4(32'hbb3fd583),
	.w5(32'hba4809bd),
	.w6(32'hb9862833),
	.w7(32'hbae1b954),
	.w8(32'hba9aa2cd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7ded7),
	.w1(32'h3b1dcc58),
	.w2(32'hb9c55d58),
	.w3(32'h3ae67fb9),
	.w4(32'h3aa4036a),
	.w5(32'hba5daf51),
	.w6(32'h3b0dead8),
	.w7(32'h3a9a464e),
	.w8(32'hba981e51),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377bf6c3),
	.w1(32'h387de22e),
	.w2(32'hba51d313),
	.w3(32'hb98c0b04),
	.w4(32'h37122590),
	.w5(32'hbad333a8),
	.w6(32'hb93413c3),
	.w7(32'hb9a0a335),
	.w8(32'hbac13760),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe8efc),
	.w1(32'h39f341df),
	.w2(32'h3a0c416e),
	.w3(32'h39976de7),
	.w4(32'h3a143152),
	.w5(32'h38c1318e),
	.w6(32'hb86f9e51),
	.w7(32'h3a03decc),
	.w8(32'hb6e89421),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04cf47),
	.w1(32'h39970193),
	.w2(32'hb849939a),
	.w3(32'h38e9f5ec),
	.w4(32'hb940cc9f),
	.w5(32'h3a483e59),
	.w6(32'h3a72593b),
	.w7(32'h39f0efb5),
	.w8(32'h3a24761a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba197615),
	.w1(32'hba9b922c),
	.w2(32'hba44140a),
	.w3(32'h3a2488c9),
	.w4(32'hbaa24520),
	.w5(32'h39ec7e2d),
	.w6(32'h3ad13302),
	.w7(32'hba26078e),
	.w8(32'hb9933b92),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2de4bd),
	.w1(32'hb9859f6e),
	.w2(32'hb9cd678b),
	.w3(32'h3b240b22),
	.w4(32'h3aea1164),
	.w5(32'h3a0fa2df),
	.w6(32'h3a5f22f8),
	.w7(32'h3a3635fd),
	.w8(32'hb9b3f3fc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d40410),
	.w1(32'hba35937e),
	.w2(32'hb9dc6128),
	.w3(32'h3adb88c7),
	.w4(32'h39969203),
	.w5(32'hba05cbe6),
	.w6(32'h3b3a09c6),
	.w7(32'h3b06ec76),
	.w8(32'hba7fcc6d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a1860f),
	.w1(32'hba1aef6a),
	.w2(32'hb9ca724f),
	.w3(32'hb9db9844),
	.w4(32'hb9b534a8),
	.w5(32'hba36c377),
	.w6(32'hb9e13bb5),
	.w7(32'hba5d0a35),
	.w8(32'hba761412),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8c836),
	.w1(32'hbacba344),
	.w2(32'hbb58b864),
	.w3(32'hbad7437f),
	.w4(32'hbaee487d),
	.w5(32'hbb406f95),
	.w6(32'hb8bea593),
	.w7(32'hbaa92b1b),
	.w8(32'hbb256317),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad41c57),
	.w1(32'h39b1ff0d),
	.w2(32'hb897061e),
	.w3(32'h3b1cb4b6),
	.w4(32'h39f0b0d0),
	.w5(32'h398201d7),
	.w6(32'h3b367a63),
	.w7(32'h3ad8a0d6),
	.w8(32'h3a254836),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb8c67),
	.w1(32'h3ae0f7ac),
	.w2(32'hbb588eaf),
	.w3(32'h3ae48f08),
	.w4(32'h3adf770e),
	.w5(32'hbb2df576),
	.w6(32'h3b062b13),
	.w7(32'h3b055d17),
	.w8(32'hbb2c8d91),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb323472),
	.w1(32'hba8820db),
	.w2(32'h392a2d6a),
	.w3(32'hbb050484),
	.w4(32'hb9b9d9fe),
	.w5(32'h3a27c3bd),
	.w6(32'hbb08fc69),
	.w7(32'hbabe8efe),
	.w8(32'hb99c56da),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0697c),
	.w1(32'hb9354dbc),
	.w2(32'h39e3d7f9),
	.w3(32'hbaae2155),
	.w4(32'hb91135b9),
	.w5(32'h39adcf7d),
	.w6(32'hbb01fa23),
	.w7(32'hba8a97d0),
	.w8(32'hba094bfc),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aa786),
	.w1(32'h3a55fd79),
	.w2(32'hbb839bbd),
	.w3(32'hb98b6db6),
	.w4(32'h3adbaefc),
	.w5(32'hbb0446f1),
	.w6(32'hbaba1d82),
	.w7(32'hba86548a),
	.w8(32'hbb18acee),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa40c2d),
	.w1(32'hbb5ec3aa),
	.w2(32'hba965de0),
	.w3(32'hbb732b45),
	.w4(32'hbba4bd98),
	.w5(32'hbb0b4832),
	.w6(32'hbb4a0c34),
	.w7(32'hbb6292fc),
	.w8(32'hbb247bd1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28d136),
	.w1(32'h3a2bb61a),
	.w2(32'hb760b22e),
	.w3(32'h3b33a398),
	.w4(32'h3abb81ec),
	.w5(32'h3a4fed54),
	.w6(32'h3abdab00),
	.w7(32'h3b116a70),
	.w8(32'h3a9c1bb2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55d12c),
	.w1(32'h3b54f5ce),
	.w2(32'h3b1a0101),
	.w3(32'h3b8deb22),
	.w4(32'h3b94fbee),
	.w5(32'h3b354817),
	.w6(32'h3bb94364),
	.w7(32'h3baaea58),
	.w8(32'h3af55758),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8cc3e),
	.w1(32'h38c709ba),
	.w2(32'hbb0b90ff),
	.w3(32'h3b0ae710),
	.w4(32'h3b17eba2),
	.w5(32'hbad14145),
	.w6(32'h3b6d71ac),
	.w7(32'h3b449fab),
	.w8(32'hb889e8e9),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b925e),
	.w1(32'hbb671b4d),
	.w2(32'hba8bed5a),
	.w3(32'hb8ae57eb),
	.w4(32'hba18dae8),
	.w5(32'hbabc34e8),
	.w6(32'hb9e3de7d),
	.w7(32'h3a0ed39d),
	.w8(32'hbab3e221),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28455c),
	.w1(32'hba8c7b81),
	.w2(32'hbb126783),
	.w3(32'hba90aa39),
	.w4(32'hba0c8183),
	.w5(32'hbb06fc2d),
	.w6(32'hba842357),
	.w7(32'h3ac9acfe),
	.w8(32'hbad0714f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d009f5),
	.w1(32'hba80ff8c),
	.w2(32'hbb54c5e2),
	.w3(32'h39daa56e),
	.w4(32'h3a4ca924),
	.w5(32'hbb082195),
	.w6(32'h3a106e98),
	.w7(32'h3a159b85),
	.w8(32'hbb05f6a9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32d503),
	.w1(32'hba803270),
	.w2(32'hba945ac0),
	.w3(32'hb8638a55),
	.w4(32'hbaa534b6),
	.w5(32'hbafd601d),
	.w6(32'h3ae3712a),
	.w7(32'h39114031),
	.w8(32'hbad20bb1),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41f0a1),
	.w1(32'hba8c0e1a),
	.w2(32'h3953c293),
	.w3(32'h3ab6a32e),
	.w4(32'h3986dad1),
	.w5(32'h3a385078),
	.w6(32'hb7fa239e),
	.w7(32'hba29681a),
	.w8(32'h38c74419),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7233f2),
	.w1(32'h3941049c),
	.w2(32'hbb0b2f76),
	.w3(32'h3adaebdb),
	.w4(32'h3ac261a1),
	.w5(32'hb9ff1f86),
	.w6(32'h39a03c17),
	.w7(32'h3a8f07e1),
	.w8(32'hb9c995ea),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e11e55),
	.w1(32'h399f6afd),
	.w2(32'h3a9c8040),
	.w3(32'hb9daa258),
	.w4(32'hb98fa798),
	.w5(32'h3b1c48cc),
	.w6(32'hb7cc11d4),
	.w7(32'hb9181efe),
	.w8(32'h3a62631e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391608f6),
	.w1(32'hb9bdd48a),
	.w2(32'hbb38e00c),
	.w3(32'h3b19ceff),
	.w4(32'h3a840e1a),
	.w5(32'hbb3b72fb),
	.w6(32'h3af2a365),
	.w7(32'h3adaec4b),
	.w8(32'hbb692205),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca98c4),
	.w1(32'hbab98484),
	.w2(32'h3a52fb34),
	.w3(32'hbadabc6e),
	.w4(32'hbaa51d59),
	.w5(32'h3a82682d),
	.w6(32'hbaeed68d),
	.w7(32'hbaf37884),
	.w8(32'h3985f299),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda56ee),
	.w1(32'hba3727bf),
	.w2(32'hbaefab35),
	.w3(32'h3bd32382),
	.w4(32'hba4f74ff),
	.w5(32'hbb23c1bd),
	.w6(32'h3bf5ef8d),
	.w7(32'hba8bef08),
	.w8(32'hbb385526),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39de64),
	.w1(32'h368e6750),
	.w2(32'h3a39d3e4),
	.w3(32'h36c5d050),
	.w4(32'h3a196f06),
	.w5(32'h3a6a057e),
	.w6(32'h3ab752b0),
	.w7(32'h39d8c649),
	.w8(32'hb9d48ae2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a435f),
	.w1(32'hb9016c80),
	.w2(32'h38da21a0),
	.w3(32'h3a8aef01),
	.w4(32'hba27c61a),
	.w5(32'h38a0c1b0),
	.w6(32'h3a0a36c8),
	.w7(32'hba152bb6),
	.w8(32'h394659a5),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83232c),
	.w1(32'h3a9ce82a),
	.w2(32'h3b1c2d43),
	.w3(32'h3a2bb57b),
	.w4(32'h3a169c78),
	.w5(32'h3b080bf1),
	.w6(32'h3a58bbb9),
	.w7(32'h3a519614),
	.w8(32'h3b0ff860),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b099ac0),
	.w1(32'h3aedf6c3),
	.w2(32'h3aa29f45),
	.w3(32'h3b22a736),
	.w4(32'h3b135369),
	.w5(32'h3adb1aa1),
	.w6(32'h3b057a04),
	.w7(32'h3af4f35c),
	.w8(32'h3b11df83),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b532926),
	.w1(32'hbb155964),
	.w2(32'h39a5024e),
	.w3(32'h3b677ed4),
	.w4(32'hba88ccb6),
	.w5(32'hba4b8032),
	.w6(32'h3ba4b35e),
	.w7(32'hbb3598aa),
	.w8(32'hbae58d1c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38163ece),
	.w1(32'hbb6cdefa),
	.w2(32'hbb0e2671),
	.w3(32'h389fb441),
	.w4(32'hbb4e1297),
	.w5(32'hbaf620a6),
	.w6(32'hba837e52),
	.w7(32'hbb5cdf93),
	.w8(32'hbaf6f076),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba013697),
	.w1(32'hb958f84f),
	.w2(32'h3b65107b),
	.w3(32'h39616f9f),
	.w4(32'h395467eb),
	.w5(32'h3b75ae57),
	.w6(32'h39cadff0),
	.w7(32'h3a32df5f),
	.w8(32'h3bb00114),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3713b),
	.w1(32'h3a30ae8f),
	.w2(32'hba9a081d),
	.w3(32'h3b0c93d1),
	.w4(32'h39228a4b),
	.w5(32'hbb21983d),
	.w6(32'h3ba2e661),
	.w7(32'h3b082a04),
	.w8(32'hbb2215d3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a998e),
	.w1(32'hba409da4),
	.w2(32'hba8b9648),
	.w3(32'hb9adfc93),
	.w4(32'hb9a18053),
	.w5(32'hba8060fd),
	.w6(32'hb955eaa8),
	.w7(32'hba96ebc9),
	.w8(32'hbaaba66b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1c5bc),
	.w1(32'hbabf8e2d),
	.w2(32'hbaddf5da),
	.w3(32'hbaf8c261),
	.w4(32'hbae53e56),
	.w5(32'hbb1a8a43),
	.w6(32'hbaa7d32c),
	.w7(32'hbaabae67),
	.w8(32'hbaf152fe),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6ab25),
	.w1(32'hb9dc15c2),
	.w2(32'h3aa37098),
	.w3(32'h3ba3b54e),
	.w4(32'hbb180c91),
	.w5(32'hbb2a2a8d),
	.w6(32'h3baa8b45),
	.w7(32'hbb4c1c37),
	.w8(32'hbb967a02),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f3466),
	.w1(32'h3a7ef3b7),
	.w2(32'hbac4b24c),
	.w3(32'h3a9aa444),
	.w4(32'h3ac2cf26),
	.w5(32'hbb232c96),
	.w6(32'h3a48e6f9),
	.w7(32'h3a5eca7e),
	.w8(32'hbab6da73),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61a867),
	.w1(32'h39e659fe),
	.w2(32'h3b0cc871),
	.w3(32'hba522124),
	.w4(32'hbac63eda),
	.w5(32'h3b5ea10e),
	.w6(32'hba4e929e),
	.w7(32'hba8643ef),
	.w8(32'h3b476a7a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813c1d),
	.w1(32'hbaf66263),
	.w2(32'hbbc0e68e),
	.w3(32'hbb86ff30),
	.w4(32'hbaf45b3c),
	.w5(32'hba740c9e),
	.w6(32'hbb8fed24),
	.w7(32'hbb83ebd6),
	.w8(32'hbb280e10),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb637574),
	.w1(32'hbb7c132d),
	.w2(32'h3c2138ce),
	.w3(32'hbb7bb1f4),
	.w4(32'h3a6d274e),
	.w5(32'h3b2693c8),
	.w6(32'h3b289f91),
	.w7(32'h3c34f7f3),
	.w8(32'hbbcc9612),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe603a7),
	.w1(32'hbbb3adb2),
	.w2(32'h3b632581),
	.w3(32'hbbdf1896),
	.w4(32'hbc4bff26),
	.w5(32'h3b83e6b2),
	.w6(32'h3b917f12),
	.w7(32'hbc377c6c),
	.w8(32'h3b8fb26b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4b3ea),
	.w1(32'hbb89ac00),
	.w2(32'hbb07dc1f),
	.w3(32'hb90c5563),
	.w4(32'hbb936627),
	.w5(32'h3aa7e9bd),
	.w6(32'hb96d5860),
	.w7(32'hbb71bf0f),
	.w8(32'h3bf0b20b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5cc7b),
	.w1(32'hb8552f8d),
	.w2(32'h3b8dc759),
	.w3(32'h3c59ddd2),
	.w4(32'hbc745791),
	.w5(32'h3b9434a5),
	.w6(32'h3c31e19b),
	.w7(32'hbc03a5e1),
	.w8(32'h3c6bda57),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c870467),
	.w1(32'h3a4da6d8),
	.w2(32'hbbeb5221),
	.w3(32'h3c689fac),
	.w4(32'hbbc35399),
	.w5(32'hbbb9ff58),
	.w6(32'h3b589df7),
	.w7(32'hbc850528),
	.w8(32'hbb3ee05b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ed9f9),
	.w1(32'h399c8d80),
	.w2(32'hbbf4032d),
	.w3(32'hbb92278a),
	.w4(32'h3b1a3908),
	.w5(32'hbaaaf7dc),
	.w6(32'hbaa88275),
	.w7(32'h3ba995b2),
	.w8(32'h3c03ac8f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03f69b),
	.w1(32'hbc5a4e09),
	.w2(32'hbb02213c),
	.w3(32'hbc2f6dff),
	.w4(32'hbb05a3d7),
	.w5(32'hbb60b2e3),
	.w6(32'hbc561a3b),
	.w7(32'hbc50e24d),
	.w8(32'hbabb3f24),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e7d77),
	.w1(32'h3b0e9177),
	.w2(32'h3c4dad77),
	.w3(32'hba5f4376),
	.w4(32'h3b954d5a),
	.w5(32'h3ccf8a83),
	.w6(32'hba065dab),
	.w7(32'h3af57a85),
	.w8(32'h3c254438),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f7050),
	.w1(32'hbc5accb6),
	.w2(32'h391db74f),
	.w3(32'hbc76810a),
	.w4(32'h3c378153),
	.w5(32'hb8cc7af3),
	.w6(32'hbcac1f22),
	.w7(32'h3cc3b07c),
	.w8(32'h3a35f122),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba83c2f),
	.w1(32'h3bae120d),
	.w2(32'h3b1e2010),
	.w3(32'hbbc2de8b),
	.w4(32'h3c3f74d0),
	.w5(32'h3bcc6d38),
	.w6(32'h3ac3ec45),
	.w7(32'h3c56888e),
	.w8(32'h3c55908f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c981b),
	.w1(32'hbc3a6bf8),
	.w2(32'hbbc4ed12),
	.w3(32'h3c1b26f7),
	.w4(32'hbc8e7c6d),
	.w5(32'hbb9da82a),
	.w6(32'h3b3382cf),
	.w7(32'hbc1b03b0),
	.w8(32'hbb23f550),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc494a04),
	.w1(32'hb9ac89be),
	.w2(32'hbc18ed6f),
	.w3(32'hbc4fc92b),
	.w4(32'h3c3ba782),
	.w5(32'hbc06c48a),
	.w6(32'hbc13e120),
	.w7(32'h3b89c579),
	.w8(32'hbbd44a2a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c3397),
	.w1(32'hbbda3a74),
	.w2(32'hba62d61c),
	.w3(32'hbb68d3c7),
	.w4(32'hbb874e80),
	.w5(32'hba781778),
	.w6(32'hbba02f84),
	.w7(32'hbc04b5a1),
	.w8(32'hbb049a55),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12d700),
	.w1(32'hb9f86863),
	.w2(32'hbb77e6b9),
	.w3(32'h3b949b19),
	.w4(32'h3b3faa09),
	.w5(32'hbc168127),
	.w6(32'hba9072c8),
	.w7(32'hbb2a6d50),
	.w8(32'h3b89b077),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6e4ae),
	.w1(32'hbb4dacfe),
	.w2(32'h3b375fe5),
	.w3(32'h3beb507d),
	.w4(32'hbc536479),
	.w5(32'h3acc1c51),
	.w6(32'h3bcdcf64),
	.w7(32'hbbc562e6),
	.w8(32'hba9fc3bc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407b12),
	.w1(32'hbb4dbd53),
	.w2(32'hbc15a482),
	.w3(32'h39b8a39b),
	.w4(32'hbbe3b7bd),
	.w5(32'hbc52d446),
	.w6(32'hbb7010d7),
	.w7(32'hbc0f519d),
	.w8(32'hbc6dbf2f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba96fb5),
	.w1(32'h3ce70d24),
	.w2(32'hbb102310),
	.w3(32'h3c126e2f),
	.w4(32'h3cac6b5e),
	.w5(32'hbc3750f2),
	.w6(32'h3d0f9a10),
	.w7(32'hbadb149b),
	.w8(32'h3c2d1812),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10a257),
	.w1(32'h3be5b605),
	.w2(32'h3c0de325),
	.w3(32'h3c7efdde),
	.w4(32'hbb9daead),
	.w5(32'h3a3aa2ed),
	.w6(32'h3b73a816),
	.w7(32'hbc52a0b8),
	.w8(32'hbbcb573f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fda71),
	.w1(32'hbc30c145),
	.w2(32'hbc434198),
	.w3(32'hbba24d60),
	.w4(32'hbbfa5f57),
	.w5(32'hbc4db726),
	.w6(32'h3ab12ba7),
	.w7(32'hbb3ce8e8),
	.w8(32'hbc43dccb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e7d6b),
	.w1(32'hbbfc91b9),
	.w2(32'h3abc8ccc),
	.w3(32'hbc3a2f23),
	.w4(32'h3aeac678),
	.w5(32'hb9d2652d),
	.w6(32'h39a0a104),
	.w7(32'h3a271545),
	.w8(32'h396f4049),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3765f3f6),
	.w1(32'h3a60873b),
	.w2(32'hbb8e5a0d),
	.w3(32'h3a857bc1),
	.w4(32'h39cf6a53),
	.w5(32'hbbaaf2a7),
	.w6(32'hb8c5ad3d),
	.w7(32'hb9fe6ffd),
	.w8(32'h3be72a28),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadca530),
	.w1(32'hbb64424f),
	.w2(32'hb9a0eebd),
	.w3(32'h3bc72358),
	.w4(32'hbc2811fa),
	.w5(32'hbbab5808),
	.w6(32'hbbf7554b),
	.w7(32'hbc5ac02f),
	.w8(32'hbc1bc1b2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc821d91),
	.w1(32'hbae73ac9),
	.w2(32'hbc1207f9),
	.w3(32'hbc467315),
	.w4(32'hbb90a37c),
	.w5(32'hbc38daba),
	.w6(32'hbb24339f),
	.w7(32'hbc6ef196),
	.w8(32'hbc8dfd06),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc1d0),
	.w1(32'h3c85b602),
	.w2(32'hbbb93563),
	.w3(32'h3c44e354),
	.w4(32'hbbb2c03e),
	.w5(32'hbb8786bc),
	.w6(32'h3c12adeb),
	.w7(32'hbc7be8fd),
	.w8(32'hbc14c693),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d39cd),
	.w1(32'h3c7413bb),
	.w2(32'h3b848337),
	.w3(32'hbaab9169),
	.w4(32'h3c33016e),
	.w5(32'h3b73e47c),
	.w6(32'h3c370edd),
	.w7(32'hbb89d41c),
	.w8(32'h3b46189e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffc522),
	.w1(32'h3a82dfe1),
	.w2(32'hbc1fb9b9),
	.w3(32'h3a7f14e9),
	.w4(32'hbc067f1c),
	.w5(32'hbb3b22bf),
	.w6(32'hbb85a869),
	.w7(32'hbb98fabf),
	.w8(32'hbc317645),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded929),
	.w1(32'hbc0b5d52),
	.w2(32'hbae023c2),
	.w3(32'hbc236aa3),
	.w4(32'hbb8ee5f4),
	.w5(32'hbc546f87),
	.w6(32'hbac3842c),
	.w7(32'hb9dd1485),
	.w8(32'hbbff1b98),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6786b),
	.w1(32'hbaa3d736),
	.w2(32'h3c569224),
	.w3(32'h3ab70538),
	.w4(32'hba67325e),
	.w5(32'h3c0a3689),
	.w6(32'hbac6877f),
	.w7(32'hbc87e0aa),
	.w8(32'h3b610e84),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac63da8),
	.w1(32'hbab3a21d),
	.w2(32'hba0747d2),
	.w3(32'hbc5d8968),
	.w4(32'hbbcb56e0),
	.w5(32'hbb1f69e6),
	.w6(32'h3b099d6f),
	.w7(32'hbadc1bb5),
	.w8(32'h3b03e06e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba154e08),
	.w1(32'h3c1855ed),
	.w2(32'hbb246adf),
	.w3(32'h3a385710),
	.w4(32'h3bf9fe67),
	.w5(32'hba3801e2),
	.w6(32'h3b46d0c2),
	.w7(32'h3af23923),
	.w8(32'h3c092771),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb981afb),
	.w1(32'h3b883872),
	.w2(32'h3b19cfbe),
	.w3(32'hbba908f3),
	.w4(32'h3b9e4fe6),
	.w5(32'h3b4e7771),
	.w6(32'h3bd2214f),
	.w7(32'h3c60470b),
	.w8(32'h3ae33736),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2900ba),
	.w1(32'hbbc8aeac),
	.w2(32'hbbac4b5c),
	.w3(32'h3b637410),
	.w4(32'hbc4e26f0),
	.w5(32'hbb46c0b9),
	.w6(32'hbb9aef9e),
	.w7(32'hbc5cce1c),
	.w8(32'hbba83dfe),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2893dc),
	.w1(32'hbc0c45c6),
	.w2(32'hbbb017c6),
	.w3(32'h3b8f16a3),
	.w4(32'hbbd359a8),
	.w5(32'hbbb54831),
	.w6(32'hbb88da9d),
	.w7(32'hbc50bf75),
	.w8(32'h39331934),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c7de3),
	.w1(32'hbbfb1fd3),
	.w2(32'h3bf8afdc),
	.w3(32'hbc7ec177),
	.w4(32'hbc7419d2),
	.w5(32'h3bf7de07),
	.w6(32'hbc7bc803),
	.w7(32'hbc583642),
	.w8(32'h3c149053),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5df750),
	.w1(32'h3b3a7c55),
	.w2(32'h3b4eaef5),
	.w3(32'h3c23ca5e),
	.w4(32'hbbb2cd6d),
	.w5(32'h3a61274b),
	.w6(32'hb8d0784e),
	.w7(32'hbb9e8c2a),
	.w8(32'hbbd20950),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3436c),
	.w1(32'hba0d111a),
	.w2(32'hbb742b85),
	.w3(32'hbbdbad91),
	.w4(32'h3bba5857),
	.w5(32'h3bd02591),
	.w6(32'hbc099745),
	.w7(32'h3aca6d51),
	.w8(32'hba19b8a3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba12171),
	.w1(32'hbbbc433d),
	.w2(32'h3a6f8cea),
	.w3(32'h3bb1956a),
	.w4(32'hbc2ab928),
	.w5(32'h3ad9a7b1),
	.w6(32'hba165289),
	.w7(32'hbb9ab679),
	.w8(32'h3ae60c57),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac72f73),
	.w1(32'h3b690e13),
	.w2(32'h3bea491c),
	.w3(32'hba2a974b),
	.w4(32'h3b304a24),
	.w5(32'h3c22d290),
	.w6(32'hba7e3427),
	.w7(32'hbb23a917),
	.w8(32'h3bbec994),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba13ccb),
	.w1(32'hbb721276),
	.w2(32'hbab108f6),
	.w3(32'h3b8e1e62),
	.w4(32'hbb9403d4),
	.w5(32'hbbd1447b),
	.w6(32'h3a5bff2d),
	.w7(32'hbbbbcd63),
	.w8(32'hbc2929eb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a9c50),
	.w1(32'h3c323349),
	.w2(32'h3a5bfcff),
	.w3(32'hbb32469b),
	.w4(32'h3cd55242),
	.w5(32'h3adc8c4c),
	.w6(32'h3c904f1f),
	.w7(32'h3bf1f6a8),
	.w8(32'h3be2e62b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4fbf4),
	.w1(32'hbb758e56),
	.w2(32'h39ae16a7),
	.w3(32'hbb8a4fbd),
	.w4(32'hbaaf0d82),
	.w5(32'hba296b1f),
	.w6(32'hba789eb6),
	.w7(32'hbc06d790),
	.w8(32'hba7854a7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c555b9),
	.w1(32'hbb15b934),
	.w2(32'hbc2aed70),
	.w3(32'hba3c2b1d),
	.w4(32'hbb13d434),
	.w5(32'hbc336d89),
	.w6(32'hbb6c9d44),
	.w7(32'hbb1f67d3),
	.w8(32'hbc58ef59),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f2c46),
	.w1(32'hbb80e5fc),
	.w2(32'hbb413c40),
	.w3(32'h3c0f6191),
	.w4(32'hbb31db7d),
	.w5(32'hbacc8115),
	.w6(32'h3c60d3dc),
	.w7(32'hbba05c01),
	.w8(32'hbb6e44b0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcb969),
	.w1(32'h399da5c4),
	.w2(32'h3be4c004),
	.w3(32'hb8f4a602),
	.w4(32'h3bc48b6d),
	.w5(32'hbb04913f),
	.w6(32'h3b8c3eaa),
	.w7(32'h3b5b183b),
	.w8(32'hbc297d05),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56cb03),
	.w1(32'hbcae503d),
	.w2(32'hbb6e6f27),
	.w3(32'hbce34c1d),
	.w4(32'hbca5f676),
	.w5(32'h3b535105),
	.w6(32'hbc7fa0da),
	.w7(32'hbbc8bed3),
	.w8(32'h3bfa6b90),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e5aaf),
	.w1(32'hbbb9af62),
	.w2(32'hbb8d9f72),
	.w3(32'h3c2a800b),
	.w4(32'hbcbba7de),
	.w5(32'hbb1d5ce9),
	.w6(32'hbbb2578f),
	.w7(32'hbc86d68e),
	.w8(32'hbb4fa7a8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af63f6c),
	.w1(32'h3aea72e9),
	.w2(32'hbc0dfe6a),
	.w3(32'h3a48f60b),
	.w4(32'h3a1d5605),
	.w5(32'hbc2231cc),
	.w6(32'hba08929c),
	.w7(32'hbabaf820),
	.w8(32'hbbb813d9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11dbff),
	.w1(32'h38ac6443),
	.w2(32'hbb380cdd),
	.w3(32'hbbf8e72d),
	.w4(32'hbb77d101),
	.w5(32'h3bacc42d),
	.w6(32'hbb1843a0),
	.w7(32'h3acc1acf),
	.w8(32'h3beb49db),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f1493),
	.w1(32'hbc1d58df),
	.w2(32'h3aee9235),
	.w3(32'hbb22c6c3),
	.w4(32'hbc670f98),
	.w5(32'h3ac3c499),
	.w6(32'hbc88c4ec),
	.w7(32'hbc03d709),
	.w8(32'h3c05297c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f1ef),
	.w1(32'hbc46aaa0),
	.w2(32'hbb764041),
	.w3(32'hbb087c97),
	.w4(32'hbc91850e),
	.w5(32'h3b7d6f4b),
	.w6(32'hbc3e62fe),
	.w7(32'hbc57d8a7),
	.w8(32'hbbe5e264),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865d24),
	.w1(32'hbaac19d8),
	.w2(32'hb992f2de),
	.w3(32'hbbb2bc92),
	.w4(32'hbb540b93),
	.w5(32'hbaf34a68),
	.w6(32'h3b440551),
	.w7(32'hba598e02),
	.w8(32'h39ebca3f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30c92b),
	.w1(32'hbb59ea69),
	.w2(32'hbc031de7),
	.w3(32'hbb2b50af),
	.w4(32'hbb1084d6),
	.w5(32'hbc23b464),
	.w6(32'hbb44c2e8),
	.w7(32'hbb7096f2),
	.w8(32'hbc38fb0d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfae0f9),
	.w1(32'h3b8b7532),
	.w2(32'h3a2e4378),
	.w3(32'hbb96e9d4),
	.w4(32'h3c2718bd),
	.w5(32'h3b115f7c),
	.w6(32'h3b914906),
	.w7(32'h3b6242fe),
	.w8(32'h3b0593f3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8353db),
	.w1(32'hbba357a0),
	.w2(32'hbbb6e0ec),
	.w3(32'h3b26fe88),
	.w4(32'hbbc79a9b),
	.w5(32'hba6047ce),
	.w6(32'h39fce5b6),
	.w7(32'hbbbd40e5),
	.w8(32'h3a34792e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fc94d),
	.w1(32'hbbe80d3a),
	.w2(32'hbad347db),
	.w3(32'hbc285047),
	.w4(32'h3bd4fc00),
	.w5(32'h3b583668),
	.w6(32'hbc9850cf),
	.w7(32'h3c995186),
	.w8(32'h3b55896e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba89e5c),
	.w1(32'h3a5e89a9),
	.w2(32'h39f6c9e2),
	.w3(32'hbc097538),
	.w4(32'h3b37f417),
	.w5(32'h3bd71b8b),
	.w6(32'h3abc7611),
	.w7(32'h3c2b3c95),
	.w8(32'h3af3544d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb613500),
	.w1(32'hbc18fb80),
	.w2(32'hbc722b4b),
	.w3(32'hbc8d9b88),
	.w4(32'hbc45f6ec),
	.w5(32'hbcd95259),
	.w6(32'hbc52f0a6),
	.w7(32'hbb08f350),
	.w8(32'hbcb96319),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c346),
	.w1(32'h3bd70c55),
	.w2(32'hb9dbbf60),
	.w3(32'h3c6ac2e0),
	.w4(32'h387ed4db),
	.w5(32'hbad8c01f),
	.w6(32'h3c7f601c),
	.w7(32'hbc89e1bc),
	.w8(32'hbb6d818d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847316),
	.w1(32'hb71ffd1b),
	.w2(32'h3a9676df),
	.w3(32'hbb61e2e1),
	.w4(32'h3b043256),
	.w5(32'h3b2cbee8),
	.w6(32'h3a92ce12),
	.w7(32'h3b06bb40),
	.w8(32'h3b1ec216),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c926f),
	.w1(32'hbb5937c6),
	.w2(32'h3ad76811),
	.w3(32'h3af50a08),
	.w4(32'hbbe7c5dd),
	.w5(32'hbab9776b),
	.w6(32'hb9fde299),
	.w7(32'hbc227561),
	.w8(32'hbc04ab38),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82cb82),
	.w1(32'h3cb4316b),
	.w2(32'hbb00b680),
	.w3(32'hbac2de39),
	.w4(32'h3c9c179f),
	.w5(32'hbc2620ec),
	.w6(32'h3bf707a8),
	.w7(32'hba460fde),
	.w8(32'h3bb3c961),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b545f25),
	.w1(32'hbb3219ed),
	.w2(32'hbb775ae6),
	.w3(32'h3ba89f60),
	.w4(32'hbbbe3753),
	.w5(32'hbb6d0679),
	.w6(32'h3a86466c),
	.w7(32'hbc624f33),
	.w8(32'h3b6e29e6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a473f),
	.w1(32'h3a7023c3),
	.w2(32'h3b2a1feb),
	.w3(32'h3af0d137),
	.w4(32'hbb7879c8),
	.w5(32'h3bebea95),
	.w6(32'hbb26590e),
	.w7(32'hbc1218f3),
	.w8(32'h3c1095c4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b5f7f),
	.w1(32'hb9d58be0),
	.w2(32'hbbaf6d32),
	.w3(32'hbae980c4),
	.w4(32'h3c09c353),
	.w5(32'h3896e055),
	.w6(32'hba3f1511),
	.w7(32'h3bf9f647),
	.w8(32'h39206efe),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ce56),
	.w1(32'hbb9bea27),
	.w2(32'h3bf5740d),
	.w3(32'hbb26a200),
	.w4(32'hbb9ec88e),
	.w5(32'h3bfc8bd5),
	.w6(32'hbb68aa1b),
	.w7(32'hbbdc2283),
	.w8(32'h3b9363fb),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a721158),
	.w1(32'hbc1ff01e),
	.w2(32'h3a5a5056),
	.w3(32'h3a72ba34),
	.w4(32'hbc12ea90),
	.w5(32'h3bf81d2c),
	.w6(32'hbb70fc35),
	.w7(32'hbc259ec5),
	.w8(32'h3b31ec79),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95dee70),
	.w1(32'h3ab1daea),
	.w2(32'hbb873cc8),
	.w3(32'hb9f21f76),
	.w4(32'h3b6f0b03),
	.w5(32'hbc3ff293),
	.w6(32'h3993724d),
	.w7(32'h39d2a890),
	.w8(32'hbc049878),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15998a),
	.w1(32'h3c5c7c49),
	.w2(32'hbb8f4854),
	.w3(32'hbb420ec3),
	.w4(32'hbc0efe23),
	.w5(32'hbbad08da),
	.w6(32'h3b621fc1),
	.w7(32'hbc584c1f),
	.w8(32'hbbae8367),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3527c7),
	.w1(32'h3c1363dd),
	.w2(32'h3c33f961),
	.w3(32'hbc4765b2),
	.w4(32'h3bd37d7c),
	.w5(32'h3c8899d9),
	.w6(32'hbbe22a4a),
	.w7(32'hbbb8476d),
	.w8(32'h3c7f24d4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c616f00),
	.w1(32'h3b217be3),
	.w2(32'h3b38e069),
	.w3(32'h3cbded1e),
	.w4(32'hbbb59f4b),
	.w5(32'hbc360d25),
	.w6(32'h3c3eb6fe),
	.w7(32'hbb915365),
	.w8(32'hbc20982d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c229d),
	.w1(32'hb9f9cf01),
	.w2(32'h3b7abd3c),
	.w3(32'hbc893c4c),
	.w4(32'h3b5af04b),
	.w5(32'hbb1a36cf),
	.w6(32'hbb9bdfc3),
	.w7(32'hbb36bf91),
	.w8(32'hbb20bacb),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33e036),
	.w1(32'hbb1b34f4),
	.w2(32'hbc48fcba),
	.w3(32'h3b8ef7f5),
	.w4(32'hbb249709),
	.w5(32'hbc3b2e79),
	.w6(32'h3bbf03d1),
	.w7(32'hbbeb41a7),
	.w8(32'hbc178cdd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c7c72),
	.w1(32'hbb578470),
	.w2(32'hbb723704),
	.w3(32'h3c41a1a6),
	.w4(32'hbc42de07),
	.w5(32'hbc029725),
	.w6(32'h3c350308),
	.w7(32'hbbb86916),
	.w8(32'h3b3fdd5d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c025474),
	.w1(32'h3b98bead),
	.w2(32'h3b1bd49a),
	.w3(32'h3c21f3de),
	.w4(32'hbc26443f),
	.w5(32'h3922a0ce),
	.w6(32'h3c214049),
	.w7(32'hbb9e8caa),
	.w8(32'hbc10a672),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1649f4),
	.w1(32'h3a174c07),
	.w2(32'hbc576578),
	.w3(32'hbbebb5f2),
	.w4(32'h3bfb1384),
	.w5(32'hbc21ca4f),
	.w6(32'hbb308eb8),
	.w7(32'hba93d0a0),
	.w8(32'hbc4f10b1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bf921),
	.w1(32'hb887285c),
	.w2(32'hbcb71d21),
	.w3(32'h3b7bdf9b),
	.w4(32'hbba10da3),
	.w5(32'hbd02cc24),
	.w6(32'h3c0c8422),
	.w7(32'hbbf1acd6),
	.w8(32'hbcf8bea0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1cd5a),
	.w1(32'h3bade37c),
	.w2(32'hbbaae460),
	.w3(32'hb9caeec9),
	.w4(32'h3c37c470),
	.w5(32'hbb94a1f5),
	.w6(32'h3c03ef7b),
	.w7(32'h3c0c0983),
	.w8(32'hbc80d38b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc680128),
	.w1(32'hbacc2c4c),
	.w2(32'hbc35d81b),
	.w3(32'hbc3a9d89),
	.w4(32'h3bd01c0f),
	.w5(32'hbc167c0b),
	.w6(32'hbb36d1f2),
	.w7(32'h3c24b33f),
	.w8(32'hbc8071b0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97c11a),
	.w1(32'hbab6a072),
	.w2(32'hbbbafb5e),
	.w3(32'hbc3d990f),
	.w4(32'h3b73ece1),
	.w5(32'h3a9bba43),
	.w6(32'hbb844cb7),
	.w7(32'hbaca985d),
	.w8(32'h3b60ec7f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9be63),
	.w1(32'hbab82aed),
	.w2(32'h3bccba26),
	.w3(32'h3c39c748),
	.w4(32'hbc4cb929),
	.w5(32'h3b41ee99),
	.w6(32'h3c1782f5),
	.w7(32'hbc759bf9),
	.w8(32'hbb46a6d9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d2b45),
	.w1(32'hbc8166f0),
	.w2(32'hbb8d0278),
	.w3(32'hbc86f59e),
	.w4(32'hbc5b1b6e),
	.w5(32'hbb439aaa),
	.w6(32'hbb85348e),
	.w7(32'hbbfe4b80),
	.w8(32'h3bce848e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f7fd2),
	.w1(32'hbbab4c95),
	.w2(32'hbad09cbb),
	.w3(32'h3bc7a138),
	.w4(32'hbceb9dd9),
	.w5(32'h3b171596),
	.w6(32'h3b890624),
	.w7(32'hbcac826d),
	.w8(32'hbb8473a1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada05d3),
	.w1(32'hbada0cb3),
	.w2(32'h3c0ee6e5),
	.w3(32'h3b9b52fc),
	.w4(32'hbbcab90c),
	.w5(32'h3a99d0e8),
	.w6(32'hbaeefd2a),
	.w7(32'hbbd3629a),
	.w8(32'hbc0f3fda),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5057),
	.w1(32'hbc52d05e),
	.w2(32'hbb852828),
	.w3(32'hbc903166),
	.w4(32'h3c3afdcf),
	.w5(32'hb9ab7cd1),
	.w6(32'hbc0d5534),
	.w7(32'h3c32aefa),
	.w8(32'hba64702e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4bc7b),
	.w1(32'h3a153e6b),
	.w2(32'hbbf87a44),
	.w3(32'hbb268b32),
	.w4(32'h3b16c90d),
	.w5(32'h3996e403),
	.w6(32'hbb85ab6d),
	.w7(32'hbc2ae68d),
	.w8(32'h3be3c5de),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3778f2),
	.w1(32'h36e365eb),
	.w2(32'hbc9afb13),
	.w3(32'h3c6937bc),
	.w4(32'hbcca9799),
	.w5(32'hbc497200),
	.w6(32'h3c53207d),
	.w7(32'hbc8241ce),
	.w8(32'hbc1e12fd),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00093e),
	.w1(32'h39334bf1),
	.w2(32'h3aa98826),
	.w3(32'h3c000b43),
	.w4(32'h3bef494e),
	.w5(32'hbb4fa0bb),
	.w6(32'h3c9d5aaa),
	.w7(32'hbbb4a8ea),
	.w8(32'h3b96301b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a757e),
	.w1(32'hbb312940),
	.w2(32'hbb354e04),
	.w3(32'hbb6aaddd),
	.w4(32'hbbb7ee39),
	.w5(32'h3bcba9b9),
	.w6(32'hbaa407e9),
	.w7(32'h3b8d7ec1),
	.w8(32'h3bda3115),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a15ceb),
	.w1(32'hbbaddfe3),
	.w2(32'h3b8c3bab),
	.w3(32'hb9ba5163),
	.w4(32'hbab7de7f),
	.w5(32'hbb1770be),
	.w6(32'hbb1021ed),
	.w7(32'hba64021d),
	.w8(32'h3b1e4a26),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c1e74),
	.w1(32'hba234a49),
	.w2(32'hbaef0478),
	.w3(32'h39cb28cd),
	.w4(32'hbb9bcc4f),
	.w5(32'h3bc3681e),
	.w6(32'hbad19fc8),
	.w7(32'hbaeab03e),
	.w8(32'h3c09b2f8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c082ca2),
	.w1(32'hbab770d8),
	.w2(32'hbc1ad7c2),
	.w3(32'h3bd598f6),
	.w4(32'hbbaa5234),
	.w5(32'hbc046af2),
	.w6(32'h3c0729c4),
	.w7(32'hbbaa0749),
	.w8(32'hbb9a496f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b89091),
	.w1(32'h3b172969),
	.w2(32'hba9ab4ee),
	.w3(32'h3be744c6),
	.w4(32'hbbe5b024),
	.w5(32'hbbac6a1d),
	.w6(32'h3c1a5463),
	.w7(32'hbbbd60d3),
	.w8(32'hba4933aa),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2de7f),
	.w1(32'h3b994c43),
	.w2(32'hba99a7cd),
	.w3(32'h3bbd3237),
	.w4(32'h39e1f14d),
	.w5(32'h3a50c5e7),
	.w6(32'h3b5f7bdf),
	.w7(32'h3b342455),
	.w8(32'h3a9f9307),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad167e2),
	.w1(32'hb99e67b5),
	.w2(32'hba930879),
	.w3(32'hb9a87f22),
	.w4(32'hba86a30c),
	.w5(32'h39778ff7),
	.w6(32'hba042618),
	.w7(32'hbb2d61e5),
	.w8(32'h3b235b7a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae93e01),
	.w1(32'hba9a7df6),
	.w2(32'h3b6c6825),
	.w3(32'h3accd995),
	.w4(32'hbb2ddfc8),
	.w5(32'h3c315e0b),
	.w6(32'h3acc56ec),
	.w7(32'hbb0fa7a9),
	.w8(32'hbb61bb1e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87fe25),
	.w1(32'h3a472e9e),
	.w2(32'h3ae56c3a),
	.w3(32'hbca3974d),
	.w4(32'h3c5f1d46),
	.w5(32'hbac2c920),
	.w6(32'hbc719a56),
	.w7(32'h3c5a5f7d),
	.w8(32'hba95025b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cf8e6),
	.w1(32'h3a5561aa),
	.w2(32'hbc055408),
	.w3(32'hb9bf8e7c),
	.w4(32'hbae83cec),
	.w5(32'hbca2b094),
	.w6(32'h3b819227),
	.w7(32'hb97b3bf2),
	.w8(32'hbcb20720),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ac059),
	.w1(32'h3c83f6de),
	.w2(32'h3b24e977),
	.w3(32'hbc37cbbe),
	.w4(32'h3c8e7172),
	.w5(32'hbb538f22),
	.w6(32'hbacc9a78),
	.w7(32'h3cb47855),
	.w8(32'hbc667185),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9e077),
	.w1(32'h3b16b97a),
	.w2(32'hbb0225f1),
	.w3(32'hbb3a78d1),
	.w4(32'h3bfa0674),
	.w5(32'hbaced3e2),
	.w6(32'h3c960aad),
	.w7(32'h3bb12c70),
	.w8(32'hbc3207d6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ef09f),
	.w1(32'hb98ddc59),
	.w2(32'h3c3a3e9c),
	.w3(32'h3baf5864),
	.w4(32'h3c1c317b),
	.w5(32'h3b4ae988),
	.w6(32'h3c268e7e),
	.w7(32'h3b74e187),
	.w8(32'h3c7e8040),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule