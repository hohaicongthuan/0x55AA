module layer_10_featuremap_350(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee7229),
	.w1(32'hbadb9654),
	.w2(32'hbc0474ae),
	.w3(32'h3abb1f98),
	.w4(32'hba1d49e5),
	.w5(32'h3b007fd4),
	.w6(32'h3bade6dc),
	.w7(32'hbb031aa6),
	.w8(32'h3b1780bc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8926e),
	.w1(32'h3c19cdb2),
	.w2(32'hb9372a2f),
	.w3(32'h3b1792d4),
	.w4(32'hbc3aa3e6),
	.w5(32'hba8ac8c6),
	.w6(32'h3bad0652),
	.w7(32'hbc4c1022),
	.w8(32'hbbcfda20),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb56b54),
	.w1(32'h3c36bf60),
	.w2(32'h39bbf003),
	.w3(32'h3bbe8548),
	.w4(32'h3b99138b),
	.w5(32'hbb3ee249),
	.w6(32'h3c10e0a6),
	.w7(32'h3c3e24a8),
	.w8(32'h3ba073f0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77ecab),
	.w1(32'h3c49b90b),
	.w2(32'h3c56a14b),
	.w3(32'hbc1960dc),
	.w4(32'hbb433460),
	.w5(32'hbbcc352c),
	.w6(32'hbbb9d0b0),
	.w7(32'hbb228d8b),
	.w8(32'hbc985a5b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d06a0),
	.w1(32'hbc016da9),
	.w2(32'h3a3c2457),
	.w3(32'hb9c529fe),
	.w4(32'hbaa11537),
	.w5(32'hba4d2647),
	.w6(32'hbc62b1a9),
	.w7(32'hbc37d136),
	.w8(32'h3b3fe1cd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8114ed),
	.w1(32'h3b80a9e9),
	.w2(32'h39311d84),
	.w3(32'hbbc48b24),
	.w4(32'hbc07ddbf),
	.w5(32'hbb4368a1),
	.w6(32'hbb7e1035),
	.w7(32'hbbbac9d7),
	.w8(32'h3b7a774f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc040b6),
	.w1(32'h3cfb610c),
	.w2(32'h3b634ed7),
	.w3(32'h3b6ecf51),
	.w4(32'h3c4b4964),
	.w5(32'hbb59b2bc),
	.w6(32'h3b0bd701),
	.w7(32'h3b372cff),
	.w8(32'hbabd956b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25c02f),
	.w1(32'hbcdc7543),
	.w2(32'hbcb05353),
	.w3(32'h3c6e9f76),
	.w4(32'hb9d1f96b),
	.w5(32'hbc67a50a),
	.w6(32'hbd125c6e),
	.w7(32'h3becc134),
	.w8(32'h3b2b2038),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a8fda),
	.w1(32'h3ac1fdcd),
	.w2(32'hbadaec87),
	.w3(32'hbb15d102),
	.w4(32'hbbdf0140),
	.w5(32'hbbb27cd5),
	.w6(32'hbabb50e8),
	.w7(32'hb9c0cf53),
	.w8(32'hbab14a82),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68fa65),
	.w1(32'h3c01dbd3),
	.w2(32'h3ba69393),
	.w3(32'hbb02521e),
	.w4(32'hba448a3d),
	.w5(32'hbb213302),
	.w6(32'hbc28b232),
	.w7(32'h3aa2eec2),
	.w8(32'hbba0dbac),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba68064),
	.w1(32'h3b4cca22),
	.w2(32'h3a3e310a),
	.w3(32'hbbe18748),
	.w4(32'hbb9d8765),
	.w5(32'h3bdb33f7),
	.w6(32'hbc2f54c5),
	.w7(32'hbc043968),
	.w8(32'h3bbbec6a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c373de4),
	.w1(32'h3c8d4f30),
	.w2(32'h3c531ad6),
	.w3(32'h3c0f062d),
	.w4(32'h3cb4d67c),
	.w5(32'h3cb4d89b),
	.w6(32'h3b8b540f),
	.w7(32'h3c803721),
	.w8(32'h3c2478b2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25acaa),
	.w1(32'hbc17b708),
	.w2(32'h3affef53),
	.w3(32'h3ce3d090),
	.w4(32'h3d009602),
	.w5(32'h3bd9bc5a),
	.w6(32'h3a4a97fa),
	.w7(32'h3caab1d1),
	.w8(32'h3bfd8c1d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11a4f6),
	.w1(32'h3c111614),
	.w2(32'hbc112d64),
	.w3(32'h3c1ef5c6),
	.w4(32'h3b920968),
	.w5(32'h38958817),
	.w6(32'h3c66accd),
	.w7(32'hbb6ebc68),
	.w8(32'hbb672086),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71c792),
	.w1(32'h3b427995),
	.w2(32'h3bb4c87d),
	.w3(32'h3acfc326),
	.w4(32'hbbac46b1),
	.w5(32'h3a888b98),
	.w6(32'hba85d0b4),
	.w7(32'hbb03f059),
	.w8(32'h3c1edc11),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ed141),
	.w1(32'h3c733c06),
	.w2(32'h3bc5617a),
	.w3(32'hb9534c05),
	.w4(32'hbc8c88a4),
	.w5(32'hbbe23a59),
	.w6(32'h3c61e474),
	.w7(32'hbae94ae2),
	.w8(32'hbc4c65e4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b138ec2),
	.w1(32'h3c0e22ed),
	.w2(32'hbb2fcaad),
	.w3(32'hbc039434),
	.w4(32'hbc10c3c7),
	.w5(32'hba8ff662),
	.w6(32'h3a290614),
	.w7(32'hbc11f5a9),
	.w8(32'h3a85e7b8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2691b9),
	.w1(32'hbc530d19),
	.w2(32'hbbb53f75),
	.w3(32'h3cc4da94),
	.w4(32'h3c97865e),
	.w5(32'hbc7acbf7),
	.w6(32'hbbaf1dc5),
	.w7(32'h3cc13cf1),
	.w8(32'h3c02244f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca6da3),
	.w1(32'hbb9e8b4f),
	.w2(32'h3966f152),
	.w3(32'hbb659c8d),
	.w4(32'h3b3890e2),
	.w5(32'hbb69a05a),
	.w6(32'hbc43a43a),
	.w7(32'hb9b8fcde),
	.w8(32'h3a676c3c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3c493),
	.w1(32'hbb5428dc),
	.w2(32'hbb27f7fc),
	.w3(32'hbb049089),
	.w4(32'hbc1aa8d6),
	.w5(32'hba9a5794),
	.w6(32'h3cca18aa),
	.w7(32'hbc1c5207),
	.w8(32'hbbe0ef5c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb430948),
	.w1(32'hbb87d3be),
	.w2(32'hbbbe7105),
	.w3(32'h3abad8c6),
	.w4(32'h3bc4634d),
	.w5(32'h3ab0b7b8),
	.w6(32'h3a4f80e9),
	.w7(32'hba0bd018),
	.w8(32'h3ba885b1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3db40f),
	.w1(32'h3c067e79),
	.w2(32'h3c0cc7ff),
	.w3(32'h38a16fa2),
	.w4(32'hbc1d270f),
	.w5(32'h39584d29),
	.w6(32'hb94ee250),
	.w7(32'hbb7261f1),
	.w8(32'hbbb3c04a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a14e9),
	.w1(32'h3b14bafd),
	.w2(32'hbc0d98ed),
	.w3(32'hbb9aad13),
	.w4(32'h3c6351d9),
	.w5(32'h3c1c3f8c),
	.w6(32'h3bcb1efd),
	.w7(32'h3c3e6e2c),
	.w8(32'h3c40b01b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f005d),
	.w1(32'hbbbdd8dc),
	.w2(32'h3ad2bede),
	.w3(32'h3ba76f63),
	.w4(32'h3be14ec8),
	.w5(32'h3bd0932d),
	.w6(32'hbc428d4a),
	.w7(32'h3c01e41a),
	.w8(32'hbb453aa1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39d49d),
	.w1(32'hbbc70681),
	.w2(32'h3b777bcd),
	.w3(32'h3bdb6698),
	.w4(32'hbb43f9e1),
	.w5(32'h3a01c687),
	.w6(32'h3cf8e0df),
	.w7(32'hbbbf02b8),
	.w8(32'hbbc25bb4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43f1b),
	.w1(32'h3c3a31ac),
	.w2(32'h3b7f15e1),
	.w3(32'hbc0748d9),
	.w4(32'hbb9080b9),
	.w5(32'hb922b1cf),
	.w6(32'hbb66c3f5),
	.w7(32'hbae6d663),
	.w8(32'h3c1fddc2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ad9e3),
	.w1(32'h3c7b0a69),
	.w2(32'h3c036e6e),
	.w3(32'hbc830a3b),
	.w4(32'hbc4f6c39),
	.w5(32'hba0b6788),
	.w6(32'hbb997621),
	.w7(32'hba39df26),
	.w8(32'h3a405333),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23508f),
	.w1(32'hbac0879a),
	.w2(32'h3ca401ec),
	.w3(32'h3c5a4be0),
	.w4(32'hbc8d15bc),
	.w5(32'hbb739e4e),
	.w6(32'h3c4fb1c5),
	.w7(32'hb939b484),
	.w8(32'hbb849312),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71528f),
	.w1(32'hbb1644ca),
	.w2(32'hbb23f7c7),
	.w3(32'h3c1f7820),
	.w4(32'hbb421ee9),
	.w5(32'h3b8271e0),
	.w6(32'h3c85aabd),
	.w7(32'hb9431dab),
	.w8(32'h3b349d8f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca174f4),
	.w1(32'h3c3c4883),
	.w2(32'h3ad40474),
	.w3(32'h3c2cb01f),
	.w4(32'hbc878526),
	.w5(32'hbc9bd835),
	.w6(32'h3cbfc39a),
	.w7(32'hbbe7d7eb),
	.w8(32'hbc95b117),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41f3cb),
	.w1(32'hbc05946a),
	.w2(32'hbbba6336),
	.w3(32'hbc35a4dc),
	.w4(32'hbc1e5ea5),
	.w5(32'hbb79b759),
	.w6(32'hbb864a18),
	.w7(32'hbbfe4dd9),
	.w8(32'h3b801b91),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afca6c9),
	.w1(32'h3c17cecf),
	.w2(32'hbbc9f6b2),
	.w3(32'h3c01c460),
	.w4(32'hba44ade1),
	.w5(32'h3af86580),
	.w6(32'h3c65e77e),
	.w7(32'hbb53ef9c),
	.w8(32'h3b8c1973),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c55ff),
	.w1(32'h3c1182d8),
	.w2(32'h3b2c6639),
	.w3(32'hbb2bed7f),
	.w4(32'hbbb2d18e),
	.w5(32'hba2e2710),
	.w6(32'hbc1dae95),
	.w7(32'hbc0aa7e9),
	.w8(32'h3bdf83c1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2e052),
	.w1(32'hbbffe0a3),
	.w2(32'hbba67122),
	.w3(32'h3ba0c78a),
	.w4(32'h3bfc4cba),
	.w5(32'hba343e03),
	.w6(32'h3b57b2bb),
	.w7(32'h3b848beb),
	.w8(32'hba93d42c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb864194),
	.w1(32'hbba168cd),
	.w2(32'hba74d217),
	.w3(32'h3ba32506),
	.w4(32'hbad933f1),
	.w5(32'h3a82a2a9),
	.w6(32'h3cf87ba4),
	.w7(32'h3b9592b8),
	.w8(32'h3ac18f89),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c073c06),
	.w1(32'h3c19b597),
	.w2(32'h3aaeb4de),
	.w3(32'hbbcc1e49),
	.w4(32'h3c2bfca0),
	.w5(32'hbb526cf7),
	.w6(32'hbc15ca12),
	.w7(32'h3b164514),
	.w8(32'hbc0c700f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf5b85e),
	.w1(32'h3b3229cd),
	.w2(32'h3b32b420),
	.w3(32'hbd2184ac),
	.w4(32'h3cd13d3d),
	.w5(32'h3cab370a),
	.w6(32'hbd55e23f),
	.w7(32'h3a69c8b8),
	.w8(32'h3ce73ad5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd21693),
	.w1(32'h3c11e63c),
	.w2(32'h3c764798),
	.w3(32'h378b3ca3),
	.w4(32'hbcc7a5ad),
	.w5(32'h3b3f73a0),
	.w6(32'h3c7d380a),
	.w7(32'hbc97bcad),
	.w8(32'hbcad7cfa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc38f01),
	.w1(32'h3be6ffdf),
	.w2(32'h3c7e0e84),
	.w3(32'h3d02161e),
	.w4(32'h3ba53035),
	.w5(32'h3ba6de2f),
	.w6(32'h3d3072d7),
	.w7(32'hbc0a4f23),
	.w8(32'hbc5efcca),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3a368),
	.w1(32'hbbe5b042),
	.w2(32'h3b541206),
	.w3(32'h3bcf2c9c),
	.w4(32'hbc1ad671),
	.w5(32'hb8d81ecc),
	.w6(32'h3c3060bc),
	.w7(32'hbb25c530),
	.w8(32'hbbd2cf02),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2afbab),
	.w1(32'hbbc09c87),
	.w2(32'hba104faf),
	.w3(32'h3b92428e),
	.w4(32'h3b6e35f2),
	.w5(32'hbb5fb94b),
	.w6(32'hbc08a98f),
	.w7(32'hba838891),
	.w8(32'h3c15c1bd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb717b29d),
	.w1(32'h3c230aaf),
	.w2(32'h3a5a439f),
	.w3(32'hbc2258e0),
	.w4(32'hbbeff35e),
	.w5(32'hbbaaa664),
	.w6(32'h3b165a6c),
	.w7(32'hba6c4115),
	.w8(32'h3bb81239),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f5f3),
	.w1(32'h3c3005bc),
	.w2(32'h3c460c06),
	.w3(32'hbc4c9305),
	.w4(32'hbb0b1388),
	.w5(32'h3b9def1b),
	.w6(32'hb9e03309),
	.w7(32'h3a270e44),
	.w8(32'h3c9b9e75),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb63b47),
	.w1(32'h3ceb96bc),
	.w2(32'h3c87a1c4),
	.w3(32'hbd0b463e),
	.w4(32'hbc813c00),
	.w5(32'hbbe56fee),
	.w6(32'h3b9a21fa),
	.w7(32'h3b333a74),
	.w8(32'hbb0fd12c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adb5ea),
	.w1(32'hbb343f9a),
	.w2(32'h3be77ad1),
	.w3(32'hbc31eece),
	.w4(32'hbc40ba52),
	.w5(32'h3be6a177),
	.w6(32'hbc6e2b10),
	.w7(32'hbc71a6ea),
	.w8(32'h3b46d7a0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf329be),
	.w1(32'h3b8a4395),
	.w2(32'h3a447b02),
	.w3(32'hbc39103f),
	.w4(32'h3a1392bb),
	.w5(32'h3c084b4e),
	.w6(32'hbb1b381b),
	.w7(32'hbb073c80),
	.w8(32'h3c28ad70),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83c0cc),
	.w1(32'h3c1d6622),
	.w2(32'h3c45af8d),
	.w3(32'h3b7b2c31),
	.w4(32'hbba07a1c),
	.w5(32'h3bc6514b),
	.w6(32'h3b1951dc),
	.w7(32'h3b353484),
	.w8(32'hbb9af547),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b5a58),
	.w1(32'h3c6068ae),
	.w2(32'h3bebcab5),
	.w3(32'h3c49bddc),
	.w4(32'h3cdc2725),
	.w5(32'h3b88c5b5),
	.w6(32'hbc398900),
	.w7(32'h3cb2b978),
	.w8(32'h3c79644b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fd52a),
	.w1(32'hbc7e512e),
	.w2(32'hbbea01c2),
	.w3(32'h3c8bb43c),
	.w4(32'h3c8a4e4d),
	.w5(32'hbb77cc51),
	.w6(32'hbb29b169),
	.w7(32'h3c644c09),
	.w8(32'h3be364b0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1196cb),
	.w1(32'h3c197dea),
	.w2(32'h3b31ae5d),
	.w3(32'hbc207e41),
	.w4(32'hbc605287),
	.w5(32'hbb6421ac),
	.w6(32'hbbcceee3),
	.w7(32'hbbb09b53),
	.w8(32'hbbfbec69),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf89338),
	.w1(32'hbbb73765),
	.w2(32'hbb661aae),
	.w3(32'h3cb12156),
	.w4(32'hbbc916ef),
	.w5(32'hbb20d3f1),
	.w6(32'h3b89ba86),
	.w7(32'hbbfb55d8),
	.w8(32'h3bec4228),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6645e3),
	.w1(32'h3bdf4404),
	.w2(32'h3ba27ced),
	.w3(32'hbbb4bdeb),
	.w4(32'hbc0c77f1),
	.w5(32'h3a6ca9e2),
	.w6(32'h3a89fe3d),
	.w7(32'h3b708ba4),
	.w8(32'hbba732ff),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb08bc),
	.w1(32'h3a8d1528),
	.w2(32'hbc1adabb),
	.w3(32'hbba4c56d),
	.w4(32'hba4185e7),
	.w5(32'h3985e7ac),
	.w6(32'h3aab0694),
	.w7(32'h3ba9edb1),
	.w8(32'h3b37d018),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66b684),
	.w1(32'h3c2ee47b),
	.w2(32'hbc23ecdc),
	.w3(32'hba3cda10),
	.w4(32'h3c02cce0),
	.w5(32'h3af8e870),
	.w6(32'hbc0810f1),
	.w7(32'h3c35dfbd),
	.w8(32'h3c7d7d6b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fa491),
	.w1(32'hbc141f68),
	.w2(32'hbac56d87),
	.w3(32'h3c1284e4),
	.w4(32'h3b9f40a8),
	.w5(32'hbb1d2e3b),
	.w6(32'h3c7bcd67),
	.w7(32'hbadacd1b),
	.w8(32'h3b8353e2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9204b3),
	.w1(32'hbb16680a),
	.w2(32'hbbe719f2),
	.w3(32'h3b75db0c),
	.w4(32'hbc00e117),
	.w5(32'hba021275),
	.w6(32'h3c2dfd50),
	.w7(32'hb9d0cd4e),
	.w8(32'hbb13b35e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989c5a7),
	.w1(32'hbbc996e6),
	.w2(32'hbbd0a3f5),
	.w3(32'h3bc09d69),
	.w4(32'h3b0bad57),
	.w5(32'hbc085e51),
	.w6(32'h3a5e6c77),
	.w7(32'h3a8b2361),
	.w8(32'hb7268c6c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b339cdc),
	.w1(32'h3bbcd53f),
	.w2(32'hbbfad638),
	.w3(32'hbc127d26),
	.w4(32'hba57384d),
	.w5(32'hbb7e9bcf),
	.w6(32'hba656d01),
	.w7(32'hbb9880e3),
	.w8(32'h3bbc24f2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c023c91),
	.w1(32'h3c3bd969),
	.w2(32'h3b198d64),
	.w3(32'hbbfed692),
	.w4(32'hbc518600),
	.w5(32'h3b8d81af),
	.w6(32'hbb2394e3),
	.w7(32'hbb34d380),
	.w8(32'hbb2257f0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6db65e),
	.w1(32'hbbcef1b7),
	.w2(32'h3c2bbcdd),
	.w3(32'hbaf88264),
	.w4(32'h3b34d385),
	.w5(32'h38b0c11e),
	.w6(32'hbbda1289),
	.w7(32'h3c48459d),
	.w8(32'h3baf0493),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb2e69),
	.w1(32'h3be36cf0),
	.w2(32'h3b80e9f0),
	.w3(32'hbb87b2c7),
	.w4(32'h3b2a2a45),
	.w5(32'hb8cc6297),
	.w6(32'h3bcb30b8),
	.w7(32'h3b900bed),
	.w8(32'h3c229f9d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf5c0a),
	.w1(32'hbb86ec28),
	.w2(32'hba3e4966),
	.w3(32'hbb62e479),
	.w4(32'hbc9faae6),
	.w5(32'h3b90ae81),
	.w6(32'h3ba0601d),
	.w7(32'hbbd3807f),
	.w8(32'h3bdeb418),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6ac89),
	.w1(32'h3a52f434),
	.w2(32'h3aaf75a2),
	.w3(32'hb8587df5),
	.w4(32'h3ad2664b),
	.w5(32'h3ab615a1),
	.w6(32'h3cc83a09),
	.w7(32'hbac63f69),
	.w8(32'hbbb76688),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981e45d),
	.w1(32'hbb40959c),
	.w2(32'hbba59d8a),
	.w3(32'h3c0be944),
	.w4(32'h3ae69cf2),
	.w5(32'h3a327b3c),
	.w6(32'h3bb2ecc8),
	.w7(32'hbbb4b46e),
	.w8(32'hbadbf681),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81cfe3),
	.w1(32'hbb408cd9),
	.w2(32'hbb9d6302),
	.w3(32'h3b4b0169),
	.w4(32'hbc34da4d),
	.w5(32'hbabc59c9),
	.w6(32'h3c976a29),
	.w7(32'hbbc0dce7),
	.w8(32'h380b05e8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd48447),
	.w1(32'h3b8f973d),
	.w2(32'h3bbb3c3d),
	.w3(32'h3a8c6594),
	.w4(32'h3aee5672),
	.w5(32'hbae75029),
	.w6(32'h3cbc4019),
	.w7(32'h3b3457d2),
	.w8(32'hbba42300),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc574af7),
	.w1(32'hbcb358ca),
	.w2(32'hbb64d04e),
	.w3(32'h3d273c01),
	.w4(32'hbb977019),
	.w5(32'hbc0ae8b9),
	.w6(32'h3b96c3fb),
	.w7(32'h3c2bcf1b),
	.w8(32'hb9b36225),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0c7fa2),
	.w1(32'h3c82f2f2),
	.w2(32'h3ba4ffad),
	.w3(32'h3b81d170),
	.w4(32'h3c2e4e2d),
	.w5(32'h3b655560),
	.w6(32'hbc8314ef),
	.w7(32'hbc0590f8),
	.w8(32'hba2c90a2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905c5a2),
	.w1(32'hbbb8c90b),
	.w2(32'hbc697f30),
	.w3(32'h3c6533d3),
	.w4(32'h3c113334),
	.w5(32'h3b59bef8),
	.w6(32'h3c1d9f28),
	.w7(32'h3a919260),
	.w8(32'h3ce15acd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca96f27),
	.w1(32'h3cdb8f95),
	.w2(32'h3cb80dd2),
	.w3(32'hbcaa983b),
	.w4(32'hbd063d2a),
	.w5(32'h3b4d8c62),
	.w6(32'hbba52535),
	.w7(32'hbd18da8a),
	.w8(32'hbc30064c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c778c28),
	.w1(32'h3c76624e),
	.w2(32'h3c0636ae),
	.w3(32'hbc60f2ce),
	.w4(32'hbc06a5e7),
	.w5(32'hbb27f077),
	.w6(32'hbc0d12f2),
	.w7(32'hbbece08b),
	.w8(32'hbbd68fb1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaa91e),
	.w1(32'hbb1a719b),
	.w2(32'hba04d6fe),
	.w3(32'h3b930e03),
	.w4(32'h3b2d0520),
	.w5(32'h3b0b7af1),
	.w6(32'h3c13df49),
	.w7(32'hbb6397a7),
	.w8(32'hbb8dcb31),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae15850),
	.w1(32'hb973a0fc),
	.w2(32'hbb4037e0),
	.w3(32'h3b0dda99),
	.w4(32'h397dd53b),
	.w5(32'hbb3d5257),
	.w6(32'h3c07bed8),
	.w7(32'h3c58fe61),
	.w8(32'hbc175133),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9394ba),
	.w1(32'hbc6bf18a),
	.w2(32'hbc4d595d),
	.w3(32'h3bc4e619),
	.w4(32'h3c9b35ee),
	.w5(32'hbb96d812),
	.w6(32'hbb20f4e5),
	.w7(32'hbba2f0b7),
	.w8(32'h3b97c6f3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1011a0),
	.w1(32'h3aedc78b),
	.w2(32'hbb0231e9),
	.w3(32'hbc0e9fd7),
	.w4(32'hbbc447e3),
	.w5(32'h3b8f4e1f),
	.w6(32'h3b214448),
	.w7(32'hbb318ba5),
	.w8(32'hbc759103),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4e16d),
	.w1(32'hbd016d90),
	.w2(32'hbc088f1b),
	.w3(32'h3d221c3f),
	.w4(32'h3d0f3340),
	.w5(32'h3b3756b1),
	.w6(32'hbb530ed6),
	.w7(32'h3c9cd7a6),
	.w8(32'h3c6e1589),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c958345),
	.w1(32'hb9c2ca3d),
	.w2(32'h3c139392),
	.w3(32'h3a8c981f),
	.w4(32'h3c33757e),
	.w5(32'hbc1d7998),
	.w6(32'hbc763ed4),
	.w7(32'h3c3cab41),
	.w8(32'h3c199a3c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0693a),
	.w1(32'h3b0e2d59),
	.w2(32'h3ba64e27),
	.w3(32'hbad6a928),
	.w4(32'hbca4c4a8),
	.w5(32'h3b544ce0),
	.w6(32'hbb8e1499),
	.w7(32'hbc16809f),
	.w8(32'hbc4d1c8e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc228857),
	.w1(32'hbcb000c0),
	.w2(32'h3aea5143),
	.w3(32'h3d01b662),
	.w4(32'h3c4ac8e8),
	.w5(32'hbc004ea3),
	.w6(32'h3c4713b6),
	.w7(32'h3cb397a5),
	.w8(32'h3b2f303a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900a3e),
	.w1(32'h3b888c86),
	.w2(32'h39d51810),
	.w3(32'h3c079c0b),
	.w4(32'hb9c012e3),
	.w5(32'hbaf00d40),
	.w6(32'h3b2f6c1f),
	.w7(32'h3b86a8d5),
	.w8(32'hbc262d61),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7cfdbd),
	.w1(32'hbca3196b),
	.w2(32'hbb9513d5),
	.w3(32'h3ca2e012),
	.w4(32'h3beda53a),
	.w5(32'h3a8b8320),
	.w6(32'h3b633dd1),
	.w7(32'h3bbc97b8),
	.w8(32'hbc30f77c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53de4f),
	.w1(32'hbc1f06ff),
	.w2(32'hbba5d84e),
	.w3(32'h3c604a76),
	.w4(32'h3ca5157d),
	.w5(32'h3aa8c911),
	.w6(32'hbbf25a05),
	.w7(32'h3bf20173),
	.w8(32'h3b7d4200),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef81e0),
	.w1(32'h3af42c0b),
	.w2(32'h3b0b94cd),
	.w3(32'hba4b3797),
	.w4(32'hbbbaf3bd),
	.w5(32'h3b1f8987),
	.w6(32'hbb9a2748),
	.w7(32'hbc1c4bab),
	.w8(32'h399477c3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c492dd2),
	.w1(32'h379c7c18),
	.w2(32'hbada247a),
	.w3(32'hba481f02),
	.w4(32'hbb7965f5),
	.w5(32'h3a177625),
	.w6(32'hb7368cff),
	.w7(32'h3a5626d1),
	.w8(32'h3a007fde),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7502a1),
	.w1(32'h3b53ea48),
	.w2(32'h3acce2a5),
	.w3(32'hbb73e6b3),
	.w4(32'hbb5d1dc5),
	.w5(32'hbb9ea6e8),
	.w6(32'hbad8024b),
	.w7(32'hbbac4fae),
	.w8(32'hbb21f8d0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf490bd),
	.w1(32'h3c1bf946),
	.w2(32'hbc190e78),
	.w3(32'hbb979253),
	.w4(32'hbb35f522),
	.w5(32'hbb986e7f),
	.w6(32'h39e9efd0),
	.w7(32'hbc3f11dc),
	.w8(32'h3bed8f92),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32f188),
	.w1(32'h3cbaf002),
	.w2(32'h3abdd347),
	.w3(32'hbc5787af),
	.w4(32'hbc53fe6b),
	.w5(32'h3b6846df),
	.w6(32'h3a852e6a),
	.w7(32'hbc12711c),
	.w8(32'h3c16604c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e17a7),
	.w1(32'hba252685),
	.w2(32'h3bd80e51),
	.w3(32'h3a0b106b),
	.w4(32'h3653d8dc),
	.w5(32'h3a9abca0),
	.w6(32'h3d3f38fc),
	.w7(32'h3c959c06),
	.w8(32'h3bdb41e4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7fce3),
	.w1(32'h3c3592fb),
	.w2(32'h3b99f051),
	.w3(32'hbc401617),
	.w4(32'hbc182cc5),
	.w5(32'hbb85eda4),
	.w6(32'hbc0ec252),
	.w7(32'hbc331c1f),
	.w8(32'hbc0fad75),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60ba43),
	.w1(32'h3c0546e4),
	.w2(32'h3b160ce3),
	.w3(32'h3c8fa926),
	.w4(32'h3caf30d0),
	.w5(32'h3b20627e),
	.w6(32'hbbbeba4c),
	.w7(32'h3c6e3995),
	.w8(32'h3bef8037),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd35b),
	.w1(32'hbba3879b),
	.w2(32'h3c84569b),
	.w3(32'h3cba8bcd),
	.w4(32'h3b34b084),
	.w5(32'h3bb63ca9),
	.w6(32'h3c7aec92),
	.w7(32'h3be8901c),
	.w8(32'hbb877c20),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60521b),
	.w1(32'h3b6647fa),
	.w2(32'h3c8987df),
	.w3(32'hbc950d37),
	.w4(32'h3c1037f4),
	.w5(32'h3b2b9dd3),
	.w6(32'hbb84f5bc),
	.w7(32'h3c20dd5a),
	.w8(32'h3c8e956a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c897477),
	.w1(32'h3d262c81),
	.w2(32'h3c5702ba),
	.w3(32'hbbb87f55),
	.w4(32'hb8b8a360),
	.w5(32'h3adc6421),
	.w6(32'h3c896a79),
	.w7(32'hbc579646),
	.w8(32'hbbb135c3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d86d2),
	.w1(32'hbcbf9d6c),
	.w2(32'hbcf6b7f8),
	.w3(32'h3c767dd4),
	.w4(32'h3b934aea),
	.w5(32'hbc6faebe),
	.w6(32'h3bc10165),
	.w7(32'h3bf9154b),
	.w8(32'hbb4057ad),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45059c),
	.w1(32'h3c9b04c2),
	.w2(32'h3c84afe8),
	.w3(32'h3bc2e809),
	.w4(32'hbaf53592),
	.w5(32'hbb201b3b),
	.w6(32'h3c676675),
	.w7(32'h3ba0c6a1),
	.w8(32'h3b87a55b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce7b90a),
	.w1(32'h3c7d010a),
	.w2(32'h3c1db064),
	.w3(32'hbb48946c),
	.w4(32'hbcb96768),
	.w5(32'hbb667649),
	.w6(32'h3d027c32),
	.w7(32'h3bc04c36),
	.w8(32'hbcc90aef),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dfe8a),
	.w1(32'hbcecb591),
	.w2(32'h3b85633e),
	.w3(32'h3d04f9d5),
	.w4(32'h3c9301ec),
	.w5(32'hbbcb478d),
	.w6(32'h3c44cd33),
	.w7(32'h3ca1b0b3),
	.w8(32'h3bc00b74),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77ae99),
	.w1(32'h3abe8f1b),
	.w2(32'h3b133004),
	.w3(32'h3bdb9e53),
	.w4(32'h3c287ca8),
	.w5(32'hbb566e6f),
	.w6(32'hbc1d0afc),
	.w7(32'h3befff4f),
	.w8(32'h3b2d42b3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc695279),
	.w1(32'hbab331dc),
	.w2(32'h3c8d371f),
	.w3(32'h3c3ee50c),
	.w4(32'h3be8edc4),
	.w5(32'h3c5d3443),
	.w6(32'h3b5b51b4),
	.w7(32'h3c3fefff),
	.w8(32'hbb1c0462),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60c6b3),
	.w1(32'h3c8a17be),
	.w2(32'h3b23b39d),
	.w3(32'hbd2d728e),
	.w4(32'h3c454151),
	.w5(32'h3c7d15ef),
	.w6(32'hbd18a1c2),
	.w7(32'hbcbef5a3),
	.w8(32'h3c0ae1f7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a68d7),
	.w1(32'hbc6046d2),
	.w2(32'hbaf77223),
	.w3(32'h3b4f5742),
	.w4(32'h3a448e0c),
	.w5(32'hbb9a40c2),
	.w6(32'h3ba33a9f),
	.w7(32'hba4fcea0),
	.w8(32'hbcabaa89),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2068f),
	.w1(32'h3b1543f2),
	.w2(32'h3b9ba223),
	.w3(32'hbbb0a105),
	.w4(32'hba3cf140),
	.w5(32'h3afdeab8),
	.w6(32'h3ba3c959),
	.w7(32'hbbfa1c8b),
	.w8(32'hbc12eeab),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b618b75),
	.w1(32'h3c25bb85),
	.w2(32'h3c2615ee),
	.w3(32'hbbe29aee),
	.w4(32'h3ced2285),
	.w5(32'h3c80666c),
	.w6(32'hbc34141b),
	.w7(32'h3c5d39cd),
	.w8(32'h3c279e1e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb19f4),
	.w1(32'hbb0ee29a),
	.w2(32'h37605d0b),
	.w3(32'hba5ae2c3),
	.w4(32'hba688945),
	.w5(32'h3ace473b),
	.w6(32'h3bcb3245),
	.w7(32'h3adc6b6a),
	.w8(32'h3b66d3b6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0736d6),
	.w1(32'h3c13b555),
	.w2(32'h3bbcc463),
	.w3(32'hbc93dc13),
	.w4(32'h3b9bd8e6),
	.w5(32'h3c985f36),
	.w6(32'hbd107150),
	.w7(32'h3c28b178),
	.w8(32'hbaa9195e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab00653),
	.w1(32'h3bae3423),
	.w2(32'h3b3772e9),
	.w3(32'hbbac8e13),
	.w4(32'hbb1d0eda),
	.w5(32'h3bb8f912),
	.w6(32'hbc67896e),
	.w7(32'hbb5c20e8),
	.w8(32'h3bd8d822),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba148c7a),
	.w1(32'hba6e6e0f),
	.w2(32'h3b6d9fac),
	.w3(32'h3b17a5cc),
	.w4(32'hbabac9fa),
	.w5(32'h3abca526),
	.w6(32'hbb032cdc),
	.w7(32'hbb299242),
	.w8(32'h3a08bd58),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a9df9),
	.w1(32'h3ba32513),
	.w2(32'h3b534b78),
	.w3(32'h3a7f196c),
	.w4(32'hbb86da1c),
	.w5(32'hbad10f9e),
	.w6(32'h3bc07304),
	.w7(32'hba780527),
	.w8(32'hbbdc54ff),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f0483),
	.w1(32'h3bc80de0),
	.w2(32'h3bb04526),
	.w3(32'h3c200dac),
	.w4(32'h3c406d9a),
	.w5(32'h3a9537ec),
	.w6(32'hbad4dc89),
	.w7(32'h3c0ca34d),
	.w8(32'h3a69570e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd33c66),
	.w1(32'h3b92229b),
	.w2(32'h3b8c9648),
	.w3(32'hba350e50),
	.w4(32'hbb39831b),
	.w5(32'h3bd95969),
	.w6(32'h3b84955f),
	.w7(32'hbb3ad056),
	.w8(32'hbba5c30c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a680eda),
	.w1(32'hbb8915fa),
	.w2(32'h3b651c3e),
	.w3(32'h3c86c60a),
	.w4(32'h3a8e1371),
	.w5(32'hbafbd7d6),
	.w6(32'h3bad9884),
	.w7(32'h3b3bed64),
	.w8(32'hbb90a565),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20cd9c),
	.w1(32'hbba6fa71),
	.w2(32'hbb83bfa8),
	.w3(32'hbb4b5072),
	.w4(32'hbb9d2f4f),
	.w5(32'hbb8ed0c2),
	.w6(32'hbbb1e252),
	.w7(32'hbb98dc44),
	.w8(32'hbc0d83db),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cd3a6),
	.w1(32'h3c328eb9),
	.w2(32'h3c857bf9),
	.w3(32'hbc521378),
	.w4(32'hb9fcdff7),
	.w5(32'h3c5b79e2),
	.w6(32'hbc88e39e),
	.w7(32'hbc771cc7),
	.w8(32'h3c2fd757),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09c3d0),
	.w1(32'hba27becc),
	.w2(32'hbb58657c),
	.w3(32'h3be68f47),
	.w4(32'hbbf39918),
	.w5(32'hbc61bd93),
	.w6(32'h3beb6777),
	.w7(32'h3bb8fada),
	.w8(32'hbc54fc89),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c286430),
	.w1(32'h3b3d1f6b),
	.w2(32'hbb1b41c2),
	.w3(32'hbb397ae8),
	.w4(32'h3baa1920),
	.w5(32'h3b2c1d48),
	.w6(32'hbb16ce7e),
	.w7(32'h3b0e99ce),
	.w8(32'h3a666b80),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cebdea),
	.w1(32'h398f1869),
	.w2(32'hbafd31c5),
	.w3(32'hbad42231),
	.w4(32'h3b45c78f),
	.w5(32'hbb00dce6),
	.w6(32'hbba68441),
	.w7(32'h3af22d41),
	.w8(32'hbb017188),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2826dc),
	.w1(32'hb98b9589),
	.w2(32'h37e57608),
	.w3(32'h3a1fe32e),
	.w4(32'hbb084e0b),
	.w5(32'h3acd09bf),
	.w6(32'h3a812054),
	.w7(32'hb9f83bc9),
	.w8(32'h3b83b73b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0d28a),
	.w1(32'h3a89a00d),
	.w2(32'h3b0fc98a),
	.w3(32'hbbc90025),
	.w4(32'h3b3d9423),
	.w5(32'h3a4ab5c5),
	.w6(32'h3b864b16),
	.w7(32'hba09fc7c),
	.w8(32'hbb13eb83),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a3a5d),
	.w1(32'h3a1e741e),
	.w2(32'h3b9c758c),
	.w3(32'h3b2478c5),
	.w4(32'hbb435d59),
	.w5(32'h3a725f66),
	.w6(32'h3ae87b5e),
	.w7(32'h3ac5cbd8),
	.w8(32'hbbe4d7bd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad76554),
	.w1(32'hbc0105ca),
	.w2(32'hbaa9f89a),
	.w3(32'hb9c02207),
	.w4(32'hbb44a21d),
	.w5(32'h3a5797d3),
	.w6(32'h3b18729b),
	.w7(32'hbba9979e),
	.w8(32'hb8ea3686),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb057299),
	.w1(32'hbb43ef8e),
	.w2(32'hba220434),
	.w3(32'hbb5111f2),
	.w4(32'h3a8c5e61),
	.w5(32'hbb4bdb91),
	.w6(32'hbbc4ec36),
	.w7(32'hba81e6a9),
	.w8(32'hba9dc92c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a119e),
	.w1(32'h39ec62e4),
	.w2(32'h3a64adfb),
	.w3(32'hbba276b0),
	.w4(32'h3c08d081),
	.w5(32'h3becc4f9),
	.w6(32'hbc2a0153),
	.w7(32'hb964b36c),
	.w8(32'h3c208343),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b323234),
	.w1(32'hbc029519),
	.w2(32'hbb790185),
	.w3(32'h3c28ce40),
	.w4(32'hbc709633),
	.w5(32'hbc06dfa7),
	.w6(32'h3c56a944),
	.w7(32'hbc459a4f),
	.w8(32'hbc832b60),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb893532),
	.w1(32'hbb100f65),
	.w2(32'hba5e8a1d),
	.w3(32'hb919de0b),
	.w4(32'hbb3b6b49),
	.w5(32'h39092396),
	.w6(32'hbb188d80),
	.w7(32'hbafc6587),
	.w8(32'hbb352200),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba947c51),
	.w1(32'h39a97bdf),
	.w2(32'hbb084981),
	.w3(32'h3b1cacaa),
	.w4(32'h3a956df9),
	.w5(32'hb9ba8ffb),
	.w6(32'h3b5ff773),
	.w7(32'h3aa3aef4),
	.w8(32'h3a5db274),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7b82c),
	.w1(32'h3822ae9d),
	.w2(32'hba34f3ff),
	.w3(32'hbab4544e),
	.w4(32'h3a9b516f),
	.w5(32'hb99e6463),
	.w6(32'h3b4e77c1),
	.w7(32'h3a56b82f),
	.w8(32'h3a56aa13),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa22420),
	.w1(32'h3b1bcd61),
	.w2(32'h3aff01f5),
	.w3(32'hbadc373d),
	.w4(32'h3ad59234),
	.w5(32'hbb50c4aa),
	.w6(32'h3996f6c2),
	.w7(32'h3b062552),
	.w8(32'hba51f6c2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c01aa),
	.w1(32'h3cb53bf2),
	.w2(32'hbb235aa6),
	.w3(32'hbb25187e),
	.w4(32'h3cbe1e91),
	.w5(32'h3b1dc267),
	.w6(32'hbb7bac3a),
	.w7(32'hbb91fe65),
	.w8(32'h3b646498),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c5c67),
	.w1(32'h3b1e361d),
	.w2(32'h3ade46a3),
	.w3(32'h3b86e6c2),
	.w4(32'h3b91810f),
	.w5(32'h3abc139c),
	.w6(32'hbbbc9792),
	.w7(32'h3c14010c),
	.w8(32'h3b9afebd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810761),
	.w1(32'h3a4fbe99),
	.w2(32'h3a0e3ed7),
	.w3(32'hbb27641a),
	.w4(32'hb9d1bb64),
	.w5(32'hba8f2872),
	.w6(32'hbbdafc24),
	.w7(32'h3a314900),
	.w8(32'hba271d87),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff5dc9),
	.w1(32'hbbdf0244),
	.w2(32'h39bf9bb4),
	.w3(32'hb97a7ebf),
	.w4(32'h3b190faa),
	.w5(32'hbb1bea1f),
	.w6(32'hbbef104e),
	.w7(32'h3b99869c),
	.w8(32'h3b959cab),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99813cc),
	.w1(32'hb7b40ab3),
	.w2(32'h3a0dc6f6),
	.w3(32'h3a72a154),
	.w4(32'hbab41884),
	.w5(32'hbafc5262),
	.w6(32'h3ba5cd19),
	.w7(32'hba81f93b),
	.w8(32'hbbd9b413),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09563d),
	.w1(32'hbb73c815),
	.w2(32'hbb8107ef),
	.w3(32'h3af569f3),
	.w4(32'hbb56352b),
	.w5(32'hbb8691be),
	.w6(32'h3b211ea2),
	.w7(32'h3b3d3373),
	.w8(32'h3b1dbd8a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b5f04),
	.w1(32'hbb88ff63),
	.w2(32'h3b421e70),
	.w3(32'h3c149243),
	.w4(32'hbc2ddbea),
	.w5(32'hbb381b87),
	.w6(32'h3c554dd5),
	.w7(32'hbb30230d),
	.w8(32'hbc0348a1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ab433),
	.w1(32'h3bbd9f88),
	.w2(32'h3baf6a13),
	.w3(32'h3c12bf83),
	.w4(32'h3c8ae9ed),
	.w5(32'h3a30902e),
	.w6(32'hbb801445),
	.w7(32'h3c4eeb55),
	.w8(32'h3c223fde),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cab73),
	.w1(32'hbb86ab12),
	.w2(32'hbad02bbe),
	.w3(32'hbb93728b),
	.w4(32'hbc1455ba),
	.w5(32'hbc0ef202),
	.w6(32'hbb8c5858),
	.w7(32'hbc0f401e),
	.w8(32'hbc6cfb3e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09c35e),
	.w1(32'hbb4c02fd),
	.w2(32'h3a9e101a),
	.w3(32'hbb96c952),
	.w4(32'h3a73e4be),
	.w5(32'h3bb85ef2),
	.w6(32'hbb27a7a9),
	.w7(32'hbb23131f),
	.w8(32'h3a833c8b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c330ed7),
	.w1(32'h3c3a0709),
	.w2(32'h3c0e28fa),
	.w3(32'h3ad92dfd),
	.w4(32'h3c92b7d5),
	.w5(32'h3c06b1a0),
	.w6(32'h3ac52d66),
	.w7(32'h3c805175),
	.w8(32'h3c5cd324),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976d7a8),
	.w1(32'h3ba504c9),
	.w2(32'h3ba16c8d),
	.w3(32'hbbbabadc),
	.w4(32'h3af3fa67),
	.w5(32'h3b8ad2b4),
	.w6(32'hbb5f3146),
	.w7(32'hbbed2acd),
	.w8(32'hba0ac7b0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98eba7),
	.w1(32'hbab88471),
	.w2(32'hba9844ea),
	.w3(32'h3becb5e0),
	.w4(32'h3ba927d9),
	.w5(32'h3a56fb79),
	.w6(32'hbc182ff6),
	.w7(32'h3c1c9c68),
	.w8(32'h3b53ef45),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c185711),
	.w1(32'h3be0b882),
	.w2(32'h3adfe4c6),
	.w3(32'h3ac13de2),
	.w4(32'h3a31c1a0),
	.w5(32'h3b40042a),
	.w6(32'h3871c5d9),
	.w7(32'hbad6726c),
	.w8(32'h39bb38c4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae961a),
	.w1(32'hbbec3b32),
	.w2(32'h3bc01c1a),
	.w3(32'h3c1f73c5),
	.w4(32'hbc99b756),
	.w5(32'hbc099108),
	.w6(32'h3cac8c37),
	.w7(32'hbc3ac1d0),
	.w8(32'hbc8b6235),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94a28f),
	.w1(32'h3b45d2bb),
	.w2(32'hbabc2a83),
	.w3(32'h3b9e06df),
	.w4(32'h3a316c16),
	.w5(32'h3b05a35e),
	.w6(32'h3a373dd2),
	.w7(32'h3ac973a5),
	.w8(32'hbb7132ea),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad01c6b),
	.w1(32'hba04bfc5),
	.w2(32'h3ab819fb),
	.w3(32'hb91260bf),
	.w4(32'h3ab7abd9),
	.w5(32'hbb5f8801),
	.w6(32'h3b06f58a),
	.w7(32'h39f68880),
	.w8(32'hbacb732d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7742e7),
	.w1(32'hbb224562),
	.w2(32'hbaceb870),
	.w3(32'hba9bc87e),
	.w4(32'hba9ee3d2),
	.w5(32'hbb7ca238),
	.w6(32'hbb2fe4cc),
	.w7(32'hb983b72b),
	.w8(32'hbb66e9f3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb6104),
	.w1(32'hbb918531),
	.w2(32'h3ae30831),
	.w3(32'hbbc7626d),
	.w4(32'hba3f9e03),
	.w5(32'h3902e24d),
	.w6(32'hbbe1a664),
	.w7(32'hbb49bb32),
	.w8(32'hbbdac830),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26f9e3),
	.w1(32'hbb8b89a7),
	.w2(32'h3bd86cd1),
	.w3(32'hba73b5fb),
	.w4(32'hbb8a261a),
	.w5(32'hbae756fe),
	.w6(32'hbbc0f05f),
	.w7(32'hbc065dce),
	.w8(32'hbbe3dc56),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a3bbf),
	.w1(32'h3aab24f7),
	.w2(32'hbb479a7c),
	.w3(32'hba8e2e17),
	.w4(32'h3b54e35b),
	.w5(32'h3b83e743),
	.w6(32'hbba9b0a2),
	.w7(32'hb89bc2cf),
	.w8(32'hba69e1fe),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1442aa),
	.w1(32'h3a8dd449),
	.w2(32'h3b2403ba),
	.w3(32'h3b4cc871),
	.w4(32'hbb071c35),
	.w5(32'hbb006b47),
	.w6(32'h3b50aa1b),
	.w7(32'hba6e6cb3),
	.w8(32'hba998dc9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b802c5a),
	.w1(32'h3a7d0161),
	.w2(32'h3b87cdb1),
	.w3(32'h3c15cbaa),
	.w4(32'h3a9489a7),
	.w5(32'hb95b6830),
	.w6(32'h3a1a8552),
	.w7(32'h3be2398e),
	.w8(32'hbb779e82),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43c9f),
	.w1(32'h3ab98bf3),
	.w2(32'h3aaaa219),
	.w3(32'h3b57528c),
	.w4(32'h38858ba0),
	.w5(32'h38a336d0),
	.w6(32'hbb1ad68f),
	.w7(32'hbb3ae61a),
	.w8(32'hbbef24e1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64bd33),
	.w1(32'h3b459cf2),
	.w2(32'h3c0a65b2),
	.w3(32'h3b9d8742),
	.w4(32'h3c4187ed),
	.w5(32'h3c8b3ac7),
	.w6(32'hbb102713),
	.w7(32'h3c36593b),
	.w8(32'h3c06bdca),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb46e17),
	.w1(32'hbbab126d),
	.w2(32'h3ca274db),
	.w3(32'h3c2d8af6),
	.w4(32'hbc3592cd),
	.w5(32'h3b8cbe5d),
	.w6(32'h3d0b43dd),
	.w7(32'hbb631e42),
	.w8(32'hbbbbe105),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdda05d),
	.w1(32'h3ba7dff3),
	.w2(32'hbaa0ec5b),
	.w3(32'h3be3c2df),
	.w4(32'h3b41a30a),
	.w5(32'hbb5e684e),
	.w6(32'h3c02b6df),
	.w7(32'h3b22e1b9),
	.w8(32'hbac515d0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a326b),
	.w1(32'hbb80d914),
	.w2(32'hb6a6079e),
	.w3(32'hbb1b833f),
	.w4(32'h3ad25e56),
	.w5(32'h39580351),
	.w6(32'hbb00f1b6),
	.w7(32'h3b0a13b5),
	.w8(32'hbac04706),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f1431),
	.w1(32'hbb2ba267),
	.w2(32'h3b3f4af0),
	.w3(32'hbbb2d428),
	.w4(32'hbbb730db),
	.w5(32'h3c08e41f),
	.w6(32'hbb4ac212),
	.w7(32'hbb87716c),
	.w8(32'h3b3b3244),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba357c8),
	.w1(32'hbbe23347),
	.w2(32'h3c2420b7),
	.w3(32'h3aab87d1),
	.w4(32'hbc06a79b),
	.w5(32'hba89fc12),
	.w6(32'h3cad86ca),
	.w7(32'hbb1f55e1),
	.w8(32'hbbaeec94),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b326bb2),
	.w1(32'hba23b284),
	.w2(32'h3acc1bfb),
	.w3(32'h3b2cf6bf),
	.w4(32'h3b00303a),
	.w5(32'h3b00148b),
	.w6(32'h3afedc1b),
	.w7(32'hbb0b21eb),
	.w8(32'hbba31e71),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954edb4),
	.w1(32'hbb1b5c58),
	.w2(32'h3b009d54),
	.w3(32'h3baa5825),
	.w4(32'h3bd80dd1),
	.w5(32'h3ad66827),
	.w6(32'h3b18c777),
	.w7(32'h3c26f990),
	.w8(32'h3b53d759),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc67c3b),
	.w1(32'h3abacc51),
	.w2(32'hbb83279e),
	.w3(32'h37867af4),
	.w4(32'h398c2196),
	.w5(32'hbb6e8307),
	.w6(32'h3b46a6de),
	.w7(32'h39e90010),
	.w8(32'hbb83daa0),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcacf1c),
	.w1(32'hbae0c7cb),
	.w2(32'h3882e78a),
	.w3(32'h3ab8469e),
	.w4(32'h3b8cc179),
	.w5(32'h3aaa589f),
	.w6(32'hbbfba261),
	.w7(32'h3b86a3e8),
	.w8(32'h3998a89f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba610e0),
	.w1(32'hb9f1d16d),
	.w2(32'h3ad54714),
	.w3(32'hbbc8d831),
	.w4(32'hbb8c89dc),
	.w5(32'h3c100d76),
	.w6(32'hbb2d3f59),
	.w7(32'hbbfc26fa),
	.w8(32'hbb95381b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf36b92),
	.w1(32'hbb5909b0),
	.w2(32'h3b80c369),
	.w3(32'hbb76a8f2),
	.w4(32'hbc47b4bb),
	.w5(32'h39c36828),
	.w6(32'h3c79d2f7),
	.w7(32'hbc5b2e4e),
	.w8(32'hbac0b602),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1f880),
	.w1(32'h3b86b24e),
	.w2(32'h3b94a1d7),
	.w3(32'h3b83f8dd),
	.w4(32'h3ad9d3c7),
	.w5(32'h3bc80d1f),
	.w6(32'hbbb4a74c),
	.w7(32'h3aaf72d2),
	.w8(32'h3a927911),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65caa4),
	.w1(32'h3bdf6bf7),
	.w2(32'h3c41bde9),
	.w3(32'h3c240daf),
	.w4(32'h3be2f629),
	.w5(32'h3b1f26fb),
	.w6(32'h3ca3d90e),
	.w7(32'h3baf5fe5),
	.w8(32'h3b83a573),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d1a99),
	.w1(32'h3a8b8aea),
	.w2(32'h39522b51),
	.w3(32'h3b8098bb),
	.w4(32'h3b85d076),
	.w5(32'hbb47528a),
	.w6(32'h3ab12e5b),
	.w7(32'h3ac86b56),
	.w8(32'hbaff539c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7600ec),
	.w1(32'hbaf1983d),
	.w2(32'hbae42b81),
	.w3(32'hba864cca),
	.w4(32'hba6ce693),
	.w5(32'h3ba797ce),
	.w6(32'hba9c0e80),
	.w7(32'hbb02aaf7),
	.w8(32'hb986f12f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0126c),
	.w1(32'hbb5f28d0),
	.w2(32'hbbbf7ecc),
	.w3(32'h3b4799fb),
	.w4(32'hbbc48707),
	.w5(32'h3b127c7b),
	.w6(32'h3ca118c3),
	.w7(32'hbb3e8c08),
	.w8(32'hbb8d397f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60e3cc),
	.w1(32'h3c3335db),
	.w2(32'h3cb0749b),
	.w3(32'hbb71b65d),
	.w4(32'h3c84188d),
	.w5(32'h3beb9eda),
	.w6(32'hbc5ee41b),
	.w7(32'hbb4911e8),
	.w8(32'h3bfc3329),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2c17),
	.w1(32'h3b3ef18e),
	.w2(32'h3b4aa92d),
	.w3(32'h3b9990bf),
	.w4(32'h3acd43cc),
	.w5(32'h3b60e712),
	.w6(32'h3b77a0c6),
	.w7(32'h3b85f89d),
	.w8(32'h3bec3728),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b961c5e),
	.w1(32'h3b1bbf46),
	.w2(32'h3b6982b0),
	.w3(32'h3bd15642),
	.w4(32'h3a859f7b),
	.w5(32'hbbb5ce71),
	.w6(32'h3c4ca64b),
	.w7(32'hba53a353),
	.w8(32'hbc322910),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8a17c),
	.w1(32'hbbd8482d),
	.w2(32'h3b9cd360),
	.w3(32'h3bb4a90c),
	.w4(32'h3a02df45),
	.w5(32'hbc035616),
	.w6(32'hbaab6788),
	.w7(32'h3b7fd80d),
	.w8(32'hbc5c5034),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4652d9),
	.w1(32'hbc48dff9),
	.w2(32'hbac053b6),
	.w3(32'h39b7914e),
	.w4(32'hbbf235fa),
	.w5(32'h3bf1b522),
	.w6(32'h3bd1497d),
	.w7(32'h3b3d1a4a),
	.w8(32'h3bdef39f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c239b60),
	.w1(32'h3c18b96f),
	.w2(32'h3b4a7697),
	.w3(32'h3c242d39),
	.w4(32'h3b9f6b70),
	.w5(32'hba3da4e4),
	.w6(32'h3b987b2a),
	.w7(32'h3c50e0bc),
	.w8(32'hbb44e587),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb081d2),
	.w1(32'h3b585127),
	.w2(32'h3b6c4ba6),
	.w3(32'h3be1a717),
	.w4(32'h3c2bdc7b),
	.w5(32'hba8cfbda),
	.w6(32'hbb87c80c),
	.w7(32'h3c87fa97),
	.w8(32'h3baf299d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394606ab),
	.w1(32'hb9d03a95),
	.w2(32'hba0bd92c),
	.w3(32'hba25a556),
	.w4(32'hb7cc9b37),
	.w5(32'h3a91b4d5),
	.w6(32'hbb370df7),
	.w7(32'hba5013bb),
	.w8(32'h3b12d15f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a264e),
	.w1(32'h3abaf0c3),
	.w2(32'h3b9ddc91),
	.w3(32'h3c849404),
	.w4(32'h3a57fc2c),
	.w5(32'h3ad0edee),
	.w6(32'h3c16a09c),
	.w7(32'h3bd1c93a),
	.w8(32'hbad02c76),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e1849),
	.w1(32'hba5910de),
	.w2(32'h3b06636c),
	.w3(32'h3afb875b),
	.w4(32'hb9810b07),
	.w5(32'hbb7bb6b7),
	.w6(32'h3b623ed4),
	.w7(32'h3a83ce36),
	.w8(32'hbb110d01),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb010914),
	.w1(32'hbb189627),
	.w2(32'hbb6da3f5),
	.w3(32'hbbaf6608),
	.w4(32'h3aba3039),
	.w5(32'hba816d2d),
	.w6(32'hbbf81cda),
	.w7(32'hbb427fe9),
	.w8(32'h3bed0c8f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e67e6),
	.w1(32'hbb48532b),
	.w2(32'h3a6b23ff),
	.w3(32'h3af8cb74),
	.w4(32'h3b87fb99),
	.w5(32'hbba90a81),
	.w6(32'hba574f18),
	.w7(32'h3a476ed2),
	.w8(32'hbba4c150),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb71ff),
	.w1(32'hb90160f5),
	.w2(32'h3b220d0d),
	.w3(32'h3c596c36),
	.w4(32'hbc1270d0),
	.w5(32'hbb1d4611),
	.w6(32'h3b51eab7),
	.w7(32'hbb1dfb06),
	.w8(32'hbc4423a6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba757f25),
	.w1(32'hb90a9abf),
	.w2(32'hbb591513),
	.w3(32'hbb966dcb),
	.w4(32'hbab6df7f),
	.w5(32'hba8d2914),
	.w6(32'h3b970bb8),
	.w7(32'hbb07f048),
	.w8(32'h3b31f2f2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee80ce),
	.w1(32'h3b7122fb),
	.w2(32'hbac3d7a3),
	.w3(32'h39a70ddd),
	.w4(32'h3b1eb78d),
	.w5(32'h3b9cf407),
	.w6(32'hbab4dcf9),
	.w7(32'h3abc9160),
	.w8(32'hbb4c3deb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b6557),
	.w1(32'hbbdb1a3e),
	.w2(32'h3b83a670),
	.w3(32'hbb50aa32),
	.w4(32'hbbf4a076),
	.w5(32'h3bd8ea6e),
	.w6(32'h3c9b4c3e),
	.w7(32'hbc04b880),
	.w8(32'hbadf21e2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b132b8c),
	.w1(32'h3c6b1201),
	.w2(32'h3c1bc81a),
	.w3(32'h3bf4f79d),
	.w4(32'h3c554f20),
	.w5(32'h3c443968),
	.w6(32'h3cbe1128),
	.w7(32'h3bdad473),
	.w8(32'h3bd6e353),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b104b),
	.w1(32'h3ba6b51d),
	.w2(32'h3c367221),
	.w3(32'hbc54d11b),
	.w4(32'h3bab23f7),
	.w5(32'h3bad4789),
	.w6(32'hbc823a43),
	.w7(32'hbba02741),
	.w8(32'h3c03691d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb254e),
	.w1(32'hbb0c7558),
	.w2(32'hba4d0648),
	.w3(32'h3aaa2c49),
	.w4(32'hbb23cb94),
	.w5(32'hbc29ea35),
	.w6(32'h3b586fcf),
	.w7(32'hba045616),
	.w8(32'hbbc178fd),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c061156),
	.w1(32'h3b6acf9d),
	.w2(32'h3ac12763),
	.w3(32'hbbcdf6f5),
	.w4(32'h3c929a52),
	.w5(32'h3b49ee58),
	.w6(32'hbc9aa973),
	.w7(32'h3c4e5809),
	.w8(32'h3c0affc3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974007),
	.w1(32'hbbbbe8e2),
	.w2(32'h3c82cfb0),
	.w3(32'h3cabb961),
	.w4(32'hbc54b38c),
	.w5(32'h3bb31c5c),
	.w6(32'h3c9c6a58),
	.w7(32'hba265448),
	.w8(32'hbc241aad),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb316a5e),
	.w1(32'h3a90e007),
	.w2(32'h3bf278eb),
	.w3(32'h3b1b1c7b),
	.w4(32'h3bee58d4),
	.w5(32'h3bea3917),
	.w6(32'hbac65e48),
	.w7(32'h3c11b4b2),
	.w8(32'hbb122203),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6061cc),
	.w1(32'h3a1a85d7),
	.w2(32'h3b17d965),
	.w3(32'hbb70cd9c),
	.w4(32'hbb3ae7df),
	.w5(32'h3c2e34b5),
	.w6(32'h3a866997),
	.w7(32'hbbbac87f),
	.w8(32'h39c434f2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb24c94),
	.w1(32'hbb5dd760),
	.w2(32'h3bb2a921),
	.w3(32'hba919fb6),
	.w4(32'hbb1f8ecd),
	.w5(32'h3b628bc8),
	.w6(32'h3c8a9be0),
	.w7(32'hba89f671),
	.w8(32'h3ac8b804),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf464a),
	.w1(32'hba5d6ed0),
	.w2(32'hbb24aa75),
	.w3(32'hbbdd1fb0),
	.w4(32'hbaadaac4),
	.w5(32'hba290624),
	.w6(32'h3bad0ec8),
	.w7(32'hbb66243d),
	.w8(32'h3aace2b5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c785ddd),
	.w1(32'h3c3e2df6),
	.w2(32'h3c192fe2),
	.w3(32'h3b4fceb6),
	.w4(32'h3c71c169),
	.w5(32'h3b2fbdf0),
	.w6(32'hbc233679),
	.w7(32'h3b856ef0),
	.w8(32'h3b9c60ec),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9240489),
	.w1(32'h3a6358eb),
	.w2(32'h383a1b58),
	.w3(32'hba10ec73),
	.w4(32'h3afc744d),
	.w5(32'hbb84c0ab),
	.w6(32'hbb99323f),
	.w7(32'hb9d01f51),
	.w8(32'hbad9583c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d9d87),
	.w1(32'hbb9033de),
	.w2(32'hbb825b41),
	.w3(32'hbb87f6dd),
	.w4(32'hbbbc45ef),
	.w5(32'hbb3e29f3),
	.w6(32'hba269927),
	.w7(32'hbbf45745),
	.w8(32'hbb455d5f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beab412),
	.w1(32'h39b9c4cd),
	.w2(32'hbad3cf64),
	.w3(32'hb9c004d4),
	.w4(32'h3a7684c7),
	.w5(32'h3aefbf3b),
	.w6(32'hba084c64),
	.w7(32'hbb4eb873),
	.w8(32'h3ac7a288),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4cd44),
	.w1(32'h3be07159),
	.w2(32'h3bcca8d2),
	.w3(32'h3bc0442e),
	.w4(32'h3c512b62),
	.w5(32'h3b851770),
	.w6(32'hbc0c257f),
	.w7(32'h3c22b5c5),
	.w8(32'h3baea7c6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa936),
	.w1(32'hbb41bcdf),
	.w2(32'h3a0f3616),
	.w3(32'hbc00d0bb),
	.w4(32'hbaa52410),
	.w5(32'h3bdcff73),
	.w6(32'hbb82cc0b),
	.w7(32'h3a679c4f),
	.w8(32'h3c0a69db),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1597a9),
	.w1(32'h3b8047cd),
	.w2(32'hbb035ad7),
	.w3(32'h3b805b99),
	.w4(32'hbaa3b890),
	.w5(32'hba92dbbc),
	.w6(32'h3b0157dc),
	.w7(32'hbaa2d8e1),
	.w8(32'h3a81d681),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf189a0),
	.w1(32'hbb40da23),
	.w2(32'hbc258425),
	.w3(32'hbb9243b2),
	.w4(32'hbb82d48c),
	.w5(32'h3957669f),
	.w6(32'hb82afe10),
	.w7(32'h3b0f3cea),
	.w8(32'h3b308987),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092881),
	.w1(32'h3bf5cfca),
	.w2(32'h3b20d861),
	.w3(32'hbbf003d0),
	.w4(32'hba90c865),
	.w5(32'hb925d25f),
	.w6(32'h3b56e1c2),
	.w7(32'hbb5ca9c0),
	.w8(32'h3ab2a53b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b3664),
	.w1(32'h37f7eb93),
	.w2(32'hbac21fb8),
	.w3(32'hba58dc88),
	.w4(32'h3b4a7d26),
	.w5(32'h3b605421),
	.w6(32'hbb20721c),
	.w7(32'h3a9419d6),
	.w8(32'h3c04e69c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1110ba),
	.w1(32'hba60a94f),
	.w2(32'h3bf3ebc6),
	.w3(32'h3c18ddca),
	.w4(32'hbb916613),
	.w5(32'h3b591dd9),
	.w6(32'h3c5692d1),
	.w7(32'hbb938b63),
	.w8(32'hbb79b099),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5f93f),
	.w1(32'h3b609fd0),
	.w2(32'h3bd55b08),
	.w3(32'h3b8028f7),
	.w4(32'hbab35a7f),
	.w5(32'hbb8b3d11),
	.w6(32'hbb9fa3e5),
	.w7(32'hbba7d0ff),
	.w8(32'hbbe9c790),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75409e),
	.w1(32'hbb6a3071),
	.w2(32'hbaf5d125),
	.w3(32'h3b202a30),
	.w4(32'h39aff71e),
	.w5(32'h3b1f7ebc),
	.w6(32'h3aa164f3),
	.w7(32'h3a98840b),
	.w8(32'h3a1490a1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5307a),
	.w1(32'hbaa24fcc),
	.w2(32'h3b9be718),
	.w3(32'h3bf8d416),
	.w4(32'hbc705bc5),
	.w5(32'hbbc8527b),
	.w6(32'h3c49ccfc),
	.w7(32'hbb79a955),
	.w8(32'hbc550b8b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57838f),
	.w1(32'hbb6ca25a),
	.w2(32'hbbcaf9e8),
	.w3(32'hbb55487d),
	.w4(32'hbb7fcd58),
	.w5(32'hbbccb4e0),
	.w6(32'hbc13093f),
	.w7(32'h3a2b0a84),
	.w8(32'hbb70154a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6273bb),
	.w1(32'hbbc4fb1a),
	.w2(32'hbb65141f),
	.w3(32'hbb7af8f0),
	.w4(32'hbb6bc52b),
	.w5(32'h3b2ddbc3),
	.w6(32'hbc38e204),
	.w7(32'hbbc96346),
	.w8(32'h3ae1adac),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeadbc),
	.w1(32'h3a80c9ed),
	.w2(32'h3b686eb7),
	.w3(32'h39fcd65c),
	.w4(32'hba3a2be7),
	.w5(32'h3a788df9),
	.w6(32'h3b1dd102),
	.w7(32'hbb02f56a),
	.w8(32'hbb196a3a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b204827),
	.w1(32'hbb7f02e7),
	.w2(32'hbac085cc),
	.w3(32'h3b4df87a),
	.w4(32'hba7cd91d),
	.w5(32'hb9a39dd6),
	.w6(32'h39d693e3),
	.w7(32'hbb52fdae),
	.w8(32'h38df7a89),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c389835),
	.w1(32'h3bf4eff6),
	.w2(32'h3c0157eb),
	.w3(32'hba7cd2e3),
	.w4(32'h3ca9a5cf),
	.w5(32'h3c52d434),
	.w6(32'hbc65c720),
	.w7(32'h3b25f978),
	.w8(32'h3c192078),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2675da),
	.w1(32'h3c069fd5),
	.w2(32'hba4475be),
	.w3(32'hbb502b9f),
	.w4(32'h3c507299),
	.w5(32'h3bc657f6),
	.w6(32'hbc17b17f),
	.w7(32'h3b5df440),
	.w8(32'h3c0af3a3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd734e),
	.w1(32'h3b4ac911),
	.w2(32'h3a019c72),
	.w3(32'h3b5c903f),
	.w4(32'h3b42dc3b),
	.w5(32'h3ae51de6),
	.w6(32'h3b025f93),
	.w7(32'h3997ce02),
	.w8(32'hbafabce5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc58b7),
	.w1(32'h3b2daa53),
	.w2(32'h3c846fc6),
	.w3(32'h3c51658d),
	.w4(32'h3c071dd1),
	.w5(32'hbacdacc5),
	.w6(32'h3b118ce2),
	.w7(32'h3c0d54e9),
	.w8(32'hbc382141),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b902521),
	.w1(32'h3a239392),
	.w2(32'hbb13a049),
	.w3(32'hba11d126),
	.w4(32'h3ac444fc),
	.w5(32'hbb9e1239),
	.w6(32'hbb2ff2f8),
	.w7(32'hbaf8a421),
	.w8(32'hbb8feff6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5536f7),
	.w1(32'hb9f3b66e),
	.w2(32'hbb7ad333),
	.w3(32'hb896ad6b),
	.w4(32'hba821b32),
	.w5(32'hbbbb1040),
	.w6(32'hbb8bb3f0),
	.w7(32'hbb45c0f4),
	.w8(32'hbb905870),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc551fff),
	.w1(32'h3c7238aa),
	.w2(32'h3d10e7d9),
	.w3(32'hbd134734),
	.w4(32'h3cd2b2cc),
	.w5(32'h3d1a2b9e),
	.w6(32'hbd16ad36),
	.w7(32'hbc00b81d),
	.w8(32'h3cef4d2c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8b838),
	.w1(32'h3abb8cd9),
	.w2(32'h3a5f0314),
	.w3(32'hbb9e1946),
	.w4(32'h3c2fd7ec),
	.w5(32'hba05ad3f),
	.w6(32'hbbe53324),
	.w7(32'h3bbff5d3),
	.w8(32'h3beba676),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5d4b3),
	.w1(32'h3c0225a5),
	.w2(32'h3b9aaa8e),
	.w3(32'hbc28418f),
	.w4(32'h3ca820f5),
	.w5(32'h3beba605),
	.w6(32'hbc851949),
	.w7(32'h3ae8e55c),
	.w8(32'h3c2adefa),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a2761),
	.w1(32'hbb13dbef),
	.w2(32'h3af18c7e),
	.w3(32'hbb54f52b),
	.w4(32'hbc014a8b),
	.w5(32'h3ba32416),
	.w6(32'h3c1d08f3),
	.w7(32'hbc035c39),
	.w8(32'hbb8424a8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd57474),
	.w1(32'h3b802603),
	.w2(32'h3beac250),
	.w3(32'h3c3b5d01),
	.w4(32'hbbf313a1),
	.w5(32'h3abaf37c),
	.w6(32'h3c64fcfc),
	.w7(32'hbbce2617),
	.w8(32'hbbbe6a41),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f20021),
	.w1(32'h3a971bfe),
	.w2(32'h389e92b2),
	.w3(32'h3b538a0e),
	.w4(32'h3af998d2),
	.w5(32'hbbcec81b),
	.w6(32'h3af573a9),
	.w7(32'h3b201d28),
	.w8(32'hbb0579dd),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9911fb),
	.w1(32'hbaa44373),
	.w2(32'hbb6ecb6f),
	.w3(32'h3b52cf31),
	.w4(32'h3ac507a7),
	.w5(32'h3babbb77),
	.w6(32'hbb0a10cf),
	.w7(32'hbb72c073),
	.w8(32'h3b61aee0),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d75b9),
	.w1(32'h3c44da09),
	.w2(32'h3c3b499e),
	.w3(32'h3bfe4e2f),
	.w4(32'h3bd6a2f3),
	.w5(32'h3a4ce4ca),
	.w6(32'h3c7fedf5),
	.w7(32'h3c18e677),
	.w8(32'hbaae2c5e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b420a68),
	.w1(32'hbb47dca7),
	.w2(32'h3a452dfc),
	.w3(32'h3ae7211e),
	.w4(32'hbb1b2120),
	.w5(32'hbb1965fc),
	.w6(32'hbb2d4dcd),
	.w7(32'hbbe2c77d),
	.w8(32'hbb3a706c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e7f67),
	.w1(32'h3bc4cd7e),
	.w2(32'hb9318850),
	.w3(32'h3abe88e0),
	.w4(32'h3bd2d97b),
	.w5(32'h3ab81788),
	.w6(32'hbb8cd361),
	.w7(32'h3a96ae3c),
	.w8(32'hbae64fe8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7129ff),
	.w1(32'h3c00f5d9),
	.w2(32'hbbfa21fa),
	.w3(32'hba859099),
	.w4(32'h3c1b0ac7),
	.w5(32'h3baa2772),
	.w6(32'h39d87316),
	.w7(32'hbba5ec58),
	.w8(32'h3789ca3f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c187a48),
	.w1(32'h3c2c879d),
	.w2(32'h3bb70919),
	.w3(32'h3be366e3),
	.w4(32'h3b541f0f),
	.w5(32'hba45162b),
	.w6(32'hbc0e71fe),
	.w7(32'hbb176e28),
	.w8(32'hb9bb2589),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b330b),
	.w1(32'h3b16106c),
	.w2(32'h3a00801e),
	.w3(32'hba3712ad),
	.w4(32'h3b1619eb),
	.w5(32'hb9bfc902),
	.w6(32'h3b878130),
	.w7(32'h3bac7447),
	.w8(32'hba222b2f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf86ebb),
	.w1(32'h3c3f4c14),
	.w2(32'h3b90b84a),
	.w3(32'hbc6c9b9b),
	.w4(32'h3cec00e5),
	.w5(32'h3c335e2b),
	.w6(32'hbcdb9767),
	.w7(32'h3b8805b7),
	.w8(32'h3c7acddf),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbdf94),
	.w1(32'hbadd4214),
	.w2(32'hb942a28c),
	.w3(32'h3add5379),
	.w4(32'h3b92d87c),
	.w5(32'h3a0cd293),
	.w6(32'hba8cdcfb),
	.w7(32'h3be418fb),
	.w8(32'hba6f2463),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139739),
	.w1(32'hbae6d377),
	.w2(32'hbc110f66),
	.w3(32'hbb696e23),
	.w4(32'hbb9bf1eb),
	.w5(32'h3b75d6cc),
	.w6(32'hb9738e98),
	.w7(32'h3aecf805),
	.w8(32'h3afa4b64),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7f210),
	.w1(32'h3b06c3fc),
	.w2(32'h3ba302be),
	.w3(32'h3b820896),
	.w4(32'h3c1abfbf),
	.w5(32'h3aafe34c),
	.w6(32'hbb986169),
	.w7(32'h3b2406fb),
	.w8(32'hbb080b7d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8806b1),
	.w1(32'hbbc2c1c6),
	.w2(32'hbb9a4a22),
	.w3(32'hba8caef1),
	.w4(32'hba2a8bf1),
	.w5(32'hbb0a2ebc),
	.w6(32'hbb8a4f21),
	.w7(32'hba900aec),
	.w8(32'hbb821703),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb534c5e),
	.w1(32'hb90f257d),
	.w2(32'h3a875489),
	.w3(32'hba0b0522),
	.w4(32'h3a8b2df9),
	.w5(32'hbb96a77c),
	.w6(32'hbae39930),
	.w7(32'h3999510d),
	.w8(32'hbba24f46),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920606),
	.w1(32'hbbaaf638),
	.w2(32'hbad76db9),
	.w3(32'hbbbb5bfe),
	.w4(32'hbb9c43b1),
	.w5(32'hbb017ded),
	.w6(32'hbbbe4251),
	.w7(32'hbb18fce2),
	.w8(32'hbafaae4a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd01e3),
	.w1(32'hba004640),
	.w2(32'hba5af679),
	.w3(32'h3a76bb20),
	.w4(32'h38d324e4),
	.w5(32'hba05e730),
	.w6(32'hba61f1fa),
	.w7(32'hbac4cddb),
	.w8(32'h3a8a9f03),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ff669),
	.w1(32'h3b188023),
	.w2(32'h3b9bb0de),
	.w3(32'hbafecc1f),
	.w4(32'h3a773f7c),
	.w5(32'h39b012eb),
	.w6(32'h3b8c1e29),
	.w7(32'h399b6ca9),
	.w8(32'h3a0a676b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba49588),
	.w1(32'h3c17a0e5),
	.w2(32'h3bacbdb1),
	.w3(32'h3c8b80c7),
	.w4(32'h3b7082c0),
	.w5(32'h3ba61d21),
	.w6(32'h3bd3b4ea),
	.w7(32'h3c2c82e6),
	.w8(32'hba354546),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf14683),
	.w1(32'h3b51f822),
	.w2(32'hbb323f27),
	.w3(32'h3b729a8e),
	.w4(32'h3c184eb5),
	.w5(32'hbb9648f6),
	.w6(32'hbb5d3152),
	.w7(32'h3bccc49a),
	.w8(32'h3b6fa877),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab75be),
	.w1(32'h3b9877ef),
	.w2(32'h3bd1315f),
	.w3(32'h3b5ae155),
	.w4(32'h3ad13270),
	.w5(32'h3a45e228),
	.w6(32'hbba86e2f),
	.w7(32'h3befe488),
	.w8(32'h3c37652f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac2e8b),
	.w1(32'h3b1ff9f3),
	.w2(32'h3a0de1be),
	.w3(32'h3aeef954),
	.w4(32'h3b2d2b19),
	.w5(32'hbb84d229),
	.w6(32'h3b029c89),
	.w7(32'h3a1200c4),
	.w8(32'hba6e6469),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabed24),
	.w1(32'h39f95229),
	.w2(32'hb93cd069),
	.w3(32'hb9d1dc8d),
	.w4(32'h3b033915),
	.w5(32'hb9df31cd),
	.w6(32'h3a8427c5),
	.w7(32'h3a925cf2),
	.w8(32'hbae17c7c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397fd768),
	.w1(32'h3a9b73c9),
	.w2(32'h3a6f0a63),
	.w3(32'hb9e11e48),
	.w4(32'h3b009228),
	.w5(32'h3b9d4e2e),
	.w6(32'hbb29632d),
	.w7(32'hba104175),
	.w8(32'h3bce9068),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac25514),
	.w1(32'hba9f2351),
	.w2(32'h3a970631),
	.w3(32'h3b8acab6),
	.w4(32'hb930dc66),
	.w5(32'hbb6f3472),
	.w6(32'h3c81eb4b),
	.w7(32'h3c5a626d),
	.w8(32'h397e1210),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09e984),
	.w1(32'hbbfca8dd),
	.w2(32'hbc32ee45),
	.w3(32'h3c0b5513),
	.w4(32'hbbfa2e71),
	.w5(32'hbc051f48),
	.w6(32'h3bf04bb5),
	.w7(32'h3b803cfd),
	.w8(32'hbbb67d27),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ab542),
	.w1(32'hbb192bd5),
	.w2(32'hbbb55b35),
	.w3(32'hbb24a56e),
	.w4(32'hbb829fc8),
	.w5(32'hbb3ea997),
	.w6(32'hbc152fd7),
	.w7(32'hbb89a19f),
	.w8(32'hbb09f03e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b19a31),
	.w1(32'hb9c23446),
	.w2(32'h37b1cf85),
	.w3(32'h3b6de045),
	.w4(32'h3a51d848),
	.w5(32'hba1b6ac2),
	.w6(32'h3a805a90),
	.w7(32'hb856061d),
	.w8(32'h3b1436d1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939e9f),
	.w1(32'hbaa743ab),
	.w2(32'hbb99be4a),
	.w3(32'hbb61188f),
	.w4(32'hbbe226b5),
	.w5(32'h3a959f44),
	.w6(32'hba619cb4),
	.w7(32'hbbb4aeb0),
	.w8(32'h3bb7712e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf6002),
	.w1(32'h3b6fc433),
	.w2(32'h3bca7a1b),
	.w3(32'h3b74f9f7),
	.w4(32'h3bd2c6fb),
	.w5(32'hbaeceda9),
	.w6(32'h3b90fed6),
	.w7(32'h3b440a8f),
	.w8(32'hbb34153d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78d643),
	.w1(32'hba99e050),
	.w2(32'hbb3e9350),
	.w3(32'hb9976950),
	.w4(32'h3b2460d6),
	.w5(32'hb6ab47f0),
	.w6(32'hbbb456d4),
	.w7(32'hba8a98ce),
	.w8(32'h3bbc95bf),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf8336),
	.w1(32'h3b89cbbf),
	.w2(32'h3b1fa77d),
	.w3(32'h3b10da65),
	.w4(32'h3b7256c0),
	.w5(32'hbb76c293),
	.w6(32'h3b5b45e7),
	.w7(32'hb8b26a76),
	.w8(32'hbac2be37),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a4aad),
	.w1(32'hbc6c01d2),
	.w2(32'hbba99c5a),
	.w3(32'h3ca12abb),
	.w4(32'hbcc509af),
	.w5(32'hbc248630),
	.w6(32'h3ca429a0),
	.w7(32'h3bbd6ecd),
	.w8(32'hbc58fd2a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a79fe),
	.w1(32'h3aed43ad),
	.w2(32'hbb068f2a),
	.w3(32'hb7ade151),
	.w4(32'hbb239dab),
	.w5(32'hba996ed2),
	.w6(32'hbb9f75c4),
	.w7(32'hbbb0b5c9),
	.w8(32'hbad9b38a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973bfdf),
	.w1(32'h3b5444e5),
	.w2(32'h3ab2a531),
	.w3(32'hbc11ce74),
	.w4(32'h3aae4f10),
	.w5(32'h3be51a14),
	.w6(32'hbba28f56),
	.w7(32'h3a2e2205),
	.w8(32'h3c336241),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule