module layer_10_featuremap_491(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb8eb8),
	.w1(32'hbb1798df),
	.w2(32'hb9c34b74),
	.w3(32'hbb33b40e),
	.w4(32'hbb9e8c12),
	.w5(32'hbb428cf8),
	.w6(32'hba22144c),
	.w7(32'hbbb69fe6),
	.w8(32'hba31ef5f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb701ca7),
	.w1(32'h3b83e9f9),
	.w2(32'hbb5a600b),
	.w3(32'h38e65250),
	.w4(32'h3a12a596),
	.w5(32'hbb056a70),
	.w6(32'hbb1437bc),
	.w7(32'hbb9846d7),
	.w8(32'hbb847edd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab30550),
	.w1(32'h3af22869),
	.w2(32'hbb3fed99),
	.w3(32'hbb9f1325),
	.w4(32'h3bf2cc65),
	.w5(32'hbc401d91),
	.w6(32'hbb316c9d),
	.w7(32'h3bacbf3a),
	.w8(32'h3bcd96f5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d30f3),
	.w1(32'h3ab4e7d8),
	.w2(32'hbb485641),
	.w3(32'h3a94ac40),
	.w4(32'hba8ee480),
	.w5(32'h3aa2e312),
	.w6(32'h3abfee2b),
	.w7(32'h3984b37b),
	.w8(32'h3a8eb9b9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8284f),
	.w1(32'hbb744ad5),
	.w2(32'hbac93528),
	.w3(32'h3b0840c8),
	.w4(32'hbb425c5b),
	.w5(32'hbb9ed6f5),
	.w6(32'h3b95925e),
	.w7(32'hbbd8b1b2),
	.w8(32'hbb2765fd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2443a),
	.w1(32'hbb23acc5),
	.w2(32'hbbd0455c),
	.w3(32'h3b3e9f2e),
	.w4(32'hbbdacdc3),
	.w5(32'hbb2882a6),
	.w6(32'h3956c1a0),
	.w7(32'hbbb0a99f),
	.w8(32'hbb8cb6ec),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03b664),
	.w1(32'h3b642826),
	.w2(32'h3c00a7c5),
	.w3(32'hbb28ed36),
	.w4(32'h3b903c20),
	.w5(32'h3a84cc0c),
	.w6(32'hbb449b73),
	.w7(32'h3b549020),
	.w8(32'h37e3eeba),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c4827),
	.w1(32'hbbef46e4),
	.w2(32'hbc17c006),
	.w3(32'h3ad4311d),
	.w4(32'hbaa2152e),
	.w5(32'hbbafda98),
	.w6(32'hbbbfa8da),
	.w7(32'hbb4d9f47),
	.w8(32'h3bb41111),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8ee1c),
	.w1(32'h3ac6b9c3),
	.w2(32'hbb919e45),
	.w3(32'hba413201),
	.w4(32'hba5d004d),
	.w5(32'hbc0345b2),
	.w6(32'h3a73f8c4),
	.w7(32'h3a592cc3),
	.w8(32'hbaadf15a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae471a0),
	.w1(32'h3a01ca1f),
	.w2(32'h3b1f4c7f),
	.w3(32'h3c32d99b),
	.w4(32'h3aa519bc),
	.w5(32'hba29d8fb),
	.w6(32'h3b9a4900),
	.w7(32'hbb36fcab),
	.w8(32'hbbe39073),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aa675),
	.w1(32'h3b4d81f4),
	.w2(32'h3b05bc8a),
	.w3(32'h399cee9b),
	.w4(32'h3b28b519),
	.w5(32'hbacc146a),
	.w6(32'hbb19fef2),
	.w7(32'hbaa3dcfa),
	.w8(32'hb9127f56),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86fab4),
	.w1(32'hbb4ed3ff),
	.w2(32'h3a813878),
	.w3(32'h3c15e540),
	.w4(32'h3a0294cb),
	.w5(32'h3ba726ea),
	.w6(32'h3b1f4d53),
	.w7(32'h3b74fbbf),
	.w8(32'h3a939cf6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cabce),
	.w1(32'h3c312100),
	.w2(32'h3943af84),
	.w3(32'h3ae14d6b),
	.w4(32'h3b335b85),
	.w5(32'h3abe5c87),
	.w6(32'h39c37eaf),
	.w7(32'h3a599421),
	.w8(32'hbad6bcc2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67bf42),
	.w1(32'hba9b213f),
	.w2(32'hbbd04975),
	.w3(32'hbb03e089),
	.w4(32'hba9af3cd),
	.w5(32'h3b1b846d),
	.w6(32'h3b31f118),
	.w7(32'h3b4504ad),
	.w8(32'h3b06a2b4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36ae04),
	.w1(32'h383b39f4),
	.w2(32'hbb846692),
	.w3(32'h3ad24b7d),
	.w4(32'hbac80d38),
	.w5(32'hbc07f326),
	.w6(32'h3c0410a4),
	.w7(32'h3a03828a),
	.w8(32'hbacafdc4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadf59a),
	.w1(32'h3a882d77),
	.w2(32'hbc04091a),
	.w3(32'hbaed8c0e),
	.w4(32'hbb4af528),
	.w5(32'hbbc49659),
	.w6(32'hbbcb3bbe),
	.w7(32'hba26edf5),
	.w8(32'hbb9d7708),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93c541),
	.w1(32'hbbcfe2a5),
	.w2(32'hbbb48500),
	.w3(32'h3b9ba489),
	.w4(32'hbb9d3964),
	.w5(32'hbb49a361),
	.w6(32'h3acb2c17),
	.w7(32'hbb67b6c8),
	.w8(32'hbb0fb7dd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5eb4e9),
	.w1(32'hbc562a07),
	.w2(32'hbc44e1c9),
	.w3(32'hbc6a31c1),
	.w4(32'hbc331248),
	.w5(32'hbb94f781),
	.w6(32'hbc143afd),
	.w7(32'hbb971f90),
	.w8(32'hbabfab20),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba83cdd),
	.w1(32'hba578f12),
	.w2(32'hb98b5ada),
	.w3(32'hbb198d12),
	.w4(32'h3abcc9af),
	.w5(32'hbb5fa410),
	.w6(32'hbb757ea3),
	.w7(32'hba84bc67),
	.w8(32'hbada3078),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3e7d6),
	.w1(32'hbb90d778),
	.w2(32'hbbbdd34e),
	.w3(32'h3c1f7d41),
	.w4(32'hbbc36478),
	.w5(32'hbbcd9186),
	.w6(32'h3bea0926),
	.w7(32'hbbc2a707),
	.w8(32'hbbaac327),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0758c),
	.w1(32'h3996ccfa),
	.w2(32'hba44a9a7),
	.w3(32'h394e4c98),
	.w4(32'hbb0ae4ad),
	.w5(32'h3ac329cd),
	.w6(32'hbb56f411),
	.w7(32'hbae94997),
	.w8(32'hba527015),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b241a90),
	.w1(32'h3bb417a7),
	.w2(32'hb96252b3),
	.w3(32'h3b3a9a8a),
	.w4(32'h3bd4d397),
	.w5(32'h3af1d2e1),
	.w6(32'hb93e719f),
	.w7(32'h3bff23ee),
	.w8(32'h3b19fa92),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dc2d3),
	.w1(32'hbc9ad1cc),
	.w2(32'hbc1c4289),
	.w3(32'hbca0a099),
	.w4(32'hbbddade2),
	.w5(32'hbbff5a89),
	.w6(32'hbc9b2220),
	.w7(32'hbb95ca7f),
	.w8(32'hbc2029f6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e6201),
	.w1(32'h3b4b01dd),
	.w2(32'hbb1ac278),
	.w3(32'hbadb1049),
	.w4(32'h3b0f575f),
	.w5(32'hbac778af),
	.w6(32'hbafcb6d3),
	.w7(32'hbb28178a),
	.w8(32'hbc16dabf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163225),
	.w1(32'h3b9ed7a2),
	.w2(32'hbb4d15cf),
	.w3(32'h3b4dac4a),
	.w4(32'hba85d4e6),
	.w5(32'hbbba8f9c),
	.w6(32'hbbaa1163),
	.w7(32'hbc0aa7d9),
	.w8(32'hbc413b98),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ac89),
	.w1(32'hbb5e2241),
	.w2(32'h3969c294),
	.w3(32'hbb7a21f3),
	.w4(32'hbb2870e1),
	.w5(32'h3a97b5a6),
	.w6(32'hbbf2c4a3),
	.w7(32'hbaaf7f49),
	.w8(32'hbbe21827),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14984d),
	.w1(32'hbab66db9),
	.w2(32'h3adc499b),
	.w3(32'hbb4b6ea8),
	.w4(32'h3a9abdac),
	.w5(32'h3bcf5506),
	.w6(32'hba0664f6),
	.w7(32'h3b1b32c9),
	.w8(32'h3b72eb20),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25a7ae),
	.w1(32'h3bbdcc55),
	.w2(32'h3b54e836),
	.w3(32'h3b6a6cee),
	.w4(32'h3ba29d68),
	.w5(32'hbbdd6fbd),
	.w6(32'h3b86199e),
	.w7(32'h3b100844),
	.w8(32'hbb94a042),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfcf4e),
	.w1(32'hba8399e0),
	.w2(32'h3b4fc428),
	.w3(32'hb9c14dd8),
	.w4(32'hbad68877),
	.w5(32'h3b3e89ff),
	.w6(32'hbb0d4eab),
	.w7(32'hbb1455a0),
	.w8(32'hbba5defc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04c24e),
	.w1(32'h3c077f89),
	.w2(32'h3b1ac586),
	.w3(32'h3b0feb6b),
	.w4(32'hbb190d05),
	.w5(32'hbbcbd0ce),
	.w6(32'h3ad7d88f),
	.w7(32'hbb6de7d2),
	.w8(32'hbc12b7ae),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66c324),
	.w1(32'hbb9c5a1a),
	.w2(32'h3ac568f4),
	.w3(32'h3acb9806),
	.w4(32'hbb7a95c2),
	.w5(32'h3bf8a908),
	.w6(32'h3af58053),
	.w7(32'hba6277ba),
	.w8(32'hbb8b1dbc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4cfe3),
	.w1(32'h3c35b0a2),
	.w2(32'h3be01dc1),
	.w3(32'h3b5ba1eb),
	.w4(32'h3c5a73f1),
	.w5(32'h3b83b55f),
	.w6(32'hbb605780),
	.w7(32'h3c07609b),
	.w8(32'h3bd36862),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb729e),
	.w1(32'h3bb4312c),
	.w2(32'h3ac80a24),
	.w3(32'hbb82fbc1),
	.w4(32'h3c0f164d),
	.w5(32'h3ba0e4a3),
	.w6(32'hbb5f3d66),
	.w7(32'h3a83e780),
	.w8(32'hbb15d35c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41d0b7),
	.w1(32'h3b3f355b),
	.w2(32'h3bfd8b71),
	.w3(32'h3c0414af),
	.w4(32'h3b7df696),
	.w5(32'h3a13121b),
	.w6(32'hba6cf3c1),
	.w7(32'hbb220b8e),
	.w8(32'hbb92a69f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58c055),
	.w1(32'hbbbbf38f),
	.w2(32'hbb4ce96c),
	.w3(32'h3a5b3968),
	.w4(32'hb9863177),
	.w5(32'h3c17891d),
	.w6(32'h3a8c91a4),
	.w7(32'hb994a786),
	.w8(32'hbb702220),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaace749),
	.w1(32'h39b159a0),
	.w2(32'hbb3db872),
	.w3(32'hbb99d9db),
	.w4(32'h3b088004),
	.w5(32'h3aeda481),
	.w6(32'hbacf4821),
	.w7(32'h3b13aa73),
	.w8(32'hba7b7de6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0fac1),
	.w1(32'hbb80dca6),
	.w2(32'hbad351ec),
	.w3(32'h3bfc23e0),
	.w4(32'hbc1bacbf),
	.w5(32'hba54e459),
	.w6(32'h39918cc9),
	.w7(32'hbc3222cb),
	.w8(32'hbbe6df0a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b1715),
	.w1(32'h3c5f6d0f),
	.w2(32'hbba6de23),
	.w3(32'h3bb370fe),
	.w4(32'h3c4fc2cc),
	.w5(32'hbbf05cd3),
	.w6(32'hbb13d47a),
	.w7(32'h3ac6f8d0),
	.w8(32'hbc20ba28),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70f524),
	.w1(32'h3c2f3381),
	.w2(32'h3a8d5e55),
	.w3(32'h3bef46f6),
	.w4(32'h3c2e5468),
	.w5(32'hbbb2a899),
	.w6(32'h3be8ab9d),
	.w7(32'h3bb4cd81),
	.w8(32'h3a56308f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba460a4),
	.w1(32'hbb3a4447),
	.w2(32'hbb9b279c),
	.w3(32'h3a3321e8),
	.w4(32'h3968af8d),
	.w5(32'hbba652b5),
	.w6(32'h398156fc),
	.w7(32'hba576044),
	.w8(32'hbb8284d2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd27718),
	.w1(32'hbbf2e320),
	.w2(32'h3b2ce4c5),
	.w3(32'hbb89b565),
	.w4(32'hbc106155),
	.w5(32'h3cc7fedd),
	.w6(32'hbb10bcf8),
	.w7(32'hbaac3346),
	.w8(32'h3b7e1470),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e61902),
	.w1(32'hbb1cc5a9),
	.w2(32'h3aad6a40),
	.w3(32'hbbe1de6f),
	.w4(32'hbb13cbc1),
	.w5(32'h3b0a50b6),
	.w6(32'h3a43404a),
	.w7(32'hbb4f107a),
	.w8(32'hb9a58380),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0110c6),
	.w1(32'h3b0c85fe),
	.w2(32'hba9a447a),
	.w3(32'hbb988aa9),
	.w4(32'h3b16b3eb),
	.w5(32'h3b5e21e5),
	.w6(32'hbb61ab86),
	.w7(32'h3abfbf37),
	.w8(32'hba320e63),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb913585),
	.w1(32'hba4f87f3),
	.w2(32'hbb90bfde),
	.w3(32'hbbdca15c),
	.w4(32'hbbb4cb56),
	.w5(32'hbbb90acd),
	.w6(32'hbb574a5a),
	.w7(32'hbbc7b810),
	.w8(32'h3ae8f026),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb1c3),
	.w1(32'h3c2610b6),
	.w2(32'h3b295726),
	.w3(32'h3a822154),
	.w4(32'h3bb4c1a6),
	.w5(32'hbbd7173c),
	.w6(32'h3b5bc014),
	.w7(32'h3a2d9d83),
	.w8(32'hbc2149b0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36da5e),
	.w1(32'hbac3c80e),
	.w2(32'hbabdd10d),
	.w3(32'h3b179f39),
	.w4(32'hbba20e52),
	.w5(32'h389a7610),
	.w6(32'hba069474),
	.w7(32'hbb64de6b),
	.w8(32'hbb528fb3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd0cac),
	.w1(32'hbb34f572),
	.w2(32'h3aae33a3),
	.w3(32'h3a3d3ee6),
	.w4(32'hb8e18cd5),
	.w5(32'h3b7fc53a),
	.w6(32'hbc052137),
	.w7(32'hba4ac12f),
	.w8(32'hbafe7536),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e115c),
	.w1(32'hbc8abf36),
	.w2(32'hbc238edb),
	.w3(32'hbc9180fd),
	.w4(32'hbc221109),
	.w5(32'h3a84f9fd),
	.w6(32'hbca1bac2),
	.w7(32'hbbdffb2b),
	.w8(32'hba2e7c54),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bfff0),
	.w1(32'h3af2b95c),
	.w2(32'hbad09c0f),
	.w3(32'hb9c4512f),
	.w4(32'hba571b2f),
	.w5(32'hbb9dd2f0),
	.w6(32'hb83b7491),
	.w7(32'hbaa8ccac),
	.w8(32'hbb238dd7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad24b3),
	.w1(32'h3b739a1a),
	.w2(32'h3c1adc70),
	.w3(32'h3c23a1d0),
	.w4(32'h3c676eb9),
	.w5(32'h3c54415e),
	.w6(32'h3bb26a36),
	.w7(32'h3bf2cd4f),
	.w8(32'h3b36c7f2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49fb92),
	.w1(32'hbb7bfe24),
	.w2(32'hbaae229a),
	.w3(32'hbb9723c5),
	.w4(32'hbae84e5f),
	.w5(32'h3afd8a4a),
	.w6(32'hbc119360),
	.w7(32'hbbb7bb97),
	.w8(32'hba2cac9e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbd3b9),
	.w1(32'hbbe8d15b),
	.w2(32'hbbad86ba),
	.w3(32'hbb8246cf),
	.w4(32'hb9d570b1),
	.w5(32'hb9f7be19),
	.w6(32'hbb8d3c89),
	.w7(32'hba186551),
	.w8(32'hbb4c1151),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53e8c7),
	.w1(32'hba665d05),
	.w2(32'hba14ac35),
	.w3(32'hbb5d28f0),
	.w4(32'h3ab50dac),
	.w5(32'h3b6ab348),
	.w6(32'hbb62be63),
	.w7(32'h3a2f18bb),
	.w8(32'hbb5ac3f6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4568a0),
	.w1(32'hbc5eaed2),
	.w2(32'hbc2fddf0),
	.w3(32'hbc44a05e),
	.w4(32'hbbede0b6),
	.w5(32'h3b2afe7b),
	.w6(32'hbc446e0f),
	.w7(32'hbb64746c),
	.w8(32'hbb914e5e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c889),
	.w1(32'hbb83de29),
	.w2(32'hbbb44b53),
	.w3(32'hb805a056),
	.w4(32'hbafe61fd),
	.w5(32'hbb8f638c),
	.w6(32'h3b219fe6),
	.w7(32'hba988a02),
	.w8(32'hbb8b1301),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc4b78),
	.w1(32'hbb8cd087),
	.w2(32'hbbf8b5cc),
	.w3(32'hbbaed113),
	.w4(32'hbbbb11a3),
	.w5(32'hba4bbff5),
	.w6(32'hbb014792),
	.w7(32'hbb30c030),
	.w8(32'hbb05adb3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ec4be),
	.w1(32'hba6a330a),
	.w2(32'h3b6a7623),
	.w3(32'h3b895b97),
	.w4(32'hbb409632),
	.w5(32'h3b2440fd),
	.w6(32'h3bb3b14d),
	.w7(32'hbb8ff899),
	.w8(32'hb93d3ee8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d54f9),
	.w1(32'h39c97b9a),
	.w2(32'hbb9cd1c5),
	.w3(32'hbb377ae7),
	.w4(32'h3a428486),
	.w5(32'hbb93243f),
	.w6(32'h3a77ebca),
	.w7(32'h392380b3),
	.w8(32'hbb0bf3a3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818989),
	.w1(32'hbb3f6cda),
	.w2(32'hbbbd24d7),
	.w3(32'h3ad9b002),
	.w4(32'hbbccaf6a),
	.w5(32'hbbb18178),
	.w6(32'hba22e6e4),
	.w7(32'hbb67a23b),
	.w8(32'hbb82b260),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9704e),
	.w1(32'hbbd54c2c),
	.w2(32'hbbd3987b),
	.w3(32'hbc1d5e32),
	.w4(32'hbc31376e),
	.w5(32'hbbe61222),
	.w6(32'hbbe506fe),
	.w7(32'hbb028189),
	.w8(32'hbb884472),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ab7b8),
	.w1(32'hbc257eee),
	.w2(32'hbbb72ac0),
	.w3(32'hbbeb7fa6),
	.w4(32'hbba6a475),
	.w5(32'h3b29927f),
	.w6(32'hbb99596d),
	.w7(32'hba9fa4f4),
	.w8(32'hbb2b169b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ec13d),
	.w1(32'hbb984ba5),
	.w2(32'h3b0045c2),
	.w3(32'hbc1f934f),
	.w4(32'h3bac598a),
	.w5(32'hbb6d859c),
	.w6(32'hbb98c02f),
	.w7(32'h3b5fa3b6),
	.w8(32'h3b0ae73f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860cf4),
	.w1(32'hbb452b85),
	.w2(32'hbb63c989),
	.w3(32'h3a6386ae),
	.w4(32'hbbde2322),
	.w5(32'hb923298b),
	.w6(32'hba0a5291),
	.w7(32'hba0e0147),
	.w8(32'hbb534b31),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a8b39),
	.w1(32'hbb686d4c),
	.w2(32'h3bb8dc69),
	.w3(32'hbb849be8),
	.w4(32'hbb4a98a1),
	.w5(32'h3bb71579),
	.w6(32'hbab775a9),
	.w7(32'hbad3f9ca),
	.w8(32'h3b51abfd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacbeaf),
	.w1(32'h3bb54d5e),
	.w2(32'h3af6735f),
	.w3(32'h3ba4ce31),
	.w4(32'h3ba3b008),
	.w5(32'hba3723e4),
	.w6(32'h393dd28a),
	.w7(32'h3bd9baa6),
	.w8(32'h3b8efacd),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaa24b),
	.w1(32'h3be7699c),
	.w2(32'h3b47a2f5),
	.w3(32'h3bd14fdc),
	.w4(32'h3bd39d56),
	.w5(32'h3bb28883),
	.w6(32'h3bc2f670),
	.w7(32'h3b05261c),
	.w8(32'h3ba896ed),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d6b227),
	.w1(32'h3af21f03),
	.w2(32'h3bc12887),
	.w3(32'h3b62ce47),
	.w4(32'hbace8ab6),
	.w5(32'h3b9f677f),
	.w6(32'hbb05be29),
	.w7(32'hbb3ce032),
	.w8(32'h3a451965),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3572c6),
	.w1(32'hbbea0b6a),
	.w2(32'hb99130c4),
	.w3(32'hbb33abb1),
	.w4(32'hbbbeedd0),
	.w5(32'hbb2ee0c0),
	.w6(32'hbbf7a198),
	.w7(32'hbc3aec40),
	.w8(32'hbc193392),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32241d),
	.w1(32'hbba84ed4),
	.w2(32'hbbcc6ddf),
	.w3(32'hbc16805e),
	.w4(32'h3bf9aae6),
	.w5(32'hbbbb13ab),
	.w6(32'hbbeab288),
	.w7(32'h3b262397),
	.w8(32'hbbebc64b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cd394),
	.w1(32'h39bb8f6b),
	.w2(32'hbbb0327b),
	.w3(32'hba6965f1),
	.w4(32'h3b5de93d),
	.w5(32'hbbea0f63),
	.w6(32'hbbb42220),
	.w7(32'hbb2fa490),
	.w8(32'hbbef82fe),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80dd33),
	.w1(32'hbb6f1243),
	.w2(32'hbb24311e),
	.w3(32'hbb32a57c),
	.w4(32'hbb16d82e),
	.w5(32'hb8c3106e),
	.w6(32'hbb53e895),
	.w7(32'hbb6c629d),
	.w8(32'hbb32dbc3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab83658),
	.w1(32'hba762877),
	.w2(32'hbb045284),
	.w3(32'hb9560041),
	.w4(32'hba6343a8),
	.w5(32'h3a5bd797),
	.w6(32'hbaa2e285),
	.w7(32'hbb188e98),
	.w8(32'hbb22d687),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e25e3),
	.w1(32'hbb9258d6),
	.w2(32'hbb511052),
	.w3(32'h3aa416a0),
	.w4(32'hbb4f967d),
	.w5(32'hba6f12a0),
	.w6(32'hba784787),
	.w7(32'hbac8a62a),
	.w8(32'h3a107268),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb790303),
	.w1(32'hbb48cfb2),
	.w2(32'hbade6e90),
	.w3(32'hbb853ba3),
	.w4(32'hbb174c88),
	.w5(32'h3aca502d),
	.w6(32'hbb0ca060),
	.w7(32'hbaa4e8da),
	.w8(32'hbaa34930),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a7160),
	.w1(32'h3b95b023),
	.w2(32'h3b88a209),
	.w3(32'hbaaddc94),
	.w4(32'h3b98881d),
	.w5(32'h3b9ff886),
	.w6(32'hbae1c81d),
	.w7(32'h3a8530d6),
	.w8(32'hb9f0d85d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16d61b),
	.w1(32'hbc3d06b6),
	.w2(32'hbbac12a7),
	.w3(32'hba21366b),
	.w4(32'hbc066a74),
	.w5(32'h3ba58908),
	.w6(32'hbc098f24),
	.w7(32'hbab2b790),
	.w8(32'h3ac85eb9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c854b),
	.w1(32'hbc6c9990),
	.w2(32'hbc2775b8),
	.w3(32'hbbd45ceb),
	.w4(32'hbc8a2bc5),
	.w5(32'hbba18d75),
	.w6(32'hbc5a1b58),
	.w7(32'hbc311c32),
	.w8(32'hbaf4362e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee536a),
	.w1(32'h3a816a65),
	.w2(32'hbbba36cf),
	.w3(32'hbb4ff29c),
	.w4(32'hbbe0a4b3),
	.w5(32'hbc11a0a8),
	.w6(32'hbb0caf3c),
	.w7(32'hbbe5997b),
	.w8(32'hbc29be48),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac4c78),
	.w1(32'hbabc3a16),
	.w2(32'h3a6d2ffb),
	.w3(32'hbb8ab276),
	.w4(32'hba8b00c2),
	.w5(32'h3a586f72),
	.w6(32'hbb7af1e3),
	.w7(32'hbb5c8df8),
	.w8(32'hba2f173e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95d51a),
	.w1(32'hbb80b0e2),
	.w2(32'h3aa77427),
	.w3(32'h393faa86),
	.w4(32'hba77bd2e),
	.w5(32'h3a466d59),
	.w6(32'hbb5896f6),
	.w7(32'hb98e681d),
	.w8(32'hbb7bb45a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca276c),
	.w1(32'h3b6ce172),
	.w2(32'h3a7d87ca),
	.w3(32'hb9998091),
	.w4(32'h3b50f749),
	.w5(32'hb909b5e8),
	.w6(32'hba25f205),
	.w7(32'hba71596c),
	.w8(32'hbb7a77d1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64afd6),
	.w1(32'hbbc8e61c),
	.w2(32'hbbb52874),
	.w3(32'hbb69f58d),
	.w4(32'hbb513efa),
	.w5(32'hb91f04ba),
	.w6(32'hbb949585),
	.w7(32'hbb690094),
	.w8(32'hbaef7898),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c9423),
	.w1(32'h372675c4),
	.w2(32'hb9894fdb),
	.w3(32'hb9e5077d),
	.w4(32'hba3010d0),
	.w5(32'hb99c4a61),
	.w6(32'h3a8b6afe),
	.w7(32'hbae60a70),
	.w8(32'hba1b00ae),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9372e78),
	.w1(32'hbaf8e6e0),
	.w2(32'hbaf99803),
	.w3(32'hbaffbfc2),
	.w4(32'hbb20ded8),
	.w5(32'hbb003b2e),
	.w6(32'h3a8dce8b),
	.w7(32'hbaec2d57),
	.w8(32'hbb3787da),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf84449),
	.w1(32'hbaee5bb2),
	.w2(32'hbaaa2dd1),
	.w3(32'hba8d821b),
	.w4(32'hbaecacee),
	.w5(32'h3a268524),
	.w6(32'hbb439a89),
	.w7(32'hbafcd276),
	.w8(32'h3a4b2e36),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb046d20),
	.w1(32'hb69eb6d6),
	.w2(32'hbb88df95),
	.w3(32'hba48c7d1),
	.w4(32'hb8d011a8),
	.w5(32'hbabe55fc),
	.w6(32'hba1a97e3),
	.w7(32'hbb00bf1d),
	.w8(32'hbb16a38a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97dbad),
	.w1(32'hbb073d24),
	.w2(32'hbaa152ca),
	.w3(32'h3a180955),
	.w4(32'hbb55c7e2),
	.w5(32'hbb0040ac),
	.w6(32'hbb073330),
	.w7(32'hbbadd7b2),
	.w8(32'hbb8a1f7f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae686b4),
	.w1(32'hba2f1dc2),
	.w2(32'hbb067c08),
	.w3(32'h387c6392),
	.w4(32'hbb5af4ca),
	.w5(32'h3b423dac),
	.w6(32'h3a899e6f),
	.w7(32'hba935e0e),
	.w8(32'hbb57b2a1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb999987),
	.w1(32'hbb194cf0),
	.w2(32'hbb2af12a),
	.w3(32'hbadb7156),
	.w4(32'hbae1f871),
	.w5(32'hba4ca9a1),
	.w6(32'hbb99cc6f),
	.w7(32'hbb9a003d),
	.w8(32'hbb688fa2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51dadf),
	.w1(32'hbc23f472),
	.w2(32'hbba1b0b7),
	.w3(32'hbca9b4b9),
	.w4(32'hbbc18898),
	.w5(32'h3ba31b9f),
	.w6(32'hbca04e95),
	.w7(32'h39aeb38f),
	.w8(32'h3b0a1ade),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00b996),
	.w1(32'h3b9a6a13),
	.w2(32'hbb4a6f38),
	.w3(32'h3ba021cb),
	.w4(32'h3b76be29),
	.w5(32'hb988ffbd),
	.w6(32'h3b456ce9),
	.w7(32'h3b35a3c3),
	.w8(32'h389d75d6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bd56e),
	.w1(32'hbb4ec546),
	.w2(32'h3ac19ed5),
	.w3(32'hbb83468a),
	.w4(32'hbaa19660),
	.w5(32'h3bfc92c0),
	.w6(32'hbb37320e),
	.w7(32'h3b18e15a),
	.w8(32'h3ba7f07f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a4233),
	.w1(32'h3ac0992c),
	.w2(32'h39992e57),
	.w3(32'h3b3f54c1),
	.w4(32'h3b3d0817),
	.w5(32'hb9fea721),
	.w6(32'hb8a15236),
	.w7(32'h3a88d60c),
	.w8(32'hbac5ab76),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64d84),
	.w1(32'hba989c1b),
	.w2(32'h3a3b36ab),
	.w3(32'hbb24f96b),
	.w4(32'h3b05053a),
	.w5(32'h3b312f33),
	.w6(32'hbb1ee577),
	.w7(32'hb869c62a),
	.w8(32'h3a8745c5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84db0a),
	.w1(32'h3ac71793),
	.w2(32'h3a0463dd),
	.w3(32'hb990da18),
	.w4(32'h3b1715d9),
	.w5(32'h374c752e),
	.w6(32'hbaf285d3),
	.w7(32'h3b3d70bd),
	.w8(32'hbaa86cc7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6daf05),
	.w1(32'h3b12a9aa),
	.w2(32'hbb04c39e),
	.w3(32'hb94e4b2b),
	.w4(32'hbae87fb3),
	.w5(32'hbbb525a1),
	.w6(32'h3b3bfed4),
	.w7(32'hbb081f53),
	.w8(32'hbbaf1eef),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08137b),
	.w1(32'hbb7ace13),
	.w2(32'hbb72b218),
	.w3(32'h39cec358),
	.w4(32'hbb7f110c),
	.w5(32'hbaa7ecdd),
	.w6(32'hbb3a6a8a),
	.w7(32'hbb1068fa),
	.w8(32'hbb057d7a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b64f),
	.w1(32'hba69ad13),
	.w2(32'hbb9dff64),
	.w3(32'hbb700cde),
	.w4(32'hba808263),
	.w5(32'hbb1bdaeb),
	.w6(32'hbb8f9d07),
	.w7(32'hbb400a88),
	.w8(32'hbbcc7a31),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a9dc1),
	.w1(32'hbba3b912),
	.w2(32'hbb938c94),
	.w3(32'h3b41247a),
	.w4(32'h3aa641a0),
	.w5(32'hba5de486),
	.w6(32'h3b7a2c88),
	.w7(32'h3a524d50),
	.w8(32'hbab811d8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32e0e7),
	.w1(32'hbc6909c7),
	.w2(32'hbbdd51e0),
	.w3(32'hbc8a6c50),
	.w4(32'hbc433b35),
	.w5(32'h3b9a5ebc),
	.w6(32'hbc8badc1),
	.w7(32'hbbb34085),
	.w8(32'h3a3ee94a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba692c2c),
	.w1(32'h3b343652),
	.w2(32'hba17fa67),
	.w3(32'h3bdc7ec8),
	.w4(32'h3bb61e44),
	.w5(32'hbb69367c),
	.w6(32'h3adc6732),
	.w7(32'h39303e47),
	.w8(32'hbc3d4a52),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11458c),
	.w1(32'h3b5c6ab6),
	.w2(32'h3a9a3b3b),
	.w3(32'h3b0ba660),
	.w4(32'h39990465),
	.w5(32'hbbcfcd36),
	.w6(32'hbaa2ec8a),
	.w7(32'hbbac41ba),
	.w8(32'hbbefd4d6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0faac3),
	.w1(32'hbb92f294),
	.w2(32'hbb022b86),
	.w3(32'h3954b254),
	.w4(32'hba6cd852),
	.w5(32'h3bf228e2),
	.w6(32'hba6f0336),
	.w7(32'h3b186aed),
	.w8(32'hbb5ac728),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9a62a),
	.w1(32'hb6b94f6d),
	.w2(32'hb9c25993),
	.w3(32'hbab030d3),
	.w4(32'h39bf9dba),
	.w5(32'hba0eca65),
	.w6(32'hbaba3f5c),
	.w7(32'hbb227393),
	.w8(32'hbad3f39a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddd7c5),
	.w1(32'hbcd03273),
	.w2(32'hbc909dcc),
	.w3(32'hbc3a247d),
	.w4(32'hbc93430b),
	.w5(32'hbb798c17),
	.w6(32'hbca333fd),
	.w7(32'hbc2482db),
	.w8(32'hbac72df3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b653273),
	.w1(32'hb913ac5b),
	.w2(32'hbb99a7e5),
	.w3(32'h3bc4f46f),
	.w4(32'hba054f6d),
	.w5(32'hbbedb233),
	.w6(32'h3bcdbfc2),
	.w7(32'h3b12330d),
	.w8(32'hbb794ec9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba170695),
	.w1(32'hba1187d5),
	.w2(32'h3a78507d),
	.w3(32'h39314127),
	.w4(32'h3afd9502),
	.w5(32'h39ba6e97),
	.w6(32'h3a0e297b),
	.w7(32'hb9e98a80),
	.w8(32'hb8034d33),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a005093),
	.w1(32'h3aa0cb20),
	.w2(32'hbb0292e8),
	.w3(32'h3a0d4ce4),
	.w4(32'h3ad56eb0),
	.w5(32'h390b1f0b),
	.w6(32'hba86c3e8),
	.w7(32'hbb1d5c8c),
	.w8(32'h3a11e7b6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a9c0d),
	.w1(32'h3b80d39b),
	.w2(32'hba19348c),
	.w3(32'hb9d13df5),
	.w4(32'hba3fd061),
	.w5(32'hba8aae3b),
	.w6(32'hbb625549),
	.w7(32'hbb468f65),
	.w8(32'hbbc5aa0a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba948d76),
	.w1(32'h3b4f3907),
	.w2(32'hb8abf276),
	.w3(32'h3b4191f9),
	.w4(32'h3ac1407b),
	.w5(32'hba43b4fe),
	.w6(32'h3b296e0b),
	.w7(32'hbb0da64d),
	.w8(32'hbb62f37c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb691212),
	.w1(32'hbb9bf6f6),
	.w2(32'hbc0d9fcd),
	.w3(32'h3b1e5b8b),
	.w4(32'h3aa38e65),
	.w5(32'hbbf21b5e),
	.w6(32'h3aa68852),
	.w7(32'hbae8899d),
	.w8(32'hbbf3f953),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c0fc2),
	.w1(32'h3a6edafd),
	.w2(32'hbb0bc41c),
	.w3(32'h394e940c),
	.w4(32'hb9ed62d0),
	.w5(32'hbb82c3f0),
	.w6(32'hbafbd6f1),
	.w7(32'hbb2bb20b),
	.w8(32'hbb96454f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf366c),
	.w1(32'h3afe814a),
	.w2(32'h3b1348cf),
	.w3(32'hbb640d73),
	.w4(32'h3a0b5308),
	.w5(32'h3b7730b9),
	.w6(32'hbaa27db8),
	.w7(32'h3b09f82d),
	.w8(32'h3ac7ff16),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae98d4),
	.w1(32'hbb75d8a6),
	.w2(32'hbb421418),
	.w3(32'hbbbe7b29),
	.w4(32'hbaece8da),
	.w5(32'h3b06324d),
	.w6(32'hbb9fcb6e),
	.w7(32'hbba6c00f),
	.w8(32'hbb47a643),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3a1d),
	.w1(32'h3ae1eca3),
	.w2(32'hbb6af507),
	.w3(32'h3b0ae690),
	.w4(32'h3b3e9117),
	.w5(32'hbb714050),
	.w6(32'h39c1bf38),
	.w7(32'hbaf1af97),
	.w8(32'hbba2ea48),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a260ddc),
	.w1(32'hbae20663),
	.w2(32'h3a0a986a),
	.w3(32'hba783418),
	.w4(32'hbb4a73c9),
	.w5(32'h39fd3520),
	.w6(32'hb9be263d),
	.w7(32'hbba2b0d0),
	.w8(32'hba7680aa),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cad15),
	.w1(32'h39f4b9cd),
	.w2(32'h399e4975),
	.w3(32'hbafe4111),
	.w4(32'h3a1a2a75),
	.w5(32'h39759530),
	.w6(32'hba7d4a17),
	.w7(32'hba968f21),
	.w8(32'hb941af52),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eda8b),
	.w1(32'hbb512e75),
	.w2(32'hbafff88e),
	.w3(32'h3b35dc82),
	.w4(32'hba971865),
	.w5(32'hba978094),
	.w6(32'h3a9736f1),
	.w7(32'h39571a81),
	.w8(32'h3a2492a7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2574a),
	.w1(32'hb9c5b171),
	.w2(32'h39ddcc93),
	.w3(32'hbaf22571),
	.w4(32'hbb01784b),
	.w5(32'h3b277ffc),
	.w6(32'h3a901dac),
	.w7(32'h39ecb98f),
	.w8(32'hbae2ddac),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabefed2),
	.w1(32'h3bbe2cc4),
	.w2(32'h3adae967),
	.w3(32'h3b12afcf),
	.w4(32'h396ea783),
	.w5(32'hbb9d119e),
	.w6(32'hb999391e),
	.w7(32'hbbb19105),
	.w8(32'hbc01e27a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387e8a79),
	.w1(32'hbb0b6ca1),
	.w2(32'hba5e9af8),
	.w3(32'hb973742a),
	.w4(32'hba052cec),
	.w5(32'h3aea3e2c),
	.w6(32'hba0bdefa),
	.w7(32'hb9f8ddeb),
	.w8(32'h3a15433b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74390),
	.w1(32'hbb861b68),
	.w2(32'hbb3738db),
	.w3(32'hbaf75812),
	.w4(32'hbb4c4038),
	.w5(32'h3abfb52d),
	.w6(32'hbb6d06df),
	.w7(32'hbb87f9e1),
	.w8(32'hbb7981c8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad09e65),
	.w1(32'h3bcb4d0c),
	.w2(32'hba48a323),
	.w3(32'h39e3b61a),
	.w4(32'h3a2b9d5e),
	.w5(32'hbbb37004),
	.w6(32'hbaf48cbf),
	.w7(32'hbbc047da),
	.w8(32'hbc43bf0e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98207b2),
	.w1(32'h3b7ab702),
	.w2(32'h3b2922ef),
	.w3(32'hba4c3bad),
	.w4(32'h3b28f098),
	.w5(32'h3a9acb3c),
	.w6(32'hbb452670),
	.w7(32'h3a93f724),
	.w8(32'h3ab4e93b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ee3f),
	.w1(32'h39d608b3),
	.w2(32'h39bd1b60),
	.w3(32'h3b553a49),
	.w4(32'hbb248e5e),
	.w5(32'h3b63a16f),
	.w6(32'h3a59e608),
	.w7(32'hbb08b109),
	.w8(32'hbad96fb1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd6770),
	.w1(32'hbab4029a),
	.w2(32'hba28e1fb),
	.w3(32'h3a226610),
	.w4(32'h3aa02f22),
	.w5(32'h3b26ea72),
	.w6(32'hb943a8f2),
	.w7(32'hbabfce88),
	.w8(32'hbaee708f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1773a),
	.w1(32'h3a963182),
	.w2(32'hbb3eaa89),
	.w3(32'h3b1edfb2),
	.w4(32'h3a3a4583),
	.w5(32'hbb8df9a7),
	.w6(32'h39dd3c56),
	.w7(32'h38e04997),
	.w8(32'hbb883f36),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a697eba),
	.w1(32'h3a25ed5a),
	.w2(32'h3aa64bd7),
	.w3(32'hbb949702),
	.w4(32'h3a3395bb),
	.w5(32'h3a7a5ef9),
	.w6(32'hbba85604),
	.w7(32'hbba66395),
	.w8(32'hbb9b7baf),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1c9e),
	.w1(32'h39238915),
	.w2(32'h3a8dc9ce),
	.w3(32'hbb8009df),
	.w4(32'h39424af2),
	.w5(32'h37dca001),
	.w6(32'hbb5aeca3),
	.w7(32'hb7dff385),
	.w8(32'hbad4c914),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72bffd),
	.w1(32'hbb685292),
	.w2(32'hbb2aa426),
	.w3(32'hb9e5f2ba),
	.w4(32'hba575192),
	.w5(32'hbb005963),
	.w6(32'hbac95d2e),
	.w7(32'h366d0ea6),
	.w8(32'hba814601),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf991d),
	.w1(32'hba8f53f8),
	.w2(32'h39b79503),
	.w3(32'h3a21c3aa),
	.w4(32'hbac9eb0f),
	.w5(32'h3a949693),
	.w6(32'h3a35c3e3),
	.w7(32'hbb3b00e3),
	.w8(32'hbb2977ba),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c713e),
	.w1(32'hba7a2f0c),
	.w2(32'hbac99f25),
	.w3(32'hba08fd75),
	.w4(32'hbacc333b),
	.w5(32'hbb24fb76),
	.w6(32'hb831df45),
	.w7(32'hbb3f4191),
	.w8(32'hbad17bb5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb259bab),
	.w1(32'h3b074946),
	.w2(32'h3b1b6417),
	.w3(32'hbb6228c5),
	.w4(32'h3ae2d9c6),
	.w5(32'h3b059aca),
	.w6(32'hba8a5967),
	.w7(32'h3b1aaa05),
	.w8(32'h3ae18662),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62d69b),
	.w1(32'h3c01295a),
	.w2(32'h3befe9bd),
	.w3(32'h3a920dca),
	.w4(32'h3bb29554),
	.w5(32'h3a8eec90),
	.w6(32'h3a0c8c92),
	.w7(32'h3a9a8207),
	.w8(32'h3b30bb71),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb876fb),
	.w1(32'hbc1a247d),
	.w2(32'hbbc80cf8),
	.w3(32'hbc28ea3e),
	.w4(32'hbc1625b0),
	.w5(32'h3af68cfb),
	.w6(32'hbc1a278c),
	.w7(32'hbb9021d1),
	.w8(32'hbbba3874),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e6b87),
	.w1(32'hbb4e2df5),
	.w2(32'hbb6e23e4),
	.w3(32'h3b110116),
	.w4(32'hbb9fa502),
	.w5(32'hbbffe183),
	.w6(32'hbb5c627d),
	.w7(32'hbbd26259),
	.w8(32'hbbd4c408),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecda50),
	.w1(32'hbae1cbb0),
	.w2(32'hbb057860),
	.w3(32'hbb27ad56),
	.w4(32'hb809442a),
	.w5(32'hba1c6e77),
	.w6(32'hbbae7ae3),
	.w7(32'hbb9629e1),
	.w8(32'hbbab092e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc28277),
	.w1(32'hbc010051),
	.w2(32'hbbaeb4c8),
	.w3(32'hbc0cb45f),
	.w4(32'hbb6405d8),
	.w5(32'h3aabc3fb),
	.w6(32'hbbf6e539),
	.w7(32'hba245a06),
	.w8(32'hbac16a80),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a1a6d),
	.w1(32'h3b19e7e4),
	.w2(32'h3b6eac76),
	.w3(32'hbb158065),
	.w4(32'hba06a803),
	.w5(32'h3b144ab1),
	.w6(32'hba863bbb),
	.w7(32'hba995ca2),
	.w8(32'h3a47ef5d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9612c13),
	.w1(32'hbad800cb),
	.w2(32'hbae3ae01),
	.w3(32'h3af0246d),
	.w4(32'hbb00ccb6),
	.w5(32'hba0cc6b7),
	.w6(32'hb8ed06d7),
	.w7(32'hbad9198b),
	.w8(32'hbb0560bc),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36c2ce),
	.w1(32'hbae09c76),
	.w2(32'hbb5bf519),
	.w3(32'hb81ece74),
	.w4(32'hbadcadb9),
	.w5(32'hbb6ffe5b),
	.w6(32'h3a622b95),
	.w7(32'hbb9444ad),
	.w8(32'hbb69dabc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926e5f),
	.w1(32'h3b155779),
	.w2(32'hbaf41bc3),
	.w3(32'h39689817),
	.w4(32'hba29289e),
	.w5(32'hbbfdb2ff),
	.w6(32'h3a98e335),
	.w7(32'hbb5bdf9f),
	.w8(32'hbc0c22fc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aa19f),
	.w1(32'hbb87139d),
	.w2(32'hbb84d907),
	.w3(32'hbb920a50),
	.w4(32'hbb683327),
	.w5(32'hba00c79f),
	.w6(32'hbb84a99e),
	.w7(32'hbb7a8f93),
	.w8(32'hbab5df74),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04ae6d),
	.w1(32'hbaf13044),
	.w2(32'hba18c403),
	.w3(32'hba76c576),
	.w4(32'hbb013f7b),
	.w5(32'h3abe3038),
	.w6(32'h3a1882fa),
	.w7(32'hbb15cc45),
	.w8(32'hb971e163),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44e002),
	.w1(32'h3a5f12b6),
	.w2(32'h3a4f3f10),
	.w3(32'hb9132deb),
	.w4(32'hb9d06aff),
	.w5(32'h3b1dc511),
	.w6(32'h39c690f2),
	.w7(32'hbb110b22),
	.w8(32'hbab8ecfc),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cceae),
	.w1(32'h3ad21149),
	.w2(32'h3b0baa34),
	.w3(32'h3a9e1bb7),
	.w4(32'hbaa224ec),
	.w5(32'hbb3ade93),
	.w6(32'hbaec4fae),
	.w7(32'hba00f25b),
	.w8(32'hbb0db367),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef84a4),
	.w1(32'hba84f65c),
	.w2(32'hbb3f5948),
	.w3(32'h3a81b91a),
	.w4(32'hbbbd670d),
	.w5(32'hbb68a5a9),
	.w6(32'hbb6fccd5),
	.w7(32'hbbe7c54f),
	.w8(32'hbb34c8d2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1897f),
	.w1(32'hb90e0901),
	.w2(32'hbb7f5031),
	.w3(32'hba94dea2),
	.w4(32'hba6abcdc),
	.w5(32'hb7b327ae),
	.w6(32'hba4cf2dc),
	.w7(32'hbb3b96e9),
	.w8(32'hbb988423),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41e3d2),
	.w1(32'h3966e6cf),
	.w2(32'hba3ca6a9),
	.w3(32'hbadcec3d),
	.w4(32'h3afa65e8),
	.w5(32'h3aef8ffd),
	.w6(32'hbb1d7344),
	.w7(32'h3a9c8b3d),
	.w8(32'h3b0ffa36),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91886a),
	.w1(32'h3af90931),
	.w2(32'hbbc19f78),
	.w3(32'h3a866690),
	.w4(32'hba0c7dd0),
	.w5(32'hbb827912),
	.w6(32'h3a286744),
	.w7(32'hbb473888),
	.w8(32'hbb4183ed),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75f9be),
	.w1(32'h3abb97c6),
	.w2(32'hbb139d24),
	.w3(32'hba98c53a),
	.w4(32'hbab3d9c6),
	.w5(32'hbb769a18),
	.w6(32'h3a5a52ba),
	.w7(32'hbbbc1eb5),
	.w8(32'hbbca5e8a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb774fd),
	.w1(32'hbb93446a),
	.w2(32'hbbe64216),
	.w3(32'hbb2c1aa7),
	.w4(32'hb8ec422d),
	.w5(32'h3a3497b8),
	.w6(32'hbb8720d3),
	.w7(32'hba8efec4),
	.w8(32'hbb4d4960),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09d493),
	.w1(32'h3b82a381),
	.w2(32'hbada5e8e),
	.w3(32'hb8f3c211),
	.w4(32'h3ba15788),
	.w5(32'hbb96e894),
	.w6(32'hba983910),
	.w7(32'h39d1ccb7),
	.w8(32'hbba2cb82),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39648436),
	.w1(32'h39524f43),
	.w2(32'hbb8aa7d0),
	.w3(32'hbaa570e6),
	.w4(32'h3b5efa13),
	.w5(32'hbb8e4ef8),
	.w6(32'hbb3dda34),
	.w7(32'hba802d39),
	.w8(32'hbb5e13db),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb453cdf),
	.w1(32'hbaba2b4c),
	.w2(32'hbabfa5d4),
	.w3(32'hbb702bcb),
	.w4(32'hba54f910),
	.w5(32'h3a813fdb),
	.w6(32'hbb033a59),
	.w7(32'h39b216c1),
	.w8(32'h39e0d46c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5504bd),
	.w1(32'h3a7dc173),
	.w2(32'hbaa2ab9e),
	.w3(32'h3aacca85),
	.w4(32'h39e52fcc),
	.w5(32'hba9f5b87),
	.w6(32'h3a798390),
	.w7(32'hba5fa03f),
	.w8(32'hbb4290f7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd0c5f),
	.w1(32'hba6ddcf5),
	.w2(32'hba87b859),
	.w3(32'hba4cad28),
	.w4(32'hb897180e),
	.w5(32'hbaf0c988),
	.w6(32'hb9afe204),
	.w7(32'hbb6dbdcc),
	.w8(32'hbb9bcf9e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b280875),
	.w1(32'h3b63c14c),
	.w2(32'h3b454ce5),
	.w3(32'h3ad5a25c),
	.w4(32'h3b6ffdd3),
	.w5(32'h3a90afc3),
	.w6(32'hbb471e7e),
	.w7(32'h3b18e62b),
	.w8(32'h3a329d61),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec2926),
	.w1(32'hbba29b6c),
	.w2(32'hbb813e1a),
	.w3(32'hb915bdee),
	.w4(32'hbb3061c7),
	.w5(32'h3b6d2647),
	.w6(32'h39a7b3cb),
	.w7(32'hba0dedbf),
	.w8(32'h3a33ec6d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7316e5),
	.w1(32'h39e9700e),
	.w2(32'h395b80cd),
	.w3(32'h3b01f8d7),
	.w4(32'hba86d60c),
	.w5(32'hbb063701),
	.w6(32'hbb3ef55c),
	.w7(32'hbb34bc7e),
	.w8(32'hbaeac488),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecea52),
	.w1(32'hbab6cf96),
	.w2(32'hbb4707b5),
	.w3(32'hbb18f30b),
	.w4(32'hba3627b7),
	.w5(32'h3b7b7cb0),
	.w6(32'hba3ddfc5),
	.w7(32'hb8b52554),
	.w8(32'hbb34c2e3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69a5b7),
	.w1(32'h3adb24b3),
	.w2(32'hb9cdc64a),
	.w3(32'h3ad91214),
	.w4(32'hbab6d6b7),
	.w5(32'h3a4a776f),
	.w6(32'h3b0537bf),
	.w7(32'h3a71b088),
	.w8(32'hbb0091f1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6858fa),
	.w1(32'hbb30ded9),
	.w2(32'hbb54a963),
	.w3(32'hbb4f2ea8),
	.w4(32'hb8b5e413),
	.w5(32'hbb404c46),
	.w6(32'hbab0b498),
	.w7(32'hbb3669f7),
	.w8(32'hbb402b87),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917db6),
	.w1(32'h3a9c1636),
	.w2(32'h39d73820),
	.w3(32'hbb7b6aac),
	.w4(32'h3aaf8fc4),
	.w5(32'h3a600511),
	.w6(32'h39c6e84d),
	.w7(32'hba27c14d),
	.w8(32'hb9d16f8b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9b78a),
	.w1(32'h3b7a90c9),
	.w2(32'h3b000e98),
	.w3(32'h3b8b1c6d),
	.w4(32'h3a1059da),
	.w5(32'h3b02e4d7),
	.w6(32'h3adcb843),
	.w7(32'h3b288d6a),
	.w8(32'h3adbe0fd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5233f),
	.w1(32'hb8e0c586),
	.w2(32'hb94d2586),
	.w3(32'h3aca1acc),
	.w4(32'hbaa7db8b),
	.w5(32'hba94a6f3),
	.w6(32'hbb026b05),
	.w7(32'hb8a3f932),
	.w8(32'hba0c759f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a9530),
	.w1(32'h39d3b31d),
	.w2(32'hb8cfd65b),
	.w3(32'hba01f41b),
	.w4(32'hb7c57de6),
	.w5(32'hb8f5ce6c),
	.w6(32'hb9a5e9c5),
	.w7(32'hba154958),
	.w8(32'h3a19187e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a97ad),
	.w1(32'h3ac3e690),
	.w2(32'hbb27e11b),
	.w3(32'h3b2626b2),
	.w4(32'h3a3b376e),
	.w5(32'hbb1f38f9),
	.w6(32'h3a748082),
	.w7(32'hbafe2619),
	.w8(32'hbb373614),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb725b03),
	.w1(32'hbb8cd213),
	.w2(32'hbb83fd6e),
	.w3(32'hbb6f31f8),
	.w4(32'hbbb71270),
	.w5(32'hbb0c0ebe),
	.w6(32'hbc249ad0),
	.w7(32'hbbdd0f8e),
	.w8(32'hbbea9c04),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba708d82),
	.w1(32'h3aa889c6),
	.w2(32'h3a98e57a),
	.w3(32'hbb838182),
	.w4(32'h3a22f250),
	.w5(32'hba04295c),
	.w6(32'hbb4d111c),
	.w7(32'h3a46e12d),
	.w8(32'hb95f6664),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af5d3b),
	.w1(32'h3a018363),
	.w2(32'hbb924f3c),
	.w3(32'h3aa96099),
	.w4(32'h3967042f),
	.w5(32'hbbf31553),
	.w6(32'hba4c92d7),
	.w7(32'hbb83d33e),
	.w8(32'hbc0042ae),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb071a00),
	.w1(32'h39d3c50c),
	.w2(32'h3b0ab8f2),
	.w3(32'hba0641bc),
	.w4(32'hbb0a5f82),
	.w5(32'hba9d21fd),
	.w6(32'h3a85f12b),
	.w7(32'hbb382f49),
	.w8(32'h39161f93),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9a323),
	.w1(32'hbafa3881),
	.w2(32'hbb2c7746),
	.w3(32'hbb31f532),
	.w4(32'h3a340587),
	.w5(32'hba5ec57e),
	.w6(32'hbad83673),
	.w7(32'h3a219915),
	.w8(32'h3a943f31),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28dc1a),
	.w1(32'hbb9ca510),
	.w2(32'hbb80c647),
	.w3(32'hbabb78b0),
	.w4(32'hbaa7b832),
	.w5(32'hba67288a),
	.w6(32'hbaa1be9f),
	.w7(32'hbb1b2768),
	.w8(32'hbad31df6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba19696),
	.w1(32'hbb290f44),
	.w2(32'hbb0bdee7),
	.w3(32'hbbb885fd),
	.w4(32'hbb1e9911),
	.w5(32'hb9ac15bb),
	.w6(32'hbba3e255),
	.w7(32'hbbbe7914),
	.w8(32'hbb8a82b1),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bebb5),
	.w1(32'hbb208c99),
	.w2(32'hbaf13458),
	.w3(32'h3973db0c),
	.w4(32'hbb194fda),
	.w5(32'hbad843af),
	.w6(32'h392fb641),
	.w7(32'hba9eb530),
	.w8(32'h387a17fd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1906),
	.w1(32'h3b69357c),
	.w2(32'h3b1befc2),
	.w3(32'hbb1b759d),
	.w4(32'h3ab13bac),
	.w5(32'h39fde623),
	.w6(32'hba357772),
	.w7(32'hbad0096a),
	.w8(32'hbb56c26e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c6dd),
	.w1(32'h39fc589f),
	.w2(32'h3a2bfb16),
	.w3(32'h3b15c3bd),
	.w4(32'hba862164),
	.w5(32'hba969c6a),
	.w6(32'hbaf38886),
	.w7(32'hbb8cbf4b),
	.w8(32'hbb0b8676),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a9fb3),
	.w1(32'hbab543fa),
	.w2(32'hb942cfb6),
	.w3(32'h39c38ffd),
	.w4(32'h39cc5d30),
	.w5(32'hba0255e8),
	.w6(32'hba8e8bbe),
	.w7(32'hbb04c60d),
	.w8(32'h39b9768e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e25a7),
	.w1(32'hbb4e596d),
	.w2(32'hbba0ecbd),
	.w3(32'hba88a461),
	.w4(32'hb98550b5),
	.w5(32'hba419c2f),
	.w6(32'hba81f1e2),
	.w7(32'h38d8e88e),
	.w8(32'hbae52838),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b0b68),
	.w1(32'h3a974650),
	.w2(32'hba779348),
	.w3(32'hbb9be11a),
	.w4(32'hba522839),
	.w5(32'hba87a0b3),
	.w6(32'hbb366264),
	.w7(32'hbb825bd0),
	.w8(32'hbb8d5d98),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f59fd),
	.w1(32'hbb492fc4),
	.w2(32'hbb738527),
	.w3(32'hba1817dc),
	.w4(32'hbb759193),
	.w5(32'hbb027bcd),
	.w6(32'hbb2a5abf),
	.w7(32'hbb1a9c46),
	.w8(32'hbb156f9e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1b424),
	.w1(32'hb87eed2b),
	.w2(32'h39b59e1a),
	.w3(32'hbb71eff5),
	.w4(32'hbb1c3308),
	.w5(32'h3a8aded9),
	.w6(32'hbb50fb10),
	.w7(32'hbb51130e),
	.w8(32'h380d902f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47e38e),
	.w1(32'hbad1c6a0),
	.w2(32'hba1a6d89),
	.w3(32'hb886f695),
	.w4(32'hbb4cbd0d),
	.w5(32'hbade2ae9),
	.w6(32'hb9e9a7f8),
	.w7(32'hbb5f842f),
	.w8(32'hbb7631b0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac73e7a),
	.w1(32'hbb741db3),
	.w2(32'h3ad3a2ba),
	.w3(32'h3b0a35ab),
	.w4(32'h3aef1e9f),
	.w5(32'h3af01ec3),
	.w6(32'h3941a0ef),
	.w7(32'h394af520),
	.w8(32'hbb83a5ec),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee5948),
	.w1(32'hbb1172cd),
	.w2(32'hbb4bcede),
	.w3(32'h3b02e478),
	.w4(32'h3a5e4ca6),
	.w5(32'h3a4c29dc),
	.w6(32'hbaf98aef),
	.w7(32'hb9ba5476),
	.w8(32'h3b132964),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43e96f),
	.w1(32'hbb9a0df8),
	.w2(32'hbb32deb8),
	.w3(32'hba9079e7),
	.w4(32'h3a8b3b88),
	.w5(32'hb99847ad),
	.w6(32'h3b027fab),
	.w7(32'h3b081388),
	.w8(32'h3b386eac),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bcc22),
	.w1(32'hbb8b39c9),
	.w2(32'hbba0f232),
	.w3(32'hbb98e78f),
	.w4(32'hbadd8970),
	.w5(32'h3acf7086),
	.w6(32'h3a8ae617),
	.w7(32'h39866634),
	.w8(32'hb8355c95),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad0502),
	.w1(32'h3bb79274),
	.w2(32'hbb1eabec),
	.w3(32'hb9d2f29b),
	.w4(32'h3badb008),
	.w5(32'hbb9a6e0d),
	.w6(32'hbb26a59c),
	.w7(32'h39b97449),
	.w8(32'hbb661f71),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b8115),
	.w1(32'h3a4d0d32),
	.w2(32'h3a020f48),
	.w3(32'h39cbb88d),
	.w4(32'hba09366e),
	.w5(32'h392c7df0),
	.w6(32'hbac0730d),
	.w7(32'hbac00f3f),
	.w8(32'hb9d8297b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0be918),
	.w1(32'hb8d7a018),
	.w2(32'hba0ec049),
	.w3(32'h3a8d1e19),
	.w4(32'hbacbdd1b),
	.w5(32'hbb28013f),
	.w6(32'h37a455f0),
	.w7(32'hbb22537b),
	.w8(32'hba91d291),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10e68f),
	.w1(32'hba1e9ae2),
	.w2(32'h3a9857b7),
	.w3(32'hbaecb4f9),
	.w4(32'hbaa37db7),
	.w5(32'h3a5ee38f),
	.w6(32'h3a3e3b84),
	.w7(32'h394ebad4),
	.w8(32'h3af6a7e3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba703f34),
	.w1(32'h3ade768e),
	.w2(32'h3b816d19),
	.w3(32'hb98cd98a),
	.w4(32'h3a5ccdde),
	.w5(32'h3b06395d),
	.w6(32'h3ae3d0cd),
	.w7(32'hba1fb44d),
	.w8(32'hb9a592cd),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb898d1),
	.w1(32'h3b9b26db),
	.w2(32'h3b01da59),
	.w3(32'h3b7bbf25),
	.w4(32'h3b858995),
	.w5(32'h3aecbd50),
	.w6(32'h3a5a6a1a),
	.w7(32'h3b53fd66),
	.w8(32'hba0b4d66),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6aa90),
	.w1(32'hb994aedf),
	.w2(32'hba923503),
	.w3(32'h3b6f3da1),
	.w4(32'h3b592f35),
	.w5(32'h3b1df95c),
	.w6(32'hbb1c441f),
	.w7(32'hb9a0c646),
	.w8(32'hba96537d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b221cef),
	.w1(32'hbaa389b8),
	.w2(32'h3a52de07),
	.w3(32'h3b97ae10),
	.w4(32'hbbb15672),
	.w5(32'hbb42a30b),
	.w6(32'h3a0dccba),
	.w7(32'hbbd6179e),
	.w8(32'hbba8a57e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77aca2),
	.w1(32'hbbb04a74),
	.w2(32'hbb84cb11),
	.w3(32'hbaf58199),
	.w4(32'hbb17715b),
	.w5(32'hbb0fa1dd),
	.w6(32'hbac72dab),
	.w7(32'hbb774a12),
	.w8(32'hbac2bc7e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a0aea),
	.w1(32'h3b0c5247),
	.w2(32'hbb5d805d),
	.w3(32'hbb537c58),
	.w4(32'hbb981da1),
	.w5(32'hbb2b3ca7),
	.w6(32'hbb045fd8),
	.w7(32'hbb63bc45),
	.w8(32'hbbbac90a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb112498),
	.w1(32'hbb93e289),
	.w2(32'hbac74bbf),
	.w3(32'hbb924501),
	.w4(32'hbb6ad24b),
	.w5(32'h3b98357c),
	.w6(32'hbb8e81c1),
	.w7(32'hbb7254fc),
	.w8(32'h3a42edc1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdc014),
	.w1(32'h3b8b0d6c),
	.w2(32'hba357822),
	.w3(32'hbb7fbd31),
	.w4(32'h3b69f37d),
	.w5(32'hbab5f955),
	.w6(32'h39fee8a5),
	.w7(32'h3b86f77f),
	.w8(32'hba480319),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0ad62),
	.w1(32'hbbf44cdc),
	.w2(32'h3bc57475),
	.w3(32'h3a72c15e),
	.w4(32'hbbe3618c),
	.w5(32'h3be4da41),
	.w6(32'hbae246b5),
	.w7(32'hbaf48b83),
	.w8(32'h3bcd33c7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c4479),
	.w1(32'h3a724e40),
	.w2(32'h3bf1a6db),
	.w3(32'h3b2c3e2b),
	.w4(32'hba851dff),
	.w5(32'hbb15980d),
	.w6(32'h3b4f0734),
	.w7(32'hbab443b5),
	.w8(32'h3a011b96),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ed450),
	.w1(32'h3bda441e),
	.w2(32'h3be23c70),
	.w3(32'hbb0d92ae),
	.w4(32'hbb7f7555),
	.w5(32'hba4bcba4),
	.w6(32'hbb4f57db),
	.w7(32'hbb363fe7),
	.w8(32'h3ae420e4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a802fd8),
	.w1(32'h3b6c4021),
	.w2(32'h3b0fab14),
	.w3(32'h3b70b120),
	.w4(32'h3b3bff00),
	.w5(32'h3a34bcc0),
	.w6(32'h3be23fad),
	.w7(32'h3b2949eb),
	.w8(32'hba52ffd7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4163),
	.w1(32'h3c675f59),
	.w2(32'h3c45d74f),
	.w3(32'h3b0b0362),
	.w4(32'h3c8c2a53),
	.w5(32'hba941d46),
	.w6(32'hba608a5e),
	.w7(32'h3a970b4a),
	.w8(32'h3a953fba),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6823b1),
	.w1(32'hbaa0aaa1),
	.w2(32'h3bd9a388),
	.w3(32'h3bbf3bf0),
	.w4(32'hbab32b8d),
	.w5(32'h3a2cbcac),
	.w6(32'h3ae0aa39),
	.w7(32'hb95dabd1),
	.w8(32'hbb0694c5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d8ef7),
	.w1(32'h3ba4b6d4),
	.w2(32'hbae49fd7),
	.w3(32'h3c00a6ce),
	.w4(32'h3b9a9113),
	.w5(32'hbb93ed88),
	.w6(32'hbb589607),
	.w7(32'h3ba76c1f),
	.w8(32'hbbc28e62),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb743083),
	.w1(32'hbae56187),
	.w2(32'h3afa5fbe),
	.w3(32'hbb16ca95),
	.w4(32'hbb27e719),
	.w5(32'hbbcde74a),
	.w6(32'hbb539ceb),
	.w7(32'hbbe515cb),
	.w8(32'hbbbc0453),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a80be),
	.w1(32'h3c625ab8),
	.w2(32'h3b554614),
	.w3(32'hbb9279b9),
	.w4(32'h3c4e95db),
	.w5(32'h39c2b270),
	.w6(32'hbb54497b),
	.w7(32'h3bc4e75e),
	.w8(32'h3a31c7d8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13d290),
	.w1(32'h3a02643d),
	.w2(32'hbaf44453),
	.w3(32'h3bb53f01),
	.w4(32'hb9303651),
	.w5(32'h3a5b75d8),
	.w6(32'h3aec5299),
	.w7(32'hba8ce7ac),
	.w8(32'h3a9afbca),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b986f),
	.w1(32'h3b823ca3),
	.w2(32'hba0b0a5c),
	.w3(32'hbad3b84b),
	.w4(32'hbaf4a2ed),
	.w5(32'hbb20a59d),
	.w6(32'hbb47b487),
	.w7(32'h3a9d005a),
	.w8(32'h3b758e1f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba282dca),
	.w1(32'h3ad59a78),
	.w2(32'h3b11a92e),
	.w3(32'h3bb99a5a),
	.w4(32'hbbcb7e84),
	.w5(32'h3c3ff1ee),
	.w6(32'h3b1f6a62),
	.w7(32'hb92f842c),
	.w8(32'h3b3f5408),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe92ae),
	.w1(32'hbc0900de),
	.w2(32'hbba760f3),
	.w3(32'hbbb5507d),
	.w4(32'hba913f8a),
	.w5(32'h3b73032b),
	.w6(32'hbbba572e),
	.w7(32'hbc0825e2),
	.w8(32'hbbb23516),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc063efc),
	.w1(32'h3a285ba0),
	.w2(32'h3aa5a280),
	.w3(32'hbb558560),
	.w4(32'hb96bb499),
	.w5(32'hbb905438),
	.w6(32'hbb9247ed),
	.w7(32'h3a37f132),
	.w8(32'h3b958e18),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98bda1),
	.w1(32'h3a8de082),
	.w2(32'h3b800c80),
	.w3(32'h3ad95e71),
	.w4(32'h3bf01a71),
	.w5(32'h3bdd9aff),
	.w6(32'h3ba8382a),
	.w7(32'h3b436b66),
	.w8(32'h3a04b224),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b2aa0),
	.w1(32'h37a4061c),
	.w2(32'h3b0d8b9a),
	.w3(32'h39922159),
	.w4(32'h3aa8ef7a),
	.w5(32'hbbd9c9ef),
	.w6(32'h3aad6555),
	.w7(32'h3b0c5160),
	.w8(32'h3ba0dd66),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1f582),
	.w1(32'h3b91425c),
	.w2(32'h3bf02276),
	.w3(32'h3b1a1270),
	.w4(32'h39a74b9e),
	.w5(32'hb990bf65),
	.w6(32'h3bd0dd74),
	.w7(32'h39c3d6cb),
	.w8(32'h3b8759be),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170136),
	.w1(32'h3a575e24),
	.w2(32'hbabc9784),
	.w3(32'h3c017bf8),
	.w4(32'hbb56f3ef),
	.w5(32'h3b2d5198),
	.w6(32'hbb8107b2),
	.w7(32'hbb6bbd21),
	.w8(32'hbb355d0d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc216408),
	.w1(32'hbc4de749),
	.w2(32'hbb36a7c9),
	.w3(32'hbb9c99ae),
	.w4(32'hbc190f0e),
	.w5(32'h3b04b747),
	.w6(32'hbb1a2398),
	.w7(32'hbb9ec8c7),
	.w8(32'h3b7acc23),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b277524),
	.w1(32'hbc26fcce),
	.w2(32'hbacabd7a),
	.w3(32'hbb98b813),
	.w4(32'hbc509e4e),
	.w5(32'h39e675b9),
	.w6(32'hbc85d0e3),
	.w7(32'hbb4f55f8),
	.w8(32'h3c44a4da),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c489f),
	.w1(32'h3b820751),
	.w2(32'hb9ff0d61),
	.w3(32'h3c035e06),
	.w4(32'hbb9e5735),
	.w5(32'hbb32fb58),
	.w6(32'h3bbba7cc),
	.w7(32'hbb658e1e),
	.w8(32'hbbdcc588),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e2130),
	.w1(32'h3b9c06e3),
	.w2(32'hbaf1b2d9),
	.w3(32'hbb15b630),
	.w4(32'h3a432bd2),
	.w5(32'hbb3cd64c),
	.w6(32'hbbcfb86e),
	.w7(32'hbbb44c27),
	.w8(32'hbbf2dd73),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e6bdf),
	.w1(32'h3bdaab06),
	.w2(32'h3b31fbdc),
	.w3(32'hbb8ac8b2),
	.w4(32'hbb98eaa8),
	.w5(32'hbb4c022b),
	.w6(32'hbbdc75e8),
	.w7(32'hbc0fcbbf),
	.w8(32'h3a10238e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c30bbf),
	.w1(32'h3aa16a7d),
	.w2(32'h3b9965df),
	.w3(32'h39848b8a),
	.w4(32'h3b808533),
	.w5(32'hbb371f9e),
	.w6(32'hb8b41982),
	.w7(32'h3b9c9bc2),
	.w8(32'h3b40f48c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ea87a),
	.w1(32'h3b57d3ac),
	.w2(32'h3b650cee),
	.w3(32'h3adad5df),
	.w4(32'hbad98680),
	.w5(32'hba47eb4f),
	.w6(32'h3a7724f9),
	.w7(32'h3b2f9a72),
	.w8(32'h3c2636ff),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80b14c),
	.w1(32'h3b67a5fe),
	.w2(32'hbb28d696),
	.w3(32'h3b3859c2),
	.w4(32'hbb039788),
	.w5(32'hbc2b74ce),
	.w6(32'h3b76c3c9),
	.w7(32'hbac522c5),
	.w8(32'hbbd87c24),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfcccd),
	.w1(32'hb92f3784),
	.w2(32'hba275f76),
	.w3(32'hbb0aa77a),
	.w4(32'hbb3084c9),
	.w5(32'h3a68d4e8),
	.w6(32'hbba53fb2),
	.w7(32'hbb8eb29f),
	.w8(32'h3b2c2fc7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f10c4a),
	.w1(32'h3a34d062),
	.w2(32'h3adc1108),
	.w3(32'h3a7b6550),
	.w4(32'hbb282593),
	.w5(32'h3b739b77),
	.w6(32'h3b9ba93a),
	.w7(32'hbbb3ec03),
	.w8(32'hbc3ec31a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0559e1),
	.w1(32'h3b912b52),
	.w2(32'h3ae2f0a0),
	.w3(32'h3b913e08),
	.w4(32'hbb470602),
	.w5(32'hbbbd6576),
	.w6(32'h39f96de2),
	.w7(32'hbc049096),
	.w8(32'hbbc86ffa),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac761f),
	.w1(32'h3ac99cbc),
	.w2(32'h39f4abdf),
	.w3(32'hba0c5396),
	.w4(32'h3b166959),
	.w5(32'h3b4918df),
	.w6(32'hbb6edd43),
	.w7(32'hbb2b5ebe),
	.w8(32'h3aefdf56),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfb2e5),
	.w1(32'hbc2df0f6),
	.w2(32'hbc28c4a2),
	.w3(32'hbc0376ab),
	.w4(32'hbc35ec29),
	.w5(32'hbc46af90),
	.w6(32'hbc22e277),
	.w7(32'hbc024c80),
	.w8(32'hb90f10a1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38ab3a),
	.w1(32'hbb14f8d3),
	.w2(32'hbba52f45),
	.w3(32'hbaaaa954),
	.w4(32'hba234043),
	.w5(32'h3b6bb0be),
	.w6(32'hb9d40844),
	.w7(32'hbb933069),
	.w8(32'h3b19d9d0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fa976),
	.w1(32'h3b0e3d9c),
	.w2(32'hbb249fa7),
	.w3(32'hbbd94ea7),
	.w4(32'hba3fba2f),
	.w5(32'h3aad9f51),
	.w6(32'h3645398d),
	.w7(32'h3a52cd89),
	.w8(32'h3a9a14d0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c7ed2),
	.w1(32'h3939fad0),
	.w2(32'hba560810),
	.w3(32'hbb01bc4f),
	.w4(32'hbb0746eb),
	.w5(32'h3b13cc09),
	.w6(32'hbb48ab99),
	.w7(32'hba800ad9),
	.w8(32'h3a93c596),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37e777),
	.w1(32'h3aa2660d),
	.w2(32'h39f4267d),
	.w3(32'h3aba91c9),
	.w4(32'h3a9a4ecb),
	.w5(32'h38a1e6a1),
	.w6(32'h3aa67d54),
	.w7(32'h3b4319da),
	.w8(32'h3b0d69f8),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c0626),
	.w1(32'hbb93a25c),
	.w2(32'hbad98c4b),
	.w3(32'h3afa8df1),
	.w4(32'hbbd51348),
	.w5(32'hbb892111),
	.w6(32'h3aeb66ba),
	.w7(32'h39da2deb),
	.w8(32'hba9194e8),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24df74),
	.w1(32'h3b9503bd),
	.w2(32'h390b38c3),
	.w3(32'hbb30dfe7),
	.w4(32'h398d7cb5),
	.w5(32'h3a6ef2e4),
	.w6(32'h3b2c768b),
	.w7(32'h3b648a26),
	.w8(32'h3a3c8011),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0084ef),
	.w1(32'h3b2f1c0e),
	.w2(32'hbba2cf5f),
	.w3(32'h3b809335),
	.w4(32'h3a9e7ada),
	.w5(32'h3a00efb6),
	.w6(32'hba08fc1d),
	.w7(32'hbad0d62b),
	.w8(32'h3ac04bf7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d71c3),
	.w1(32'hb9abbf06),
	.w2(32'hbbed417e),
	.w3(32'h3ab166e9),
	.w4(32'hbb9c8279),
	.w5(32'h3b5a7b40),
	.w6(32'hbb96038f),
	.w7(32'h3c396408),
	.w8(32'h3bd0872c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99fb6a),
	.w1(32'h3bc3b07d),
	.w2(32'h3abd13ca),
	.w3(32'h39121682),
	.w4(32'hbaf99d49),
	.w5(32'hbb3f573b),
	.w6(32'h3b8d803f),
	.w7(32'hbb1fadbd),
	.w8(32'hbad2c15b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22dc1f),
	.w1(32'hbb09ed7d),
	.w2(32'h3aaa9457),
	.w3(32'hbb19539b),
	.w4(32'hbaf2ed2b),
	.w5(32'hbbddd1c2),
	.w6(32'h39a9c397),
	.w7(32'hbb9eb187),
	.w8(32'h3aa80ea0),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99801d),
	.w1(32'h3b42de49),
	.w2(32'h3c3a5433),
	.w3(32'h3aa43159),
	.w4(32'h3bd15259),
	.w5(32'h3b114a2d),
	.w6(32'hbb1b881c),
	.w7(32'h3c37837e),
	.w8(32'h3b5dde52),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43b1a),
	.w1(32'hbb13dd0e),
	.w2(32'hbb381d0f),
	.w3(32'hbb530fc2),
	.w4(32'hbb65fe83),
	.w5(32'hbb7ebb39),
	.w6(32'hba91a661),
	.w7(32'hbba7bf5e),
	.w8(32'hb9d07fe2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc60d1a),
	.w1(32'hbb4aed37),
	.w2(32'hb96b6991),
	.w3(32'hbb094b59),
	.w4(32'hbb623a32),
	.w5(32'h3bb94576),
	.w6(32'hba65308d),
	.w7(32'h3aa85292),
	.w8(32'hba0b86c2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50c8ac),
	.w1(32'hb9aee054),
	.w2(32'h3aa28f80),
	.w3(32'hba311060),
	.w4(32'hbb3a9c36),
	.w5(32'h39a72ffd),
	.w6(32'hba1b622e),
	.w7(32'hbb6985f7),
	.w8(32'h3baaaf8e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2cceb),
	.w1(32'hba23c062),
	.w2(32'h3b3278bb),
	.w3(32'h39e5958a),
	.w4(32'hbba0eaf8),
	.w5(32'hbbd6b88e),
	.w6(32'hba8a0514),
	.w7(32'hbb3ce04f),
	.w8(32'hbaacd84a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc121027),
	.w1(32'h3a25ef46),
	.w2(32'h3c0d5104),
	.w3(32'hbc03f9a2),
	.w4(32'hbb8d74cb),
	.w5(32'hbb309114),
	.w6(32'hbc09d5df),
	.w7(32'h3abab010),
	.w8(32'h3b0a3d26),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be15f),
	.w1(32'hba4594c8),
	.w2(32'hbb1aa5a3),
	.w3(32'h3b547504),
	.w4(32'hbb620a89),
	.w5(32'hbb6c77f5),
	.w6(32'h3b2f2abd),
	.w7(32'h3a088b55),
	.w8(32'h3b9b23b1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b3ade),
	.w1(32'h3ba51272),
	.w2(32'h3c123496),
	.w3(32'h3ad620ce),
	.w4(32'h3bb31895),
	.w5(32'h3bf4790d),
	.w6(32'h3bb2de0f),
	.w7(32'h3b565699),
	.w8(32'h3b953c17),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e630f),
	.w1(32'hbbb1160b),
	.w2(32'hbb52290f),
	.w3(32'h3be8eb8c),
	.w4(32'hbb7e974e),
	.w5(32'hbb4e9a93),
	.w6(32'hb9ea703f),
	.w7(32'h39332bb0),
	.w8(32'h3a8e82c4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7c869),
	.w1(32'h3b1131ac),
	.w2(32'h3700c08b),
	.w3(32'h3b134c6f),
	.w4(32'h3a2fc733),
	.w5(32'h3929c91a),
	.w6(32'hbb6baee7),
	.w7(32'h3aeef49c),
	.w8(32'h3b67031b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b766e7d),
	.w1(32'h3a9d88e4),
	.w2(32'hbb657750),
	.w3(32'h3b1a2e62),
	.w4(32'hbb7467e8),
	.w5(32'hbaf88d48),
	.w6(32'h3b3360d1),
	.w7(32'hbc01e64f),
	.w8(32'hb9984bb7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23acee),
	.w1(32'h3b95a928),
	.w2(32'h38d39d6a),
	.w3(32'hb8dc15d3),
	.w4(32'hbb1e9c9e),
	.w5(32'hbad999ea),
	.w6(32'hb963f4db),
	.w7(32'hbb02e327),
	.w8(32'hbb90a60e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc446239),
	.w1(32'hbbabbd92),
	.w2(32'hbae55c7d),
	.w3(32'hbb7fd328),
	.w4(32'hbb6f16ba),
	.w5(32'hbb6f302e),
	.w6(32'hbc22098c),
	.w7(32'hbb02cd40),
	.w8(32'hba078bcf),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe8841),
	.w1(32'hba101d47),
	.w2(32'hbaf28082),
	.w3(32'hba80d52f),
	.w4(32'hbb4fae92),
	.w5(32'hbb6ba302),
	.w6(32'h3865d3f7),
	.w7(32'hbb8c093e),
	.w8(32'h38892414),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b533d),
	.w1(32'h3a3c4d7e),
	.w2(32'h3baaee57),
	.w3(32'hbb7d3ab3),
	.w4(32'h3a868e84),
	.w5(32'h3a98185b),
	.w6(32'h39cee0e8),
	.w7(32'h3bcecce6),
	.w8(32'h3b1b71bb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule