module layer_10_featuremap_425(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3bf30),
	.w1(32'hb9289b27),
	.w2(32'hb94001b8),
	.w3(32'h39228226),
	.w4(32'hba2467a3),
	.w5(32'hb9d6299c),
	.w6(32'hb8b299ea),
	.w7(32'hb9966d84),
	.w8(32'hb91688cd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6a971),
	.w1(32'hb9a52ec1),
	.w2(32'hb964cbd5),
	.w3(32'hba414a44),
	.w4(32'hb95f4c78),
	.w5(32'hba03a35f),
	.w6(32'hb8df3101),
	.w7(32'h385989c6),
	.w8(32'hb8336b33),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba264cec),
	.w1(32'hbaa60f5a),
	.w2(32'hb970edcd),
	.w3(32'hb9a848f5),
	.w4(32'hbac0afa1),
	.w5(32'hba8c7b26),
	.w6(32'hba007adf),
	.w7(32'hba4824f0),
	.w8(32'hba4d7771),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9872f9b),
	.w1(32'h3a962ca9),
	.w2(32'h3a5878a7),
	.w3(32'hb8cbca1b),
	.w4(32'h3a7d3cc5),
	.w5(32'h3a7c99f2),
	.w6(32'hb90cb4a5),
	.w7(32'h39a8ec00),
	.w8(32'h39024067),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b312e),
	.w1(32'hb92c6c71),
	.w2(32'hb9807eda),
	.w3(32'h3a013c81),
	.w4(32'hb989d3d0),
	.w5(32'hb97dc949),
	.w6(32'h391057f7),
	.w7(32'hb816e04c),
	.w8(32'hb9b26095),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfecaa),
	.w1(32'hba6da862),
	.w2(32'hba7228f3),
	.w3(32'h39fc46bb),
	.w4(32'hba7a78ed),
	.w5(32'hba24e40b),
	.w6(32'hb822192e),
	.w7(32'hba2232d8),
	.w8(32'hb9e4c175),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba844460),
	.w1(32'hb9aa0142),
	.w2(32'h38edcbd8),
	.w3(32'hbaa9163e),
	.w4(32'h39f139a6),
	.w5(32'h3898e658),
	.w6(32'hba90ed57),
	.w7(32'h3a22c347),
	.w8(32'h3ab30d94),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39078235),
	.w1(32'h3a679579),
	.w2(32'hb9d94c35),
	.w3(32'h3a8aef83),
	.w4(32'h3a86d737),
	.w5(32'h3a32916d),
	.w6(32'h3a8b5e66),
	.w7(32'h3ad33804),
	.w8(32'h3979ab9f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98120f4),
	.w1(32'hba9ec1e6),
	.w2(32'hba120d98),
	.w3(32'h3a0655ec),
	.w4(32'hba07f7a6),
	.w5(32'hba2b3d2a),
	.w6(32'h3a64a4c3),
	.w7(32'hb9004fc8),
	.w8(32'hba6386e4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39924b62),
	.w1(32'h3ab6fc89),
	.w2(32'h3b0d43ae),
	.w3(32'h3ab2a9fb),
	.w4(32'h3b03ee3e),
	.w5(32'h3af5f2c4),
	.w6(32'hb98c22d1),
	.w7(32'h3ab5244c),
	.w8(32'h3b114d0b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91827e),
	.w1(32'h39772b64),
	.w2(32'h39debd3d),
	.w3(32'hba9408b7),
	.w4(32'hb9af1824),
	.w5(32'hba484fdc),
	.w6(32'hba798756),
	.w7(32'hb9aad8d0),
	.w8(32'h36448d62),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fd30e),
	.w1(32'hb914c80d),
	.w2(32'h3a0460e8),
	.w3(32'h3a10ac6b),
	.w4(32'hba9a6037),
	.w5(32'h39df4146),
	.w6(32'h390ed2f1),
	.w7(32'hbae2cd6f),
	.w8(32'hba37faff),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e546b),
	.w1(32'h39a32741),
	.w2(32'hba20dd67),
	.w3(32'hba2d25f1),
	.w4(32'h3a796106),
	.w5(32'hb7a1c4b8),
	.w6(32'hba897741),
	.w7(32'h39aa839b),
	.w8(32'hb988e097),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba841d2f),
	.w1(32'h391cea7e),
	.w2(32'h3aa73040),
	.w3(32'hba2ba3fe),
	.w4(32'hb96b246a),
	.w5(32'hb94c4073),
	.w6(32'hba32e976),
	.w7(32'hb9ee3ae4),
	.w8(32'hb901d443),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad588c6),
	.w1(32'h3869c505),
	.w2(32'h36e37ae0),
	.w3(32'h3af25da3),
	.w4(32'h3ac30a4d),
	.w5(32'h391361de),
	.w6(32'h392a4185),
	.w7(32'h3a5c4d4c),
	.w8(32'h3a638988),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d4419),
	.w1(32'h3b07e0ae),
	.w2(32'h3af71ae2),
	.w3(32'h3ade5666),
	.w4(32'h3b0b5f2b),
	.w5(32'h3ab68360),
	.w6(32'h3a50a426),
	.w7(32'h3ad93669),
	.w8(32'h3a949c09),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a3ee3),
	.w1(32'hb919e3ab),
	.w2(32'h38d8737f),
	.w3(32'h38895b5c),
	.w4(32'hbadbb3c7),
	.w5(32'hbaaf9dc5),
	.w6(32'hb96ee58f),
	.w7(32'hbae4f16b),
	.w8(32'hbaf328da),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37dc6b),
	.w1(32'h3af2b453),
	.w2(32'h3a9024d5),
	.w3(32'hbaa48566),
	.w4(32'h3a543f77),
	.w5(32'h3a0b0886),
	.w6(32'hbad8196c),
	.w7(32'h3a11b08d),
	.w8(32'h3926edb9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0faf06),
	.w1(32'h3aa94323),
	.w2(32'h3aaf4b1e),
	.w3(32'h3adfcbdd),
	.w4(32'h3ab50f5b),
	.w5(32'h3a277aaa),
	.w6(32'h3adb98bd),
	.w7(32'h3a41d69b),
	.w8(32'h3a07517b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375f9242),
	.w1(32'hb9c685af),
	.w2(32'hba6b3197),
	.w3(32'h39985eff),
	.w4(32'hb9aca86a),
	.w5(32'h397ae455),
	.w6(32'h395b2500),
	.w7(32'hb8ac03ba),
	.w8(32'h3939a1fb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d59fe),
	.w1(32'hba3ac1be),
	.w2(32'hba4180b6),
	.w3(32'hb951a103),
	.w4(32'hba16b3f0),
	.w5(32'hb9dedcff),
	.w6(32'h3929c81c),
	.w7(32'h3984ad36),
	.w8(32'h38b33bbc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a784ec3),
	.w1(32'h3a67f5f2),
	.w2(32'h3a5cdbb8),
	.w3(32'h39188ff3),
	.w4(32'h3a4d1223),
	.w5(32'h3a6c48e5),
	.w6(32'h39c64f7b),
	.w7(32'h3a476745),
	.w8(32'h39f2a97f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28a98f),
	.w1(32'hba88f2c6),
	.w2(32'h3adc5bc1),
	.w3(32'h3b2730be),
	.w4(32'h3a8cc97f),
	.w5(32'h3ac40872),
	.w6(32'h3ad8a2b9),
	.w7(32'h3a17eb7d),
	.w8(32'h3ad0894c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395be15f),
	.w1(32'h3a8a5e16),
	.w2(32'h3ab0200d),
	.w3(32'h3a7775e8),
	.w4(32'h3a5ed86a),
	.w5(32'h3a749c3e),
	.w6(32'hba07547e),
	.w7(32'hb90aa08e),
	.w8(32'h3a00241b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab413d3),
	.w1(32'hba51f806),
	.w2(32'h3a95dfe0),
	.w3(32'hba8f6120),
	.w4(32'hb92cb7ca),
	.w5(32'h3a2ddfa3),
	.w6(32'hba214ab5),
	.w7(32'hb9acc98a),
	.w8(32'h3a79fbc6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a809338),
	.w1(32'hbaa3b087),
	.w2(32'hbaa022f2),
	.w3(32'h3a2eeaa5),
	.w4(32'hba99398a),
	.w5(32'hb98c393f),
	.w6(32'h3a06dd48),
	.w7(32'hba87d6be),
	.w8(32'hb95e326e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015271),
	.w1(32'h399b0b65),
	.w2(32'h3a79f0e0),
	.w3(32'hbad569ac),
	.w4(32'h3a66a78e),
	.w5(32'h39939504),
	.w6(32'hbac6702a),
	.w7(32'h3a01d7d4),
	.w8(32'h3a127565),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389453f5),
	.w1(32'h392fb34e),
	.w2(32'h39955c1c),
	.w3(32'h391773e4),
	.w4(32'h39f83266),
	.w5(32'hb9832e9a),
	.w6(32'h3692b8af),
	.w7(32'h3a183e8e),
	.w8(32'h397940bb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a3398),
	.w1(32'h3a0db4ed),
	.w2(32'h3a98e670),
	.w3(32'hba187e66),
	.w4(32'hbaa464c6),
	.w5(32'hb9802206),
	.w6(32'hb93f3613),
	.w7(32'hba5c4967),
	.w8(32'hb8f9b225),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c3e73),
	.w1(32'h3ada9a73),
	.w2(32'h3ab4e7b9),
	.w3(32'h3ab1c56d),
	.w4(32'h3b073989),
	.w5(32'h3ae02672),
	.w6(32'h3a79c839),
	.w7(32'h3b0b2c43),
	.w8(32'h3ae7898d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22e2a0),
	.w1(32'h3abeb867),
	.w2(32'h3aa9c17d),
	.w3(32'h398525a4),
	.w4(32'h3a8f15ef),
	.w5(32'h3a84a3dd),
	.w6(32'h39c5a8f1),
	.w7(32'h3a31f3c7),
	.w8(32'h3ac9da86),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a629d0b),
	.w1(32'h39b8ecd5),
	.w2(32'h39848f16),
	.w3(32'h3960b45b),
	.w4(32'h390921ce),
	.w5(32'hb9201138),
	.w6(32'h3aa7912e),
	.w7(32'h39d6acd5),
	.w8(32'h3974685c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb2044),
	.w1(32'h39d1602e),
	.w2(32'h3a411803),
	.w3(32'h3a8b5a9d),
	.w4(32'h38aa6ac9),
	.w5(32'hba0d4f2a),
	.w6(32'h3a0ea268),
	.w7(32'h398b97dd),
	.w8(32'hb934d809),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f0a41),
	.w1(32'hb9f75b2c),
	.w2(32'hb900ce80),
	.w3(32'h3892f211),
	.w4(32'h39c1e718),
	.w5(32'h3889ccac),
	.w6(32'hba3dae59),
	.w7(32'h39b76ccc),
	.w8(32'h39473170),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6714),
	.w1(32'h3a381720),
	.w2(32'h3a19bbd6),
	.w3(32'hbaab603d),
	.w4(32'h3a3a46c9),
	.w5(32'h3a272200),
	.w6(32'hba98d391),
	.w7(32'h3a6dae95),
	.w8(32'h3989798e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d9fbe),
	.w1(32'h3a9d1856),
	.w2(32'h3a9165f3),
	.w3(32'h3a440f7a),
	.w4(32'h3a7377e2),
	.w5(32'h3a6cc3de),
	.w6(32'h39922a16),
	.w7(32'h3a7da1f0),
	.w8(32'h39a9c3ec),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b3b32),
	.w1(32'h3ae268f1),
	.w2(32'h3b132b51),
	.w3(32'h3a730196),
	.w4(32'h3a5c43e2),
	.w5(32'h3a560c68),
	.w6(32'h3a1012d4),
	.w7(32'h3a65e4b9),
	.w8(32'h3b034598),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3f064),
	.w1(32'hbaeb54b7),
	.w2(32'h391c7590),
	.w3(32'hbb041aff),
	.w4(32'hbb2fe08f),
	.w5(32'hba7e53b4),
	.w6(32'hb9b42892),
	.w7(32'hb9d3e119),
	.w8(32'h39aecbf8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04022f),
	.w1(32'hbae8861d),
	.w2(32'h3a4a5f0d),
	.w3(32'hbb06d026),
	.w4(32'hbb30029d),
	.w5(32'hb996e408),
	.w6(32'hba9c3f66),
	.w7(32'hbb1e595a),
	.w8(32'hb9e70535),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eefd36),
	.w1(32'h380c668d),
	.w2(32'hb9ad49c5),
	.w3(32'hba07fc87),
	.w4(32'hb6c905dd),
	.w5(32'hb9788073),
	.w6(32'hb9fc8a90),
	.w7(32'h396f055d),
	.w8(32'h38c21848),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0002a),
	.w1(32'hba3a751c),
	.w2(32'hba8ab5d9),
	.w3(32'hb990174e),
	.w4(32'hb8907403),
	.w5(32'hb88cc6db),
	.w6(32'hb9d9c3d4),
	.w7(32'hba8e4f70),
	.w8(32'hba8049aa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b7786),
	.w1(32'h3901c4a2),
	.w2(32'hb93a0931),
	.w3(32'hba20c692),
	.w4(32'h39ff0562),
	.w5(32'hb6a15df7),
	.w6(32'hbaa51169),
	.w7(32'h3947bce2),
	.w8(32'h398dba1d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fc6658),
	.w1(32'h39371081),
	.w2(32'h3a490373),
	.w3(32'h3a060203),
	.w4(32'hb9be90b3),
	.w5(32'h3a35fd65),
	.w6(32'h3a0e4850),
	.w7(32'hba1cda14),
	.w8(32'hb96a8f31),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1150be),
	.w1(32'h3a40fe1a),
	.w2(32'h3a2bb804),
	.w3(32'h3abdd0f8),
	.w4(32'h3add116f),
	.w5(32'h3a6c86fd),
	.w6(32'h39a8b18a),
	.w7(32'h3a4f8dd0),
	.w8(32'h3a8a3610),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d6bc8),
	.w1(32'h3a945a56),
	.w2(32'h3aaefa64),
	.w3(32'h3a1405c3),
	.w4(32'h3b007bac),
	.w5(32'h3adb2246),
	.w6(32'hb9fa4c89),
	.w7(32'h3ad9a128),
	.w8(32'h3b059880),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b380e9),
	.w1(32'h3a925c92),
	.w2(32'h3b0ae89b),
	.w3(32'h3ab80f0a),
	.w4(32'h3b25a8e3),
	.w5(32'h3b2b441a),
	.w6(32'h39a82406),
	.w7(32'h3ae615d3),
	.w8(32'h3b0b32b1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1fbca),
	.w1(32'h3b1f2bd1),
	.w2(32'h3ae33f5c),
	.w3(32'h3a9e7504),
	.w4(32'h3b148bf5),
	.w5(32'h3a6487bd),
	.w6(32'h3a40b276),
	.w7(32'h3b01226e),
	.w8(32'h3abc7928),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9999257),
	.w1(32'hba3490de),
	.w2(32'hbabcda97),
	.w3(32'h39466a8c),
	.w4(32'h39dc3527),
	.w5(32'h3891b76f),
	.w6(32'hba4cb322),
	.w7(32'hba1cb521),
	.w8(32'hba6b3d8f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997cac5),
	.w1(32'h3a44a2d9),
	.w2(32'h3a8c9428),
	.w3(32'hba0e1497),
	.w4(32'h3aa0bb55),
	.w5(32'h3a6f4a0e),
	.w6(32'hb99504a6),
	.w7(32'h3ab36c33),
	.w8(32'h3a603c20),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b017e8f),
	.w1(32'h3b1bf4c4),
	.w2(32'h3b273295),
	.w3(32'h3acd3064),
	.w4(32'h3b1ed648),
	.w5(32'h3ae45749),
	.w6(32'h3a9b641a),
	.w7(32'h3b3ba38d),
	.w8(32'h3ad90a53),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa131e8),
	.w1(32'hb95a4ef1),
	.w2(32'h3a0e5701),
	.w3(32'h38cf94bc),
	.w4(32'hb89d2660),
	.w5(32'h3a681fb4),
	.w6(32'h3a9919e3),
	.w7(32'hb9a82cd6),
	.w8(32'h39c59651),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be857e),
	.w1(32'hb8d1db9a),
	.w2(32'hb992bb00),
	.w3(32'hb965a4b1),
	.w4(32'hba23dce0),
	.w5(32'hba21e423),
	.w6(32'h38933258),
	.w7(32'hba250b11),
	.w8(32'hba08f7fb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab568cd),
	.w1(32'h398b2d9c),
	.w2(32'h3a1c60cc),
	.w3(32'hba839bf5),
	.w4(32'h3a736fe9),
	.w5(32'h3a46c943),
	.w6(32'hba37cd4f),
	.w7(32'h3ab3c2fb),
	.w8(32'h3a24887d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9454854),
	.w1(32'hb9064d22),
	.w2(32'hb970a877),
	.w3(32'h3a5fca3d),
	.w4(32'h3a8a084f),
	.w5(32'h39f21a82),
	.w6(32'h3a01896a),
	.w7(32'h3a8020e3),
	.w8(32'hb9a829e9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38640f16),
	.w1(32'h3a807b05),
	.w2(32'h39370f75),
	.w3(32'hb8a0036a),
	.w4(32'h3a843ba5),
	.w5(32'h391b8fbe),
	.w6(32'hb8a350b9),
	.w7(32'h3a701f31),
	.w8(32'h39a5f64f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02be99),
	.w1(32'hba167b8e),
	.w2(32'hb9a73017),
	.w3(32'h3a103170),
	.w4(32'hb98876a0),
	.w5(32'hba242a75),
	.w6(32'h39c7e323),
	.w7(32'hb90bf41f),
	.w8(32'h3940df00),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ab86a),
	.w1(32'hba473c36),
	.w2(32'hba40f4a4),
	.w3(32'hb9aae0d7),
	.w4(32'hba0f0918),
	.w5(32'h38df4c4b),
	.w6(32'hb921a699),
	.w7(32'hba1f50b6),
	.w8(32'h3468cb62),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19c603),
	.w1(32'hbab22781),
	.w2(32'hba8797fa),
	.w3(32'hb988bb72),
	.w4(32'hbab9ab40),
	.w5(32'hba8c568f),
	.w6(32'hb97de16e),
	.w7(32'hbaa98e06),
	.w8(32'hbad5cd90),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a1956),
	.w1(32'hb9ffcdd0),
	.w2(32'hba07c801),
	.w3(32'hb924e168),
	.w4(32'hba142b45),
	.w5(32'h3831f4aa),
	.w6(32'hbaa448de),
	.w7(32'hba1ef4e3),
	.w8(32'hba35beb0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e7fe2),
	.w1(32'hba238a53),
	.w2(32'hb90648ab),
	.w3(32'hba889442),
	.w4(32'hba5f3160),
	.w5(32'hb9f56b9a),
	.w6(32'hba90cff1),
	.w7(32'hbaa29836),
	.w8(32'hbaa58487),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c28bb7),
	.w1(32'hb98da964),
	.w2(32'hb982b768),
	.w3(32'h3a1a3413),
	.w4(32'hba1a0b55),
	.w5(32'hb9d75202),
	.w6(32'hb9a001e6),
	.w7(32'hba14fa67),
	.w8(32'h39904dc3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84bff7),
	.w1(32'h387c25c6),
	.w2(32'h38b49edb),
	.w3(32'hba56bc55),
	.w4(32'h39e9916f),
	.w5(32'hb909a9eb),
	.w6(32'hba1d9ee0),
	.w7(32'h39e5f290),
	.w8(32'h3a04fe27),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4f586),
	.w1(32'hb4ed70dc),
	.w2(32'h394d703f),
	.w3(32'h39eb0235),
	.w4(32'hb990da51),
	.w5(32'hb7f10a17),
	.w6(32'h39db3ebc),
	.w7(32'hb9ca1536),
	.w8(32'hb8d0746b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36b0df),
	.w1(32'hba6d95cf),
	.w2(32'hba432ff0),
	.w3(32'h3a83d819),
	.w4(32'hba923ead),
	.w5(32'hba5203f0),
	.w6(32'h3a5a9f4e),
	.w7(32'hbabc0d85),
	.w8(32'hbad79ca5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65acbb),
	.w1(32'h3a9c8d52),
	.w2(32'h3a735452),
	.w3(32'hbaa6f0f1),
	.w4(32'h3a3a8a5f),
	.w5(32'h3a31f573),
	.w6(32'hbaa62680),
	.w7(32'h3a41a520),
	.w8(32'h3a075384),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dc2f0),
	.w1(32'h39ceefd8),
	.w2(32'h3a10c341),
	.w3(32'h39e4c2f6),
	.w4(32'h3a0a7681),
	.w5(32'h39b5b3b3),
	.w6(32'h39f5224c),
	.w7(32'h3a74f93a),
	.w8(32'h3a75f4fe),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7557b8),
	.w1(32'hbabd1e10),
	.w2(32'hbb021003),
	.w3(32'h3a8037d3),
	.w4(32'hbaa48c9e),
	.w5(32'hbadb7948),
	.w6(32'h3a92ac3d),
	.w7(32'hbaa17e39),
	.w8(32'hbae21183),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadb386),
	.w1(32'hba00007c),
	.w2(32'h39a8c00f),
	.w3(32'hba175e6a),
	.w4(32'h39b2c91e),
	.w5(32'h38e3d7c0),
	.w6(32'hbaa0dca3),
	.w7(32'hb794ca26),
	.w8(32'h3a184510),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba829b40),
	.w1(32'hba431278),
	.w2(32'h395bb936),
	.w3(32'hbaa05c57),
	.w4(32'hb9d80adf),
	.w5(32'h3a169aac),
	.w6(32'hba99d9da),
	.w7(32'hb9cdd052),
	.w8(32'hb9c57f02),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89a73b),
	.w1(32'h39f69314),
	.w2(32'h38964d3c),
	.w3(32'h39d73227),
	.w4(32'hba2277ac),
	.w5(32'h3ac9a637),
	.w6(32'h3987de26),
	.w7(32'hba9dfdff),
	.w8(32'h3b2f4d53),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba894bfb),
	.w1(32'hbaf9a050),
	.w2(32'hbaae70dc),
	.w3(32'hbaf8b98a),
	.w4(32'hbaaf07a5),
	.w5(32'hbaf7bf4c),
	.w6(32'hba7d7687),
	.w7(32'hbb34d811),
	.w8(32'hbb11d745),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68d7a2),
	.w1(32'hbb104380),
	.w2(32'hba517d4f),
	.w3(32'hbb97249a),
	.w4(32'hba7e542f),
	.w5(32'h3ab668e7),
	.w6(32'hbb8f1110),
	.w7(32'h3b95c864),
	.w8(32'h3b8ca95b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7fa95),
	.w1(32'h3b307ead),
	.w2(32'h3a8b6f35),
	.w3(32'hbafcc2d0),
	.w4(32'h3af96899),
	.w5(32'h37db324d),
	.w6(32'h3abac465),
	.w7(32'hb7a23198),
	.w8(32'h3896f2e1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6412df),
	.w1(32'hba86b9a5),
	.w2(32'h398ba55f),
	.w3(32'h3ba7b581),
	.w4(32'hb992272c),
	.w5(32'hb927aaf4),
	.w6(32'h3b94814a),
	.w7(32'hba1d74c4),
	.w8(32'hbaf3b8fd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e40141),
	.w1(32'hbaa94cab),
	.w2(32'h3b52b88a),
	.w3(32'h3a8a1b65),
	.w4(32'hbb44b33f),
	.w5(32'hbbaf6cd2),
	.w6(32'hbb95bac5),
	.w7(32'hb9612244),
	.w8(32'hba40d156),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa45c1d),
	.w1(32'hba93a74c),
	.w2(32'hba9e0d00),
	.w3(32'hbb6f76d3),
	.w4(32'h3b03a18e),
	.w5(32'h3b066fdf),
	.w6(32'hb94c14f1),
	.w7(32'hba3a7096),
	.w8(32'hb81d50fd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af853f6),
	.w1(32'h3b15f39d),
	.w2(32'hbb42ce78),
	.w3(32'h3b502491),
	.w4(32'hbb25acbd),
	.w5(32'hbba62a21),
	.w6(32'hb9e65a6f),
	.w7(32'hbb70139c),
	.w8(32'hbb99c5ca),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85f512),
	.w1(32'hbb4d5ebf),
	.w2(32'hbb528cd7),
	.w3(32'hbaff64fc),
	.w4(32'hbb015079),
	.w5(32'hbb459429),
	.w6(32'hbb4902cf),
	.w7(32'hba9c352a),
	.w8(32'hba59d9d1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3c6dd),
	.w1(32'h3ad658e2),
	.w2(32'h3a0e14cf),
	.w3(32'hbbc2ef49),
	.w4(32'h3a944d82),
	.w5(32'h3a95abe4),
	.w6(32'hbb340c37),
	.w7(32'h3b11b0b7),
	.w8(32'h3ad74f6b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4f4aa),
	.w1(32'hbb10c47f),
	.w2(32'hb9af446f),
	.w3(32'hbb1a7550),
	.w4(32'hbb5f5984),
	.w5(32'hbae249c8),
	.w6(32'hbae03ab0),
	.w7(32'hbb4b8545),
	.w8(32'h3809d665),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9919e69),
	.w1(32'h3be5ca85),
	.w2(32'h3c238d5c),
	.w3(32'hba6680a8),
	.w4(32'h3bfd74d4),
	.w5(32'h3be52ce5),
	.w6(32'h3a084d12),
	.w7(32'h3bdffb98),
	.w8(32'h3bcd4ed5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074dc5),
	.w1(32'h3a6b08f0),
	.w2(32'hb96750a9),
	.w3(32'h3bd21e9d),
	.w4(32'hba75cd82),
	.w5(32'h39cd90c9),
	.w6(32'h3bc34a9d),
	.w7(32'hb9f3df18),
	.w8(32'h3a086d55),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2369d0),
	.w1(32'h3b35b8b3),
	.w2(32'h3b23aad8),
	.w3(32'h3a393c84),
	.w4(32'h3ab1d24e),
	.w5(32'h3b13ca91),
	.w6(32'h3b0dbfb1),
	.w7(32'h3ad14edf),
	.w8(32'h3a691d6e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd62db),
	.w1(32'hb99dcaaa),
	.w2(32'hbb27f846),
	.w3(32'h3b5077f0),
	.w4(32'hbac958bb),
	.w5(32'hbb568c95),
	.w6(32'h3b9d848c),
	.w7(32'hbb31e178),
	.w8(32'hba815233),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25783c),
	.w1(32'hbb91e26e),
	.w2(32'hbb714c34),
	.w3(32'hbb7ed071),
	.w4(32'hbb9b0aa1),
	.w5(32'hbb196ec7),
	.w6(32'hba56d030),
	.w7(32'hbb38761e),
	.w8(32'h39a79046),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d0c4f4),
	.w1(32'hbb22962a),
	.w2(32'hbaf08151),
	.w3(32'hb9e2c745),
	.w4(32'hba36a4b7),
	.w5(32'hba7958c5),
	.w6(32'h3a7df909),
	.w7(32'h3a347d45),
	.w8(32'hbbd22e74),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62e603),
	.w1(32'hbae55c47),
	.w2(32'hbb077d9c),
	.w3(32'hbb71ce6f),
	.w4(32'hbaf06d25),
	.w5(32'hbb216bec),
	.w6(32'hbbbc8b6d),
	.w7(32'h3a0df212),
	.w8(32'h3ac29b8f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ca219),
	.w1(32'hbb25950c),
	.w2(32'hbb9ff799),
	.w3(32'hbb5c95d9),
	.w4(32'hbb13a537),
	.w5(32'hbbf2e9b5),
	.w6(32'hba6da06c),
	.w7(32'hba2175ce),
	.w8(32'hbaa88eab),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb968f),
	.w1(32'hbb046758),
	.w2(32'hbad55786),
	.w3(32'hbb3fe341),
	.w4(32'hb85916b5),
	.w5(32'h391eb2be),
	.w6(32'hba5e7a51),
	.w7(32'hbb8920bb),
	.w8(32'hbb5b231b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf86ee8),
	.w1(32'h3a650b08),
	.w2(32'h39163cec),
	.w3(32'h393d913f),
	.w4(32'h3b00d17d),
	.w5(32'h3b346ad0),
	.w6(32'hb9ba90ab),
	.w7(32'h37d40873),
	.w8(32'h3a68e060),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2031a),
	.w1(32'hbb5e565a),
	.w2(32'hba83ae71),
	.w3(32'hbb1bcf16),
	.w4(32'hbb9cdb41),
	.w5(32'h3a3d8f84),
	.w6(32'hba331a35),
	.w7(32'hbb5e3993),
	.w8(32'h3aaa1992),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ca1de),
	.w1(32'hbb689e1a),
	.w2(32'hbb9c069e),
	.w3(32'hb984f4fc),
	.w4(32'hbad7cb3e),
	.w5(32'hbb6ba784),
	.w6(32'h3a80fb73),
	.w7(32'hba6ac259),
	.w8(32'hba615dd4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34daa2),
	.w1(32'h3b3a0f44),
	.w2(32'h3b12cffc),
	.w3(32'hba1c5025),
	.w4(32'h3a9bda52),
	.w5(32'hb9dd59f5),
	.w6(32'hbb29d669),
	.w7(32'h3b67bf64),
	.w8(32'h3b3a39f2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b86c1),
	.w1(32'h3981a435),
	.w2(32'h39d140df),
	.w3(32'h3ab3909d),
	.w4(32'h3aebb7ae),
	.w5(32'h3b5c8ab1),
	.w6(32'h3b417ed4),
	.w7(32'h3b646551),
	.w8(32'h3b4c70cb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab97a00),
	.w1(32'hba354eff),
	.w2(32'h3a97378f),
	.w3(32'h3a2f1d3e),
	.w4(32'h3a2be4e4),
	.w5(32'h3b1d39c2),
	.w6(32'hb99176df),
	.w7(32'hbb512a58),
	.w8(32'hba1da2ab),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab89dbf),
	.w1(32'hbb7f904b),
	.w2(32'hbbae7272),
	.w3(32'h3ac0851f),
	.w4(32'hbaf57c30),
	.w5(32'hba368ffb),
	.w6(32'hbadab935),
	.w7(32'hbacfec66),
	.w8(32'hba2143a8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f1ef4),
	.w1(32'hbb57749c),
	.w2(32'hbb100c24),
	.w3(32'hb8ea78cb),
	.w4(32'hbb54dcba),
	.w5(32'h3a08f7e7),
	.w6(32'hba358985),
	.w7(32'hba37e09f),
	.w8(32'h37ad27aa),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3222f2),
	.w1(32'h3ba4bde3),
	.w2(32'h3bf12732),
	.w3(32'h38405006),
	.w4(32'h3bfa1b08),
	.w5(32'h3c09992a),
	.w6(32'hbadddb43),
	.w7(32'h3c32d597),
	.w8(32'h3bfa943b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7f04d),
	.w1(32'h394ec404),
	.w2(32'hbaef987c),
	.w3(32'h3b72a71f),
	.w4(32'hb9366de4),
	.w5(32'h38d513e7),
	.w6(32'h3b135d57),
	.w7(32'h3b376a1f),
	.w8(32'h3b0267d5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4ba89),
	.w1(32'hba9bdadf),
	.w2(32'hbb5c983e),
	.w3(32'hbab52a55),
	.w4(32'h3ac782b8),
	.w5(32'h3aad9261),
	.w6(32'h3b0d227b),
	.w7(32'hbb824e3d),
	.w8(32'hbb06ac43),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54c009),
	.w1(32'hbbca1bc7),
	.w2(32'hbb1a38f3),
	.w3(32'hbb11da38),
	.w4(32'h3a8f8942),
	.w5(32'h3ae5f586),
	.w6(32'hbb8f7516),
	.w7(32'h3ace97c8),
	.w8(32'hbaa964f7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3a7b9),
	.w1(32'hbb00b366),
	.w2(32'hba9bbc96),
	.w3(32'h3b8c989e),
	.w4(32'h3a9ed366),
	.w5(32'h3b267a49),
	.w6(32'hb790e51a),
	.w7(32'hb9e5e40b),
	.w8(32'h392bb550),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1b6d),
	.w1(32'hbb3d0007),
	.w2(32'hbba23089),
	.w3(32'hbb92e303),
	.w4(32'hbaa83261),
	.w5(32'hbb007349),
	.w6(32'hbb0d62ca),
	.w7(32'hbb630340),
	.w8(32'hbb84bc67),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a042586),
	.w1(32'hba61913e),
	.w2(32'hba49e3b9),
	.w3(32'h3a8ba131),
	.w4(32'hbae498fe),
	.w5(32'h3b009cb5),
	.w6(32'h3833b433),
	.w7(32'hba717818),
	.w8(32'hba876333),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b3561),
	.w1(32'h3b039428),
	.w2(32'hba35615e),
	.w3(32'hbb53e4b1),
	.w4(32'h3a4d1804),
	.w5(32'hbbbe3243),
	.w6(32'hbb685a52),
	.w7(32'h3a8d7af5),
	.w8(32'hbb69f4c2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d76b6),
	.w1(32'h394ffcef),
	.w2(32'h3a5e2d58),
	.w3(32'hbb8ecd54),
	.w4(32'hb9f5921d),
	.w5(32'h3b42e6ed),
	.w6(32'hb8fcc126),
	.w7(32'h3aaf89a9),
	.w8(32'h3a879289),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7eec3),
	.w1(32'h3b1cba77),
	.w2(32'h3a7374ed),
	.w3(32'h3a025d17),
	.w4(32'h3adb0951),
	.w5(32'hba246a3b),
	.w6(32'hba03dc1b),
	.w7(32'h3a68ccbb),
	.w8(32'hba6123d0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b312d20),
	.w1(32'hbb55630b),
	.w2(32'hb7fb49a8),
	.w3(32'h398afe44),
	.w4(32'hbb5b5f14),
	.w5(32'hbaa0e37d),
	.w6(32'h3b1d1f17),
	.w7(32'hbb3b3394),
	.w8(32'hbb515d86),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b701333),
	.w1(32'h3b8afdd8),
	.w2(32'h3ba2395e),
	.w3(32'h3b2c28c1),
	.w4(32'h3c1cb91d),
	.w5(32'h3b8e0c56),
	.w6(32'h3ac2587b),
	.w7(32'h3ba49c95),
	.w8(32'h3b6f2a5c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33f176),
	.w1(32'hbb72d3bc),
	.w2(32'hbb1410d6),
	.w3(32'h3bbefbda),
	.w4(32'hbada0b84),
	.w5(32'hbba151ac),
	.w6(32'h3bb9953d),
	.w7(32'h3b86f98f),
	.w8(32'h3b9f2e52),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9e3aa),
	.w1(32'hbaebeec7),
	.w2(32'hba5a4243),
	.w3(32'hbba6fe89),
	.w4(32'hba7a763a),
	.w5(32'hbad090db),
	.w6(32'h3af4be28),
	.w7(32'hbade30af),
	.w8(32'hbb64ab81),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56f244),
	.w1(32'hbb6e1b1d),
	.w2(32'hbaacf3e5),
	.w3(32'hbb0084fd),
	.w4(32'hbaedb7a6),
	.w5(32'h3b475857),
	.w6(32'hba2d82c4),
	.w7(32'h397d6551),
	.w8(32'h3ae11ce4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3293e2),
	.w1(32'hbb7f6318),
	.w2(32'hbb37acdc),
	.w3(32'hbb84b3c2),
	.w4(32'hbba06cb1),
	.w5(32'hbb4f057e),
	.w6(32'hbb2e3b69),
	.w7(32'hbba974ca),
	.w8(32'hbb7e5794),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b034713),
	.w1(32'hba7e7688),
	.w2(32'hba824320),
	.w3(32'h3b30872c),
	.w4(32'h3a7364ca),
	.w5(32'hb95ededc),
	.w6(32'h3abdfd3d),
	.w7(32'h3afa28fb),
	.w8(32'h39c7ab41),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90130e),
	.w1(32'h3a7296d3),
	.w2(32'h39e4307e),
	.w3(32'h3aeea403),
	.w4(32'hba968d5e),
	.w5(32'h3abae6bf),
	.w6(32'hbaec3b4f),
	.w7(32'h3b885300),
	.w8(32'h3ada2d24),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ade42),
	.w1(32'hbaad86a0),
	.w2(32'hba549e74),
	.w3(32'hbae6872a),
	.w4(32'hbaadae8d),
	.w5(32'h39aa7e7d),
	.w6(32'hbb5068a5),
	.w7(32'hba5cc7ca),
	.w8(32'hba8a8c65),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4adf9f),
	.w1(32'hbb0ec746),
	.w2(32'hbb85c9d3),
	.w3(32'hbabb876f),
	.w4(32'hbae5d472),
	.w5(32'hbb31a054),
	.w6(32'hba68483a),
	.w7(32'h3a0f4768),
	.w8(32'h3a38b6a1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d4203),
	.w1(32'h3b0b704b),
	.w2(32'h3ac2058f),
	.w3(32'h3aa2b265),
	.w4(32'h3b0cd74c),
	.w5(32'h3b1c077e),
	.w6(32'h3b0b8b2a),
	.w7(32'h3b80e0bd),
	.w8(32'h3abc3d97),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96f38a),
	.w1(32'hbb204aff),
	.w2(32'hb8df9975),
	.w3(32'h3b1e3874),
	.w4(32'hbb3b73ed),
	.w5(32'hbbba8b4f),
	.w6(32'h3b19f86f),
	.w7(32'hbb7ca5f6),
	.w8(32'hbb498224),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbfeba),
	.w1(32'hb8fb1c40),
	.w2(32'hbb02d0c7),
	.w3(32'hbb027955),
	.w4(32'hbae7f04c),
	.w5(32'h3ae86cf0),
	.w6(32'hbb24125e),
	.w7(32'hbb1500dd),
	.w8(32'hba6c775f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53e957),
	.w1(32'hb9e61dd7),
	.w2(32'hbb260cbe),
	.w3(32'hbb030e5f),
	.w4(32'hbb755d2c),
	.w5(32'hbb4514c7),
	.w6(32'hba28739f),
	.w7(32'hbb7ad0f1),
	.w8(32'hbb688013),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949e2a3),
	.w1(32'hb9129dfc),
	.w2(32'hba440025),
	.w3(32'h3aa9e3e3),
	.w4(32'h3ab1a191),
	.w5(32'h3a20289e),
	.w6(32'h3ae85cf5),
	.w7(32'hbba7612f),
	.w8(32'hbad2defd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd8345),
	.w1(32'h39611f87),
	.w2(32'hbaca14dc),
	.w3(32'hbb999190),
	.w4(32'hba546b5b),
	.w5(32'hb90f25d6),
	.w6(32'hbadc426a),
	.w7(32'hba2719d2),
	.w8(32'hba39d4ff),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86f27e),
	.w1(32'hbb15c5df),
	.w2(32'hba835d82),
	.w3(32'hba657fa6),
	.w4(32'hb9ab138a),
	.w5(32'h3b2b8a56),
	.w6(32'hbb1399ce),
	.w7(32'hbb2b1958),
	.w8(32'hbb3636bc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38d377),
	.w1(32'hbab0a5ac),
	.w2(32'hba8d0190),
	.w3(32'h39a9f3d7),
	.w4(32'h3ad7f7a0),
	.w5(32'hba414405),
	.w6(32'hbb552c15),
	.w7(32'h3b02af03),
	.w8(32'h3a5e7b97),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba1adf),
	.w1(32'h3ad5e012),
	.w2(32'h3b41ecbd),
	.w3(32'h3b105214),
	.w4(32'h3a84c186),
	.w5(32'hb9c21640),
	.w6(32'h3b1a5972),
	.w7(32'h3b6ab120),
	.w8(32'h3ad62d13),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9986651),
	.w1(32'h3aee1574),
	.w2(32'h39fac030),
	.w3(32'hbae0898a),
	.w4(32'hbaa7e4e5),
	.w5(32'hb962902a),
	.w6(32'h3a93821f),
	.w7(32'hbab07a73),
	.w8(32'hbb221ba7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba338d75),
	.w1(32'hb96457b9),
	.w2(32'hb9dc243a),
	.w3(32'h37f501b9),
	.w4(32'h3b3873a2),
	.w5(32'hb8ae68d4),
	.w6(32'hbb08b0d0),
	.w7(32'h3956170e),
	.w8(32'hbb69a76b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebda8d),
	.w1(32'hb935ac62),
	.w2(32'hbae68b52),
	.w3(32'h3aafdd4d),
	.w4(32'h3b317c0d),
	.w5(32'hba6b56c8),
	.w6(32'hbae78a39),
	.w7(32'h3aa9fe06),
	.w8(32'h38b6cec5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b22da),
	.w1(32'hbae7ea08),
	.w2(32'hbade56f9),
	.w3(32'hbb232b3f),
	.w4(32'hbb005b02),
	.w5(32'h3a9988b5),
	.w6(32'hb9bd00ff),
	.w7(32'h3a57f3a6),
	.w8(32'hb9a7a38c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10eafa),
	.w1(32'h3ad3350f),
	.w2(32'hba8696ca),
	.w3(32'hbb2d51c0),
	.w4(32'h3bec6c4c),
	.w5(32'h378fa866),
	.w6(32'hbaafd526),
	.w7(32'h3b871102),
	.w8(32'h3b36a0a5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91c2b3),
	.w1(32'h3b8aa237),
	.w2(32'h3a8bbadf),
	.w3(32'h3b28459a),
	.w4(32'h3b7a3d20),
	.w5(32'h3b8ec6d5),
	.w6(32'hba80e174),
	.w7(32'h3b1141a4),
	.w8(32'h3b79c9de),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7144b3),
	.w1(32'hbb023fa2),
	.w2(32'hbabe6583),
	.w3(32'h3b15ad37),
	.w4(32'h3a700ef0),
	.w5(32'h3ae50662),
	.w6(32'hb97be516),
	.w7(32'hba3d9485),
	.w8(32'hbaade070),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9634669),
	.w1(32'hbab3f591),
	.w2(32'h3958311c),
	.w3(32'hbaa33864),
	.w4(32'h3a7e75e0),
	.w5(32'h3b491977),
	.w6(32'hbad9966c),
	.w7(32'h3b231801),
	.w8(32'hba76b7fb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4eaa05),
	.w1(32'h38baa64c),
	.w2(32'h3a89862b),
	.w3(32'hba536455),
	.w4(32'h3a1bdcef),
	.w5(32'hba8c25c1),
	.w6(32'hbab68af6),
	.w7(32'hbb4ee814),
	.w8(32'hbaf1c96e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab62db2),
	.w1(32'h3af93ea8),
	.w2(32'h398ef022),
	.w3(32'hbb324613),
	.w4(32'h3b151eda),
	.w5(32'h3ad42a06),
	.w6(32'hbb85214d),
	.w7(32'h3bc80fda),
	.w8(32'h3b55d6b4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36baa3),
	.w1(32'hbaa24aa9),
	.w2(32'hba505aee),
	.w3(32'hba11426a),
	.w4(32'hba8474bd),
	.w5(32'h3ade5b60),
	.w6(32'hbac54b40),
	.w7(32'h3a8518bf),
	.w8(32'h3b0a97af),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3737f6),
	.w1(32'h3b874447),
	.w2(32'h393a5564),
	.w3(32'h3a22982a),
	.w4(32'hba296089),
	.w5(32'hbb54de12),
	.w6(32'hbb271d28),
	.w7(32'hbb24fb01),
	.w8(32'hbb74ed41),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d7267),
	.w1(32'hbacb807c),
	.w2(32'hbaeff4d1),
	.w3(32'hbb6bfbb2),
	.w4(32'h3a880f5a),
	.w5(32'h3a7f0e9f),
	.w6(32'hbb3a6423),
	.w7(32'h3a907729),
	.w8(32'h3ad8325e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a802cc4),
	.w1(32'h3b235ef4),
	.w2(32'h3a67d6fc),
	.w3(32'h3b7b77e6),
	.w4(32'hbafc7c0e),
	.w5(32'hb8631215),
	.w6(32'h3b56f204),
	.w7(32'hbaa982b0),
	.w8(32'hbad79bfb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a405c1a),
	.w1(32'h3ac0baaa),
	.w2(32'hbb44c727),
	.w3(32'hb887c8d6),
	.w4(32'hb99c4b74),
	.w5(32'hba7c24b7),
	.w6(32'hbb0151c4),
	.w7(32'hb82ae63a),
	.w8(32'hbb830a4d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932b6d),
	.w1(32'hbab6b53f),
	.w2(32'h3a27b291),
	.w3(32'hbb8530c1),
	.w4(32'h36d0a257),
	.w5(32'h3a843c41),
	.w6(32'hb86e85d2),
	.w7(32'h393c6d5f),
	.w8(32'h39aaa243),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39109fc9),
	.w1(32'hbb119c31),
	.w2(32'hbb448013),
	.w3(32'h3b217c85),
	.w4(32'hbaaa2fcc),
	.w5(32'h3a0ea0b1),
	.w6(32'h3b18a0c0),
	.w7(32'hba88578a),
	.w8(32'h3a80ebb2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d6a0b),
	.w1(32'hb9f887b7),
	.w2(32'h39b4f634),
	.w3(32'h3943c4ce),
	.w4(32'hba54f2f1),
	.w5(32'h3ace3cc1),
	.w6(32'h3b2b0717),
	.w7(32'h39fd400b),
	.w8(32'h3b81d445),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f2e67),
	.w1(32'hbb7c5239),
	.w2(32'hbadd3864),
	.w3(32'h3a9b4330),
	.w4(32'hbb5b50c6),
	.w5(32'hbba75583),
	.w6(32'h3b4def0e),
	.w7(32'hbb0d2331),
	.w8(32'hbb3f675b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fde989),
	.w1(32'h3a448fb4),
	.w2(32'hba24a840),
	.w3(32'hbb3e5695),
	.w4(32'hbaff9b7f),
	.w5(32'hbb8d35fa),
	.w6(32'hbb2918d2),
	.w7(32'hbb5c28bb),
	.w8(32'hbb4077de),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05f0e7),
	.w1(32'hbaf6d418),
	.w2(32'hba8e9609),
	.w3(32'hbb6480dd),
	.w4(32'hbb0dfe4b),
	.w5(32'h3a92c379),
	.w6(32'hbb2867c5),
	.w7(32'hbaf40610),
	.w8(32'h39b2c93d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac53f21),
	.w1(32'hbb36f162),
	.w2(32'hbb02855c),
	.w3(32'hba9a5b76),
	.w4(32'hbb9a7c36),
	.w5(32'hbb5dc9f0),
	.w6(32'hbaed9744),
	.w7(32'hbb1b4bf2),
	.w8(32'hbbbcfd6d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb370476),
	.w1(32'h3ad85836),
	.w2(32'h3b15f3c2),
	.w3(32'hbac47b2b),
	.w4(32'hba942297),
	.w5(32'h3a3fd3c6),
	.w6(32'hbb3e87bf),
	.w7(32'hb96f0afa),
	.w8(32'hbb3555ea),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac329fe),
	.w1(32'hbb222b3b),
	.w2(32'h3a38435f),
	.w3(32'h3a1ad380),
	.w4(32'hbb24a551),
	.w5(32'h3a028c55),
	.w6(32'hbae4b572),
	.w7(32'h3a1756e0),
	.w8(32'hba0ee71c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e1f12),
	.w1(32'hbaefd386),
	.w2(32'hbb3e97a5),
	.w3(32'h38e4af45),
	.w4(32'h394ce7a9),
	.w5(32'h39e20aa8),
	.w6(32'hbac036c2),
	.w7(32'h3aafcab9),
	.w8(32'h3aaf42c0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e7aa8),
	.w1(32'h3b90200a),
	.w2(32'h3abccdaa),
	.w3(32'h3a396746),
	.w4(32'h38af7b97),
	.w5(32'hbb261965),
	.w6(32'hbae09a7d),
	.w7(32'h38856419),
	.w8(32'hbb2935d2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fe145),
	.w1(32'h3b2ecdbf),
	.w2(32'hbaf38e6f),
	.w3(32'hbb872b67),
	.w4(32'hbaaaad4f),
	.w5(32'h39e8db04),
	.w6(32'hbb19aa11),
	.w7(32'hbb515e9e),
	.w8(32'h3b2d5af1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb424ba8),
	.w1(32'h3a8b2ef4),
	.w2(32'hb99ae6a4),
	.w3(32'hbb025ea9),
	.w4(32'hb9c8536b),
	.w5(32'hbb01ea14),
	.w6(32'hbb727dbc),
	.w7(32'hbb062b6c),
	.w8(32'hbbab7b59),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65523f),
	.w1(32'h3b93042f),
	.w2(32'h3bb34abf),
	.w3(32'h3a6eb179),
	.w4(32'h3c237452),
	.w5(32'h3bda1715),
	.w6(32'hbb879945),
	.w7(32'h3bc66298),
	.w8(32'h39b1d169),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde80bf),
	.w1(32'h3a271072),
	.w2(32'hb932897c),
	.w3(32'h3b75684a),
	.w4(32'h3a4b0ea3),
	.w5(32'h3aa29c85),
	.w6(32'h3abc55c9),
	.w7(32'h3a91c5f0),
	.w8(32'h3b10ebb6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a787ac),
	.w1(32'hbb997900),
	.w2(32'hbb491e7c),
	.w3(32'hba184568),
	.w4(32'hbb39e828),
	.w5(32'hbae84659),
	.w6(32'h399d7f05),
	.w7(32'h3a03f6e7),
	.w8(32'hbaff4d27),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aadc1),
	.w1(32'h3b04604f),
	.w2(32'h3b52ecb4),
	.w3(32'hbb76017e),
	.w4(32'hb959bf37),
	.w5(32'h3af9f9d8),
	.w6(32'hb91ded84),
	.w7(32'h3a340588),
	.w8(32'hb9339730),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39b580),
	.w1(32'hba5f1bbf),
	.w2(32'h3b8f075f),
	.w3(32'h3a8298e2),
	.w4(32'hba2f8b39),
	.w5(32'h3b47be06),
	.w6(32'h3b214b7d),
	.w7(32'h3a365868),
	.w8(32'hbab8253f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31c137),
	.w1(32'h3b38839a),
	.w2(32'hba80ecae),
	.w3(32'hb8bce76d),
	.w4(32'h3a6dc483),
	.w5(32'hb9a4f587),
	.w6(32'h398f03d4),
	.w7(32'h3b1b967d),
	.w8(32'h3ae85d6c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01aef7),
	.w1(32'h3a2e24f3),
	.w2(32'h3b064d68),
	.w3(32'hb8d84b18),
	.w4(32'h3b596351),
	.w5(32'h39aa4738),
	.w6(32'h3a29097d),
	.w7(32'h3a81a80a),
	.w8(32'h3b1fb2f6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d69ba),
	.w1(32'hbb39ad28),
	.w2(32'hbb61cd44),
	.w3(32'hbb02010d),
	.w4(32'hba919004),
	.w5(32'hbb12042a),
	.w6(32'hbad91df3),
	.w7(32'hbb7953c8),
	.w8(32'hba9e27ee),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a453dda),
	.w1(32'h3ac71817),
	.w2(32'hb9071130),
	.w3(32'h3a6f016b),
	.w4(32'hbaa84f98),
	.w5(32'h3b3b87fc),
	.w6(32'hbaa2a2d3),
	.w7(32'hb949aa73),
	.w8(32'h3a16e1bd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe6202),
	.w1(32'h3bd22993),
	.w2(32'h3bacff95),
	.w3(32'h3aed3297),
	.w4(32'h3a415691),
	.w5(32'h38cb50db),
	.w6(32'h3b663c03),
	.w7(32'h3adbadff),
	.w8(32'h3a9fb839),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9561db),
	.w1(32'hba089f88),
	.w2(32'hb804fa03),
	.w3(32'hb9f25eda),
	.w4(32'hbab3e226),
	.w5(32'h3ae990c8),
	.w6(32'h398efba5),
	.w7(32'hbb528b73),
	.w8(32'h3a3f435d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4035b),
	.w1(32'h39863511),
	.w2(32'hbba41538),
	.w3(32'h39baf9a2),
	.w4(32'hba09aae2),
	.w5(32'hb9c114a3),
	.w6(32'h39b47488),
	.w7(32'h388f88ff),
	.w8(32'hbaf1ba91),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34072e),
	.w1(32'h39a25da8),
	.w2(32'hba4e853e),
	.w3(32'hbb72c891),
	.w4(32'h3a0486c5),
	.w5(32'h3b14f850),
	.w6(32'hbae4c7eb),
	.w7(32'h3b6ec04c),
	.w8(32'h3b6a651c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30cffd),
	.w1(32'hbabc2942),
	.w2(32'hbb437c43),
	.w3(32'h3b46687c),
	.w4(32'hbac62eba),
	.w5(32'hba158ce0),
	.w6(32'h3b6923e8),
	.w7(32'hba8b7484),
	.w8(32'hba984a2f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984be3a),
	.w1(32'h3b4589bf),
	.w2(32'h3ac75a9e),
	.w3(32'h3b07d862),
	.w4(32'h3bc43d20),
	.w5(32'h3b776451),
	.w6(32'hb85d596a),
	.w7(32'h3adc01f7),
	.w8(32'hbb3651eb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a025af1),
	.w1(32'hba0e3d86),
	.w2(32'hbb21d1cb),
	.w3(32'hb9c54fcd),
	.w4(32'hbaa8b40d),
	.w5(32'h3a58f036),
	.w6(32'h3a543bde),
	.w7(32'hb9422f10),
	.w8(32'hbae12483),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba609b55),
	.w1(32'h3baa0902),
	.w2(32'h3a03a6bc),
	.w3(32'hb8c879d9),
	.w4(32'h3b4ec73d),
	.w5(32'h3b4af702),
	.w6(32'h3a54cf91),
	.w7(32'h3b26c2f8),
	.w8(32'h3b1cd404),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8edc67),
	.w1(32'hb9018c64),
	.w2(32'hbb7c82cf),
	.w3(32'hba9487c4),
	.w4(32'h3ae792e5),
	.w5(32'h3a3b90b5),
	.w6(32'hb9a0cd8b),
	.w7(32'h3b87db24),
	.w8(32'h3b59ee7d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b9ac1),
	.w1(32'hb950ed96),
	.w2(32'h39ffa5fb),
	.w3(32'h3b259814),
	.w4(32'h3a5a9e31),
	.w5(32'h3abb3990),
	.w6(32'h3af0920b),
	.w7(32'hb9158513),
	.w8(32'h3a9d22af),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392eeb05),
	.w1(32'hbabcc665),
	.w2(32'hba8e96e4),
	.w3(32'h3937b87e),
	.w4(32'hbb4ec080),
	.w5(32'hba2eecc3),
	.w6(32'hbb1e9438),
	.w7(32'hba870a2b),
	.w8(32'h3b2403cb),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f1516),
	.w1(32'h3b568535),
	.w2(32'h3b1d6887),
	.w3(32'h3a98d252),
	.w4(32'h3b86a075),
	.w5(32'hbaeb0efb),
	.w6(32'h39ecef6c),
	.w7(32'h3c165684),
	.w8(32'h3bbf2fbb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10e652),
	.w1(32'hbb33747b),
	.w2(32'hba8cc5e9),
	.w3(32'hbac2e0a9),
	.w4(32'hbaee9cac),
	.w5(32'h3ab861de),
	.w6(32'h3b0b6e62),
	.w7(32'hbb129a5b),
	.w8(32'h3b271c72),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a41f4c),
	.w1(32'hbb1246dc),
	.w2(32'h3b395df3),
	.w3(32'hba8371b1),
	.w4(32'hbb6fb04c),
	.w5(32'h39b6d8f8),
	.w6(32'h3a85f4ad),
	.w7(32'h3af5364a),
	.w8(32'h3b8d2eee),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a693754),
	.w1(32'h3bbce31d),
	.w2(32'h3baef754),
	.w3(32'hb9bd9bd7),
	.w4(32'hb912d3df),
	.w5(32'h396a0a65),
	.w6(32'h392c6a50),
	.w7(32'h3b691edb),
	.w8(32'h3b82c7ad),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06be90),
	.w1(32'hb97e7f16),
	.w2(32'hbac8552f),
	.w3(32'h3b1fb745),
	.w4(32'hba92d033),
	.w5(32'hba6c4cee),
	.w6(32'h3ba44aa3),
	.w7(32'h39e9d58d),
	.w8(32'hbb2638e5),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f8e07),
	.w1(32'hba3ecf7c),
	.w2(32'hbb07820b),
	.w3(32'hbae3de40),
	.w4(32'hbaefb2c4),
	.w5(32'hbb13fa21),
	.w6(32'h39549367),
	.w7(32'hba860816),
	.w8(32'h3a613368),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9fb3e),
	.w1(32'hbb1b84dc),
	.w2(32'hba071da9),
	.w3(32'hba72cfd5),
	.w4(32'hbb30c14a),
	.w5(32'hba63a894),
	.w6(32'hbac678cc),
	.w7(32'hbac885a7),
	.w8(32'hba9bab13),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb083563),
	.w1(32'hbac3747d),
	.w2(32'hbbab92ee),
	.w3(32'hbb43423a),
	.w4(32'hbb4a80c4),
	.w5(32'hbb1d9ac2),
	.w6(32'hbb41f81a),
	.w7(32'hbaaa8eb6),
	.w8(32'hba7284f9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc010dd1),
	.w1(32'hba29f4d0),
	.w2(32'hbafeb5d5),
	.w3(32'hbb886e8e),
	.w4(32'hbb4e67b6),
	.w5(32'hb9c008aa),
	.w6(32'hbb5f3283),
	.w7(32'hbb078796),
	.w8(32'hbb20270a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964583c),
	.w1(32'h3b1e619b),
	.w2(32'h3ac73f97),
	.w3(32'h3a81ce77),
	.w4(32'hba1ef20a),
	.w5(32'h3b240911),
	.w6(32'h3a5d5d8a),
	.w7(32'hba157960),
	.w8(32'h3b5b3776),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb125b59),
	.w1(32'h394bd40c),
	.w2(32'hba137d29),
	.w3(32'hbb90d236),
	.w4(32'h3b388e25),
	.w5(32'h3b1a536a),
	.w6(32'hba8ec09e),
	.w7(32'h39a3bdc2),
	.w8(32'hba146ab4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904ccd),
	.w1(32'hba8e4331),
	.w2(32'hba014cf0),
	.w3(32'hbaeeca5b),
	.w4(32'hbae195a2),
	.w5(32'h3aefe3ed),
	.w6(32'hba3b83e2),
	.w7(32'hbb47894c),
	.w8(32'hba4373ee),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399eae30),
	.w1(32'h378ad26a),
	.w2(32'hbb80ac6c),
	.w3(32'hba3ad8d1),
	.w4(32'h39b3ea24),
	.w5(32'hbb1d52a7),
	.w6(32'hba9e7131),
	.w7(32'hba1a117a),
	.w8(32'hbb457297),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e87d6),
	.w1(32'h39fa3ecb),
	.w2(32'h399bf3df),
	.w3(32'h3b972934),
	.w4(32'hba990f12),
	.w5(32'hbb5b38cb),
	.w6(32'h3aa4e7ec),
	.w7(32'hb9c5c42d),
	.w8(32'hbace8387),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3799d539),
	.w1(32'h3b4b9fab),
	.w2(32'h3aa7d82c),
	.w3(32'h3a94522e),
	.w4(32'h3aefeeda),
	.w5(32'hbb2992a0),
	.w6(32'hbb1cc442),
	.w7(32'h3b7924b2),
	.w8(32'h3ae2876b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aefc6),
	.w1(32'hbb341de4),
	.w2(32'hbac1c20e),
	.w3(32'hba15068c),
	.w4(32'hbb18a8c7),
	.w5(32'hba11c44e),
	.w6(32'h3a6896cd),
	.w7(32'hbb2e9e60),
	.w8(32'hb8c0b1ad),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32adf7),
	.w1(32'h3b55d9be),
	.w2(32'hb9809387),
	.w3(32'h3ae61b12),
	.w4(32'hbb361509),
	.w5(32'hb9e83854),
	.w6(32'h3b119d81),
	.w7(32'hbaf68a84),
	.w8(32'h39e34289),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdbec7),
	.w1(32'hba5f4bb4),
	.w2(32'hbabe9bb7),
	.w3(32'hbae7856d),
	.w4(32'hbb0ef293),
	.w5(32'hbaf0e49e),
	.w6(32'hbad1ea0d),
	.w7(32'hbb58104d),
	.w8(32'hbb70dc36),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba962088),
	.w1(32'h3ba32a98),
	.w2(32'h3bb6c042),
	.w3(32'hbb208389),
	.w4(32'h3bb95321),
	.w5(32'h3b6c5a44),
	.w6(32'hbb034912),
	.w7(32'h3baeed59),
	.w8(32'h3b6da315),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97d62c),
	.w1(32'h3a4d7907),
	.w2(32'h3af8af08),
	.w3(32'h3b8fc1b3),
	.w4(32'hbab7364a),
	.w5(32'h3b4fb6a1),
	.w6(32'h3ba51316),
	.w7(32'h3a49c373),
	.w8(32'h3b502fc7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8174f7),
	.w1(32'hba8abcdc),
	.w2(32'hba0e31a2),
	.w3(32'h3bae33c5),
	.w4(32'hb9542103),
	.w5(32'h397ce7fc),
	.w6(32'h3bb8f408),
	.w7(32'h3a6589ef),
	.w8(32'hba4746d0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad34ebe),
	.w1(32'h3b2fa87c),
	.w2(32'h3a68450f),
	.w3(32'h3a767319),
	.w4(32'hb9050886),
	.w5(32'hb9f772b4),
	.w6(32'hba9d6e61),
	.w7(32'h3b90f1fc),
	.w8(32'h3bbfdf44),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d10152),
	.w1(32'hbbdb8db2),
	.w2(32'hbba0ea2a),
	.w3(32'hba82acc4),
	.w4(32'hbbab9096),
	.w5(32'hba58875a),
	.w6(32'h3bad1c9c),
	.w7(32'hbb45668b),
	.w8(32'hb8b21113),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc6195),
	.w1(32'hbae8ba71),
	.w2(32'h3bc0386f),
	.w3(32'hbb85b523),
	.w4(32'h3b42a91e),
	.w5(32'h3c1cd79e),
	.w6(32'hbb1957c2),
	.w7(32'h3bb7e8f5),
	.w8(32'h3bd33878),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad22764),
	.w1(32'hbaff0085),
	.w2(32'hb958d078),
	.w3(32'hbb2e0cc2),
	.w4(32'hbbe055ac),
	.w5(32'hbb08fc2a),
	.w6(32'hba0d024b),
	.w7(32'hbbe722ff),
	.w8(32'hbaf832ff),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c710b),
	.w1(32'hba508e60),
	.w2(32'h3ba2ff32),
	.w3(32'hbafff837),
	.w4(32'hbb1c5592),
	.w5(32'hbb08a6e1),
	.w6(32'hbade1678),
	.w7(32'hbbb7a432),
	.w8(32'h39c4094f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1661fd),
	.w1(32'hbb10fa0d),
	.w2(32'hbb97d592),
	.w3(32'hbb934f8b),
	.w4(32'hb86579d2),
	.w5(32'hbbb86aea),
	.w6(32'h3c179ea8),
	.w7(32'h3a821fe9),
	.w8(32'hbbfadaed),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d19cb),
	.w1(32'h39c8fa50),
	.w2(32'h3af5ea9b),
	.w3(32'hbc237b90),
	.w4(32'h3b3c2de8),
	.w5(32'h3bce5282),
	.w6(32'hbbfadda8),
	.w7(32'h3ac786af),
	.w8(32'hbb30e5a4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43a440),
	.w1(32'hba89d385),
	.w2(32'h393e5f1a),
	.w3(32'hbb34f231),
	.w4(32'hbac52d1b),
	.w5(32'h3ad83aac),
	.w6(32'hbb55e78f),
	.w7(32'hba57ce6a),
	.w8(32'hbace6896),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a45925),
	.w1(32'hbb041788),
	.w2(32'hb978a3af),
	.w3(32'h3b53d512),
	.w4(32'h3aa55e41),
	.w5(32'h3b859aff),
	.w6(32'hbb20ae50),
	.w7(32'h3b1ca75b),
	.w8(32'h3b1251b5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2387d4),
	.w1(32'h3acf2e65),
	.w2(32'hbb1d02ca),
	.w3(32'h3a8e258e),
	.w4(32'h3b125c19),
	.w5(32'hbb301903),
	.w6(32'h39d274e2),
	.w7(32'h3ab31bd3),
	.w8(32'hbb1e0028),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6dac4),
	.w1(32'hbb951dcb),
	.w2(32'hbaa2b9fe),
	.w3(32'hb9bfeae2),
	.w4(32'hbbc71f70),
	.w5(32'hbb4886e2),
	.w6(32'hbbf5e54a),
	.w7(32'h3adf5016),
	.w8(32'h3984873f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaca69f),
	.w1(32'h3b83ece1),
	.w2(32'h3b222bab),
	.w3(32'h3be03be6),
	.w4(32'h3b4b3c28),
	.w5(32'hbbac6275),
	.w6(32'h3ba40d83),
	.w7(32'h3bf050d3),
	.w8(32'hbabe64d5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7aef3),
	.w1(32'h3b123535),
	.w2(32'hba8b91e1),
	.w3(32'h3bbf153e),
	.w4(32'h3b88043e),
	.w5(32'h3a339b5c),
	.w6(32'h3b9cdcf1),
	.w7(32'h3b904661),
	.w8(32'h3b9cf7e5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fbf72),
	.w1(32'h3c6e2d9a),
	.w2(32'h3c2009a8),
	.w3(32'h3b7512c9),
	.w4(32'h3cb01edd),
	.w5(32'h3c720106),
	.w6(32'hba2bd6a6),
	.w7(32'h3c874b40),
	.w8(32'h3c3a28a2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b123806),
	.w1(32'h3b96056d),
	.w2(32'hbb727c97),
	.w3(32'h3b275b70),
	.w4(32'h3c08f2ad),
	.w5(32'h3bbc1fb2),
	.w6(32'hb9cc451e),
	.w7(32'h3b89d189),
	.w8(32'h3b2f76d5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00cc53),
	.w1(32'h3ac5866e),
	.w2(32'h3ae952aa),
	.w3(32'h3ae49305),
	.w4(32'h3af86537),
	.w5(32'h39502923),
	.w6(32'hbb7e2a4b),
	.w7(32'hbaece816),
	.w8(32'h3afafc1e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96db497),
	.w1(32'hbb5d222a),
	.w2(32'h39301365),
	.w3(32'h3af910ea),
	.w4(32'h3b1ac151),
	.w5(32'h3a94888f),
	.w6(32'h3a9da0b9),
	.w7(32'h3b7f08fc),
	.w8(32'h3aedb907),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ed97b),
	.w1(32'h3b48a533),
	.w2(32'hbb403419),
	.w3(32'h3bb9f5da),
	.w4(32'h3b4ac102),
	.w5(32'h3bc00891),
	.w6(32'h3bc7f486),
	.w7(32'h3abbc494),
	.w8(32'hba449804),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71c765),
	.w1(32'h3bc9cb51),
	.w2(32'h3a669bd1),
	.w3(32'hbb4972bf),
	.w4(32'h3ba58135),
	.w5(32'hbb904885),
	.w6(32'h3a913ece),
	.w7(32'hbaf99185),
	.w8(32'h38b1e656),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcd39e),
	.w1(32'hbc094930),
	.w2(32'hbb23dd37),
	.w3(32'h3b154ed5),
	.w4(32'hbc444fed),
	.w5(32'hbb9bb8cd),
	.w6(32'hbb1d1d3a),
	.w7(32'hbbde5449),
	.w8(32'h3a135ae6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1334fa),
	.w1(32'hba050e56),
	.w2(32'h3a1e76d8),
	.w3(32'hbb09670b),
	.w4(32'hbbb58332),
	.w5(32'h3b2cb0c9),
	.w6(32'h3921b25f),
	.w7(32'hb8eb34f5),
	.w8(32'h3b7b0b03),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1edf1),
	.w1(32'h3a5fe126),
	.w2(32'hba676fe5),
	.w3(32'h3c232eb3),
	.w4(32'h3ad4ce7e),
	.w5(32'hba506e80),
	.w6(32'h3b4f306f),
	.w7(32'h3aad9283),
	.w8(32'hbb3d599f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baef780),
	.w1(32'h3b5c1357),
	.w2(32'hb9c782af),
	.w3(32'h3bfc5420),
	.w4(32'hbafbc0e2),
	.w5(32'h3a177de1),
	.w6(32'h3bc6a8c0),
	.w7(32'hbb423f54),
	.w8(32'hba8b73b3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07bf00),
	.w1(32'hba0d312c),
	.w2(32'hba81c518),
	.w3(32'hbb33aa9f),
	.w4(32'hbb9029f2),
	.w5(32'h3b038ee0),
	.w6(32'hb936c577),
	.w7(32'hbb1f4beb),
	.w8(32'h3a0fbef6),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fd8bd),
	.w1(32'hbbc9ae32),
	.w2(32'hba7909f1),
	.w3(32'hbbb7fe1a),
	.w4(32'hbb948106),
	.w5(32'hbb62e021),
	.w6(32'hba9c8527),
	.w7(32'h3b2f8277),
	.w8(32'h3be1b866),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29b1a6),
	.w1(32'h3bce0cea),
	.w2(32'h3a5278ce),
	.w3(32'hb9b3e4a5),
	.w4(32'h3c2aeea2),
	.w5(32'h3b5d9091),
	.w6(32'h39fe9b2c),
	.w7(32'h3c06de9b),
	.w8(32'h3c21be5c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9148440),
	.w1(32'h3b371a74),
	.w2(32'h3b07ca38),
	.w3(32'hbb9c523b),
	.w4(32'h3bf65e8c),
	.w5(32'h3ba6c8ba),
	.w6(32'h3b484ac0),
	.w7(32'h3c1d36f9),
	.w8(32'h3c248f1d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ede4b6),
	.w1(32'hbb6dd113),
	.w2(32'h3b73c950),
	.w3(32'hbade632a),
	.w4(32'hbb9c6ca6),
	.w5(32'hba6c63d5),
	.w6(32'h3a3c78dd),
	.w7(32'h3bb088c8),
	.w8(32'h3ac7cb51),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14e030),
	.w1(32'hbad37ff2),
	.w2(32'hb9f124a7),
	.w3(32'h3acc80bc),
	.w4(32'h3a606c2d),
	.w5(32'h3bed19bf),
	.w6(32'hbb489619),
	.w7(32'hb96f1ecc),
	.w8(32'hba2ee370),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee9e49),
	.w1(32'hbb7befe4),
	.w2(32'hbc0f6608),
	.w3(32'hbc2e29f2),
	.w4(32'hbb40cca8),
	.w5(32'h3c0b8261),
	.w6(32'hbbf43278),
	.w7(32'hb9a2371b),
	.w8(32'h3abf04c1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e5c657),
	.w1(32'h3a973176),
	.w2(32'h3b7398f2),
	.w3(32'h3c4fcf02),
	.w4(32'hbb2a0eda),
	.w5(32'hbbc908cb),
	.w6(32'h3b0d307d),
	.w7(32'hba2b33bc),
	.w8(32'hbbc9481e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31ff30),
	.w1(32'h3bbe2030),
	.w2(32'hbaa4ee9c),
	.w3(32'hbb7e8768),
	.w4(32'hbaa77297),
	.w5(32'hbb84c020),
	.w6(32'hbb832547),
	.w7(32'h3a494fa6),
	.w8(32'hbac1c47d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5988d1),
	.w1(32'h3b9f8099),
	.w2(32'h3c085b1e),
	.w3(32'hbb8c4749),
	.w4(32'h3b19cf8e),
	.w5(32'h3b712cb8),
	.w6(32'hbb65f681),
	.w7(32'h3a3fbfd9),
	.w8(32'h3afd7375),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba753cd5),
	.w1(32'h3a186201),
	.w2(32'hbb35fd77),
	.w3(32'h3b0a1f3c),
	.w4(32'hbb64a1ad),
	.w5(32'hbb5520fc),
	.w6(32'h3c5e037d),
	.w7(32'hbb105612),
	.w8(32'hbba8422a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2bc62),
	.w1(32'hbbd936b1),
	.w2(32'hbb4387b8),
	.w3(32'h3b3856fc),
	.w4(32'hbb17a4d5),
	.w5(32'h3b3325d0),
	.w6(32'hbb975fba),
	.w7(32'hbc0e751c),
	.w8(32'hbb674ec6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb576f83),
	.w1(32'hba82c320),
	.w2(32'hbb8df19e),
	.w3(32'h3bb9d1cd),
	.w4(32'hbba7f272),
	.w5(32'hbafbf54c),
	.w6(32'hba1b723d),
	.w7(32'h3b1360bb),
	.w8(32'hba1c853b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75b1d),
	.w1(32'hb8616528),
	.w2(32'hb8d5b2c2),
	.w3(32'hbb2add82),
	.w4(32'hbb17ecb9),
	.w5(32'hba980fb5),
	.w6(32'h3aa95ee2),
	.w7(32'hbb1ef56e),
	.w8(32'hbbd8c7fc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6cd9d),
	.w1(32'h3b976f00),
	.w2(32'hba0a4ebb),
	.w3(32'hbbe51cbd),
	.w4(32'hb7a9c96d),
	.w5(32'hbb20fc98),
	.w6(32'hbb9f20ba),
	.w7(32'hbb92d1cc),
	.w8(32'h3ab38a50),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891c4ed),
	.w1(32'hbb0df4a9),
	.w2(32'hbb43eccf),
	.w3(32'hb81fcedd),
	.w4(32'hbae061d8),
	.w5(32'hbb3ccb0a),
	.w6(32'h3a704f1a),
	.w7(32'hbb42f7da),
	.w8(32'hbb73e3c8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6378c),
	.w1(32'h3b37ce10),
	.w2(32'h3b1363cf),
	.w3(32'h3a0d7f54),
	.w4(32'h3bd6db56),
	.w5(32'h3c0879c4),
	.w6(32'hbb9f0ba6),
	.w7(32'h3b953e81),
	.w8(32'h3c3153dd),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe4f24),
	.w1(32'h3af85a4a),
	.w2(32'h3c03f493),
	.w3(32'h3c5346b4),
	.w4(32'h3b8fa989),
	.w5(32'h3c4161ea),
	.w6(32'h3c02b0a0),
	.w7(32'h3bc14907),
	.w8(32'h3c2dd7ea),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db1c7b),
	.w1(32'h3bb0b237),
	.w2(32'hb919dfe5),
	.w3(32'h39b538ca),
	.w4(32'h3b34697a),
	.w5(32'h3bd19016),
	.w6(32'h3b0a6abb),
	.w7(32'hbbf9e1c3),
	.w8(32'hbbc161ee),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba773f36),
	.w1(32'hba8911a8),
	.w2(32'hbb106856),
	.w3(32'h3b6f5688),
	.w4(32'hbaa33d90),
	.w5(32'hbb1ff9c6),
	.w6(32'h390ca50c),
	.w7(32'hba72d54e),
	.w8(32'h3b68760d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23dbb6),
	.w1(32'hb9ecee35),
	.w2(32'h3afdb07f),
	.w3(32'hbc27cec4),
	.w4(32'hbb6551bb),
	.w5(32'h3be0fe88),
	.w6(32'hbb97d89e),
	.w7(32'hbb8ec6df),
	.w8(32'hbab9bfac),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc54ff4),
	.w1(32'hbbf40096),
	.w2(32'hbbb69d32),
	.w3(32'h3ba6b199),
	.w4(32'hbc06e710),
	.w5(32'h3b5773cc),
	.w6(32'h3a770467),
	.w7(32'hbbf4c2ec),
	.w8(32'hba6247f9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf15eb3),
	.w1(32'h3a922d04),
	.w2(32'hbade088e),
	.w3(32'h3c3ad57b),
	.w4(32'h3b9b8c69),
	.w5(32'h3b6d1614),
	.w6(32'h3c1233c0),
	.w7(32'h3b9a7454),
	.w8(32'hb893b378),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54d84c),
	.w1(32'hb9896bf8),
	.w2(32'h3b210153),
	.w3(32'hb9aaed13),
	.w4(32'h3b9aa92e),
	.w5(32'h3ba66f94),
	.w6(32'hbb40ae18),
	.w7(32'h3ae1440c),
	.w8(32'h3a9ae05a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba456dff),
	.w1(32'h3873e7a4),
	.w2(32'h3b2c5d78),
	.w3(32'hbb831949),
	.w4(32'h3b0d4428),
	.w5(32'hbc6d5644),
	.w6(32'hb9878f8d),
	.w7(32'hb951e335),
	.w8(32'hbc391baa),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c075d0e),
	.w1(32'hbbf0dd03),
	.w2(32'hbbf5e16e),
	.w3(32'hb9095363),
	.w4(32'hbc08f737),
	.w5(32'hbba7cdb5),
	.w6(32'h3ab38051),
	.w7(32'hbc2299f6),
	.w8(32'hbc1a4474),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2303ec),
	.w1(32'h3b58982f),
	.w2(32'hbbf70841),
	.w3(32'hbc12fae2),
	.w4(32'h3bf30069),
	.w5(32'hb9d93b26),
	.w6(32'hbc5652fb),
	.w7(32'h3b7e8550),
	.w8(32'hba3ab7a3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3723b),
	.w1(32'hbc364f9a),
	.w2(32'hbc4ebd16),
	.w3(32'hbc27a31d),
	.w4(32'hbb45551f),
	.w5(32'hbbd93b98),
	.w6(32'hbb89327b),
	.w7(32'h3b264631),
	.w8(32'h3bf1d8fd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8398c6),
	.w1(32'h3b8825d3),
	.w2(32'h3afe8f49),
	.w3(32'hbb9ad5ed),
	.w4(32'h3b1ed957),
	.w5(32'hbadceab4),
	.w6(32'h3be49320),
	.w7(32'h3c013fbf),
	.w8(32'hbaced1ca),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b7976),
	.w1(32'hbab258ef),
	.w2(32'hba08bc55),
	.w3(32'hbc122ae7),
	.w4(32'h3a85f281),
	.w5(32'hbb3ddf2a),
	.w6(32'hbbe82f33),
	.w7(32'hbace65c6),
	.w8(32'hbaaa872b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d1e72),
	.w1(32'h3bb8fc2f),
	.w2(32'hba37e89d),
	.w3(32'hbb65fa2b),
	.w4(32'h3be80872),
	.w5(32'hbbddd55d),
	.w6(32'hbacbf0d6),
	.w7(32'h3b12c749),
	.w8(32'hbb967eca),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9851b0),
	.w1(32'h3b57891b),
	.w2(32'h3bc670f0),
	.w3(32'h3b81fb2c),
	.w4(32'h3b254fb5),
	.w5(32'h3c8af5bc),
	.w6(32'h3b2fe25e),
	.w7(32'h3ade300a),
	.w8(32'h3bf26662),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa193bc),
	.w1(32'hbb4cf07b),
	.w2(32'hbb911c5a),
	.w3(32'h3b973fbf),
	.w4(32'hbb6c2f6e),
	.w5(32'hb967a5b2),
	.w6(32'h3b1d7696),
	.w7(32'hb9b387b2),
	.w8(32'hba373afc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a098f3a),
	.w1(32'h3b92c4eb),
	.w2(32'h3b5ccbc2),
	.w3(32'h3ba732a3),
	.w4(32'h3c3e8e54),
	.w5(32'h3c946fe4),
	.w6(32'hba5a3ae5),
	.w7(32'h3b62367a),
	.w8(32'h3bb00d0d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15c911),
	.w1(32'hbbe7279b),
	.w2(32'hbb032fd9),
	.w3(32'h3c15f680),
	.w4(32'hbb3b1dae),
	.w5(32'h3bf5f2bf),
	.w6(32'h3baf1397),
	.w7(32'hbb925908),
	.w8(32'h3bc2bfdf),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3676c),
	.w1(32'hbb8e725f),
	.w2(32'hb8a46c74),
	.w3(32'h3b4526ab),
	.w4(32'hbb6b6f3e),
	.w5(32'hbbc2a9c9),
	.w6(32'h3c2c53a4),
	.w7(32'hbba5581f),
	.w8(32'hbb25514c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf19de),
	.w1(32'hbba8feab),
	.w2(32'hbab728f7),
	.w3(32'hbb6ee108),
	.w4(32'hbbb334f6),
	.w5(32'hbbd68a8b),
	.w6(32'h3a953a3f),
	.w7(32'hb9d202c8),
	.w8(32'hbaa60168),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a93ff),
	.w1(32'h3a541f6d),
	.w2(32'hba176805),
	.w3(32'h3b84251c),
	.w4(32'hbae5b60d),
	.w5(32'hba56f1ef),
	.w6(32'h3bee554d),
	.w7(32'hbb43e038),
	.w8(32'hbbc1c643),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule