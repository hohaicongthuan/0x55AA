module layer_8_featuremap_193(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeed560),
	.w1(32'hbb7628df),
	.w2(32'h3c18016d),
	.w3(32'hbc900890),
	.w4(32'hbbdd5fcd),
	.w5(32'h3b424beb),
	.w6(32'hbb08aec5),
	.w7(32'h3a631748),
	.w8(32'hba81ab40),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99a189),
	.w1(32'hbaa8f7c4),
	.w2(32'hba1245d5),
	.w3(32'hbbc13b3a),
	.w4(32'h3acb08ec),
	.w5(32'h3a47ae15),
	.w6(32'hba582a6d),
	.w7(32'h37505b67),
	.w8(32'h39c875a5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d239b6),
	.w1(32'hbb0d1d5c),
	.w2(32'hbb65ad0d),
	.w3(32'h3b59b880),
	.w4(32'h3b09423b),
	.w5(32'h394b55b7),
	.w6(32'h38430d3c),
	.w7(32'hbafaeea6),
	.w8(32'hbafc68fe),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be21297),
	.w1(32'h3c003b50),
	.w2(32'h3bb30df9),
	.w3(32'hba4553d9),
	.w4(32'h3ba4185d),
	.w5(32'h3bc77f29),
	.w6(32'hbb63f59d),
	.w7(32'hbb431197),
	.w8(32'hbabb7cd6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ba6d8),
	.w1(32'h370e9584),
	.w2(32'h3b634ecc),
	.w3(32'h3aa659ab),
	.w4(32'hb9c48639),
	.w5(32'h3b3f783c),
	.w6(32'h3a0fd118),
	.w7(32'h3b300269),
	.w8(32'h3b50e89b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becdf86),
	.w1(32'h3bfa447a),
	.w2(32'hbbcb3d81),
	.w3(32'h3bade110),
	.w4(32'h3bce62e7),
	.w5(32'hbbec0dbf),
	.w6(32'h3afed4a4),
	.w7(32'hbbcf0912),
	.w8(32'hbc0e7f0e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac50c17),
	.w1(32'h3a01e05a),
	.w2(32'h3a284a21),
	.w3(32'hbacdc0b6),
	.w4(32'hba390eef),
	.w5(32'hb9eb41b2),
	.w6(32'h3a710fc8),
	.w7(32'h3a243f29),
	.w8(32'h3b22b985),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c4f8),
	.w1(32'hbb5fe5cb),
	.w2(32'h3be9fd01),
	.w3(32'hbaaaa535),
	.w4(32'h3af6a1c8),
	.w5(32'h3c04ab17),
	.w6(32'h3b982b59),
	.w7(32'h3b9b309a),
	.w8(32'h3bff8f8d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba877cf5),
	.w1(32'hbba63300),
	.w2(32'h3b4ce263),
	.w3(32'h3b98b0c3),
	.w4(32'hbba1ba32),
	.w5(32'h3b6a4292),
	.w6(32'hbbf60be4),
	.w7(32'hbb8bb302),
	.w8(32'hba9e62a7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc105b00),
	.w1(32'h3c07a25e),
	.w2(32'h3c3d6fd4),
	.w3(32'h3a6c6940),
	.w4(32'h3c224933),
	.w5(32'h3c3721c6),
	.w6(32'h3b895a72),
	.w7(32'h3bd79194),
	.w8(32'h3c000209),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39d9a9),
	.w1(32'h3a4a4cf4),
	.w2(32'h3bd01b86),
	.w3(32'hbb5b8764),
	.w4(32'hbc5c6a6a),
	.w5(32'hba3f9e5a),
	.w6(32'hbb291c2d),
	.w7(32'hbb87501d),
	.w8(32'h3bba0037),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09c7f5),
	.w1(32'hbaa25ff9),
	.w2(32'h3c2bf3e2),
	.w3(32'hbc25e162),
	.w4(32'h3ca4bd12),
	.w5(32'h3cd78b03),
	.w6(32'h3ba99f48),
	.w7(32'h3bc41d64),
	.w8(32'h3c0f4cb4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2c09a),
	.w1(32'h3aa8697f),
	.w2(32'hbb31b3bb),
	.w3(32'h3d19e584),
	.w4(32'hba0a73e7),
	.w5(32'hbb7d03ab),
	.w6(32'hbac8cdb4),
	.w7(32'hbba3152f),
	.w8(32'hbb5c9d7e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba809d18),
	.w1(32'hbacb3afa),
	.w2(32'hbb75ec9d),
	.w3(32'h39ac1c0e),
	.w4(32'h3b9e3720),
	.w5(32'h3af53db3),
	.w6(32'hbb85f8e1),
	.w7(32'hbb3b64dd),
	.w8(32'h3b02b18e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97665c6),
	.w1(32'h3a07ef52),
	.w2(32'h3ad3174a),
	.w3(32'h3b1d4f02),
	.w4(32'h3ac6877b),
	.w5(32'h3b406439),
	.w6(32'h3aab1969),
	.w7(32'h3a80ff1a),
	.w8(32'h3b21532b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea258),
	.w1(32'hba52a95d),
	.w2(32'h3bb5d0ce),
	.w3(32'h3b91e34e),
	.w4(32'h39c69265),
	.w5(32'h3ba57331),
	.w6(32'hbbaf49d6),
	.w7(32'h3ae01351),
	.w8(32'hb954f187),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907631b),
	.w1(32'hbaaaf339),
	.w2(32'hbbac7a96),
	.w3(32'hbc02d87c),
	.w4(32'hbbb516a0),
	.w5(32'hbbe44c4a),
	.w6(32'hbc009363),
	.w7(32'hbc0af2bb),
	.w8(32'hbbe52b94),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb98053),
	.w1(32'hbb877a84),
	.w2(32'hbb3d2018),
	.w3(32'hbb2780d7),
	.w4(32'h3b314000),
	.w5(32'hba7ca02f),
	.w6(32'hbb2d7bfa),
	.w7(32'h3a1676da),
	.w8(32'h3bf41921),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc363a98),
	.w1(32'h3b89b240),
	.w2(32'h3c9bb3cc),
	.w3(32'hbbd0efa6),
	.w4(32'hbc666d6a),
	.w5(32'h3c612852),
	.w6(32'h3be5b3dc),
	.w7(32'h3c36cf92),
	.w8(32'h3c0069be),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02c964),
	.w1(32'hbb67b978),
	.w2(32'hbb93761e),
	.w3(32'hbace7280),
	.w4(32'h3aaf0175),
	.w5(32'hbb4e8ba1),
	.w6(32'hbbd1224c),
	.w7(32'hbb5c5bf0),
	.w8(32'hbb9cd01a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad96ee),
	.w1(32'hbac83ac6),
	.w2(32'hbb2b4696),
	.w3(32'h3ba1bf46),
	.w4(32'hbb929f1d),
	.w5(32'hbb6136a6),
	.w6(32'hbac22dc5),
	.w7(32'hbbc404fd),
	.w8(32'hbb052aff),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add4628),
	.w1(32'hbbfa581f),
	.w2(32'hbc2680b5),
	.w3(32'h3aca0946),
	.w4(32'hbbc9ed83),
	.w5(32'hbc48b515),
	.w6(32'hbbc30dba),
	.w7(32'hbc1b9543),
	.w8(32'hbbee75d9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a2059),
	.w1(32'hbb92cb28),
	.w2(32'h3d010d5d),
	.w3(32'hbc8599b7),
	.w4(32'hbc1ca8dc),
	.w5(32'h3ccae39e),
	.w6(32'hbc46e9b6),
	.w7(32'hba8b9532),
	.w8(32'h3c35e3d9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f23b8),
	.w1(32'hbc378bb1),
	.w2(32'hbc481ecf),
	.w3(32'h3c12bcdf),
	.w4(32'hbc1a6466),
	.w5(32'hbc176c22),
	.w6(32'hbbfcf0a6),
	.w7(32'hbc19db1a),
	.w8(32'hbc140546),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc243901),
	.w1(32'hbaf84c83),
	.w2(32'hbb8dfc8e),
	.w3(32'hbc2d2832),
	.w4(32'hbbee5ff3),
	.w5(32'hbc0ac774),
	.w6(32'hbb8474d5),
	.w7(32'hbbd85038),
	.w8(32'hbbf3a659),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc050ea8),
	.w1(32'hbc17b133),
	.w2(32'h3ab61a3f),
	.w3(32'hbc1694a7),
	.w4(32'hbb6ff490),
	.w5(32'hb9e6781b),
	.w6(32'hbb11d1d4),
	.w7(32'hb7c0b48c),
	.w8(32'h3a96ba34),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8748f),
	.w1(32'h3ba9f812),
	.w2(32'h3b97eb2b),
	.w3(32'hbabae88f),
	.w4(32'h3a88c283),
	.w5(32'h3bc97f12),
	.w6(32'h3b2e78b2),
	.w7(32'h3b72e43e),
	.w8(32'h3b197944),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf5034b),
	.w1(32'h3c18a7ec),
	.w2(32'h3c49b67d),
	.w3(32'hbbca190f),
	.w4(32'hbd1608ae),
	.w5(32'hbd0022c7),
	.w6(32'hbc059240),
	.w7(32'hbcfa1a61),
	.w8(32'hbc90382c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf01cc3),
	.w1(32'h39238952),
	.w2(32'hbbe6ed76),
	.w3(32'hbb995c86),
	.w4(32'h3b06de55),
	.w5(32'hbbdcc26d),
	.w6(32'h3bd98c9e),
	.w7(32'hbb93f193),
	.w8(32'h3b5f7ae6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae22f6e),
	.w1(32'hbaf1f284),
	.w2(32'h39aa70a4),
	.w3(32'h3a9d6100),
	.w4(32'h39aef9bb),
	.w5(32'h3c1fc880),
	.w6(32'h39953cfe),
	.w7(32'hba2624d5),
	.w8(32'h3a2af4f9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24d4dc),
	.w1(32'hbb94decf),
	.w2(32'hbb48fe09),
	.w3(32'h3cc37835),
	.w4(32'h3a9be883),
	.w5(32'h3b4c8c16),
	.w6(32'h3afcf9a5),
	.w7(32'h3923469b),
	.w8(32'h3aefb2e9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c604a),
	.w1(32'hbb6b308c),
	.w2(32'hbb0d0bec),
	.w3(32'h3b27f26d),
	.w4(32'hbbddbbc5),
	.w5(32'hbbad7dab),
	.w6(32'hba10dfca),
	.w7(32'hba15c004),
	.w8(32'hbc0a8749),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8ec69),
	.w1(32'hbaf43c74),
	.w2(32'h3b9360dd),
	.w3(32'hbbbf2835),
	.w4(32'h3a8ef66a),
	.w5(32'h3c6db4fc),
	.w6(32'hbb966876),
	.w7(32'hbb1ffeef),
	.w8(32'h3a146111),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066094),
	.w1(32'hba27c475),
	.w2(32'hbb50cadd),
	.w3(32'h3c26d8e9),
	.w4(32'hbae28933),
	.w5(32'hbab7c21a),
	.w6(32'h3abe4366),
	.w7(32'h3b2934d7),
	.w8(32'h39e344e0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe09c77),
	.w1(32'h3a8f65f8),
	.w2(32'hbba89da5),
	.w3(32'hbbaefb8c),
	.w4(32'h3bae205b),
	.w5(32'h3a9d9b85),
	.w6(32'hbb513742),
	.w7(32'hbaaf1aaf),
	.w8(32'hbb77533f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcebf44),
	.w1(32'hbc0539d7),
	.w2(32'h3a74345d),
	.w3(32'hb945b852),
	.w4(32'hbc2b9531),
	.w5(32'hbbc0009e),
	.w6(32'hbb4d00d9),
	.w7(32'hbaa4143d),
	.w8(32'h3aa418d7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab90092),
	.w1(32'h39c98ed5),
	.w2(32'h3b09a770),
	.w3(32'hb9c60d38),
	.w4(32'h3b276e00),
	.w5(32'h3bf76732),
	.w6(32'hb9886eee),
	.w7(32'h397dd9bf),
	.w8(32'hbb180a81),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a23ff),
	.w1(32'hbb9523a8),
	.w2(32'hbb38ee8c),
	.w3(32'h3b711960),
	.w4(32'hbb8c997f),
	.w5(32'hbb3671e9),
	.w6(32'hbb9b6a04),
	.w7(32'hbb815a57),
	.w8(32'hbbaf46f5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9571e),
	.w1(32'hbc13b175),
	.w2(32'hbb2ec0a6),
	.w3(32'hbb975e34),
	.w4(32'hbc167fed),
	.w5(32'hbb955fd6),
	.w6(32'hbc164027),
	.w7(32'hbabc9364),
	.w8(32'h3aec4c93),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b3aca),
	.w1(32'hb9a93bc1),
	.w2(32'hba3b38b7),
	.w3(32'h3af9b22d),
	.w4(32'hbb9e49bb),
	.w5(32'hbb4e4e81),
	.w6(32'h39ba907a),
	.w7(32'hb95bc0cc),
	.w8(32'hbb068684),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45abc7),
	.w1(32'h3c4d012f),
	.w2(32'h3c97e4b9),
	.w3(32'h3b0f2517),
	.w4(32'h3ca0a630),
	.w5(32'h3c8b2c22),
	.w6(32'h3c48e444),
	.w7(32'h3c347686),
	.w8(32'hb990b14c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a1359),
	.w1(32'hbc6d9831),
	.w2(32'h3b5cf9ce),
	.w3(32'h39901473),
	.w4(32'hbc2c34a5),
	.w5(32'h3c06b27e),
	.w6(32'hbc262069),
	.w7(32'h3a2960fc),
	.w8(32'hbbf5d12f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00b4f0),
	.w1(32'hba2f7f1f),
	.w2(32'hbba412f8),
	.w3(32'hbc0798e5),
	.w4(32'hbbd6eb5e),
	.w5(32'hbbdfcbfe),
	.w6(32'h3a84b778),
	.w7(32'hbb1275b6),
	.w8(32'hbae6460d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4e936),
	.w1(32'hbc1ba607),
	.w2(32'hba9a7baf),
	.w3(32'hbb17cc7d),
	.w4(32'hbc420731),
	.w5(32'hbbd98799),
	.w6(32'hbc210fab),
	.w7(32'hbbb03648),
	.w8(32'hbc07e183),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0a76b),
	.w1(32'hbb28793c),
	.w2(32'h3c4b3763),
	.w3(32'hbbf91253),
	.w4(32'hbbd6e7d3),
	.w5(32'h3c6a1d53),
	.w6(32'h39908f62),
	.w7(32'hba9bfebe),
	.w8(32'h399d6024),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f6e80),
	.w1(32'hbbdc8225),
	.w2(32'h39bb9d9f),
	.w3(32'hbbc0efff),
	.w4(32'hbb9622d7),
	.w5(32'h39203433),
	.w6(32'hbbb97027),
	.w7(32'hbb8bc700),
	.w8(32'h3b3b673f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0f5c),
	.w1(32'hbbca778f),
	.w2(32'hbb57a1f3),
	.w3(32'h3b860b0b),
	.w4(32'hbc1f08d0),
	.w5(32'hbbffd457),
	.w6(32'h39244bad),
	.w7(32'h3b5e9b5d),
	.w8(32'hbae77629),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc479c1a),
	.w1(32'hbc737772),
	.w2(32'hb88f4ccb),
	.w3(32'hbcb52120),
	.w4(32'hbccf6f2e),
	.w5(32'hbb6559e0),
	.w6(32'hbc4c7324),
	.w7(32'hbc11da83),
	.w8(32'hbbe6d814),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb978e),
	.w1(32'hbbb1b1f9),
	.w2(32'hbbbbebe8),
	.w3(32'hbc1c9da0),
	.w4(32'hbb9df677),
	.w5(32'hbb8d5a53),
	.w6(32'hbb3443d7),
	.w7(32'hbbe6a98b),
	.w8(32'hbc056310),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb741b0e),
	.w1(32'h3ae404ea),
	.w2(32'h3c006686),
	.w3(32'hbb47d018),
	.w4(32'h3bde27cf),
	.w5(32'h3c55b146),
	.w6(32'h3bd98644),
	.w7(32'h3a26ad16),
	.w8(32'h3b031786),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53aa6e),
	.w1(32'hbc1bdf7f),
	.w2(32'hbbf48f28),
	.w3(32'h3bc7517c),
	.w4(32'h3a94a859),
	.w5(32'hba116244),
	.w6(32'h3b445dfc),
	.w7(32'h3ac75304),
	.w8(32'hbbb3f032),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd89644),
	.w1(32'hbb2f853f),
	.w2(32'h3c17bb3b),
	.w3(32'hbbed9147),
	.w4(32'hbbb3c250),
	.w5(32'h3c7c4cab),
	.w6(32'h3b97806d),
	.w7(32'h3bdddd91),
	.w8(32'h3b7c0b26),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb587caf),
	.w1(32'h3b8f2ef2),
	.w2(32'h3c04b97f),
	.w3(32'hba9c890e),
	.w4(32'h3b7cd450),
	.w5(32'h3bf0b0c8),
	.w6(32'h3b94d776),
	.w7(32'h3b98d948),
	.w8(32'h3bf6b248),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515ad9),
	.w1(32'hbb8b20fc),
	.w2(32'h3c0df7e6),
	.w3(32'h3b5bda24),
	.w4(32'h3a8744cb),
	.w5(32'h3c145685),
	.w6(32'h3ac627c7),
	.w7(32'h3c0b3b51),
	.w8(32'h3bafbe65),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5d1a1),
	.w1(32'hbb80be74),
	.w2(32'h39acb6a9),
	.w3(32'h3b056958),
	.w4(32'hb8b9ee6a),
	.w5(32'h3b7b2284),
	.w6(32'hbbc25462),
	.w7(32'hb92000c3),
	.w8(32'h3aae48d1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0e5d8),
	.w1(32'hbcd2a24b),
	.w2(32'h3b7d10ef),
	.w3(32'hbc09d327),
	.w4(32'hbcd94ac2),
	.w5(32'hbb9f949b),
	.w6(32'hbc50788f),
	.w7(32'h3b10c11e),
	.w8(32'h3b9b7867),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fe78e),
	.w1(32'hbb4d01c5),
	.w2(32'hbba37121),
	.w3(32'hbba36241),
	.w4(32'h3a602df0),
	.w5(32'hbb67007a),
	.w6(32'hbbd0b357),
	.w7(32'hbc43088d),
	.w8(32'h3b0688b8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd10c9d),
	.w1(32'hba7f0b43),
	.w2(32'h3b96a350),
	.w3(32'hbbc0342d),
	.w4(32'hbb9e29d4),
	.w5(32'h3be2f24b),
	.w6(32'h3b0d86b4),
	.w7(32'hbab37574),
	.w8(32'hbadce9b1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb145743),
	.w1(32'hbb574818),
	.w2(32'h3b447d69),
	.w3(32'hbb80a12b),
	.w4(32'hbb8682fc),
	.w5(32'h3b988b3d),
	.w6(32'hbb4a9721),
	.w7(32'hbb8e77fc),
	.w8(32'h3c0c786f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00b0ac),
	.w1(32'hba9dd0a1),
	.w2(32'hbad8c2a9),
	.w3(32'h3c4d4b5e),
	.w4(32'hbb6bb0fa),
	.w5(32'hbb2b45d0),
	.w6(32'hbbe33d31),
	.w7(32'hbbc6aa60),
	.w8(32'hbb2b786a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfb3b0),
	.w1(32'h3b34d2fb),
	.w2(32'h3b2d707e),
	.w3(32'hbc44c112),
	.w4(32'hbaca9b17),
	.w5(32'hb853c2f8),
	.w6(32'h399c5abf),
	.w7(32'h3b910dde),
	.w8(32'h3baea171),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396992bb),
	.w1(32'hbb247918),
	.w2(32'hbb29b1e5),
	.w3(32'h3b170f21),
	.w4(32'h3baa021c),
	.w5(32'h3bf2b3a6),
	.w6(32'h3b69f1a3),
	.w7(32'h3b9ba390),
	.w8(32'h3a948938),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c1ee6),
	.w1(32'h3b3eea4f),
	.w2(32'h3bf63d5f),
	.w3(32'h3bb24215),
	.w4(32'h3b987761),
	.w5(32'h3bb26259),
	.w6(32'h3c3f3967),
	.w7(32'h3c36f192),
	.w8(32'h3bc8f5f9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2053a3),
	.w1(32'hbba501bd),
	.w2(32'h3b8fed97),
	.w3(32'hbb572279),
	.w4(32'h3c2dbc04),
	.w5(32'h3c977daf),
	.w6(32'hbb6d26b3),
	.w7(32'h3b413428),
	.w8(32'h3c842da3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85f8ab),
	.w1(32'hba054cf7),
	.w2(32'hbaf7ff55),
	.w3(32'h3d05181b),
	.w4(32'h3b57fa9a),
	.w5(32'h3ababa5d),
	.w6(32'h3b5aa6a4),
	.w7(32'h3a9b63fc),
	.w8(32'h3b74cde8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6eb03),
	.w1(32'hbb985f46),
	.w2(32'h388c2124),
	.w3(32'h3ab6afa1),
	.w4(32'hbbf7a58b),
	.w5(32'hbbd7a0fe),
	.w6(32'h393b8af0),
	.w7(32'hbb05793b),
	.w8(32'h38133f9c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30ac19),
	.w1(32'h3addc13f),
	.w2(32'h3b4e4a3d),
	.w3(32'hbbb101b9),
	.w4(32'h39bb5fa6),
	.w5(32'h3bbce269),
	.w6(32'hbb04cef4),
	.w7(32'h3b1c1368),
	.w8(32'hbaaadcc1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc263dd),
	.w1(32'hbc12bbcd),
	.w2(32'hbb2e04b5),
	.w3(32'hbbf88609),
	.w4(32'hbc0efea0),
	.w5(32'hbbd63dce),
	.w6(32'h3b076a08),
	.w7(32'h3b79781d),
	.w8(32'hbb9385a7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ddfb8),
	.w1(32'hbb659826),
	.w2(32'hbb93dd6b),
	.w3(32'hbb3cc913),
	.w4(32'hbc1b0f6b),
	.w5(32'hbbc9fffa),
	.w6(32'hbbba7e14),
	.w7(32'hbb9051bf),
	.w8(32'hbbfd55a9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae52c2),
	.w1(32'h3c5fbb96),
	.w2(32'h3caad279),
	.w3(32'hbc7ce9d8),
	.w4(32'hbc79b422),
	.w5(32'h3b5edd8e),
	.w6(32'hbba3b177),
	.w7(32'hbc3861a7),
	.w8(32'h3b62d5d0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a5cb4),
	.w1(32'h3bc8c524),
	.w2(32'hbc017c15),
	.w3(32'h39e3b5a8),
	.w4(32'h3a4b87c7),
	.w5(32'hbc69269c),
	.w6(32'h34507cab),
	.w7(32'hbc3c6a39),
	.w8(32'h3bf4312c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a1565),
	.w1(32'hbb503f3e),
	.w2(32'h3b53269c),
	.w3(32'h3acec4cc),
	.w4(32'h3b9c733b),
	.w5(32'h3a93edda),
	.w6(32'hbc0e30e2),
	.w7(32'hbbc9faec),
	.w8(32'h3a9c056a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48da26),
	.w1(32'hbc03455d),
	.w2(32'hbba0d556),
	.w3(32'h3b4aa713),
	.w4(32'hba9d2236),
	.w5(32'hbb623d43),
	.w6(32'hbc106a62),
	.w7(32'hbc31444e),
	.w8(32'hbbf971e4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f00f0),
	.w1(32'h3b98357b),
	.w2(32'h3c0b81d9),
	.w3(32'hb9f2ebf0),
	.w4(32'h3c2599db),
	.w5(32'h3b8f8d65),
	.w6(32'h3b493de0),
	.w7(32'h3ba7bc5c),
	.w8(32'h3be5f998),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee2493),
	.w1(32'h3b6fe8df),
	.w2(32'h3b919605),
	.w3(32'h3ae38249),
	.w4(32'h3be83a8e),
	.w5(32'h3bbab11c),
	.w6(32'hba3b0d21),
	.w7(32'h3b1abcc4),
	.w8(32'h3c4d4353),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19374d),
	.w1(32'hb9e50394),
	.w2(32'h3b811a2f),
	.w3(32'h3c529b27),
	.w4(32'h3b876a66),
	.w5(32'h3ba0a291),
	.w6(32'hbb3db835),
	.w7(32'hbb73f661),
	.w8(32'h3b2e94b5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b336766),
	.w1(32'hbb7d1e19),
	.w2(32'hbb6bc093),
	.w3(32'h3c0530b4),
	.w4(32'h3aa55333),
	.w5(32'h39d94902),
	.w6(32'hba7d121c),
	.w7(32'hba91aec0),
	.w8(32'h3b9aab53),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bbbc8),
	.w1(32'hba843a1a),
	.w2(32'h3c3b4e50),
	.w3(32'h3b854e64),
	.w4(32'hbc2442e9),
	.w5(32'h3bd1ac60),
	.w6(32'hbb24cf0c),
	.w7(32'h3b913103),
	.w8(32'h3b9238a8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc348c52),
	.w1(32'hbb5a758a),
	.w2(32'h3c29a729),
	.w3(32'hbb4eb688),
	.w4(32'hbbd038a1),
	.w5(32'h3b705f31),
	.w6(32'hbc3210e8),
	.w7(32'hbbbc9e36),
	.w8(32'h3b3b70ac),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be84ae4),
	.w1(32'hbbb21f42),
	.w2(32'h379f25ad),
	.w3(32'h3c01b877),
	.w4(32'hbbe065c8),
	.w5(32'hba6fd861),
	.w6(32'hbbe423c7),
	.w7(32'hbb1b4eaa),
	.w8(32'h3afc6db3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c8828),
	.w1(32'h3ba23ee1),
	.w2(32'h3bbffd15),
	.w3(32'h3ae95a81),
	.w4(32'h3b91e17a),
	.w5(32'hba8b2eec),
	.w6(32'h3aaae2e2),
	.w7(32'hbb77be1a),
	.w8(32'h3b5aebfc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b311d),
	.w1(32'hbb7b12f5),
	.w2(32'hbc0e32a5),
	.w3(32'h3c05fc03),
	.w4(32'hbbd01308),
	.w5(32'hbb89581a),
	.w6(32'hbc80b703),
	.w7(32'hbc896c6c),
	.w8(32'hbc13e6ac),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56f3b7),
	.w1(32'hbb03541d),
	.w2(32'h3b855959),
	.w3(32'hbc6cbbe6),
	.w4(32'h3b841f79),
	.w5(32'h3c24553a),
	.w6(32'hb81efb84),
	.w7(32'hba4ebe71),
	.w8(32'h3b58be05),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7525e4),
	.w1(32'h3c01bbc0),
	.w2(32'h3c090e19),
	.w3(32'h3c9d07cc),
	.w4(32'h3c871184),
	.w5(32'h3c15664c),
	.w6(32'h3b9dd30a),
	.w7(32'h3c995f0d),
	.w8(32'hbb8073ce),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb049c7),
	.w1(32'h38b79660),
	.w2(32'h3cbc4eb8),
	.w3(32'hbb939651),
	.w4(32'hbb5e0d84),
	.w5(32'h3c55028d),
	.w6(32'h3bbce9e7),
	.w7(32'h3bc77588),
	.w8(32'h3c2ec5a0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c345c0b),
	.w1(32'h3c6cb63c),
	.w2(32'h3c2c2901),
	.w3(32'h3c4ff70e),
	.w4(32'h3c11c82f),
	.w5(32'h3be0d08d),
	.w6(32'h38e3f740),
	.w7(32'h3a843511),
	.w8(32'h3b5ebed3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aac0c),
	.w1(32'h3b85a8be),
	.w2(32'h3b89a0a6),
	.w3(32'hbbf0b517),
	.w4(32'h39272b51),
	.w5(32'h3ae2b68c),
	.w6(32'hbb1d8380),
	.w7(32'hbb8797b5),
	.w8(32'h3a985539),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10a80a),
	.w1(32'hb96c0bda),
	.w2(32'h3b30083d),
	.w3(32'h3b814513),
	.w4(32'hba69f538),
	.w5(32'h3a7bbec3),
	.w6(32'hbbe4078a),
	.w7(32'hbc09f558),
	.w8(32'hbc0383bc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b0698),
	.w1(32'h3b122e35),
	.w2(32'h3b407f33),
	.w3(32'h3a443a39),
	.w4(32'h3a981035),
	.w5(32'h3bb2d5df),
	.w6(32'hbb85a2a2),
	.w7(32'hbbc80d26),
	.w8(32'hbbf5e747),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07f237),
	.w1(32'hbbe0492e),
	.w2(32'hbb92ea5f),
	.w3(32'h3b2b25c4),
	.w4(32'h3ae3d6ae),
	.w5(32'h3beb2817),
	.w6(32'hbb3cdfaa),
	.w7(32'hbba046cb),
	.w8(32'h3a0e9289),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d05da),
	.w1(32'hbaf0eddf),
	.w2(32'hbaac0b90),
	.w3(32'h3c287e24),
	.w4(32'h3b719e9e),
	.w5(32'h3b5971ab),
	.w6(32'hbb7bf7f5),
	.w7(32'hbbad18af),
	.w8(32'hbb94866a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb762a0f),
	.w1(32'hbb3e2a64),
	.w2(32'hbb88b2da),
	.w3(32'h3b64e3a7),
	.w4(32'hbb9ca742),
	.w5(32'hbb8cfe61),
	.w6(32'hbaeb82a0),
	.w7(32'hbab3120e),
	.w8(32'hbbc0ba07),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1664a0),
	.w1(32'h3aea2041),
	.w2(32'hbb0d1965),
	.w3(32'hbba4579a),
	.w4(32'h3b346096),
	.w5(32'h3a97dad2),
	.w6(32'hbb2b6740),
	.w7(32'h3a36d5e0),
	.w8(32'h3ae01c17),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10450b),
	.w1(32'hbb420fe1),
	.w2(32'hb95b2be7),
	.w3(32'h3b75cd1a),
	.w4(32'hbb49adbe),
	.w5(32'hbb008dc3),
	.w6(32'hbb162595),
	.w7(32'hba3cef1b),
	.w8(32'hba2d62ee),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda7de1),
	.w1(32'hbbe3ae96),
	.w2(32'hbb828cfd),
	.w3(32'hbb91836a),
	.w4(32'hbb9cc27b),
	.w5(32'hbb58c4e6),
	.w6(32'hbb07fa88),
	.w7(32'hbb5f41c1),
	.w8(32'hbc1af563),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a4ccc),
	.w1(32'hbbd3242f),
	.w2(32'h3b61679a),
	.w3(32'hbc318d2f),
	.w4(32'hbbf610de),
	.w5(32'hb9c720a5),
	.w6(32'hbb43a6b4),
	.w7(32'h37b38971),
	.w8(32'h3a6be8cc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9871ec),
	.w1(32'h39787932),
	.w2(32'h3b8944f9),
	.w3(32'hbbacff69),
	.w4(32'h3bb8d2e3),
	.w5(32'h3be6430c),
	.w6(32'h3ab92443),
	.w7(32'hb99ff27a),
	.w8(32'h3b0fbc9c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af815ab),
	.w1(32'hbbf4d2d8),
	.w2(32'hbaac80eb),
	.w3(32'h3b30eff9),
	.w4(32'hbb1b4bc2),
	.w5(32'hb9e2f279),
	.w6(32'hbc0ee541),
	.w7(32'hba4e5a4e),
	.w8(32'h3c03b8fc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cfc21),
	.w1(32'hbbf8bb81),
	.w2(32'hbc0d8ed0),
	.w3(32'h3c3b2bfe),
	.w4(32'hbc1f4236),
	.w5(32'hbc4dd10b),
	.w6(32'hbc26100b),
	.w7(32'hbc1dce63),
	.w8(32'hb9e04a5f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbe73d),
	.w1(32'h3c36cba4),
	.w2(32'h3b852acf),
	.w3(32'h3ab18e97),
	.w4(32'h3b0c5df1),
	.w5(32'h3b6de6ed),
	.w6(32'h3b1f536c),
	.w7(32'h3ae8a062),
	.w8(32'h3b6856f1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b6c16),
	.w1(32'h3ae62834),
	.w2(32'h3a8870e8),
	.w3(32'h3ae138e8),
	.w4(32'hbaedf12a),
	.w5(32'hbadfd420),
	.w6(32'h3b2ae15f),
	.w7(32'hbb4efaab),
	.w8(32'hb98538fb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c1bdc),
	.w1(32'hbb5470e0),
	.w2(32'hbb794eb7),
	.w3(32'h3ad25a4c),
	.w4(32'hba2fadd2),
	.w5(32'hbbd1665e),
	.w6(32'hbbfc1520),
	.w7(32'hbc07147e),
	.w8(32'hbb50d208),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8236),
	.w1(32'hbc03c691),
	.w2(32'hbc0164dd),
	.w3(32'hbb5f0a7e),
	.w4(32'hbc4ce20d),
	.w5(32'hbc33e78a),
	.w6(32'hbc4aaea0),
	.w7(32'hbc17347c),
	.w8(32'hbc0d97e3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31215a),
	.w1(32'hbb555e8b),
	.w2(32'hbbdb91de),
	.w3(32'hbbd686dc),
	.w4(32'h3916d87a),
	.w5(32'hbbbd6954),
	.w6(32'hbbbe09c1),
	.w7(32'hbb97d8e1),
	.w8(32'h3a04732d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaff50c),
	.w1(32'hbba85846),
	.w2(32'h38a2f2fd),
	.w3(32'h3b21ea6d),
	.w4(32'hbb7fe346),
	.w5(32'h3bf80162),
	.w6(32'hbbc0bd6a),
	.w7(32'hbb9d3195),
	.w8(32'h3c3337e0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde6374),
	.w1(32'h3b2946ab),
	.w2(32'h3be7c746),
	.w3(32'h3b33d971),
	.w4(32'hbbd5eddc),
	.w5(32'h3a798723),
	.w6(32'h3b0c9563),
	.w7(32'hbb981309),
	.w8(32'h3bd35006),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab77205),
	.w1(32'h3a8c5a45),
	.w2(32'h3bd9ea58),
	.w3(32'h3a537e45),
	.w4(32'hbaa99c14),
	.w5(32'h3abd4af7),
	.w6(32'hbc057036),
	.w7(32'hbbbbb1f3),
	.w8(32'hbb95022a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0eb2f),
	.w1(32'hba17f23a),
	.w2(32'h3aefe8e2),
	.w3(32'hbb477674),
	.w4(32'h3b4d173a),
	.w5(32'h3c246ceb),
	.w6(32'hbb26f8ff),
	.w7(32'hba2158b8),
	.w8(32'hbbabdec9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae0d9d),
	.w1(32'hb9cebf70),
	.w2(32'hbb4aa451),
	.w3(32'h3c44c2e1),
	.w4(32'hba118abf),
	.w5(32'hbbb0b437),
	.w6(32'h3b993682),
	.w7(32'h3906d604),
	.w8(32'h3b5a8320),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0c7c5),
	.w1(32'hbb15ab5e),
	.w2(32'hba91f62b),
	.w3(32'hba637e45),
	.w4(32'hbb286712),
	.w5(32'hba999c0c),
	.w6(32'hbb2d1b79),
	.w7(32'hbb1ca76e),
	.w8(32'hba667306),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd41516),
	.w1(32'hbc35f4d9),
	.w2(32'hbc48623f),
	.w3(32'hbb7904ea),
	.w4(32'hbc422fc0),
	.w5(32'hbc44e9db),
	.w6(32'hbbbc91ae),
	.w7(32'hbbb4b6e5),
	.w8(32'hbc259f46),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42cfae),
	.w1(32'hbbd0ab69),
	.w2(32'hbc22d218),
	.w3(32'hbbfa70c9),
	.w4(32'hbba83335),
	.w5(32'hbc0e6f57),
	.w6(32'hbb609c8c),
	.w7(32'hbbd94a82),
	.w8(32'hbbdb2e6a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb881509),
	.w1(32'hbbfeccbd),
	.w2(32'hbc311cd9),
	.w3(32'hbb3cefb7),
	.w4(32'hbc1d774e),
	.w5(32'hbc04ae7e),
	.w6(32'hbc2c38f1),
	.w7(32'hbb8e8e70),
	.w8(32'hbc408f6b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bae95),
	.w1(32'h399925ae),
	.w2(32'h3a2cf7e8),
	.w3(32'hbc606e81),
	.w4(32'h3ab159f9),
	.w5(32'hbb9109e4),
	.w6(32'hbbe6631e),
	.w7(32'hbc295408),
	.w8(32'hbb8988a2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841c48),
	.w1(32'hbb424077),
	.w2(32'hb9cc60e7),
	.w3(32'hbba65629),
	.w4(32'h3a56bbe9),
	.w5(32'h3bf2834f),
	.w6(32'hbabf9e5a),
	.w7(32'h398aea06),
	.w8(32'hbbf1581a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d239a),
	.w1(32'hba872493),
	.w2(32'hba80c4f4),
	.w3(32'hbb1b8917),
	.w4(32'hba075c55),
	.w5(32'hba6846df),
	.w6(32'h3a6c6fef),
	.w7(32'hb969e2e9),
	.w8(32'hba1036c8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1c20b),
	.w1(32'h3ba4c10a),
	.w2(32'hbafeb72a),
	.w3(32'hbb13fe42),
	.w4(32'hb8946680),
	.w5(32'hbb062089),
	.w6(32'h3bb2520c),
	.w7(32'hbb160b6c),
	.w8(32'h3c0cfda7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda7698),
	.w1(32'hbab8dc1b),
	.w2(32'hbb6ed5b6),
	.w3(32'h3be24796),
	.w4(32'hbbb33191),
	.w5(32'hbbec87bc),
	.w6(32'h3aaa2acc),
	.w7(32'hbb40cdb7),
	.w8(32'hbb67929f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0fd2f),
	.w1(32'hb8d836a8),
	.w2(32'h3bb15c27),
	.w3(32'hbc02e663),
	.w4(32'h3b19d1ce),
	.w5(32'h3b94e7ac),
	.w6(32'h399adfc0),
	.w7(32'h3b046847),
	.w8(32'hbb1b941b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b609daf),
	.w1(32'hbb06f318),
	.w2(32'h3ab09360),
	.w3(32'hbaae7f64),
	.w4(32'hb7dfb28b),
	.w5(32'h3b19590e),
	.w6(32'hb764bb94),
	.w7(32'h3abbc880),
	.w8(32'h39cb68dc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ec0c3),
	.w1(32'hbc05f623),
	.w2(32'hbb93f93d),
	.w3(32'h3bd546b8),
	.w4(32'hbba4b527),
	.w5(32'hbb9feb8f),
	.w6(32'hbc5f9710),
	.w7(32'hbc1b7eb1),
	.w8(32'hbc144eef),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41a4f1),
	.w1(32'h397f2b0c),
	.w2(32'h3bbef015),
	.w3(32'hbc7cf2a7),
	.w4(32'h3b72f4ba),
	.w5(32'h3c065104),
	.w6(32'hbacf1cd0),
	.w7(32'h3ab7099f),
	.w8(32'hbb9ba208),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070b40),
	.w1(32'hbb0bd763),
	.w2(32'hba03834e),
	.w3(32'h39b3b76b),
	.w4(32'hba536594),
	.w5(32'hb96e515d),
	.w6(32'hba6c467e),
	.w7(32'h3a117a72),
	.w8(32'h3b16ae59),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e110e),
	.w1(32'hbc2d1987),
	.w2(32'hbc194dd9),
	.w3(32'h3b533b82),
	.w4(32'hbc2b413c),
	.w5(32'hbc154382),
	.w6(32'hbbe1d66d),
	.w7(32'hbbe06552),
	.w8(32'hbbefe5a0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2365c2),
	.w1(32'h3abeeb32),
	.w2(32'hbad48b68),
	.w3(32'hbc205b01),
	.w4(32'h3bca03c7),
	.w5(32'h3b984ed5),
	.w6(32'hba393970),
	.w7(32'hbb3e1f4f),
	.w8(32'hbb394ff4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fdcee),
	.w1(32'hbc5ad822),
	.w2(32'hbc5daad0),
	.w3(32'h3ba50fa5),
	.w4(32'hbc5192af),
	.w5(32'hbc6650d0),
	.w6(32'hbbfb9070),
	.w7(32'hbc3e8dbf),
	.w8(32'hbba49ea9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4035f0),
	.w1(32'hb99163e1),
	.w2(32'h3aee43dd),
	.w3(32'hbc6e835a),
	.w4(32'hba28145c),
	.w5(32'h3a3dbebb),
	.w6(32'hbb2baa31),
	.w7(32'hbab05e49),
	.w8(32'hbb37d06b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a98a),
	.w1(32'h3c04446d),
	.w2(32'h3cc22836),
	.w3(32'hbbf8b879),
	.w4(32'hbb2baa36),
	.w5(32'h3b649541),
	.w6(32'h3c0a5722),
	.w7(32'h3ca6ccb7),
	.w8(32'h3cd46569),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule