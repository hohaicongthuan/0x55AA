module layer_10_featuremap_309(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18977f),
	.w1(32'hb8a2cedd),
	.w2(32'hb9dbe610),
	.w3(32'hb800c265),
	.w4(32'hba4eb061),
	.w5(32'h3a4d1de2),
	.w6(32'h3ab894a0),
	.w7(32'hb635ccb7),
	.w8(32'h3a04bb1a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b827b7f),
	.w1(32'h3aa1b552),
	.w2(32'hbb061770),
	.w3(32'h3bb1c226),
	.w4(32'hba546025),
	.w5(32'hbb041852),
	.w6(32'h3bb5cef3),
	.w7(32'hba4b7624),
	.w8(32'hbb4fd12f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90519b1),
	.w1(32'hb96f4c1c),
	.w2(32'hbae73ca2),
	.w3(32'h3a74a3c9),
	.w4(32'hba703da8),
	.w5(32'hb89cc376),
	.w6(32'h3b5178bd),
	.w7(32'h392e094a),
	.w8(32'h392b7d59),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0571c4),
	.w1(32'h3b185d34),
	.w2(32'h3bb03885),
	.w3(32'hbb45e67c),
	.w4(32'hb8bbb0e0),
	.w5(32'h3a0310ba),
	.w6(32'hbad32675),
	.w7(32'h3b5066dd),
	.w8(32'h3ab4700a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba972f68),
	.w1(32'hbb112bb1),
	.w2(32'hba144a49),
	.w3(32'hba016c84),
	.w4(32'h3ab5b18d),
	.w5(32'h3a28be51),
	.w6(32'hbb631ef1),
	.w7(32'hba89d735),
	.w8(32'h3a8efc68),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e45b92),
	.w1(32'hba1115b8),
	.w2(32'h391f28a3),
	.w3(32'h3aaad951),
	.w4(32'h3a9e1610),
	.w5(32'h3b352bf2),
	.w6(32'h3a4c4bc6),
	.w7(32'h3a0c1922),
	.w8(32'h3b0995ec),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b910b71),
	.w1(32'h3c6080f7),
	.w2(32'h3c845e08),
	.w3(32'h3ad1a590),
	.w4(32'h3beb0f3b),
	.w5(32'h3b81ecc3),
	.w6(32'h3c19ecb3),
	.w7(32'h3c330965),
	.w8(32'h3bca6f9a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fc54f),
	.w1(32'h3a862a24),
	.w2(32'hbc22cc19),
	.w3(32'hbc430db9),
	.w4(32'hbc325791),
	.w5(32'hbc12d537),
	.w6(32'hbc4016f6),
	.w7(32'hbbae8ef8),
	.w8(32'hbb9b77e0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9b68b),
	.w1(32'hba43b039),
	.w2(32'hbaa7440a),
	.w3(32'hba14c77a),
	.w4(32'h3a0cb49a),
	.w5(32'hb98dfe2d),
	.w6(32'h38aa3ad8),
	.w7(32'hb96a5699),
	.w8(32'hba08e593),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d0cd),
	.w1(32'hb9785b81),
	.w2(32'h3a2ef2f0),
	.w3(32'hbb8c4138),
	.w4(32'hbae4601e),
	.w5(32'hbb860a26),
	.w6(32'h3c1b8c0c),
	.w7(32'h3c0a58f5),
	.w8(32'h3bb72e4a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6e6f4),
	.w1(32'hba8ac7c1),
	.w2(32'hb658d5c0),
	.w3(32'hb9bb3b50),
	.w4(32'h39341e48),
	.w5(32'h3b0aac41),
	.w6(32'hbabbe7c5),
	.w7(32'h39433a6b),
	.w8(32'h3a95101f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4886dc),
	.w1(32'h3c79f1e8),
	.w2(32'h3c8c2116),
	.w3(32'h3a81ee09),
	.w4(32'h3bfbe2e6),
	.w5(32'h3b338407),
	.w6(32'h3c2d927b),
	.w7(32'h3c82a8e9),
	.w8(32'h3c426b00),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd780a0),
	.w1(32'hb957c76d),
	.w2(32'hba0c6a6b),
	.w3(32'hbbbf24b0),
	.w4(32'hbb02adc9),
	.w5(32'hbb3dafb0),
	.w6(32'h3c0d6503),
	.w7(32'h3c149042),
	.w8(32'h3b904a85),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9231605),
	.w1(32'h3a952752),
	.w2(32'hbb498b20),
	.w3(32'hbb7ef54c),
	.w4(32'hbb77a72a),
	.w5(32'hbb9ac19c),
	.w6(32'hb963ad7e),
	.w7(32'hbb1ef35c),
	.w8(32'hbb3b0e36),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21c97f),
	.w1(32'hbb8262ee),
	.w2(32'hbbd567ed),
	.w3(32'h3badd8df),
	.w4(32'h3b0aed91),
	.w5(32'hbb842cff),
	.w6(32'h3b87ab3b),
	.w7(32'h3b087969),
	.w8(32'hbb2d3150),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97a292),
	.w1(32'hba4555d1),
	.w2(32'hbbf0f1d9),
	.w3(32'hbb4c2b09),
	.w4(32'hbb91d47b),
	.w5(32'hbbc7e5d9),
	.w6(32'h3baa7c63),
	.w7(32'h3ad0273b),
	.w8(32'h3b3ea750),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaa98f),
	.w1(32'h394f6641),
	.w2(32'h39cdedcb),
	.w3(32'h3b19e5df),
	.w4(32'h3b086e59),
	.w5(32'h387f3f2b),
	.w6(32'h3aeb5bb6),
	.w7(32'h3ad969d5),
	.w8(32'h3887ed54),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc923f8c),
	.w1(32'hbc1130e4),
	.w2(32'hbc219f4f),
	.w3(32'hbb8f0c66),
	.w4(32'hbb1774c5),
	.w5(32'hbc2e529a),
	.w6(32'h3c06194f),
	.w7(32'h3bc63123),
	.w8(32'h3b065f7a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d07f2),
	.w1(32'hbae41c87),
	.w2(32'hba9c7f9c),
	.w3(32'hbb9aa678),
	.w4(32'h394f5832),
	.w5(32'hbb0141de),
	.w6(32'h3b97f714),
	.w7(32'h3c1570a5),
	.w8(32'h3b991b6b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb809b693),
	.w1(32'hba8b2c3b),
	.w2(32'hbac022e8),
	.w3(32'h39e0a18a),
	.w4(32'hba879548),
	.w5(32'hbaa9fdf0),
	.w6(32'hba67c4d4),
	.w7(32'hbac6a774),
	.w8(32'hba3a88c0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64ee7b),
	.w1(32'hbb52c712),
	.w2(32'hbb13f0cc),
	.w3(32'hbae61aa8),
	.w4(32'hba947563),
	.w5(32'h3ab8bdb7),
	.w6(32'hba7341fb),
	.w7(32'hb9b51782),
	.w8(32'h3b023b8f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf40bc5),
	.w1(32'h3b8ff999),
	.w2(32'h3ae9ccbf),
	.w3(32'h3b9e1e22),
	.w4(32'h3b3bb9bc),
	.w5(32'h3a0845cc),
	.w6(32'h3adebfe4),
	.w7(32'h3b03587f),
	.w8(32'hba8d31ee),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f5906),
	.w1(32'hbb81f3c1),
	.w2(32'hbc284933),
	.w3(32'hbb93b62f),
	.w4(32'h3c5681cf),
	.w5(32'h3a8d1f4c),
	.w6(32'h3c703963),
	.w7(32'h3c88c046),
	.w8(32'h3c1fbd8f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dd0ee),
	.w1(32'hbb4cc200),
	.w2(32'hbac066bc),
	.w3(32'h3b4d706d),
	.w4(32'h3b272ded),
	.w5(32'h3a9d4f41),
	.w6(32'h3c465cff),
	.w7(32'h3bfc36b0),
	.w8(32'h3be92ee8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9051f3),
	.w1(32'h3baa813b),
	.w2(32'hbb62c108),
	.w3(32'h3c8d05c5),
	.w4(32'h3b592014),
	.w5(32'hbb5244e5),
	.w6(32'h3c6463f1),
	.w7(32'h3b544fa4),
	.w8(32'hba4ff174),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23213e),
	.w1(32'h39ff3abe),
	.w2(32'h3ac33cc9),
	.w3(32'h3aecdac1),
	.w4(32'h3b48b9c9),
	.w5(32'h3a9f1cf2),
	.w6(32'h3ade8870),
	.w7(32'h3af0b529),
	.w8(32'h3b1e9d10),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cdbb90),
	.w1(32'h3a848567),
	.w2(32'h3b10363f),
	.w3(32'h3acc1da0),
	.w4(32'h3ac6c69f),
	.w5(32'h3914e238),
	.w6(32'h3b23ea57),
	.w7(32'h3b1ef1c8),
	.w8(32'h3ab5760a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bfa07),
	.w1(32'h3c15004a),
	.w2(32'h39938303),
	.w3(32'h3c1e15d9),
	.w4(32'hb9d4e46c),
	.w5(32'hbb24a5c6),
	.w6(32'h3bc0b63f),
	.w7(32'hbc094743),
	.w8(32'hba3a1888),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61c517),
	.w1(32'h3ac14059),
	.w2(32'h3996cf0b),
	.w3(32'h3b7e6676),
	.w4(32'h3b115ea3),
	.w5(32'h38ad3754),
	.w6(32'hb96446ac),
	.w7(32'h3a99e160),
	.w8(32'h3a63c584),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ecf5b),
	.w1(32'h3c461930),
	.w2(32'h3bf0d5d6),
	.w3(32'h3c57ff30),
	.w4(32'h3c0868bf),
	.w5(32'h3b1aaca4),
	.w6(32'h3c745806),
	.w7(32'h3b8180c2),
	.w8(32'h3b6c8fb5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b012c50),
	.w1(32'h3b4bb902),
	.w2(32'h3b22d574),
	.w3(32'h395491e8),
	.w4(32'hba8d728f),
	.w5(32'h3abbd188),
	.w6(32'h3b2d810d),
	.w7(32'h3a1b6a75),
	.w8(32'h3aa7a7d2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cd5f1),
	.w1(32'hbae77693),
	.w2(32'h392fd4ba),
	.w3(32'h3acabb5b),
	.w4(32'h3ac712ab),
	.w5(32'h37984c64),
	.w6(32'h39c79a53),
	.w7(32'h39b156ce),
	.w8(32'h3b0389fc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8cefc),
	.w1(32'hba293f14),
	.w2(32'hba6310df),
	.w3(32'hbb7af755),
	.w4(32'hbb80b428),
	.w5(32'hbb735fd7),
	.w6(32'h3b839e47),
	.w7(32'h3b3cf992),
	.w8(32'h3a0da54d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60a037),
	.w1(32'hb9754e2e),
	.w2(32'hbb25345a),
	.w3(32'h3af6d30a),
	.w4(32'hba891f0f),
	.w5(32'hba225e19),
	.w6(32'h3a604bfe),
	.w7(32'hbb0c5b6f),
	.w8(32'h3981e121),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6c903),
	.w1(32'h3aae589a),
	.w2(32'h3b2cdc6c),
	.w3(32'hbb14a33c),
	.w4(32'hbad03231),
	.w5(32'h39baf335),
	.w6(32'hbb177907),
	.w7(32'hba9c1d59),
	.w8(32'hba9a42fe),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96c2d0),
	.w1(32'hba882b7b),
	.w2(32'h3ac00e8e),
	.w3(32'hbb9d1ea1),
	.w4(32'h39cab6f5),
	.w5(32'hba957088),
	.w6(32'hb8d9de28),
	.w7(32'h3b79859a),
	.w8(32'h3ae0ee4d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b531b),
	.w1(32'hbc25839e),
	.w2(32'h3b38398e),
	.w3(32'hbb2175be),
	.w4(32'hbb3218d4),
	.w5(32'h3c6fdbf2),
	.w6(32'h3c27e86c),
	.w7(32'h3cb43a2f),
	.w8(32'h3ca9f746),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a3dca),
	.w1(32'h3b72910c),
	.w2(32'hb9dcf95e),
	.w3(32'h3ca1c93c),
	.w4(32'h3c3a4300),
	.w5(32'h3b89338c),
	.w6(32'h3c3f509a),
	.w7(32'h3bc1a80c),
	.w8(32'hbabefe33),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccd407),
	.w1(32'h3c99c4b2),
	.w2(32'h3c27fd93),
	.w3(32'h3ca6aa53),
	.w4(32'h3c7698e2),
	.w5(32'h3be3d6a4),
	.w6(32'h3c3f0e13),
	.w7(32'h3bb3e69d),
	.w8(32'h3b2ea06d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e7c81),
	.w1(32'hba8ea365),
	.w2(32'hbb40785a),
	.w3(32'h3b11c218),
	.w4(32'hba109d3d),
	.w5(32'h38beec41),
	.w6(32'h398bd875),
	.w7(32'hbae0a5fb),
	.w8(32'h38e8750b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa27b19),
	.w1(32'h375497fd),
	.w2(32'h3ab6c8aa),
	.w3(32'hbae8fc87),
	.w4(32'hba3b6324),
	.w5(32'h3b199139),
	.w6(32'h3a240d73),
	.w7(32'h39ee7740),
	.w8(32'h3b116518),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae799b2),
	.w1(32'h3a84a16a),
	.w2(32'h3af1c9df),
	.w3(32'h3b8c02f3),
	.w4(32'h3b4f12be),
	.w5(32'hbb0cb33a),
	.w6(32'h3b2f047a),
	.w7(32'h3b1ebe7c),
	.w8(32'hbb029ed0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2244fe),
	.w1(32'hbb039710),
	.w2(32'h38d9ffa1),
	.w3(32'hbb08e707),
	.w4(32'h3b0e6f44),
	.w5(32'hbb3e2ed9),
	.w6(32'hba946e80),
	.w7(32'h3b235e18),
	.w8(32'hba61d1a5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46f08f),
	.w1(32'hbb2498df),
	.w2(32'hbb8d248a),
	.w3(32'hbc5db69c),
	.w4(32'h3ada46e0),
	.w5(32'hbbacebd7),
	.w6(32'h3c2785fb),
	.w7(32'h3c4f54e6),
	.w8(32'h3bd55ad1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba919c93),
	.w1(32'hba7f6dc3),
	.w2(32'hbb113614),
	.w3(32'h3b99dbfc),
	.w4(32'h3b5ad5e3),
	.w5(32'h3b17df60),
	.w6(32'h3c2402f9),
	.w7(32'h3c05b4a7),
	.w8(32'h3bc43fc6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1967de),
	.w1(32'hbb8c83ca),
	.w2(32'hba51fc07),
	.w3(32'h3b8424b0),
	.w4(32'h3b14544c),
	.w5(32'h3a7ab7e5),
	.w6(32'h3c50ddc7),
	.w7(32'h3c2f2991),
	.w8(32'h3c0538bd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace8ed3),
	.w1(32'h3b93ac3b),
	.w2(32'h3a2a2031),
	.w3(32'h3aa8f464),
	.w4(32'h3ab7eaed),
	.w5(32'h3a9a6882),
	.w6(32'h3bce14d7),
	.w7(32'h3b95d8fa),
	.w8(32'h3b8b0a56),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02e679),
	.w1(32'h3b0e8b9f),
	.w2(32'h3a89860d),
	.w3(32'hbc11262a),
	.w4(32'h3b8b28f8),
	.w5(32'hbb8db0bf),
	.w6(32'h3c1bcddb),
	.w7(32'h3cbeb47c),
	.w8(32'h3c2b8cd9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cbc54),
	.w1(32'hbb155a88),
	.w2(32'hbb08ee90),
	.w3(32'hbb788d13),
	.w4(32'hbb4e738b),
	.w5(32'h3a877af4),
	.w6(32'hbb224f32),
	.w7(32'hbab1aed8),
	.w8(32'h395163f2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82c999),
	.w1(32'hba3694b8),
	.w2(32'hba23715f),
	.w3(32'hb96904ff),
	.w4(32'h39a06059),
	.w5(32'hbaf8bf33),
	.w6(32'hba722b30),
	.w7(32'hbaec5400),
	.w8(32'hbb3a94d8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83e9545),
	.w1(32'hba0a45a5),
	.w2(32'hbb2033cd),
	.w3(32'hb90c864a),
	.w4(32'hba4e428e),
	.w5(32'hbb0c1840),
	.w6(32'h395b8a15),
	.w7(32'h3a1f1e9a),
	.w8(32'hbaf9d9a3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d338e),
	.w1(32'hbadc61a3),
	.w2(32'hbb8b25e3),
	.w3(32'hb96738f7),
	.w4(32'h3a20fe2b),
	.w5(32'hba3e82de),
	.w6(32'h3b804398),
	.w7(32'h3b73e1df),
	.w8(32'h3b171ecc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae95cd1),
	.w1(32'h39b1b9d2),
	.w2(32'hbadf3a0c),
	.w3(32'hba67a6ac),
	.w4(32'hb7d5014e),
	.w5(32'hba683ea1),
	.w6(32'h3b156338),
	.w7(32'h3ab888fe),
	.w8(32'hba097436),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04289a),
	.w1(32'h3ad01669),
	.w2(32'h3b77a720),
	.w3(32'hbc484485),
	.w4(32'hba6bbd03),
	.w5(32'hb9d0748a),
	.w6(32'h3c37c317),
	.w7(32'h3ca43135),
	.w8(32'h3c4aaf50),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e2442),
	.w1(32'hb9fcf63b),
	.w2(32'hbae7652c),
	.w3(32'h3b2482bf),
	.w4(32'h3b61c169),
	.w5(32'h3ab82c5a),
	.w6(32'h3ac8efca),
	.w7(32'h3ad4f146),
	.w8(32'h3b1f94b3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4acbd4),
	.w1(32'hba2cfc5d),
	.w2(32'hb96bba6f),
	.w3(32'h3980e748),
	.w4(32'h3abec394),
	.w5(32'hb986de37),
	.w6(32'hba681dc0),
	.w7(32'h3924c240),
	.w8(32'hb83513d9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83d5c5),
	.w1(32'h39a3afca),
	.w2(32'h3a0f9dea),
	.w3(32'hb9457268),
	.w4(32'h3a4844d5),
	.w5(32'h3a89e7c9),
	.w6(32'hba6d6a45),
	.w7(32'hb91b0f3b),
	.w8(32'h3b5dbb38),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3089cd),
	.w1(32'h3b1c9876),
	.w2(32'h3b5ba108),
	.w3(32'h3b73e0fe),
	.w4(32'h3b156174),
	.w5(32'h3b071f4a),
	.w6(32'h3bc5efac),
	.w7(32'h3b2a15ab),
	.w8(32'h3aa77d41),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b404acb),
	.w1(32'h3b087ece),
	.w2(32'h3b1d05ba),
	.w3(32'h3b3b48a0),
	.w4(32'h3b413ea6),
	.w5(32'h3b301957),
	.w6(32'hb7ccef4c),
	.w7(32'h3acf0156),
	.w8(32'h3add2ad4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b833ad3),
	.w1(32'h3bcb5e13),
	.w2(32'h3bbd2dff),
	.w3(32'h3a5137bc),
	.w4(32'h3b25e21f),
	.w5(32'h3a3324c1),
	.w6(32'h39a159b2),
	.w7(32'h37b8ad09),
	.w8(32'hba9e33fe),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a01b),
	.w1(32'hba93485e),
	.w2(32'hbac5915a),
	.w3(32'hbb875cea),
	.w4(32'hb909fbd1),
	.w5(32'hba802731),
	.w6(32'h3b07a915),
	.w7(32'h3af71c27),
	.w8(32'h3a7142bf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc244b1a),
	.w1(32'hbb9ed24d),
	.w2(32'hbbe1da40),
	.w3(32'hba27b25a),
	.w4(32'hbb359a9b),
	.w5(32'hbb1cdd06),
	.w6(32'h3b3a89d2),
	.w7(32'hbbe416f7),
	.w8(32'hbb39ba7d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17a84d),
	.w1(32'hbabab4f3),
	.w2(32'hba9f0913),
	.w3(32'hba0d54f1),
	.w4(32'hba446ddc),
	.w5(32'hba4c77c0),
	.w6(32'hba071358),
	.w7(32'hbabca5bf),
	.w8(32'hba03a703),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d19eb8),
	.w1(32'hb9a96208),
	.w2(32'h39f5223e),
	.w3(32'hba330371),
	.w4(32'h3a5955dc),
	.w5(32'hbb04e207),
	.w6(32'hba53394b),
	.w7(32'h3906916c),
	.w8(32'hbab82560),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf73b86),
	.w1(32'hba8d853c),
	.w2(32'h39d70379),
	.w3(32'hbac4f528),
	.w4(32'h399f252f),
	.w5(32'h3ac40661),
	.w6(32'hbb0f0cba),
	.w7(32'hb956b7dc),
	.w8(32'hba90d896),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1ded7),
	.w1(32'h3a51dce3),
	.w2(32'h3a19d9de),
	.w3(32'h3a5c95ed),
	.w4(32'h3ad77ae4),
	.w5(32'h3a56f5c2),
	.w6(32'h39ef2cb4),
	.w7(32'h392b4d21),
	.w8(32'h3a44c98d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf57476),
	.w1(32'h3b8db721),
	.w2(32'hba973459),
	.w3(32'hbbd8c411),
	.w4(32'hbc33675c),
	.w5(32'hbc299f97),
	.w6(32'h3b74f9a4),
	.w7(32'h3abbc6e8),
	.w8(32'h3b937a49),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadac2e9),
	.w1(32'hbb5d82af),
	.w2(32'hbb839131),
	.w3(32'h3b4bbc8e),
	.w4(32'hbaf5bb8b),
	.w5(32'hbb9f4924),
	.w6(32'h3b493598),
	.w7(32'h3c0d8b25),
	.w8(32'h3a035254),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb90577),
	.w1(32'hbbdcc4c6),
	.w2(32'hbc6530ff),
	.w3(32'h3a435e7f),
	.w4(32'h390aba04),
	.w5(32'hbc4efe3d),
	.w6(32'h3a3fc48e),
	.w7(32'hbb3a3cc3),
	.w8(32'hbbeb8a88),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeb25c),
	.w1(32'hbb993de0),
	.w2(32'hbba02053),
	.w3(32'h3c53d5d0),
	.w4(32'h3baa5134),
	.w5(32'h3b3563ca),
	.w6(32'h3c219374),
	.w7(32'h3bfbaeaa),
	.w8(32'h3bccf277),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc82f5),
	.w1(32'h394d7209),
	.w2(32'h3a9cb5bf),
	.w3(32'h396328f6),
	.w4(32'h3ad512b4),
	.w5(32'h39e037f4),
	.w6(32'h3a99f603),
	.w7(32'h3b0f6fbd),
	.w8(32'hba33f15a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba903c13),
	.w1(32'hbaa27a55),
	.w2(32'h3a0a072b),
	.w3(32'hba1f34d8),
	.w4(32'hb9a897bd),
	.w5(32'h3a43600c),
	.w6(32'hba22272c),
	.w7(32'h38d552da),
	.w8(32'hba66b6ad),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc201b),
	.w1(32'hba3e335a),
	.w2(32'hba1a30b0),
	.w3(32'h3aadc61e),
	.w4(32'h39a89616),
	.w5(32'hbaf1fae1),
	.w6(32'hbab21ae6),
	.w7(32'hbb42ec40),
	.w8(32'hbb22dc08),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825d32),
	.w1(32'hbad83e9e),
	.w2(32'hbb1e0c16),
	.w3(32'hb9f75802),
	.w4(32'hb9804098),
	.w5(32'hb91756ef),
	.w6(32'h3a835134),
	.w7(32'h3a2a6c1a),
	.w8(32'hb90e29d8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82cbd6),
	.w1(32'hb8626134),
	.w2(32'h37ad983f),
	.w3(32'h3a2f7536),
	.w4(32'h39842dbb),
	.w5(32'hbb18a745),
	.w6(32'h3ab4ffc1),
	.w7(32'h3a98ca90),
	.w8(32'hbb40f123),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6e365),
	.w1(32'hbb5fa2de),
	.w2(32'hbab7369b),
	.w3(32'hbc22cbe2),
	.w4(32'hbb8d7226),
	.w5(32'h3b00cfe0),
	.w6(32'hbb1ea85a),
	.w7(32'h3b64ab15),
	.w8(32'h3b9e4357),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856748),
	.w1(32'hbaad2eab),
	.w2(32'hbb52e384),
	.w3(32'hbba61daf),
	.w4(32'hbbce5dd4),
	.w5(32'hbbc38004),
	.w6(32'h38ee09ee),
	.w7(32'h3bc2e799),
	.w8(32'h3afe5471),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5be16),
	.w1(32'h3af6b229),
	.w2(32'hbb741ddb),
	.w3(32'h3c19598b),
	.w4(32'h3b171ec0),
	.w5(32'hbaead395),
	.w6(32'h3c3f76c9),
	.w7(32'h3bd00113),
	.w8(32'h3b844644),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a1d4c),
	.w1(32'hbb5a3e8f),
	.w2(32'hbbe50a57),
	.w3(32'hb8e05e58),
	.w4(32'hbba89c0c),
	.w5(32'hbb8bb9b3),
	.w6(32'h3b663281),
	.w7(32'hba9836c5),
	.w8(32'hb9e9aa5c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b890e21),
	.w1(32'h3b1fbd71),
	.w2(32'h3bdeab4b),
	.w3(32'h3a5b02d8),
	.w4(32'h39c9a8ad),
	.w5(32'h3a3a6465),
	.w6(32'h3b62f996),
	.w7(32'h3b3c8d87),
	.w8(32'h3b26dbe3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a953f02),
	.w1(32'h3ac76607),
	.w2(32'hbad1fe4f),
	.w3(32'h3ae5432f),
	.w4(32'h39ca6111),
	.w5(32'hbb1f000f),
	.w6(32'h3b5c8e3e),
	.w7(32'h3b76e5a9),
	.w8(32'hbb03ece7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe67f43),
	.w1(32'hbb33e2c4),
	.w2(32'hbb7c7c8d),
	.w3(32'hbb33e947),
	.w4(32'hb94247f4),
	.w5(32'hbaee8d3f),
	.w6(32'h3abf4a70),
	.w7(32'h3bb19037),
	.w8(32'h3a4bd8c6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e4463),
	.w1(32'h3b13792d),
	.w2(32'h3b251d68),
	.w3(32'hbac990d4),
	.w4(32'hb8b2eef6),
	.w5(32'h3aacf5f0),
	.w6(32'h3a70bb70),
	.w7(32'h3b261685),
	.w8(32'h3a929033),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f4643),
	.w1(32'hbb1208ff),
	.w2(32'hba2d52af),
	.w3(32'hb9dbd9de),
	.w4(32'h3a20debf),
	.w5(32'h3a2a8ba7),
	.w6(32'hbb02efc0),
	.w7(32'hb66382e5),
	.w8(32'hba59f08b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f8c72),
	.w1(32'h3b01c7d7),
	.w2(32'h3af4f2e6),
	.w3(32'hb77f143d),
	.w4(32'h3a16b481),
	.w5(32'hb93027ca),
	.w6(32'h3b0f4cb3),
	.w7(32'h3b021f09),
	.w8(32'h3a0dd467),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d648b),
	.w1(32'h3b19f07b),
	.w2(32'h3acf0e69),
	.w3(32'h3b165f06),
	.w4(32'h3ac6dc7b),
	.w5(32'h3a07b638),
	.w6(32'h3b1f78f2),
	.w7(32'h3a5ad1cd),
	.w8(32'h39fd9ab4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c2b55),
	.w1(32'hba27aad8),
	.w2(32'hbabd9a28),
	.w3(32'h3b4df231),
	.w4(32'hba768f65),
	.w5(32'h399313ad),
	.w6(32'h3b841fe8),
	.w7(32'h3a9ab1a9),
	.w8(32'h39681ae9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acad4b1),
	.w1(32'h3ac568fd),
	.w2(32'h3abdd2b5),
	.w3(32'hb8f25fac),
	.w4(32'hb994e705),
	.w5(32'h3b0c817f),
	.w6(32'hba877bc0),
	.w7(32'hba9e5e76),
	.w8(32'h3adf6f4e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae55ac4),
	.w1(32'hbb7387f5),
	.w2(32'h39b17cc0),
	.w3(32'h3b13cd7a),
	.w4(32'h3ac0813b),
	.w5(32'hbb2732d5),
	.w6(32'h3b6d1c51),
	.w7(32'h3b71a7bb),
	.w8(32'h3b245310),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded140),
	.w1(32'hbb7f5651),
	.w2(32'hbbe1ca85),
	.w3(32'hbc222e48),
	.w4(32'hbbc26de2),
	.w5(32'hbc06acae),
	.w6(32'hbae111ae),
	.w7(32'hb93b51be),
	.w8(32'hb955b4e1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf24cce),
	.w1(32'h3bf31781),
	.w2(32'h3b34db43),
	.w3(32'h3b786ad7),
	.w4(32'h3b92eaa2),
	.w5(32'h3b586cba),
	.w6(32'h3aebc77b),
	.w7(32'h3b87fa00),
	.w8(32'h3bc8eaf4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f364e),
	.w1(32'h3a85170e),
	.w2(32'h3b615de4),
	.w3(32'hbc6128c7),
	.w4(32'h3b95fa81),
	.w5(32'h3bc0f7bf),
	.w6(32'h3bf40891),
	.w7(32'h3c9f69f3),
	.w8(32'h3c57f9bf),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8c09f),
	.w1(32'h3b96d51a),
	.w2(32'h3b1a3c35),
	.w3(32'h3c3827c7),
	.w4(32'h3c1fee08),
	.w5(32'h3b6d797a),
	.w6(32'h3c39e34d),
	.w7(32'h3c0fb9f1),
	.w8(32'h3be1b042),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe262d5),
	.w1(32'hbc06b0ea),
	.w2(32'hbc271e98),
	.w3(32'hb8339eea),
	.w4(32'hbbcb5ae5),
	.w5(32'hbc211556),
	.w6(32'h3c0a2638),
	.w7(32'h3a91a69b),
	.w8(32'hba979c96),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7a0c8),
	.w1(32'h3b9d29f1),
	.w2(32'h3a97adcb),
	.w3(32'h3b2ca9d6),
	.w4(32'h3a83846d),
	.w5(32'h3a3c3273),
	.w6(32'h3bdc7451),
	.w7(32'h3b737892),
	.w8(32'h3b72aac9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d1b60),
	.w1(32'h3b3d9aaf),
	.w2(32'hbb04820f),
	.w3(32'h3bf890fe),
	.w4(32'h3a8e12a8),
	.w5(32'hbb82bfbd),
	.w6(32'h3c0f888e),
	.w7(32'h3b5d5fcc),
	.w8(32'hb8842305),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7abbcb),
	.w1(32'h3add3849),
	.w2(32'hbb422e3d),
	.w3(32'hbadf7234),
	.w4(32'hbb331565),
	.w5(32'h39d1272f),
	.w6(32'hbafc210d),
	.w7(32'hbb93e222),
	.w8(32'hb9cdbe32),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf19c45),
	.w1(32'h3adf96d3),
	.w2(32'hbae59995),
	.w3(32'hbba9bf5b),
	.w4(32'h3967e04d),
	.w5(32'hbb7c85fa),
	.w6(32'h3c580a79),
	.w7(32'h3c26387f),
	.w8(32'h3b8e8b4a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c1b6),
	.w1(32'h3c07166f),
	.w2(32'h3c32a195),
	.w3(32'hbbc7696f),
	.w4(32'h3ae6819e),
	.w5(32'h3bf4b757),
	.w6(32'h3c16daad),
	.w7(32'h3c22c2ca),
	.w8(32'h3c5680da),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc313d09),
	.w1(32'hbc807975),
	.w2(32'hbcadd90f),
	.w3(32'hb8cd07c5),
	.w4(32'h3a06a8e8),
	.w5(32'hbba493e3),
	.w6(32'hbc4fca77),
	.w7(32'h3bc51fb0),
	.w8(32'h3b90e428),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf37d18),
	.w1(32'h3b139a5f),
	.w2(32'h3b24d8f8),
	.w3(32'h3b8515bb),
	.w4(32'h3ba476f4),
	.w5(32'h3ad005ea),
	.w6(32'h3b046efa),
	.w7(32'hba413cce),
	.w8(32'hbbaf72bf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838310),
	.w1(32'h3ad0fb50),
	.w2(32'h3b6d111a),
	.w3(32'h3c5a03b0),
	.w4(32'h3c052f31),
	.w5(32'h3b6c60f9),
	.w6(32'h3c7d0a09),
	.w7(32'h3bb9a9df),
	.w8(32'h3bb7b8f9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf22a2),
	.w1(32'h3b6c7dc1),
	.w2(32'h3c24a5e5),
	.w3(32'hbc48158b),
	.w4(32'h3c2b2cae),
	.w5(32'h3c4a58c6),
	.w6(32'h3be9d1bb),
	.w7(32'h3cd351a2),
	.w8(32'h3cb15711),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e78d0),
	.w1(32'hbb40d040),
	.w2(32'hb9eb5af4),
	.w3(32'hbb87a74a),
	.w4(32'h3a011622),
	.w5(32'hbabefae1),
	.w6(32'hbba510ce),
	.w7(32'h3a47e403),
	.w8(32'hbb994990),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd148da2),
	.w1(32'hbd05bc24),
	.w2(32'hbcd1fb8f),
	.w3(32'hbc9435e3),
	.w4(32'hbc86e477),
	.w5(32'hbca350d8),
	.w6(32'hbbfe368b),
	.w7(32'h3c325e0b),
	.w8(32'hbb938f0b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc210f22),
	.w1(32'hb9b88c5d),
	.w2(32'h3ba8202c),
	.w3(32'hbc18869a),
	.w4(32'hb8fcbd56),
	.w5(32'h3b2061c9),
	.w6(32'hbb83c495),
	.w7(32'h3bedf4b4),
	.w8(32'h3c1c1938),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c76da),
	.w1(32'hbb23021c),
	.w2(32'hba2cacf2),
	.w3(32'hbb29e626),
	.w4(32'hba826741),
	.w5(32'h383cadd8),
	.w6(32'hbab46e70),
	.w7(32'hbacd3b79),
	.w8(32'h3a704d27),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e077),
	.w1(32'h3afffe0f),
	.w2(32'hbb7d7add),
	.w3(32'h396ace2c),
	.w4(32'hba4349db),
	.w5(32'hbb846201),
	.w6(32'h3b1d9168),
	.w7(32'h398c657d),
	.w8(32'h3a2dce9a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb093c91),
	.w1(32'h3b580d32),
	.w2(32'h3b43f772),
	.w3(32'h3976ecf8),
	.w4(32'hba76bca8),
	.w5(32'hbaf4ef47),
	.w6(32'h3c5c0fa9),
	.w7(32'h3c0f5b7a),
	.w8(32'h3b327f3a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa05dbd),
	.w1(32'h3adb25b9),
	.w2(32'hb9915dc8),
	.w3(32'h3b663db5),
	.w4(32'h3abcc33f),
	.w5(32'hb87e8f14),
	.w6(32'h3bbd2e75),
	.w7(32'h3a91c635),
	.w8(32'hb9537e37),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39848884),
	.w1(32'hbb4eadb4),
	.w2(32'hbc0d0110),
	.w3(32'h3b72092b),
	.w4(32'h38209566),
	.w5(32'hba01d6c0),
	.w6(32'h3b23bad5),
	.w7(32'hbb325b86),
	.w8(32'hbb1a448b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac16a13),
	.w1(32'hbae6cd69),
	.w2(32'hbb2353fa),
	.w3(32'h3a9184b8),
	.w4(32'h3952634e),
	.w5(32'h3ace8e6b),
	.w6(32'h3aac883a),
	.w7(32'h3abb7fe2),
	.w8(32'h3aa4270c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9befe2),
	.w1(32'h3b80ad39),
	.w2(32'h3c2601a0),
	.w3(32'hb9f00dd0),
	.w4(32'h3b710fee),
	.w5(32'h3b8f103d),
	.w6(32'h3bbd9b9b),
	.w7(32'h3c1fc944),
	.w8(32'h3c35543a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9705351),
	.w1(32'hba45ea35),
	.w2(32'hbbfcef23),
	.w3(32'hbbed1f14),
	.w4(32'hbb817604),
	.w5(32'hbc1ffc84),
	.w6(32'hba58c4b6),
	.w7(32'h3a104ca1),
	.w8(32'hbb3cc4c4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb400d7e),
	.w1(32'hbb090bf5),
	.w2(32'hb8db0072),
	.w3(32'h3ad1127f),
	.w4(32'h3b346445),
	.w5(32'h3b3de52e),
	.w6(32'h3bdb356e),
	.w7(32'h3b9a5838),
	.w8(32'h3b9a5f6b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3969de0d),
	.w1(32'hba0ee4f2),
	.w2(32'hba9cbc98),
	.w3(32'h3a9ea2f2),
	.w4(32'h3924be2c),
	.w5(32'h39b300d4),
	.w6(32'hb9d85327),
	.w7(32'hbab3f4d1),
	.w8(32'h3a736aa6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a633ec1),
	.w1(32'hba546bcf),
	.w2(32'hb906815c),
	.w3(32'hb8e35d26),
	.w4(32'hb88d49a9),
	.w5(32'hba5e9ddd),
	.w6(32'h3ace2454),
	.w7(32'h3a912879),
	.w8(32'hbb1bbdb2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba329603),
	.w1(32'hb9ad8891),
	.w2(32'hbaa0a052),
	.w3(32'hbb1659c7),
	.w4(32'hba7c8555),
	.w5(32'h3b38f5ab),
	.w6(32'hbb0221af),
	.w7(32'hbb598637),
	.w8(32'h3afde33f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0a240),
	.w1(32'h3a1c7241),
	.w2(32'h3aaa1d2d),
	.w3(32'h3a12f5d1),
	.w4(32'h3a8c1c0d),
	.w5(32'hbacbd0fc),
	.w6(32'h3a375c43),
	.w7(32'h3aa38a08),
	.w8(32'hba103bdb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafddb54),
	.w1(32'hbb971c88),
	.w2(32'hbb322585),
	.w3(32'h3a8b3077),
	.w4(32'h3ab7413c),
	.w5(32'h3b1a9ef6),
	.w6(32'h3c372d17),
	.w7(32'h3bad8e3c),
	.w8(32'h3bae6db3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac68a61),
	.w1(32'hbae46e49),
	.w2(32'hbaebd257),
	.w3(32'hba852bba),
	.w4(32'hba50a90b),
	.w5(32'h3990bd10),
	.w6(32'h38e6cc46),
	.w7(32'hb9df3532),
	.w8(32'h37e4e2a9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1fd3c),
	.w1(32'h3b9483f4),
	.w2(32'h3be8a84b),
	.w3(32'hbb629276),
	.w4(32'h3b9e2af6),
	.w5(32'h3bc2ae31),
	.w6(32'h3a459284),
	.w7(32'h3bf4e609),
	.w8(32'h3c2c0f11),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c013b),
	.w1(32'h3b485c13),
	.w2(32'hbb617791),
	.w3(32'h3c2b7e1d),
	.w4(32'h3928b802),
	.w5(32'hbb3547b9),
	.w6(32'h3c1c3c65),
	.w7(32'h3a2a3c2a),
	.w8(32'hbb8cf206),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989315a),
	.w1(32'h3ae8d28e),
	.w2(32'h3a8485bb),
	.w3(32'h39482703),
	.w4(32'hba37ea9c),
	.w5(32'hba9f2248),
	.w6(32'h3a252a63),
	.w7(32'h3a1bdde3),
	.w8(32'h3934e1f4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee89ac),
	.w1(32'h3a5cb631),
	.w2(32'hb9e0802f),
	.w3(32'h38bd3ed8),
	.w4(32'h3a168153),
	.w5(32'h3a9edb65),
	.w6(32'h3a88bfa4),
	.w7(32'h3a4606f3),
	.w8(32'hba08c8b3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e2595),
	.w1(32'hba37e87f),
	.w2(32'h38fe35dd),
	.w3(32'h3a3fa7e2),
	.w4(32'h3924bf1c),
	.w5(32'h3a16eb7c),
	.w6(32'h399247d6),
	.w7(32'h39f7f0d4),
	.w8(32'h3a31ed32),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cfdff),
	.w1(32'h3aa7412d),
	.w2(32'h3a859518),
	.w3(32'h3ab12ee0),
	.w4(32'h3ae059c1),
	.w5(32'h3aaff876),
	.w6(32'h3ad49867),
	.w7(32'h3ac56107),
	.w8(32'h3b1f8433),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c810e),
	.w1(32'h3b8d18f1),
	.w2(32'h3b0c8394),
	.w3(32'h3b38d6a5),
	.w4(32'hbbbdb733),
	.w5(32'hbc1695aa),
	.w6(32'h3bb1ad9f),
	.w7(32'h3c228e74),
	.w8(32'h3bb64513),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987067),
	.w1(32'hba043c63),
	.w2(32'h3aea0d48),
	.w3(32'hbc18dae0),
	.w4(32'hbb906903),
	.w5(32'hbb60c8ff),
	.w6(32'h3aef5bcb),
	.w7(32'h3b891f88),
	.w8(32'h3ad298ec),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a094a),
	.w1(32'hba134213),
	.w2(32'hbabf01d6),
	.w3(32'hbad39a17),
	.w4(32'hba4334d8),
	.w5(32'hba0ff171),
	.w6(32'hb77ddfa9),
	.w7(32'h3abb04ae),
	.w8(32'h3a2c4dc4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb438413),
	.w1(32'hbb86d6e5),
	.w2(32'hbae37452),
	.w3(32'h3a16df91),
	.w4(32'hba4b2b46),
	.w5(32'hbb23e653),
	.w6(32'hbb1feff2),
	.w7(32'hba921790),
	.w8(32'h3a91bfb2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15a2e2),
	.w1(32'h3ae846bd),
	.w2(32'h393abc81),
	.w3(32'h3b16cbe4),
	.w4(32'h39027810),
	.w5(32'h3a91b0ef),
	.w6(32'h3bfd9b02),
	.w7(32'h3b4a6deb),
	.w8(32'hb8de5b5e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa91b6b),
	.w1(32'hbaab5c07),
	.w2(32'hbb41d941),
	.w3(32'h3ac0da51),
	.w4(32'hbb3a17e3),
	.w5(32'hbb969c08),
	.w6(32'h3b73f4b3),
	.w7(32'hba592aae),
	.w8(32'hbaa5f8c1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ee456),
	.w1(32'hbb68bce8),
	.w2(32'hbbe6d93c),
	.w3(32'h3b2a87ae),
	.w4(32'hbbcce9ba),
	.w5(32'hbb8424a0),
	.w6(32'h3b5770fa),
	.w7(32'hbae97766),
	.w8(32'hb96c131c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc275655),
	.w1(32'h3acd8915),
	.w2(32'h391a148c),
	.w3(32'hbc3b9bc0),
	.w4(32'hbb04679c),
	.w5(32'hbb3d1282),
	.w6(32'h3baacf96),
	.w7(32'h3c2487e6),
	.w8(32'h3bed45d5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9ef1c),
	.w1(32'h3aba0216),
	.w2(32'hba8556bc),
	.w3(32'h3b6e5b0e),
	.w4(32'h3ae36932),
	.w5(32'hba979cf7),
	.w6(32'h3b9a2d0a),
	.w7(32'h3a78fdc6),
	.w8(32'hb9f19282),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fda3a),
	.w1(32'h3a211158),
	.w2(32'hbb62693e),
	.w3(32'hbb8d4ffd),
	.w4(32'h39e12479),
	.w5(32'hbb252fe1),
	.w6(32'h3b5c152b),
	.w7(32'h3bd80cb0),
	.w8(32'h3b168c13),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb854ca1),
	.w1(32'h3b662dbd),
	.w2(32'h3b358988),
	.w3(32'hbc08a366),
	.w4(32'h3af67c22),
	.w5(32'h3b94253c),
	.w6(32'h3bfea2e9),
	.w7(32'h3c7981e3),
	.w8(32'h3c56186a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59c8f1),
	.w1(32'hbb860749),
	.w2(32'hbbca6add),
	.w3(32'h3a404129),
	.w4(32'hbabfe537),
	.w5(32'hbaf10242),
	.w6(32'h3b8444ab),
	.w7(32'h3a9267af),
	.w8(32'h3b26f23b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812436),
	.w1(32'hbb8fdb1f),
	.w2(32'h391153e8),
	.w3(32'hbb9c68cf),
	.w4(32'hbae3b063),
	.w5(32'hba589811),
	.w6(32'h3b5d1cb6),
	.w7(32'h3b856c09),
	.w8(32'h3ab882ef),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993cdc8),
	.w1(32'hba04d14b),
	.w2(32'hba46537b),
	.w3(32'h39fb7cd4),
	.w4(32'h3ae4b03b),
	.w5(32'hba476b3a),
	.w6(32'h3b1e1410),
	.w7(32'h3afd3126),
	.w8(32'hba438855),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c3222),
	.w1(32'h3bb7fca5),
	.w2(32'h3b098c3f),
	.w3(32'h3c31253a),
	.w4(32'h393052f1),
	.w5(32'hbb0a4c04),
	.w6(32'h3bf3f32a),
	.w7(32'hb9ef61d3),
	.w8(32'h3b1d0013),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f8d86),
	.w1(32'hbb26dba8),
	.w2(32'hbb579c13),
	.w3(32'hbac4b375),
	.w4(32'hbacf32fb),
	.w5(32'hb9f68c3a),
	.w6(32'h3b57c3cf),
	.w7(32'h3ad8c0e7),
	.w8(32'h3a281a20),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03998c),
	.w1(32'h3a6eba68),
	.w2(32'h399ca602),
	.w3(32'h39f4fb2d),
	.w4(32'hb9288f3b),
	.w5(32'hba897367),
	.w6(32'h39eeedc7),
	.w7(32'h3a009ea9),
	.w8(32'hb91143f4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b058c),
	.w1(32'hb7b90f2c),
	.w2(32'hba1234b9),
	.w3(32'hba661591),
	.w4(32'hbaadeec0),
	.w5(32'hbaa4610e),
	.w6(32'h395f12d2),
	.w7(32'h3a037111),
	.w8(32'hb999cbae),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1605d),
	.w1(32'hbad8d05c),
	.w2(32'h3b310e79),
	.w3(32'hbbda4af4),
	.w4(32'hbb88bbca),
	.w5(32'hba2b61ab),
	.w6(32'hba0351f7),
	.w7(32'h3a345410),
	.w8(32'h3b279f4c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb478550),
	.w1(32'hbbbc13fa),
	.w2(32'hbb3020f1),
	.w3(32'hbb25a428),
	.w4(32'hbb82bc87),
	.w5(32'hbb9c3e25),
	.w6(32'h39f634ad),
	.w7(32'hbae804ed),
	.w8(32'hbb413943),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab90796),
	.w1(32'h3a144a3e),
	.w2(32'h39eeac3f),
	.w3(32'h3aebecba),
	.w4(32'h3a2ee92a),
	.w5(32'h3ae8d8eb),
	.w6(32'h3c1641f5),
	.w7(32'h3c07234f),
	.w8(32'h3bfb1b64),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab68b34),
	.w1(32'h3a1f58d5),
	.w2(32'h3ab287d5),
	.w3(32'h3a834d1c),
	.w4(32'h3a727640),
	.w5(32'h3a1c30b0),
	.w6(32'h3a8de683),
	.w7(32'h3a8cb5f3),
	.w8(32'h3a98034f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9641b98),
	.w1(32'h39edb08d),
	.w2(32'h3aa43ee7),
	.w3(32'hbb2485dc),
	.w4(32'hbb15045b),
	.w5(32'hbb4e6920),
	.w6(32'h3c0515e3),
	.w7(32'h3ba9f302),
	.w8(32'h3ad5f8b8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b276259),
	.w1(32'hb8d4f216),
	.w2(32'h3a815d5f),
	.w3(32'h3a8ed064),
	.w4(32'hbb087da9),
	.w5(32'hbb007088),
	.w6(32'h3b8a0dff),
	.w7(32'h3a84a057),
	.w8(32'hb9adcf6a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafaa558),
	.w1(32'h3b078415),
	.w2(32'hbaf51b85),
	.w3(32'h3a548429),
	.w4(32'h3c0da4f7),
	.w5(32'h3c1fcec6),
	.w6(32'h3c484e35),
	.w7(32'h3c8f4fd2),
	.w8(32'h3c634c96),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc91086),
	.w1(32'hb87c027a),
	.w2(32'hbab7c908),
	.w3(32'h3c51b1d4),
	.w4(32'h3ad6c98d),
	.w5(32'h3a874d91),
	.w6(32'h3c60b930),
	.w7(32'hb973de98),
	.w8(32'h3b9ead70),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afef4a3),
	.w1(32'h3a745eb6),
	.w2(32'hbab3ecd7),
	.w3(32'h3ad13961),
	.w4(32'hbb14624d),
	.w5(32'hbb1ceae2),
	.w6(32'h3b29e008),
	.w7(32'hbb2fd632),
	.w8(32'hbb8c98d7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c5d64),
	.w1(32'hbab349e9),
	.w2(32'hba8f45b3),
	.w3(32'hbb1bfd55),
	.w4(32'hba164314),
	.w5(32'h3adc1267),
	.w6(32'hb9e15831),
	.w7(32'hba3d0a35),
	.w8(32'h3799732b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6eef2),
	.w1(32'hb907321c),
	.w2(32'h3ac12840),
	.w3(32'h3901f2fa),
	.w4(32'h3a0f13dc),
	.w5(32'h3b4fa60c),
	.w6(32'h3ad35847),
	.w7(32'h3b016dc4),
	.w8(32'h3b8d1f9f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7586f),
	.w1(32'hbaf7ac81),
	.w2(32'hbb4d2294),
	.w3(32'h3692b5e1),
	.w4(32'hbb2e6aa5),
	.w5(32'hba647f6b),
	.w6(32'h3abae05c),
	.w7(32'hbafa6d66),
	.w8(32'h39874f6a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3940e),
	.w1(32'h3b91d9ee),
	.w2(32'h3b14a5b8),
	.w3(32'h3b9e34dc),
	.w4(32'h3b263880),
	.w5(32'h3afffabd),
	.w6(32'h3ae0f307),
	.w7(32'h38e73eb2),
	.w8(32'hbb3b9175),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0871f7),
	.w1(32'h385bb3c9),
	.w2(32'h3ae19b34),
	.w3(32'hba69ae4b),
	.w4(32'h3b419374),
	.w5(32'h391d4087),
	.w6(32'h3a89eda0),
	.w7(32'h3b199e9d),
	.w8(32'hb9fdee9f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88d625),
	.w1(32'hb9a37515),
	.w2(32'h3b11fb85),
	.w3(32'h3a97269f),
	.w4(32'h3b69aad0),
	.w5(32'hba571a80),
	.w6(32'hb9f54035),
	.w7(32'h3a67ad96),
	.w8(32'hb6e0cb31),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd2adc),
	.w1(32'hbb5078e7),
	.w2(32'h3a1486e3),
	.w3(32'hbbad0b5a),
	.w4(32'hbb9b2e6f),
	.w5(32'hba899d75),
	.w6(32'h3b52b9e9),
	.w7(32'h3b9b5d05),
	.w8(32'h3b4e3589),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba244ca3),
	.w1(32'hb91df4e4),
	.w2(32'h3b16a126),
	.w3(32'hbb123e1f),
	.w4(32'hba4300c7),
	.w5(32'hba21edf5),
	.w6(32'hba59772e),
	.w7(32'h3a76f411),
	.w8(32'h3b069645),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf9453),
	.w1(32'hbb02346e),
	.w2(32'hbaef9e84),
	.w3(32'hb9f77930),
	.w4(32'hba56cd1a),
	.w5(32'hb9db1496),
	.w6(32'h3abbbfc6),
	.w7(32'hba0f317b),
	.w8(32'h3b0e12f9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba148d04),
	.w1(32'hbacb7da2),
	.w2(32'hb9259f81),
	.w3(32'hb99eb6ac),
	.w4(32'h3a101c58),
	.w5(32'h3ac32a45),
	.w6(32'hbadd3cd6),
	.w7(32'h3a5232bd),
	.w8(32'h38f085d1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c116beb),
	.w1(32'h3c0ae782),
	.w2(32'h3b9aa2bc),
	.w3(32'h3b9d1da4),
	.w4(32'hba3da89b),
	.w5(32'hbbad90d1),
	.w6(32'h3b546f07),
	.w7(32'hba6b9f74),
	.w8(32'hbb96aeb3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa25e36),
	.w1(32'hbaaa8035),
	.w2(32'hba28bf7f),
	.w3(32'hbad087c2),
	.w4(32'hbad6f93c),
	.w5(32'hba2acfb9),
	.w6(32'hb8ed1201),
	.w7(32'hba9c5110),
	.w8(32'h36d85769),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f34d07),
	.w1(32'hba3dd38a),
	.w2(32'hba52419d),
	.w3(32'h39f669ce),
	.w4(32'hbacc09d9),
	.w5(32'hba2f6f0e),
	.w6(32'h3a22bb3f),
	.w7(32'hba18ac15),
	.w8(32'h3a10ebf2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afec2eb),
	.w1(32'hbb4dccc1),
	.w2(32'hba21c6b2),
	.w3(32'hba5b4e5e),
	.w4(32'h3a1d6806),
	.w5(32'h396bbf31),
	.w6(32'h3ad8f120),
	.w7(32'h3b639b73),
	.w8(32'h3a4c3124),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97362f),
	.w1(32'h3a4487f3),
	.w2(32'h3baa626d),
	.w3(32'hbb5c099e),
	.w4(32'h3a548b20),
	.w5(32'hba1bb7e6),
	.w6(32'hbb170295),
	.w7(32'h3bfdc65c),
	.w8(32'h3b9e0d20),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96d9ac),
	.w1(32'h3a7a75bd),
	.w2(32'hb9b97c7e),
	.w3(32'h3ac01553),
	.w4(32'h386e2a8c),
	.w5(32'hbac10f24),
	.w6(32'h3b22612b),
	.w7(32'h3aac000a),
	.w8(32'h39f5a4e6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc016b5),
	.w1(32'h3b563ee3),
	.w2(32'hb814a406),
	.w3(32'h3b3617e8),
	.w4(32'hba5175ca),
	.w5(32'hbba05cfe),
	.w6(32'h3c55b706),
	.w7(32'h3bc4d75f),
	.w8(32'hbb0be746),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f6601),
	.w1(32'h39a59d4d),
	.w2(32'hbaf4b379),
	.w3(32'hbb147c85),
	.w4(32'hbbb2a200),
	.w5(32'h39bc0216),
	.w6(32'hbaae1899),
	.w7(32'hbb6ad22a),
	.w8(32'h3b87d0d8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44758),
	.w1(32'h3b83bfaf),
	.w2(32'hb78453b2),
	.w3(32'hba80d917),
	.w4(32'h3b87d165),
	.w5(32'h3bcbd689),
	.w6(32'h3c5b72ca),
	.w7(32'h3c442305),
	.w8(32'h3c5f87e2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fc419),
	.w1(32'h39c0059f),
	.w2(32'hbb196615),
	.w3(32'h3b1854c0),
	.w4(32'h3a85acad),
	.w5(32'hbb5fb12c),
	.w6(32'h3bf49eec),
	.w7(32'h3c026fc3),
	.w8(32'h3bba9ee8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a785),
	.w1(32'hb7b4034e),
	.w2(32'h3a5c3526),
	.w3(32'hbbbcd70a),
	.w4(32'h3a2fbbfe),
	.w5(32'hbb0322d9),
	.w6(32'h3bb9f5de),
	.w7(32'h3c120be8),
	.w8(32'h3b23fc97),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfc3dc),
	.w1(32'h3ac925b4),
	.w2(32'h3a556670),
	.w3(32'h3b14f63a),
	.w4(32'h3b1f0674),
	.w5(32'h3a6a293b),
	.w6(32'h3b23f421),
	.w7(32'h3b57b4cc),
	.w8(32'h3b276340),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a526e),
	.w1(32'hbac0d254),
	.w2(32'hbb249dbc),
	.w3(32'hbb24e19c),
	.w4(32'hbadc6d14),
	.w5(32'hba4416f9),
	.w6(32'h3b3a78e5),
	.w7(32'h3ab29f9a),
	.w8(32'h3b5ee112),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4faa9b),
	.w1(32'h390037c6),
	.w2(32'h3a86bee3),
	.w3(32'h3a046e8d),
	.w4(32'h3abf91d0),
	.w5(32'hbb09c591),
	.w6(32'h3b052e6d),
	.w7(32'h3b07d718),
	.w8(32'hbb90f18c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb429ec),
	.w1(32'hba3abf0b),
	.w2(32'h3a54a35f),
	.w3(32'hb9e325ca),
	.w4(32'h3a59a3a3),
	.w5(32'hb98a5902),
	.w6(32'hb8dd65d0),
	.w7(32'hb982cbea),
	.w8(32'hbb1b7e70),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad995e0),
	.w1(32'hbb739c5d),
	.w2(32'hbb5b7c21),
	.w3(32'hbb02d572),
	.w4(32'hbb0a59d0),
	.w5(32'hbb58f69b),
	.w6(32'hbaf526ea),
	.w7(32'hbb3b5f96),
	.w8(32'hbb291ab3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39127028),
	.w1(32'h395b748e),
	.w2(32'hbb940216),
	.w3(32'hbb8b35bb),
	.w4(32'hbb7dc3aa),
	.w5(32'hbbc22b00),
	.w6(32'h3ac3851e),
	.w7(32'h3a0b6970),
	.w8(32'h3a171913),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2abe2),
	.w1(32'hbb66fbd7),
	.w2(32'hbaccde82),
	.w3(32'hbb3760dc),
	.w4(32'hba89190e),
	.w5(32'hbaa06768),
	.w6(32'hbb72d448),
	.w7(32'hba28ac9a),
	.w8(32'hbb00ed0a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06f70a),
	.w1(32'hbaccdeee),
	.w2(32'hba519fe2),
	.w3(32'hbac70df8),
	.w4(32'hbac4816f),
	.w5(32'hba224b79),
	.w6(32'hbae6d5a8),
	.w7(32'hba54a200),
	.w8(32'hba2dc054),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4de635),
	.w1(32'h3a1ae91d),
	.w2(32'hba1a90d2),
	.w3(32'h3af69a35),
	.w4(32'h3a9e4190),
	.w5(32'h3ad5e04b),
	.w6(32'h3afb24ac),
	.w7(32'hb98a3e96),
	.w8(32'h3b243b34),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f0e00),
	.w1(32'h3bb4d19d),
	.w2(32'h3b5a26a8),
	.w3(32'h3a962ab6),
	.w4(32'h3bd421fb),
	.w5(32'h3bbd5da7),
	.w6(32'h3bd10fe5),
	.w7(32'h3c352e0f),
	.w8(32'h3c423680),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39701282),
	.w1(32'h3ba63427),
	.w2(32'h3c106b18),
	.w3(32'hbb8a17c8),
	.w4(32'h3ac4830d),
	.w5(32'h3b87db42),
	.w6(32'h3a84bf49),
	.w7(32'h3c040c15),
	.w8(32'h3c013026),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e81e8),
	.w1(32'hbb2c47db),
	.w2(32'hbb0fb04d),
	.w3(32'hba03431b),
	.w4(32'hba9ae954),
	.w5(32'hbab0d6b0),
	.w6(32'h38da1ed5),
	.w7(32'hba7fabdd),
	.w8(32'hbaffe042),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49fcff),
	.w1(32'h3b3e4bba),
	.w2(32'hbb9e6642),
	.w3(32'hba0cbdd6),
	.w4(32'h3bbad960),
	.w5(32'hbbe04e51),
	.w6(32'h3c6fd631),
	.w7(32'h3c4e017c),
	.w8(32'h3ae2a490),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933aa94),
	.w1(32'hb98339df),
	.w2(32'hbb4e02ca),
	.w3(32'h3aea1a81),
	.w4(32'hbb89428b),
	.w5(32'h3aae3a0b),
	.w6(32'h3c13fa00),
	.w7(32'h3ba2ad86),
	.w8(32'h3c0a7eff),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393227d7),
	.w1(32'h3b25f6b0),
	.w2(32'h3b8822f5),
	.w3(32'hbb1c8f2c),
	.w4(32'hb888d113),
	.w5(32'h3ae811bc),
	.w6(32'h3ad50c82),
	.w7(32'h3b567ff3),
	.w8(32'h3a7145e2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c471b0),
	.w1(32'h3995f0a2),
	.w2(32'hba00c896),
	.w3(32'h3a4a12e8),
	.w4(32'h3ac16c90),
	.w5(32'hba4166af),
	.w6(32'hb93cb118),
	.w7(32'h376ec0e5),
	.w8(32'hba140210),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafc95f),
	.w1(32'hba9f386a),
	.w2(32'hb8a51ec4),
	.w3(32'hbae07be8),
	.w4(32'hba8772ce),
	.w5(32'hbade4ac3),
	.w6(32'hbb2fe7b1),
	.w7(32'hb9a25de0),
	.w8(32'hbadbfd4a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84b42e),
	.w1(32'hba8d34dc),
	.w2(32'hb9bfde18),
	.w3(32'hbafa283c),
	.w4(32'hb98b1d10),
	.w5(32'hba7199ba),
	.w6(32'hbb0ab918),
	.w7(32'hba6226d2),
	.w8(32'hbaf352f4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9511e2),
	.w1(32'h3bfb1429),
	.w2(32'h3c1059a0),
	.w3(32'hbb71dcd9),
	.w4(32'h386ddb24),
	.w5(32'h3b90e0bf),
	.w6(32'h3b1355b3),
	.w7(32'h3ba61008),
	.w8(32'h3bc6ef20),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6852c9),
	.w1(32'hba8be846),
	.w2(32'hbb350f00),
	.w3(32'h3a94ab04),
	.w4(32'h3a891255),
	.w5(32'h3b0debbb),
	.w6(32'h3b56f140),
	.w7(32'h3a8d6121),
	.w8(32'h3b762785),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c187642),
	.w1(32'h3ba9d72b),
	.w2(32'hbb0295b0),
	.w3(32'h3c4d04c9),
	.w4(32'h3bb339bc),
	.w5(32'hba7a736f),
	.w6(32'h3c60580f),
	.w7(32'h3be850d1),
	.w8(32'h3a06d65a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb79e),
	.w1(32'hbabe5c72),
	.w2(32'h3917e830),
	.w3(32'h3a9e99a7),
	.w4(32'hb859c9cd),
	.w5(32'h3aecd65c),
	.w6(32'h3a2acde7),
	.w7(32'h3a74a8b7),
	.w8(32'h3b343e31),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8378a9),
	.w1(32'h3b5cd93e),
	.w2(32'h3a09c4ca),
	.w3(32'hba13c925),
	.w4(32'h3b60f796),
	.w5(32'hbb248467),
	.w6(32'h3c50ef7b),
	.w7(32'h3c575a52),
	.w8(32'h3bc5fcf1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc450),
	.w1(32'hbab90b82),
	.w2(32'h3a272fec),
	.w3(32'hbba65c0f),
	.w4(32'h39d3d8d9),
	.w5(32'h3b93a503),
	.w6(32'h3b47e38a),
	.w7(32'h3b8e10c0),
	.w8(32'h3bfedec8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39604a20),
	.w1(32'h3ad6d3c3),
	.w2(32'h39ba177b),
	.w3(32'h3aa7f85f),
	.w4(32'h3a6c780b),
	.w5(32'hb9bd2c1d),
	.w6(32'h3b0ed7bd),
	.w7(32'h3a67f6a5),
	.w8(32'h397f491f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38771257),
	.w1(32'h38bc3bbc),
	.w2(32'hbb6a6dc3),
	.w3(32'h3a8a1e3f),
	.w4(32'h398d4b8c),
	.w5(32'hbac6a723),
	.w6(32'h39d600c4),
	.w7(32'h3a51eda5),
	.w8(32'hbb3e934a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed9015),
	.w1(32'hbb3c6393),
	.w2(32'hbb13b851),
	.w3(32'hbb1b091b),
	.w4(32'hba896b17),
	.w5(32'hba026687),
	.w6(32'hbb6a1bae),
	.w7(32'hbb2250fc),
	.w8(32'hb8b973ff),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ebe5b),
	.w1(32'h3b0438a4),
	.w2(32'hba16c1dc),
	.w3(32'hb9a7c8b6),
	.w4(32'h3885ccc6),
	.w5(32'hbab627ca),
	.w6(32'h3b355c89),
	.w7(32'h3b97c172),
	.w8(32'h3b1e787e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48c11d),
	.w1(32'hbbc639e5),
	.w2(32'hbba3b285),
	.w3(32'h3b18937d),
	.w4(32'hba80a3c4),
	.w5(32'h3a5844e7),
	.w6(32'h3a81be3e),
	.w7(32'hbad87401),
	.w8(32'hbaa224f8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b035e8d),
	.w1(32'hb966985c),
	.w2(32'hb9fb9450),
	.w3(32'h3b89d936),
	.w4(32'h3b3befb0),
	.w5(32'h3b28356a),
	.w6(32'h3bcd590c),
	.w7(32'h3b9950da),
	.w8(32'h3bb993c4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3863e8),
	.w1(32'h3b74bc72),
	.w2(32'h3b689cec),
	.w3(32'h3aa4038a),
	.w4(32'h3ab8810a),
	.w5(32'h3a00adac),
	.w6(32'h3b847678),
	.w7(32'h3b51f8bf),
	.w8(32'h3843baff),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12ff4b),
	.w1(32'h3b5b2cea),
	.w2(32'hbac71c5b),
	.w3(32'h3c3ecb95),
	.w4(32'h3b14d824),
	.w5(32'h3a1b7ad4),
	.w6(32'h3c437c9b),
	.w7(32'h3ba4efe7),
	.w8(32'h3b89e2dd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbecdf0),
	.w1(32'hbb81dc30),
	.w2(32'hbb3c3399),
	.w3(32'hbb6bae0e),
	.w4(32'hbb5af1f9),
	.w5(32'hbb75ba3c),
	.w6(32'h3b05269a),
	.w7(32'h3ae86e7d),
	.w8(32'h38c04884),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ca284f),
	.w1(32'h3a04ab74),
	.w2(32'hba2b00bb),
	.w3(32'hb9cb7b40),
	.w4(32'h3ad0ffde),
	.w5(32'hbaf57f73),
	.w6(32'h3c095fcb),
	.w7(32'h3bda50b7),
	.w8(32'h3b9c88b5),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ad35f),
	.w1(32'hba4d8485),
	.w2(32'hbaa5a800),
	.w3(32'hbae02764),
	.w4(32'hbaba9710),
	.w5(32'h3918e5e7),
	.w6(32'hb8839c71),
	.w7(32'hba9c717e),
	.w8(32'h38f6fb58),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d45c4c),
	.w1(32'hba856e13),
	.w2(32'hb9bb38a3),
	.w3(32'h39fdb47f),
	.w4(32'hb9784996),
	.w5(32'hbba75228),
	.w6(32'hb9812d65),
	.w7(32'hba638fdd),
	.w8(32'hbb5429cf),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ec86f),
	.w1(32'hbc173097),
	.w2(32'hbb467615),
	.w3(32'hbb3a03b7),
	.w4(32'hbb7932f7),
	.w5(32'h3ba1c682),
	.w6(32'h3ab8717e),
	.w7(32'h3bdeede6),
	.w8(32'h3c10a6b8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22ceb1),
	.w1(32'h3aea04ca),
	.w2(32'hbaab5068),
	.w3(32'h3a34d44f),
	.w4(32'h3b8b13d8),
	.w5(32'h390261ae),
	.w6(32'h3b288f0a),
	.w7(32'h3ba06b18),
	.w8(32'h3adbb75c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7d2c),
	.w1(32'hbb6fa8c1),
	.w2(32'hbb01f709),
	.w3(32'h3b918d36),
	.w4(32'h3b801925),
	.w5(32'hbae939a4),
	.w6(32'h3c1d73b4),
	.w7(32'h3bd0a264),
	.w8(32'h3b9b085f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28d4d0),
	.w1(32'h3c1d7dd6),
	.w2(32'h3c27685c),
	.w3(32'hbc025802),
	.w4(32'hbb136d5f),
	.w5(32'h3b589346),
	.w6(32'h3baeb22a),
	.w7(32'h3c407ab4),
	.w8(32'h3bfba6c7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c95a70),
	.w1(32'hba1809d8),
	.w2(32'hb8020246),
	.w3(32'h3a137477),
	.w4(32'h3a3bd203),
	.w5(32'hbac2a005),
	.w6(32'hba2919bd),
	.w7(32'hb9a7b66f),
	.w8(32'hbaf57cd0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad94fdd),
	.w1(32'hbafdd7cb),
	.w2(32'hbab2307f),
	.w3(32'hbb24cbff),
	.w4(32'hbb0f4c94),
	.w5(32'hb942f116),
	.w6(32'hb9c46c99),
	.w7(32'hb92575e3),
	.w8(32'h3978d871),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10d986),
	.w1(32'h3b78531a),
	.w2(32'h3c2e2193),
	.w3(32'hbbbe06fc),
	.w4(32'h3b4ab843),
	.w5(32'h3c1faff7),
	.w6(32'hbbdc347d),
	.w7(32'h3c99ecfa),
	.w8(32'h3c96dc63),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47536c),
	.w1(32'hbac21c62),
	.w2(32'h3b119f8c),
	.w3(32'hbc09d59e),
	.w4(32'hba29bc9b),
	.w5(32'hbafd4cbe),
	.w6(32'h3b80be8f),
	.w7(32'h3c182f60),
	.w8(32'h3bac8c4a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc203056),
	.w1(32'hba0ebdc2),
	.w2(32'h3b8f66a0),
	.w3(32'hbc5258df),
	.w4(32'h3a752354),
	.w5(32'h3ba7fd0f),
	.w6(32'hbb75515f),
	.w7(32'h3c663a98),
	.w8(32'h3c1704b7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad65b),
	.w1(32'h3aae1536),
	.w2(32'h3aeb7e60),
	.w3(32'h3b7d8c35),
	.w4(32'h3b275944),
	.w5(32'h3b18b5c8),
	.w6(32'hb9a23031),
	.w7(32'h3aa2e366),
	.w8(32'h39d6eca4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd6c59),
	.w1(32'h3b53fabf),
	.w2(32'hbab2408d),
	.w3(32'h3c208b9c),
	.w4(32'h3b13df4b),
	.w5(32'h3a1dc2b2),
	.w6(32'h3bc74ac9),
	.w7(32'h3ac98b66),
	.w8(32'h3a08c563),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33f864),
	.w1(32'h3937ac63),
	.w2(32'h39ad3be6),
	.w3(32'h39b02b14),
	.w4(32'h3a0b4cc9),
	.w5(32'hb9d4c63f),
	.w6(32'h38d2436d),
	.w7(32'h3a707ecf),
	.w8(32'hba4a93d7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c33af),
	.w1(32'hbacb9dd7),
	.w2(32'h397611de),
	.w3(32'h3b0d30b2),
	.w4(32'hba8af693),
	.w5(32'h3ad9bdeb),
	.w6(32'h3aa45619),
	.w7(32'hbab0dd50),
	.w8(32'h3a609267),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac105cc),
	.w1(32'h3b6e6e7c),
	.w2(32'h3bb1b206),
	.w3(32'hbb40902d),
	.w4(32'h3a83f197),
	.w5(32'hbb2bda6f),
	.w6(32'hba99322b),
	.w7(32'h3ac4d6c3),
	.w8(32'hba885a71),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12fcbd),
	.w1(32'hba865a78),
	.w2(32'hba2481aa),
	.w3(32'h38904f96),
	.w4(32'hba0b98e2),
	.w5(32'hbb51dfe4),
	.w6(32'hbb0dc924),
	.w7(32'hb9c0e00d),
	.w8(32'hbb90f180),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a05b9),
	.w1(32'h3a835e40),
	.w2(32'h3bc6a56c),
	.w3(32'hbbb8b0db),
	.w4(32'hb8bc6964),
	.w5(32'hb5c3be60),
	.w6(32'hbbd4e396),
	.w7(32'h3a1a152f),
	.w8(32'h3b0edb44),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cb216),
	.w1(32'hbad12b5a),
	.w2(32'hbb186282),
	.w3(32'h3b9f3d11),
	.w4(32'h3b4c2c41),
	.w5(32'hbb6b1d40),
	.w6(32'h3c31a415),
	.w7(32'h3c0c3ca4),
	.w8(32'hbb2ec09d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9799fac),
	.w1(32'h3adac88d),
	.w2(32'h3b1f9e17),
	.w3(32'h39a66d21),
	.w4(32'h3b5c13fa),
	.w5(32'hbb1348bf),
	.w6(32'h3b396ed5),
	.w7(32'h3bd7a6f5),
	.w8(32'h3aa5d033),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7f24),
	.w1(32'hbb53f931),
	.w2(32'hbb47fd2e),
	.w3(32'hbad06ab1),
	.w4(32'hba845069),
	.w5(32'hbb86978e),
	.w6(32'hbae4f9eb),
	.w7(32'h3a087cac),
	.w8(32'hbb8c6105),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc980080),
	.w1(32'hbb198df9),
	.w2(32'h3b8cfed5),
	.w3(32'hbc6b83e1),
	.w4(32'h3b35f774),
	.w5(32'h3bf57be2),
	.w6(32'hba9440af),
	.w7(32'h3cbc48c0),
	.w8(32'h3c94914a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7d45),
	.w1(32'hbaaa265e),
	.w2(32'hb6811094),
	.w3(32'h3ad666fa),
	.w4(32'hb9b84b1c),
	.w5(32'h3ac8666e),
	.w6(32'h3b72aca1),
	.w7(32'h3b3d526c),
	.w8(32'h3c0e8097),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d49b8),
	.w1(32'h3b06aad6),
	.w2(32'h3b9ff6fc),
	.w3(32'h3c04c437),
	.w4(32'h3c29b8f8),
	.w5(32'h3a8212ed),
	.w6(32'h3c6b8681),
	.w7(32'h3c71c981),
	.w8(32'hba7fd467),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6bbad),
	.w1(32'hbb6b7f1c),
	.w2(32'hb8e7a9a2),
	.w3(32'hbbf7643f),
	.w4(32'hbb2bc074),
	.w5(32'h3aef7884),
	.w6(32'h3a2f9b8a),
	.w7(32'h3aaefa19),
	.w8(32'h3b893237),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b813658),
	.w1(32'hba30979f),
	.w2(32'h3b809bdd),
	.w3(32'hba247f57),
	.w4(32'h3b4c96ab),
	.w5(32'h3b49bb03),
	.w6(32'h3b79e01d),
	.w7(32'h3b6270dc),
	.w8(32'h3a970d6e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0783a),
	.w1(32'h3b6475da),
	.w2(32'h3bae0667),
	.w3(32'h3b7aa5d7),
	.w4(32'h3bc55980),
	.w5(32'h3ad388c1),
	.w6(32'h3b47a112),
	.w7(32'h3bb06eed),
	.w8(32'h3a60185f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac26131),
	.w1(32'hba622b40),
	.w2(32'h3be0ba98),
	.w3(32'hba9009c4),
	.w4(32'h3bcaf953),
	.w5(32'h3af456a1),
	.w6(32'hbb503b70),
	.w7(32'h3b682ab6),
	.w8(32'h3b03c600),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab26f94),
	.w1(32'h3b63e322),
	.w2(32'h3c12e370),
	.w3(32'h3b81af52),
	.w4(32'h3c17bd80),
	.w5(32'h39e91301),
	.w6(32'h3ba6293b),
	.w7(32'h3c3e2db7),
	.w8(32'h3b411725),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac173a),
	.w1(32'h3b6e2d22),
	.w2(32'h3bb05522),
	.w3(32'h3b37170c),
	.w4(32'h3b9d0ac8),
	.w5(32'h3b8677a3),
	.w6(32'h3bbbbc66),
	.w7(32'h3ba6ed11),
	.w8(32'h3b3c0f97),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15ecb4),
	.w1(32'h3b2e1076),
	.w2(32'hbafc2371),
	.w3(32'hbb956984),
	.w4(32'hbb4df835),
	.w5(32'hbbfb1562),
	.w6(32'h3b95fdfe),
	.w7(32'h3b974dcc),
	.w8(32'h3b466f62),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fccb1),
	.w1(32'hbbd12992),
	.w2(32'hbac8e7d3),
	.w3(32'hbc11dfc8),
	.w4(32'hbac6a963),
	.w5(32'hba852d8e),
	.w6(32'h3b51fb82),
	.w7(32'h3c103f68),
	.w8(32'h3bcb05d5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8377a6),
	.w1(32'h3bb3cff1),
	.w2(32'h3bc03ea7),
	.w3(32'hbc016d3d),
	.w4(32'hba5afb82),
	.w5(32'hb8b6b416),
	.w6(32'h3baac894),
	.w7(32'h3bd0d884),
	.w8(32'h3c38f926),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75ca9b),
	.w1(32'h3b956fb8),
	.w2(32'hb8431c46),
	.w3(32'h3b2db92a),
	.w4(32'h3bc4156c),
	.w5(32'hb741775a),
	.w6(32'h3b8cfb13),
	.w7(32'hbb46433f),
	.w8(32'hbb29b27f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc732ae),
	.w1(32'hbb4621dc),
	.w2(32'hba8880e3),
	.w3(32'hbb255c1a),
	.w4(32'hbb62eef7),
	.w5(32'hb9b934b8),
	.w6(32'hbaeebb14),
	.w7(32'hbad28447),
	.w8(32'hbb2b7c3b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf4e7b),
	.w1(32'hba91b09c),
	.w2(32'hba4a4a33),
	.w3(32'hb9c336bc),
	.w4(32'hb9dcc1a4),
	.w5(32'hba916e0d),
	.w6(32'hbb7c506c),
	.w7(32'hbb48f29a),
	.w8(32'h39828145),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029da1),
	.w1(32'hbb367136),
	.w2(32'hbaccbbc0),
	.w3(32'hb9847191),
	.w4(32'hbaab2f51),
	.w5(32'hbbb305f1),
	.w6(32'h3a899d3d),
	.w7(32'hbaa14f1b),
	.w8(32'hbbc5e935),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f080),
	.w1(32'hbc3058e1),
	.w2(32'hbc05427c),
	.w3(32'hbc1c8f49),
	.w4(32'hbbdc0db8),
	.w5(32'hbc101fda),
	.w6(32'hbb1cfe1b),
	.w7(32'hbab6a523),
	.w8(32'hbbc663d0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf410b0),
	.w1(32'hbc140052),
	.w2(32'hbb8785ce),
	.w3(32'hba98b2e9),
	.w4(32'hba377e88),
	.w5(32'h3b858f04),
	.w6(32'hbbf6ff4a),
	.w7(32'hbb844ef6),
	.w8(32'h3b86bead),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac01929),
	.w1(32'h391c2db6),
	.w2(32'h3b0936be),
	.w3(32'h3b618a5b),
	.w4(32'h3abae268),
	.w5(32'h3b0aa00a),
	.w6(32'h3b7d6c78),
	.w7(32'h3afe5417),
	.w8(32'h3b2e49cc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa07a70),
	.w1(32'hba1cf875),
	.w2(32'hbbc4f18d),
	.w3(32'hba615797),
	.w4(32'hba8e0be7),
	.w5(32'hbc09bccd),
	.w6(32'hba26f73f),
	.w7(32'hba833e1f),
	.w8(32'hbb3b15c7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f5657),
	.w1(32'hbabbd438),
	.w2(32'hba1b6b27),
	.w3(32'hbc1157d6),
	.w4(32'hbbe1825c),
	.w5(32'hbba809a7),
	.w6(32'h3983ca8d),
	.w7(32'h3ab4ab54),
	.w8(32'hbae06429),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398953cb),
	.w1(32'hba113f46),
	.w2(32'hbb2b10a1),
	.w3(32'hbb66e0dd),
	.w4(32'h3a8f54a3),
	.w5(32'hb8f6577c),
	.w6(32'h3b9b0141),
	.w7(32'h3b9832de),
	.w8(32'h3b1f753a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa65d19),
	.w1(32'h3b14ae37),
	.w2(32'h3b12b037),
	.w3(32'hba089c85),
	.w4(32'hbb047475),
	.w5(32'hbb8f8d64),
	.w6(32'h3b5be710),
	.w7(32'h3aefb9de),
	.w8(32'hbae0f0dd),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d1712),
	.w1(32'hbbd8fce3),
	.w2(32'hbcb5ce70),
	.w3(32'hbc02c023),
	.w4(32'hbc2632ce),
	.w5(32'hbc963f99),
	.w6(32'hba1c620d),
	.w7(32'hbbcfd37e),
	.w8(32'hbba806fb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb658581),
	.w1(32'hbb540a78),
	.w2(32'hbad0f46d),
	.w3(32'hbb0eb66d),
	.w4(32'h3a2bbd97),
	.w5(32'hb9df26f9),
	.w6(32'hbb2705d0),
	.w7(32'hbaa0e1f3),
	.w8(32'hba0515c7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e0479),
	.w1(32'hbb8fdfc6),
	.w2(32'h3aade141),
	.w3(32'h3b128e77),
	.w4(32'h3bb18c41),
	.w5(32'h3c0027bf),
	.w6(32'hba400c2f),
	.w7(32'h3bdfca65),
	.w8(32'h3c17da2e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule