module layer_6_featuremap_58(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc3bbb),
	.w1(32'hbbfa6ba0),
	.w2(32'hbb64daa8),
	.w3(32'h3b27f6fa),
	.w4(32'h3c2e8be4),
	.w5(32'h3c4de7ae),
	.w6(32'hbb83eece),
	.w7(32'h3c09ae16),
	.w8(32'h3c9b95ac),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c248e3e),
	.w1(32'hba180f92),
	.w2(32'h3ba606d0),
	.w3(32'h3b76f70a),
	.w4(32'hbabb3062),
	.w5(32'hba67faca),
	.w6(32'h3a37a782),
	.w7(32'h3ad4fdfb),
	.w8(32'hbbe626c3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68ff06),
	.w1(32'h3b67c2bb),
	.w2(32'hbd153489),
	.w3(32'hbc10a892),
	.w4(32'h3b88ae9a),
	.w5(32'h3d082bf2),
	.w6(32'hbb89d874),
	.w7(32'hbcd0bb57),
	.w8(32'h3d43f844),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8abe6b),
	.w1(32'hbb81cf58),
	.w2(32'hbb77cdd1),
	.w3(32'hbb40d80a),
	.w4(32'hbc04eeb5),
	.w5(32'hbc3bcdc4),
	.w6(32'hbb378787),
	.w7(32'hbb63675c),
	.w8(32'hbbf4f5fb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a266c3e),
	.w1(32'h3c29670a),
	.w2(32'hbc92a86a),
	.w3(32'hbbc655fc),
	.w4(32'h3bd6391f),
	.w5(32'h3c0b9032),
	.w6(32'hbc3339c7),
	.w7(32'hbca912da),
	.w8(32'h3d1bdeee),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6128c),
	.w1(32'hbb31d0f3),
	.w2(32'hbafc8156),
	.w3(32'hbb132608),
	.w4(32'h3a36432d),
	.w5(32'hb79e9d9d),
	.w6(32'hbb4515f2),
	.w7(32'h3ac0e334),
	.w8(32'h3b8c67f6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8021a7),
	.w1(32'hbab45902),
	.w2(32'h3b2ce4e2),
	.w3(32'hba3a6ecb),
	.w4(32'hbb90bba1),
	.w5(32'hbba7699e),
	.w6(32'h3a259c3e),
	.w7(32'h39ab8909),
	.w8(32'hbc1f885c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83148c),
	.w1(32'hbc19e18a),
	.w2(32'hbb636fae),
	.w3(32'hbcb29aa6),
	.w4(32'h3c86a530),
	.w5(32'h3cbec168),
	.w6(32'hbcea522d),
	.w7(32'h3a618cb7),
	.w8(32'h3cf69a2e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bb2e4),
	.w1(32'hbb7ced99),
	.w2(32'h3c6c5542),
	.w3(32'h3c10f8f4),
	.w4(32'h3b747db6),
	.w5(32'hbc634bd5),
	.w6(32'h3b4f486e),
	.w7(32'h3c7c9392),
	.w8(32'hbc628172),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33af5a),
	.w1(32'h3a9a5c52),
	.w2(32'hbba35ee6),
	.w3(32'hbb3bcdc5),
	.w4(32'hbba16244),
	.w5(32'hbb5598f8),
	.w6(32'hb993a9d5),
	.w7(32'hbbdd9530),
	.w8(32'hbba5adb4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc70f87),
	.w1(32'h3c54af96),
	.w2(32'hbb484f7d),
	.w3(32'h3b798ada),
	.w4(32'h3b3349c8),
	.w5(32'h3b593eea),
	.w6(32'h3c7af48a),
	.w7(32'h3b59df2d),
	.w8(32'h3b52c602),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac0d32),
	.w1(32'h3aae4f91),
	.w2(32'hbb47e3f7),
	.w3(32'hbba1c1f3),
	.w4(32'hba85e379),
	.w5(32'h3c887852),
	.w6(32'hbbc87d92),
	.w7(32'hbbe1b126),
	.w8(32'h3c1f03e6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14b8b3),
	.w1(32'hbb5a2a0b),
	.w2(32'h3a8a4d24),
	.w3(32'hbbcd0cb0),
	.w4(32'hbb00275c),
	.w5(32'hbbc316a1),
	.w6(32'hbb6d3a93),
	.w7(32'h3a85def1),
	.w8(32'hbbc40811),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ad66f),
	.w1(32'h3952d5bc),
	.w2(32'h3c537581),
	.w3(32'h393a4fd6),
	.w4(32'h3c899302),
	.w5(32'h39b6e0cf),
	.w6(32'h3a4191ba),
	.w7(32'h3c7be4cf),
	.w8(32'h3c6af65b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1fb02),
	.w1(32'hbbcbdfd0),
	.w2(32'h3b880cce),
	.w3(32'h3aa7a572),
	.w4(32'h3b8d27c0),
	.w5(32'h3b1f7081),
	.w6(32'hba239e63),
	.w7(32'h3c077f30),
	.w8(32'h3b027cba),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b042716),
	.w1(32'hbab1fbe7),
	.w2(32'h3aff95d9),
	.w3(32'h3baa4145),
	.w4(32'h3a44089f),
	.w5(32'h3a53b817),
	.w6(32'h3b834267),
	.w7(32'h3bc97a2a),
	.w8(32'h3bdfc8e4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5415bc),
	.w1(32'hbbf89661),
	.w2(32'hbcd7e2d8),
	.w3(32'hbc271cb2),
	.w4(32'hba919111),
	.w5(32'h3c7ff8d8),
	.w6(32'hbc1c98dd),
	.w7(32'hbc959d86),
	.w8(32'h3d1e85d8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f1a27),
	.w1(32'h3b7d9e04),
	.w2(32'h3b7c67a2),
	.w3(32'h3ac224e8),
	.w4(32'hba8b66a8),
	.w5(32'h3bd36a1a),
	.w6(32'h3b812c6a),
	.w7(32'h3b921dbd),
	.w8(32'h3bf5e923),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc26405),
	.w1(32'h3bb347a7),
	.w2(32'hba944c36),
	.w3(32'hbb6c0b88),
	.w4(32'hbc60f71a),
	.w5(32'hbc67904c),
	.w6(32'h38c522f5),
	.w7(32'hbc02949c),
	.w8(32'hbc49744b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19284d),
	.w1(32'hbcbfa2f1),
	.w2(32'hbcb3124a),
	.w3(32'hbc7035f0),
	.w4(32'hbc2f0d7b),
	.w5(32'hbc5a29d1),
	.w6(32'hbcb4b959),
	.w7(32'hbc77c1ef),
	.w8(32'hbc4f26a9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4f7b9),
	.w1(32'hbb302051),
	.w2(32'h39abe359),
	.w3(32'hbb0dbffc),
	.w4(32'hbb4975aa),
	.w5(32'hbb958524),
	.w6(32'hbb32cc09),
	.w7(32'h3b2af396),
	.w8(32'hbb8651a2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c3ef6),
	.w1(32'hbc1210b2),
	.w2(32'h3bc9e379),
	.w3(32'hbb3a7274),
	.w4(32'h3c38a3da),
	.w5(32'h3bad2137),
	.w6(32'hbb6b3acd),
	.w7(32'h3c852fc7),
	.w8(32'h3c5e4060),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44c668),
	.w1(32'hbc546e06),
	.w2(32'hbc99e5ab),
	.w3(32'hbc10b30e),
	.w4(32'h3c4961d2),
	.w5(32'h3c045945),
	.w6(32'hbce5a63f),
	.w7(32'h3c2e6954),
	.w8(32'h3d61cc43),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d192998),
	.w1(32'hbbe46869),
	.w2(32'h3d612ac4),
	.w3(32'h3ac35b28),
	.w4(32'h3c33a128),
	.w5(32'hbcf6b34e),
	.w6(32'h3b9cab68),
	.w7(32'h3d39f4f7),
	.w8(32'hbd0fffd3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfeb31),
	.w1(32'hbd0d100b),
	.w2(32'hbc720566),
	.w3(32'hba93feff),
	.w4(32'hbbca00af),
	.w5(32'hbc77db51),
	.w6(32'hbc2fc318),
	.w7(32'h3c154f7e),
	.w8(32'h3c42b1f3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed0c6),
	.w1(32'hbca63a70),
	.w2(32'hbcc73127),
	.w3(32'hbd0ca5b7),
	.w4(32'hbcbd66e2),
	.w5(32'hbc94f531),
	.w6(32'hbd0bcaef),
	.w7(32'hbcc52ff5),
	.w8(32'hbbe1a2b4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d28516),
	.w1(32'hbb0644cd),
	.w2(32'h3bb4ec72),
	.w3(32'h3a53058b),
	.w4(32'hbbe51686),
	.w5(32'hbc114cef),
	.w6(32'h3a98309b),
	.w7(32'h3b92cb6f),
	.w8(32'hbb9aeb95),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47b74d),
	.w1(32'h3adca993),
	.w2(32'h3a27d8f8),
	.w3(32'h3b014717),
	.w4(32'hbbf106d7),
	.w5(32'hbc05bba9),
	.w6(32'h3b854b7f),
	.w7(32'hbab94b3b),
	.w8(32'hbc2a214e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbada6a1),
	.w1(32'hb981f14c),
	.w2(32'h3ada66a8),
	.w3(32'h3b57f97f),
	.w4(32'h3b0197d6),
	.w5(32'h3ac33204),
	.w6(32'h3b16719e),
	.w7(32'h3ae8b1d8),
	.w8(32'h3955da40),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c195853),
	.w1(32'hbcc193ae),
	.w2(32'hbca5e958),
	.w3(32'hbd0eeeab),
	.w4(32'hbc8babff),
	.w5(32'hbca498b2),
	.w6(32'hbd4f8a90),
	.w7(32'hbb5bf888),
	.w8(32'h3c4ba913),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bdf1a),
	.w1(32'hbc4cbc49),
	.w2(32'hbc843fcc),
	.w3(32'h3b8a6f43),
	.w4(32'hbbf208b9),
	.w5(32'h3c0a1c46),
	.w6(32'h3bb96cec),
	.w7(32'h3bb1bf61),
	.w8(32'h3c5cffbd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99c39c),
	.w1(32'h3c912bdd),
	.w2(32'hbb21d158),
	.w3(32'h3bd9f7a7),
	.w4(32'h3aecd09a),
	.w5(32'h3c92ad14),
	.w6(32'h3b13b154),
	.w7(32'hbcb26269),
	.w8(32'h3b416d5a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd044568),
	.w1(32'hbc84e583),
	.w2(32'h3aa2f8c4),
	.w3(32'hbc946242),
	.w4(32'h3c8314d5),
	.w5(32'hbc541d8b),
	.w6(32'hbc41ce57),
	.w7(32'h3c82e189),
	.w8(32'h3c87af19),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce49094),
	.w1(32'hbc529d1f),
	.w2(32'hbd0327ed),
	.w3(32'hbc3a3314),
	.w4(32'h3c5cd87e),
	.w5(32'h3c1ed35f),
	.w6(32'hbcf51547),
	.w7(32'hbb932d81),
	.w8(32'h3cf068ee),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdaf4e),
	.w1(32'hbae93471),
	.w2(32'h3a5b9f58),
	.w3(32'h3a320398),
	.w4(32'h3b9c21a2),
	.w5(32'h3ad26db4),
	.w6(32'hbb2b8be6),
	.w7(32'h3b29873d),
	.w8(32'h3b29afe3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c41a7),
	.w1(32'h3c255392),
	.w2(32'h3b8b8a54),
	.w3(32'hbb9f9038),
	.w4(32'hbc28767b),
	.w5(32'h3c839bc1),
	.w6(32'h3a616b78),
	.w7(32'hbcb8cf5d),
	.w8(32'hbc3c6283),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9aa763),
	.w1(32'hbba8453c),
	.w2(32'hbc095999),
	.w3(32'h3a21706e),
	.w4(32'h3b2d4c5f),
	.w5(32'hbb18dd40),
	.w6(32'hba9daa2b),
	.w7(32'hb89f3b7b),
	.w8(32'h3bd1517d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc95cf),
	.w1(32'hba302579),
	.w2(32'hb92d3b80),
	.w3(32'hbb631f29),
	.w4(32'hbc005ee7),
	.w5(32'hbbe75d15),
	.w6(32'h3a8c2da2),
	.w7(32'hbb48a6b6),
	.w8(32'hbbd44af0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f04c),
	.w1(32'h3c0a6652),
	.w2(32'h3c32c023),
	.w3(32'h3bf259ad),
	.w4(32'h3c82e02f),
	.w5(32'hbc148973),
	.w6(32'h3c3b0aea),
	.w7(32'h3c43606b),
	.w8(32'h3aba6cec),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e42f5),
	.w1(32'h3c1344cc),
	.w2(32'h3c83ebd3),
	.w3(32'h3cc161a4),
	.w4(32'h3c958c9f),
	.w5(32'h3c419525),
	.w6(32'hbb39f3f0),
	.w7(32'h3cd55a16),
	.w8(32'hb9a919a6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82c481),
	.w1(32'hbc629d38),
	.w2(32'h3c9b2ec7),
	.w3(32'hbb5d6820),
	.w4(32'hbcb9bea3),
	.w5(32'hbcf52e4e),
	.w6(32'h3c505aee),
	.w7(32'h3c802456),
	.w8(32'hbd148f3d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d66fa),
	.w1(32'hbbaa31d3),
	.w2(32'hb8ac2a4f),
	.w3(32'hbbb4a62b),
	.w4(32'hbbd2adb6),
	.w5(32'hbbf048a6),
	.w6(32'hbb96fa75),
	.w7(32'hbb5cc08e),
	.w8(32'hbbf1f3f4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5e450),
	.w1(32'hbc67e4c1),
	.w2(32'hbc6ba908),
	.w3(32'hbb401005),
	.w4(32'h39ac8147),
	.w5(32'h3b479e00),
	.w6(32'hbc3bf3c3),
	.w7(32'hbc0e1bd8),
	.w8(32'h3c1c072d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13cf06),
	.w1(32'hbcdd097f),
	.w2(32'hbc6a3433),
	.w3(32'hbcb9e8f3),
	.w4(32'hbd080aec),
	.w5(32'hbcd6591a),
	.w6(32'hbc49e420),
	.w7(32'hbc9dc057),
	.w8(32'hbb0e63f6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccf041),
	.w1(32'hbb7a841e),
	.w2(32'hb99f912b),
	.w3(32'hbb49945f),
	.w4(32'h3ab7ce74),
	.w5(32'hba6b55ec),
	.w6(32'hbb718cd6),
	.w7(32'hb8b284f5),
	.w8(32'h3a0722c8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc54b89),
	.w1(32'h3b44700f),
	.w2(32'h3be3907d),
	.w3(32'h3b283bce),
	.w4(32'h3b2d9f38),
	.w5(32'hbc217bf7),
	.w6(32'h3ba350a3),
	.w7(32'h3c9ca0ba),
	.w8(32'hbc8bfc65),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c0d05),
	.w1(32'h3b4982c2),
	.w2(32'h3c452557),
	.w3(32'h3bf03068),
	.w4(32'h3aa327e6),
	.w5(32'hbbc7d0f7),
	.w6(32'h3be9f144),
	.w7(32'h3c2922e6),
	.w8(32'hbc2c819e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce74e37),
	.w1(32'hbc619782),
	.w2(32'hbc565446),
	.w3(32'hbc362a94),
	.w4(32'h3cb3bdf1),
	.w5(32'h3ca5303d),
	.w6(32'hbcd6106f),
	.w7(32'h3cc4ec34),
	.w8(32'h3d826d6d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1939cf),
	.w1(32'h3ac3b5ba),
	.w2(32'h3b40af6b),
	.w3(32'hbaddb85b),
	.w4(32'hb9e25f01),
	.w5(32'hb9054c81),
	.w6(32'h3ac4b2d0),
	.w7(32'h3b2c4818),
	.w8(32'h3a481f48),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e1af7),
	.w1(32'h3be2f34b),
	.w2(32'hbbe49ff5),
	.w3(32'h3c8963d3),
	.w4(32'h3c7bd24f),
	.w5(32'hbb2b4580),
	.w6(32'h3c9de0cb),
	.w7(32'h3cbb2cbb),
	.w8(32'h3c9dd990),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c679d38),
	.w1(32'hbb79f61b),
	.w2(32'hb98dc1a0),
	.w3(32'hbb2281db),
	.w4(32'hbbc1bd8b),
	.w5(32'hbb991cff),
	.w6(32'hbb91856e),
	.w7(32'hbac3e9af),
	.w8(32'hbb56217f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8239d),
	.w1(32'hbc5e6193),
	.w2(32'hbb802350),
	.w3(32'hbc1dd924),
	.w4(32'hbc305a1d),
	.w5(32'hbc2eb777),
	.w6(32'hbbb9da6a),
	.w7(32'hbb02305a),
	.w8(32'hbbc40702),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5effa),
	.w1(32'hbaf84f85),
	.w2(32'h3c4f25f1),
	.w3(32'hba814552),
	.w4(32'h3b8f69fa),
	.w5(32'h3b2b9705),
	.w6(32'hbaa2a3b2),
	.w7(32'h3c1cdfa6),
	.w8(32'h3be80235),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be61b83),
	.w1(32'hbbfc85c7),
	.w2(32'hb9337482),
	.w3(32'h3be35d28),
	.w4(32'h3c227d01),
	.w5(32'h3abf503d),
	.w6(32'hbadfa5f1),
	.w7(32'h3c3c12ae),
	.w8(32'h3bc155bf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dcc05),
	.w1(32'h3bb11065),
	.w2(32'h3c037d69),
	.w3(32'h3bd18552),
	.w4(32'h3bd62ad6),
	.w5(32'h3b666a9e),
	.w6(32'hb875adb4),
	.w7(32'h3bb032f2),
	.w8(32'hbaff7110),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c0b2c),
	.w1(32'h3bead0a2),
	.w2(32'h39fddd90),
	.w3(32'h3bb3592a),
	.w4(32'hbbaca0bb),
	.w5(32'hbbd1354a),
	.w6(32'h3af3a76a),
	.w7(32'hbc477bc1),
	.w8(32'hbc66881d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb37dc),
	.w1(32'h3b9638be),
	.w2(32'h3cea3631),
	.w3(32'hbbae56ee),
	.w4(32'h3c890dfb),
	.w5(32'h3cbb2e7b),
	.w6(32'h3bd15a4f),
	.w7(32'h3d096136),
	.w8(32'h3d1d24fb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02032a),
	.w1(32'h3bad82b1),
	.w2(32'h3c705bd5),
	.w3(32'h3b5da07e),
	.w4(32'h3bf8427c),
	.w5(32'h3bceacdb),
	.w6(32'h3c446c25),
	.w7(32'h3c8a64f9),
	.w8(32'h3c33e733),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad6910),
	.w1(32'hbb741f98),
	.w2(32'hbc4c875b),
	.w3(32'h3abd8a6e),
	.w4(32'hbb8dcce2),
	.w5(32'hbbd4a28a),
	.w6(32'hbb8511aa),
	.w7(32'hbc3d4e4b),
	.w8(32'hbc46bc51),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbde0e6),
	.w1(32'hbca7b93e),
	.w2(32'hbc323028),
	.w3(32'hbc8e0121),
	.w4(32'hbc5d8e39),
	.w5(32'hbbcf2e55),
	.w6(32'hbc481f13),
	.w7(32'hbb75e226),
	.w8(32'hbb41cdd7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b7d1d),
	.w1(32'hbbc9bb5c),
	.w2(32'hbc016d3c),
	.w3(32'h3af12bc9),
	.w4(32'hba5d41e2),
	.w5(32'hbb989e0d),
	.w6(32'h368ed217),
	.w7(32'hbbc7ab51),
	.w8(32'hbc10912d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049de6),
	.w1(32'hbb101e77),
	.w2(32'hbb143d54),
	.w3(32'h3ae0981c),
	.w4(32'hbb97b619),
	.w5(32'hbc13ecb1),
	.w6(32'h3ab74432),
	.w7(32'h3b444051),
	.w8(32'h3b82d528),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d019224),
	.w1(32'h3c856107),
	.w2(32'hbc16b99b),
	.w3(32'h3c0a42e7),
	.w4(32'hb8496ade),
	.w5(32'hbb1ccdf7),
	.w6(32'hbbc0e4a9),
	.w7(32'hbc8f6ab0),
	.w8(32'hbbe80362),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3cfb6),
	.w1(32'hbc97285b),
	.w2(32'hbd685593),
	.w3(32'hbb0b8fd7),
	.w4(32'hbd0a8316),
	.w5(32'hbd25145a),
	.w6(32'hbcd0715d),
	.w7(32'hbd8b2937),
	.w8(32'hbd99178f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule