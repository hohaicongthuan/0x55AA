module layer_8_featuremap_106(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfca8c),
	.w1(32'h3b40db6c),
	.w2(32'h3a68c9cb),
	.w3(32'hbb9ac64a),
	.w4(32'h3b3ed6b6),
	.w5(32'hbaf7d8e6),
	.w6(32'h3b8f4b19),
	.w7(32'h3c441497),
	.w8(32'hbcba880a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fbd65),
	.w1(32'h3b845a1f),
	.w2(32'hbb56d079),
	.w3(32'h3b21a336),
	.w4(32'h3b93bde6),
	.w5(32'hbbe719a7),
	.w6(32'h3b1865b5),
	.w7(32'hb9ce6c85),
	.w8(32'hbbafce74),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823caa),
	.w1(32'h3b65bc0c),
	.w2(32'hbc646a90),
	.w3(32'hbc5a58ea),
	.w4(32'hbba30bf5),
	.w5(32'hbbc478e2),
	.w6(32'hba1fc252),
	.w7(32'h3ae4ebb8),
	.w8(32'hbc1d0f35),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81aa87),
	.w1(32'hbbe1ad89),
	.w2(32'h3bcc8894),
	.w3(32'hbbb7f92c),
	.w4(32'hbb3cc09e),
	.w5(32'h3c2b8dcb),
	.w6(32'hbb9a1e19),
	.w7(32'hbb810b6b),
	.w8(32'h3cdba890),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15f54a),
	.w1(32'h3a88e427),
	.w2(32'h3a1ce03d),
	.w3(32'h3b989da2),
	.w4(32'hbbed49c9),
	.w5(32'h3bc75645),
	.w6(32'hbc7e6d01),
	.w7(32'hbaf0af6a),
	.w8(32'hbc7a65ae),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c2e41),
	.w1(32'hbc1ae4e2),
	.w2(32'hbc23a1ad),
	.w3(32'hbc2e5439),
	.w4(32'hbc602baa),
	.w5(32'h3cc44f7f),
	.w6(32'hbc607a8e),
	.w7(32'h3bb3c053),
	.w8(32'h3c89e98d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95699f),
	.w1(32'hbb221295),
	.w2(32'hbc59fa43),
	.w3(32'hbbbbda7e),
	.w4(32'h3bc505e0),
	.w5(32'hbc7fce9b),
	.w6(32'hbc463e53),
	.w7(32'hbc7a83d3),
	.w8(32'h3c950edf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc303d98),
	.w1(32'h3bab399b),
	.w2(32'h3b52e336),
	.w3(32'hbb223b06),
	.w4(32'h3c74b76f),
	.w5(32'hbcc07ab2),
	.w6(32'hbc13331d),
	.w7(32'hbcb7c8c2),
	.w8(32'hbba960cc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b477876),
	.w1(32'hbc3e5438),
	.w2(32'h382abf9f),
	.w3(32'h3b260088),
	.w4(32'hbace3eed),
	.w5(32'hbc704330),
	.w6(32'hbb86ecc9),
	.w7(32'hbc1c5ed6),
	.w8(32'h3b525839),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6be3f),
	.w1(32'h3b3b4266),
	.w2(32'hbba807d5),
	.w3(32'h3c53caaf),
	.w4(32'h3b9e6607),
	.w5(32'hbb783868),
	.w6(32'hbc5de738),
	.w7(32'hbc83587d),
	.w8(32'h3d828f61),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5631b1),
	.w1(32'hbada8faf),
	.w2(32'hbc6a29c8),
	.w3(32'hb9c79fc9),
	.w4(32'hbc4b9bac),
	.w5(32'hbc48a0ff),
	.w6(32'hbb4f73cd),
	.w7(32'h3bd76eb0),
	.w8(32'hbcb99c21),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38686e),
	.w1(32'hbbe1fe58),
	.w2(32'h3c139d64),
	.w3(32'hbc0529c0),
	.w4(32'hbc2fac4b),
	.w5(32'h3c121a94),
	.w6(32'hbb3da809),
	.w7(32'hbc09749b),
	.w8(32'h3b750dda),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52ff56),
	.w1(32'hb9b6f99d),
	.w2(32'hba93b2ff),
	.w3(32'hbb56eb19),
	.w4(32'hbb30a1dd),
	.w5(32'hbb417257),
	.w6(32'hbd0163a7),
	.w7(32'hbae999f3),
	.w8(32'hbafddc5d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9cab5),
	.w1(32'hbb76200e),
	.w2(32'hba8506c0),
	.w3(32'hbb193a28),
	.w4(32'hba552f2a),
	.w5(32'hba4b5e60),
	.w6(32'h39c375b6),
	.w7(32'hbac1a103),
	.w8(32'hbafa5d15),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35674f),
	.w1(32'hba50acc0),
	.w2(32'h37b9358b),
	.w3(32'hbb59afdd),
	.w4(32'hbaf2bc73),
	.w5(32'hbb4bd31b),
	.w6(32'hbb0e4668),
	.w7(32'hbaff8981),
	.w8(32'hbb1dd7b4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd334a),
	.w1(32'h3a201b4b),
	.w2(32'h3b97f228),
	.w3(32'hbb460d7f),
	.w4(32'h3bb2e306),
	.w5(32'h3a9b4f0e),
	.w6(32'hbb0c044b),
	.w7(32'h3abf0856),
	.w8(32'h3b18e51a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb76f07),
	.w1(32'h3b23f32f),
	.w2(32'hbb85d680),
	.w3(32'hbb4832fa),
	.w4(32'h3a28da28),
	.w5(32'hba2d1d12),
	.w6(32'h3bba5bc6),
	.w7(32'hb93c1bc3),
	.w8(32'hbb65baea),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8290d),
	.w1(32'hbb23d413),
	.w2(32'hbbc30f64),
	.w3(32'hbb676f51),
	.w4(32'hbc233e26),
	.w5(32'hbc05315c),
	.w6(32'hbb255596),
	.w7(32'hbb802bb2),
	.w8(32'hb915dd12),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c70f7),
	.w1(32'h3a81931b),
	.w2(32'h3ab4f20a),
	.w3(32'hbbddf58e),
	.w4(32'h3bf4e9b0),
	.w5(32'h3b891c77),
	.w6(32'hbb4fd444),
	.w7(32'h3b27a04b),
	.w8(32'hba81bec4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbee9e4),
	.w1(32'h3bea542a),
	.w2(32'h3bddfafd),
	.w3(32'hbbcc9ee4),
	.w4(32'h3b0fef25),
	.w5(32'hbbad67a9),
	.w6(32'h3b326c22),
	.w7(32'h3b346dce),
	.w8(32'hbac07ccb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0afc1a),
	.w1(32'h3c07036b),
	.w2(32'hbbb25b7e),
	.w3(32'h39dc0512),
	.w4(32'h3b869c97),
	.w5(32'hbbd07866),
	.w6(32'h3c43c815),
	.w7(32'h3a02f638),
	.w8(32'hbb2d53cc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb449b84),
	.w1(32'hba70f648),
	.w2(32'hbc1c81a4),
	.w3(32'hbb6455d3),
	.w4(32'hbb714a92),
	.w5(32'hbb0138d1),
	.w6(32'hbbb581c2),
	.w7(32'hb6ab031c),
	.w8(32'hbbf36102),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe21bd5),
	.w1(32'hbbaf30b0),
	.w2(32'hbbb5b931),
	.w3(32'hbb36ab74),
	.w4(32'hbb281587),
	.w5(32'hbb3f6203),
	.w6(32'hbc1112eb),
	.w7(32'hbc1d01ea),
	.w8(32'hbc6e2dec),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49f03d),
	.w1(32'hba42bce5),
	.w2(32'h3ad70bb2),
	.w3(32'hbbcc08e2),
	.w4(32'hbc1a23c8),
	.w5(32'hbbab5b7d),
	.w6(32'hbc130bac),
	.w7(32'hbb6bda5d),
	.w8(32'hba890f6c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3450e),
	.w1(32'h3a22dc09),
	.w2(32'h3bfb5783),
	.w3(32'h3a13304c),
	.w4(32'h39642f5f),
	.w5(32'hbb54a002),
	.w6(32'h39d5dbce),
	.w7(32'h3c224987),
	.w8(32'h3c4a409f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5a4e1),
	.w1(32'h3c05bb6f),
	.w2(32'hbb8eea33),
	.w3(32'hb9cfe9eb),
	.w4(32'h3b6372fd),
	.w5(32'hbb68c600),
	.w6(32'h3c2ab9a4),
	.w7(32'h3b35cb1f),
	.w8(32'hbc7be111),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891ea7),
	.w1(32'h3c333557),
	.w2(32'h3b81a5c2),
	.w3(32'hbc2d348f),
	.w4(32'hbb74c445),
	.w5(32'hbb9ca391),
	.w6(32'hbbc52ba6),
	.w7(32'h3bc852b0),
	.w8(32'h3bacc5c2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75179c),
	.w1(32'hbadd51ef),
	.w2(32'h3b7f199f),
	.w3(32'hbc04367f),
	.w4(32'h3b842e08),
	.w5(32'hbac51603),
	.w6(32'hbaf74800),
	.w7(32'hbc287978),
	.w8(32'hbbc8f9ac),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a446119),
	.w1(32'hbb5839cd),
	.w2(32'h3b904d8d),
	.w3(32'hbb19707b),
	.w4(32'h3bddeddf),
	.w5(32'hba69d85e),
	.w6(32'hbc7e9b04),
	.w7(32'h3b1cbaed),
	.w8(32'hbb19e902),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a772f),
	.w1(32'hba795d88),
	.w2(32'hbc100fcc),
	.w3(32'hba3d270a),
	.w4(32'h3c288dae),
	.w5(32'h3c1b31bb),
	.w6(32'hbc039180),
	.w7(32'h3a2a0c21),
	.w8(32'h3bbcb995),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56c518),
	.w1(32'hbc920567),
	.w2(32'h39df78bc),
	.w3(32'hbb7f57ce),
	.w4(32'hbb4a391f),
	.w5(32'hbb7fc02a),
	.w6(32'hbc090666),
	.w7(32'hbba0429d),
	.w8(32'hbba4976b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcd63c),
	.w1(32'h3a0707a8),
	.w2(32'h37e833cd),
	.w3(32'hbb82fad8),
	.w4(32'hbb72a63b),
	.w5(32'hbab65e09),
	.w6(32'hbbbf90ce),
	.w7(32'h3afc75fd),
	.w8(32'h3b93864b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79d9c1),
	.w1(32'hb97ec7ae),
	.w2(32'h3c584965),
	.w3(32'h3abb5d0b),
	.w4(32'h3c395c6b),
	.w5(32'h3c749ac5),
	.w6(32'h3bebe626),
	.w7(32'h3cba22d4),
	.w8(32'h3cda3126),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4faa9f),
	.w1(32'h3be96431),
	.w2(32'hbb95dc50),
	.w3(32'h3c9716c5),
	.w4(32'hbb64d950),
	.w5(32'hbb87b4bf),
	.w6(32'h3cf3b068),
	.w7(32'hbbc01245),
	.w8(32'h3b3e2129),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafc34b),
	.w1(32'hbbcc5294),
	.w2(32'h3b171a6d),
	.w3(32'hbafcd7ed),
	.w4(32'h3b21ce57),
	.w5(32'h3a8ba48d),
	.w6(32'hbb81eb76),
	.w7(32'h3a5eb19a),
	.w8(32'hbb3eb1b7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aced1ed),
	.w1(32'h3bb8973b),
	.w2(32'h38f06679),
	.w3(32'h3ad15515),
	.w4(32'h3b1cf3ce),
	.w5(32'h3be3cf73),
	.w6(32'hbaeeab20),
	.w7(32'h3c6ecfca),
	.w8(32'h3c37ec5a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe09009),
	.w1(32'hbb64f2fd),
	.w2(32'hba21c4f5),
	.w3(32'h3bfb2698),
	.w4(32'h39a7e348),
	.w5(32'h3b45383e),
	.w6(32'h3c1f2f68),
	.w7(32'h3c52c5ef),
	.w8(32'h3c1db69e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbec78f),
	.w1(32'h3c905eea),
	.w2(32'h3c0450a7),
	.w3(32'h38bb2d01),
	.w4(32'hbb48b489),
	.w5(32'hbbc5310b),
	.w6(32'h3c6eaa4a),
	.w7(32'hba89543b),
	.w8(32'h3809e49b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c065105),
	.w1(32'h3b3c7766),
	.w2(32'h3bb19789),
	.w3(32'h3aa73738),
	.w4(32'h3ab641f6),
	.w5(32'h3bb3d84f),
	.w6(32'hba88c98a),
	.w7(32'h3b8e2140),
	.w8(32'h3a8fda12),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee8d9),
	.w1(32'h3bb423b9),
	.w2(32'h3b291720),
	.w3(32'h3b7f2590),
	.w4(32'hba622048),
	.w5(32'hba387b7b),
	.w6(32'h3a7fdc09),
	.w7(32'hbc0ba0c5),
	.w8(32'hbbd0e1a0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a954a10),
	.w1(32'h3b1443f8),
	.w2(32'h3b23d238),
	.w3(32'hba1d27ea),
	.w4(32'h39f07d1f),
	.w5(32'hb9b7359c),
	.w6(32'hbc0ca63b),
	.w7(32'hbb0d6c24),
	.w8(32'h3afa0b7a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9b543),
	.w1(32'h3a9d743c),
	.w2(32'h3b836070),
	.w3(32'h3b44f3e0),
	.w4(32'h3b8b4de1),
	.w5(32'h3aa3f625),
	.w6(32'h3a1d918b),
	.w7(32'h3ab8baf9),
	.w8(32'hbae1fcc0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccd978),
	.w1(32'h3b3f6e7f),
	.w2(32'h3ae2c57a),
	.w3(32'h39a00341),
	.w4(32'hba8156c9),
	.w5(32'hbaaddef3),
	.w6(32'h3aa67f66),
	.w7(32'hbafc1411),
	.w8(32'h3becfbaf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48bf28),
	.w1(32'hb8ff9be2),
	.w2(32'hb9a30ecc),
	.w3(32'hba22960e),
	.w4(32'hba5b9577),
	.w5(32'h39b49835),
	.w6(32'h3b6164a5),
	.w7(32'hba809d80),
	.w8(32'hb9fee333),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc53728),
	.w1(32'hbb7cba68),
	.w2(32'hbbae9c87),
	.w3(32'hb9044538),
	.w4(32'h3aee4c16),
	.w5(32'hbb2d0421),
	.w6(32'h39c798a4),
	.w7(32'h3b6d9ff2),
	.w8(32'hbb715c7b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfed73a),
	.w1(32'hbbfef87d),
	.w2(32'h3bb44dea),
	.w3(32'hbbb93885),
	.w4(32'hbba3fe67),
	.w5(32'h3a0655b0),
	.w6(32'hbc01c1fe),
	.w7(32'h3afc5420),
	.w8(32'h3c2ade7a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b8917),
	.w1(32'hba2a2c1d),
	.w2(32'h3b105014),
	.w3(32'h3a20d450),
	.w4(32'h3932fc3e),
	.w5(32'hbbf25257),
	.w6(32'h3c3a777b),
	.w7(32'hbabd3f39),
	.w8(32'hbc3c1fb8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b64950),
	.w1(32'hbb80a213),
	.w2(32'hbaf85574),
	.w3(32'hbb45168a),
	.w4(32'hbb208307),
	.w5(32'hbb015bc3),
	.w6(32'hbbdcabec),
	.w7(32'h3ae66c02),
	.w8(32'hbc036961),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b56f7),
	.w1(32'hbb9b36c5),
	.w2(32'h3bea6484),
	.w3(32'h3932c8f2),
	.w4(32'hbb51d399),
	.w5(32'hbbe6b347),
	.w6(32'hbc1e3857),
	.w7(32'hbb8070df),
	.w8(32'hbbb73fbf),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b006b06),
	.w1(32'hba83110b),
	.w2(32'h3c6c0375),
	.w3(32'hbbcdcb06),
	.w4(32'h3ba502d0),
	.w5(32'h3bac64cb),
	.w6(32'hbb0f1cd3),
	.w7(32'h3bb4fbff),
	.w8(32'h3be607cd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45d3ed),
	.w1(32'h3c1dd1e7),
	.w2(32'hbad3d41a),
	.w3(32'h3bb2b1d6),
	.w4(32'h3b51e9a8),
	.w5(32'hbae3f948),
	.w6(32'h3bd2da77),
	.w7(32'hbb685f11),
	.w8(32'hbc681f99),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f35af),
	.w1(32'hbc9a7884),
	.w2(32'h3ad67bf0),
	.w3(32'hbabbff73),
	.w4(32'hbc3985f5),
	.w5(32'hbc21db2b),
	.w6(32'hbc8fc6a4),
	.w7(32'hbb8b320e),
	.w8(32'hbc206004),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb3f6c),
	.w1(32'hbb218caf),
	.w2(32'hbaf6c81f),
	.w3(32'hbbdb9686),
	.w4(32'h3af5262d),
	.w5(32'h3ac41308),
	.w6(32'hbc4c9c14),
	.w7(32'hbae115f6),
	.w8(32'h3a96a7a2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba14263),
	.w1(32'h3a8ad3b6),
	.w2(32'h382f4d6a),
	.w3(32'h3bee74ca),
	.w4(32'hb7f53dc4),
	.w5(32'h3aafb92b),
	.w6(32'hbac1676c),
	.w7(32'hba1ac196),
	.w8(32'h3aeb648a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2305d9),
	.w1(32'hbad3c42c),
	.w2(32'hbb0e2b26),
	.w3(32'hb92cae64),
	.w4(32'h3a892d3b),
	.w5(32'h3af60af6),
	.w6(32'h3a64fa4c),
	.w7(32'h3bb1208e),
	.w8(32'h3a2bfe25),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1eb1c),
	.w1(32'h3ab9ce31),
	.w2(32'h3b953dfa),
	.w3(32'hbbfdf464),
	.w4(32'h3a875c99),
	.w5(32'hba2bdc5c),
	.w6(32'hbc023e33),
	.w7(32'h3b199abb),
	.w8(32'hbb3bfab1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ed737),
	.w1(32'hbb0d13cf),
	.w2(32'hb8ab6c99),
	.w3(32'h3aec84ee),
	.w4(32'h3b26a97f),
	.w5(32'hb880199b),
	.w6(32'hbae89814),
	.w7(32'hbc18f6f0),
	.w8(32'hbbcb8e29),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39466b8b),
	.w1(32'h3b691da4),
	.w2(32'hbb7f044a),
	.w3(32'hbaa16c95),
	.w4(32'h3c03f97d),
	.w5(32'h3ba5ed0d),
	.w6(32'hbbdf14f4),
	.w7(32'hbc47c92b),
	.w8(32'hbc00861b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9fcf3),
	.w1(32'hbc75bbfc),
	.w2(32'hb8c7bcac),
	.w3(32'hbb7ad95a),
	.w4(32'hb92858e3),
	.w5(32'h3a9b3d3c),
	.w6(32'hbc811d51),
	.w7(32'hba867907),
	.w8(32'h39f01772),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc28f),
	.w1(32'hbb3d7e6b),
	.w2(32'hbb608647),
	.w3(32'h395584ba),
	.w4(32'hbb1804ea),
	.w5(32'hbb66d622),
	.w6(32'hb88aaf3f),
	.w7(32'hba535b07),
	.w8(32'hbb739fa8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd82a),
	.w1(32'h3c14962c),
	.w2(32'hbb355c2a),
	.w3(32'hbbdbb81e),
	.w4(32'h3b3dfca8),
	.w5(32'h3baa1ede),
	.w6(32'h3ac02d20),
	.w7(32'h3c260f43),
	.w8(32'h3b73442d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc726062),
	.w1(32'hbc268043),
	.w2(32'h3be90b85),
	.w3(32'h3bdbd301),
	.w4(32'h3c22ca7d),
	.w5(32'h3b851db1),
	.w6(32'hbb0f31e6),
	.w7(32'h3c72f09a),
	.w8(32'h3c995589),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0f965),
	.w1(32'h3c6d4309),
	.w2(32'h3a5094f7),
	.w3(32'h3ad914aa),
	.w4(32'hbb6a082c),
	.w5(32'hbba0bb5f),
	.w6(32'h3c6e3fec),
	.w7(32'h3a1cc84d),
	.w8(32'hbc04dfe0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba120ded),
	.w1(32'hbb1d8a2a),
	.w2(32'h3a754d7b),
	.w3(32'hbbc1cb29),
	.w4(32'hbb4975c8),
	.w5(32'hbbdc3090),
	.w6(32'hbbc3046a),
	.w7(32'h3b27a77a),
	.w8(32'h3bf247b5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2dbbce),
	.w1(32'hbb13369a),
	.w2(32'h3c4e934a),
	.w3(32'hbbaf601d),
	.w4(32'h3b24984f),
	.w5(32'hb9cdc1c1),
	.w6(32'h3bb1c9b5),
	.w7(32'h3b4b1ef5),
	.w8(32'h3b1962a1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ef485),
	.w1(32'h3cb4a918),
	.w2(32'hbb48f963),
	.w3(32'hba5efb58),
	.w4(32'hba23bb46),
	.w5(32'hb9a44d7d),
	.w6(32'h3bd134e8),
	.w7(32'hbb9d1f55),
	.w8(32'hbbc75270),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d8719),
	.w1(32'hbade45df),
	.w2(32'hbb3fc7cf),
	.w3(32'hba76566b),
	.w4(32'hba0afc5d),
	.w5(32'h3b2a6849),
	.w6(32'hbb76e331),
	.w7(32'hbb8b8194),
	.w8(32'hbbd664aa),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a911245),
	.w1(32'hbb0cd537),
	.w2(32'hbbf71064),
	.w3(32'h3a8c6bc8),
	.w4(32'h3c02708f),
	.w5(32'h3c278f56),
	.w6(32'hbb4f277d),
	.w7(32'h3c1161fd),
	.w8(32'h3c840307),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae790b6),
	.w1(32'h3c37c242),
	.w2(32'hb948b4d4),
	.w3(32'h3c2babec),
	.w4(32'hbb5053bb),
	.w5(32'hbaf4eb31),
	.w6(32'h3ca36eb4),
	.w7(32'h3b3124da),
	.w8(32'hbb2a780d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa44919),
	.w1(32'h3ac3ebff),
	.w2(32'h3a54037e),
	.w3(32'hbbdf5a8f),
	.w4(32'h3c204134),
	.w5(32'h3bc32825),
	.w6(32'hbb9d1e57),
	.w7(32'hbb95674b),
	.w8(32'h3b8506fe),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8455b0),
	.w1(32'hbbff31ed),
	.w2(32'hbbc6e27a),
	.w3(32'h3c0e9be7),
	.w4(32'h3bca7a7b),
	.w5(32'hb959273b),
	.w6(32'h3af55728),
	.w7(32'hbc55e051),
	.w8(32'hbbfd1c34),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99327c),
	.w1(32'h3b4a3e04),
	.w2(32'h3b6c81c7),
	.w3(32'h3a291045),
	.w4(32'h3a689900),
	.w5(32'h3a2e67d2),
	.w6(32'hbbbc5375),
	.w7(32'h3bca1d1b),
	.w8(32'h3c0d2cb3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43211f),
	.w1(32'hbbae3fde),
	.w2(32'h3c3af94d),
	.w3(32'h3ba57197),
	.w4(32'hbad5be9d),
	.w5(32'hba8da70b),
	.w6(32'h3b8fb76f),
	.w7(32'h3c089908),
	.w8(32'h3c9cded5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c351b20),
	.w1(32'h3c84d39a),
	.w2(32'hbb61bd04),
	.w3(32'h3b9cabd0),
	.w4(32'h3aadb6f9),
	.w5(32'h3b173e33),
	.w6(32'h3ccd1753),
	.w7(32'hbc2f0482),
	.w8(32'hbbbe4935),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d5518),
	.w1(32'hbb7e98f0),
	.w2(32'h3aabb497),
	.w3(32'hba8729d2),
	.w4(32'hbbe65653),
	.w5(32'hbb86945d),
	.w6(32'hbb0639ea),
	.w7(32'h3b6c538b),
	.w8(32'hbb987331),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac73928),
	.w1(32'hbb6201c4),
	.w2(32'h3b4e476f),
	.w3(32'h3a07f324),
	.w4(32'hb987256c),
	.w5(32'h3b76c45c),
	.w6(32'hbb91ba56),
	.w7(32'h3a4a28f5),
	.w8(32'h3b245f38),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f518b),
	.w1(32'h3b870bad),
	.w2(32'hbb28e0cd),
	.w3(32'h3c0a6063),
	.w4(32'hbb2235f4),
	.w5(32'h3c093557),
	.w6(32'h3b189a6a),
	.w7(32'hbbf9152a),
	.w8(32'hba85c411),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf5496),
	.w1(32'h3bb29b25),
	.w2(32'hbb0d4ce6),
	.w3(32'h3b31a9e0),
	.w4(32'hba0c5bb1),
	.w5(32'hbb900808),
	.w6(32'hbb82a77e),
	.w7(32'h38ed8581),
	.w8(32'hbb61ac7a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e0e8a),
	.w1(32'hbc1e36d0),
	.w2(32'hbb48b3b3),
	.w3(32'h3b0e6e6a),
	.w4(32'hba99babf),
	.w5(32'hbb5d8834),
	.w6(32'h3b671220),
	.w7(32'h3a52c59e),
	.w8(32'hbbb82977),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31300c),
	.w1(32'hbc4262ca),
	.w2(32'hbbdd7607),
	.w3(32'hb9e6424f),
	.w4(32'h3a09f770),
	.w5(32'hbaf3bef9),
	.w6(32'hba15741b),
	.w7(32'hbcd4bbcf),
	.w8(32'hbc7bbd01),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6876a3),
	.w1(32'hbcaa67c8),
	.w2(32'h3b4bb18b),
	.w3(32'hbb70a67b),
	.w4(32'hbbf8f2ed),
	.w5(32'hbc6f4ae6),
	.w6(32'hbc06f669),
	.w7(32'hbc5ded97),
	.w8(32'hbc907c92),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26d84d),
	.w1(32'h3cb5d1e3),
	.w2(32'hbcb25ac9),
	.w3(32'hbc61f8b8),
	.w4(32'hbb76043e),
	.w5(32'h3abca42c),
	.w6(32'hbc5ab7f7),
	.w7(32'h3b6ad43d),
	.w8(32'hbcb066f5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2399a),
	.w1(32'h3ca1667f),
	.w2(32'hbc611814),
	.w3(32'hbb5a0cbf),
	.w4(32'h3c0e8f72),
	.w5(32'hbbb00e2c),
	.w6(32'hbc619744),
	.w7(32'hbb2f758a),
	.w8(32'hbc89ace4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58a025),
	.w1(32'h3cf1b1fd),
	.w2(32'h3ba018d8),
	.w3(32'hbc81e826),
	.w4(32'hbc526edb),
	.w5(32'hbc60b634),
	.w6(32'hbc9dfd5c),
	.w7(32'hbcc5da57),
	.w8(32'h3c4a5fde),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc3daa),
	.w1(32'hbbf4e108),
	.w2(32'h3bd41e06),
	.w3(32'hbbf98f66),
	.w4(32'hbb92a321),
	.w5(32'hbba2f5f6),
	.w6(32'hbba20a22),
	.w7(32'h3bdcebcc),
	.w8(32'h3c77f011),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44b5ca),
	.w1(32'hbc08dca7),
	.w2(32'hbbb56892),
	.w3(32'hbbe68467),
	.w4(32'hbb8776be),
	.w5(32'h3a83c31e),
	.w6(32'hbaab402b),
	.w7(32'hbbcbf9ad),
	.w8(32'h3c855e90),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11fb79),
	.w1(32'h3a9b6e26),
	.w2(32'hbc260ba9),
	.w3(32'hbbeefb11),
	.w4(32'hbc5c3891),
	.w5(32'hbb871341),
	.w6(32'h3bf5a0a4),
	.w7(32'hbbf5fe0b),
	.w8(32'h3c08d6cf),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc504f2f),
	.w1(32'hbc8814ab),
	.w2(32'h3c481c02),
	.w3(32'hbc2758a6),
	.w4(32'h3c15d76e),
	.w5(32'hbb005fe8),
	.w6(32'h3b9b6742),
	.w7(32'h3c2b81ac),
	.w8(32'hbb20307a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0f08b),
	.w1(32'h3c19646b),
	.w2(32'h3c0c4763),
	.w3(32'hbbcaa7bf),
	.w4(32'hbb9db751),
	.w5(32'h38c7f29c),
	.w6(32'hbb84a144),
	.w7(32'h3baef261),
	.w8(32'hbb0ead18),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba46cfe),
	.w1(32'hbb727111),
	.w2(32'h3c276545),
	.w3(32'hbbcd568f),
	.w4(32'hbba37695),
	.w5(32'h3c82c85a),
	.w6(32'hbc088236),
	.w7(32'hbbb4d33d),
	.w8(32'h3be3c564),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6062c),
	.w1(32'hbbb93c01),
	.w2(32'h3c583913),
	.w3(32'h3b9ec850),
	.w4(32'hbc4996cb),
	.w5(32'hbcc7b9f1),
	.w6(32'hbb8c2627),
	.w7(32'hbcd582ae),
	.w8(32'hbc9fad05),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d498be7),
	.w1(32'hbc1220f6),
	.w2(32'h3c0fb024),
	.w3(32'hbc36db14),
	.w4(32'hbc3bdb2b),
	.w5(32'h39b20390),
	.w6(32'hbca5d02f),
	.w7(32'hbb945da4),
	.w8(32'h3c7a1ea1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b4369),
	.w1(32'hbcacdcc7),
	.w2(32'hbc827918),
	.w3(32'hbc2f3480),
	.w4(32'h3a83922a),
	.w5(32'h3c0e24c9),
	.w6(32'hbc8f7171),
	.w7(32'hbc11b535),
	.w8(32'hbbb78740),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98eb5a),
	.w1(32'h3b223250),
	.w2(32'h3bcbe4f1),
	.w3(32'h3b80ab2d),
	.w4(32'hbbc74892),
	.w5(32'hbb9f2568),
	.w6(32'h3c218667),
	.w7(32'hbb69d8bc),
	.w8(32'hbbc6cec6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccb836),
	.w1(32'hbbc51377),
	.w2(32'hbbad96b6),
	.w3(32'hbbca9996),
	.w4(32'h3b23607d),
	.w5(32'h3b327ffb),
	.w6(32'hbbe287d2),
	.w7(32'hbae924dc),
	.w8(32'hbb4f0f9d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe21069),
	.w1(32'hbb6dcdb0),
	.w2(32'h3ca2cbb4),
	.w3(32'h3ba01cde),
	.w4(32'hbc621113),
	.w5(32'hbc971df7),
	.w6(32'hb956533d),
	.w7(32'hbb280a50),
	.w8(32'hbc1b191f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d14fc99),
	.w1(32'hbc99194d),
	.w2(32'hbc6e87f9),
	.w3(32'hbc5d51bc),
	.w4(32'h3bd23ac5),
	.w5(32'h3c47a158),
	.w6(32'hbc179418),
	.w7(32'h3bb63ca7),
	.w8(32'hbc24e230),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6fbc0c),
	.w1(32'h3d275b2f),
	.w2(32'h3b9d31ae),
	.w3(32'hbc80519e),
	.w4(32'h3aec6e13),
	.w5(32'hbb97b100),
	.w6(32'h3bdd2cc6),
	.w7(32'hbb38dcee),
	.w8(32'hbcc51a1f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33df9d),
	.w1(32'h3d0c867f),
	.w2(32'hbab1c47e),
	.w3(32'hbc432900),
	.w4(32'h3cad7e95),
	.w5(32'h3c50df21),
	.w6(32'hbc865ef6),
	.w7(32'h3ca21da2),
	.w8(32'h3c605cdb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7ccef),
	.w1(32'hbbf779ec),
	.w2(32'hbc19a61e),
	.w3(32'h3c19edee),
	.w4(32'hbc03b36e),
	.w5(32'h3baa0aa2),
	.w6(32'h3ba36227),
	.w7(32'hbb80412b),
	.w8(32'h3d01b5d6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf353a6),
	.w1(32'h3a63d079),
	.w2(32'h3bc986ef),
	.w3(32'h3aac63a2),
	.w4(32'hbad0e830),
	.w5(32'hbba200b1),
	.w6(32'h3cd43ad7),
	.w7(32'hbc09da49),
	.w8(32'h3c0d8fbc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf768c5),
	.w1(32'h3b6a8e04),
	.w2(32'h3c656c07),
	.w3(32'hbc4faf8e),
	.w4(32'hbb67d663),
	.w5(32'hbc2c30a6),
	.w6(32'hbc388ae8),
	.w7(32'h3b6451df),
	.w8(32'hbcc3d971),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76c382),
	.w1(32'h3b521e5f),
	.w2(32'h3b9fab50),
	.w3(32'hbc6905f4),
	.w4(32'hbbb2c421),
	.w5(32'hbc868ff6),
	.w6(32'hbc8bfd54),
	.w7(32'hbca80fe9),
	.w8(32'hbce0998b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9eb58),
	.w1(32'h3cabe7a2),
	.w2(32'hbc4b1a44),
	.w3(32'hbcbd81cb),
	.w4(32'h394acad2),
	.w5(32'h3a890f22),
	.w6(32'hbc543902),
	.w7(32'hbcacdaef),
	.w8(32'hbc925b43),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8e6b2),
	.w1(32'hbcb90d89),
	.w2(32'hbade6118),
	.w3(32'hba58b092),
	.w4(32'hbb8419d4),
	.w5(32'h3956b9d0),
	.w6(32'hbc66e9a1),
	.w7(32'hbc935696),
	.w8(32'hbc529afe),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8abaea),
	.w1(32'hbb99f31c),
	.w2(32'h3c41beb0),
	.w3(32'hbbfe5b7f),
	.w4(32'h3ab518e1),
	.w5(32'h3c97d56f),
	.w6(32'hbcb596ba),
	.w7(32'h3c6c030d),
	.w8(32'h3cc4a3f3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6aca7),
	.w1(32'hbcb205e8),
	.w2(32'hbb557192),
	.w3(32'h3c2d8dca),
	.w4(32'hbb3de6bb),
	.w5(32'h3a95351f),
	.w6(32'h3c3b0169),
	.w7(32'hbaf7a75e),
	.w8(32'hb9d8a038),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e4cde),
	.w1(32'h3cc48009),
	.w2(32'hbbb60b57),
	.w3(32'hbaaf3326),
	.w4(32'hbab28e0a),
	.w5(32'h3c362a0e),
	.w6(32'h3c264e4e),
	.w7(32'hbc2c2a9e),
	.w8(32'hba461133),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b60189),
	.w1(32'h3bd3a6b6),
	.w2(32'h3b9c1cea),
	.w3(32'h3b28183e),
	.w4(32'h3ac23808),
	.w5(32'h3a0e46ae),
	.w6(32'hbbb273fd),
	.w7(32'hbb074ba9),
	.w8(32'h3c2b89e5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3bb87),
	.w1(32'hbc680b87),
	.w2(32'h3b98c43c),
	.w3(32'hbc0cdf52),
	.w4(32'hbc118b4f),
	.w5(32'h39cefd09),
	.w6(32'h3bc518af),
	.w7(32'hbbe0fe46),
	.w8(32'h3bb915eb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223200),
	.w1(32'h3c07e7ef),
	.w2(32'hbbba3eeb),
	.w3(32'hbbb97745),
	.w4(32'h3c272361),
	.w5(32'h3c289491),
	.w6(32'h3c9192f0),
	.w7(32'hbc44edf8),
	.w8(32'hbb244f9f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa683e),
	.w1(32'h3c0c452d),
	.w2(32'h3b9fa20a),
	.w3(32'hbb037747),
	.w4(32'hbc9da1e8),
	.w5(32'hbc836876),
	.w6(32'h3bfb3a61),
	.w7(32'hbc99a187),
	.w8(32'hbc16d225),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c278471),
	.w1(32'h3bea792d),
	.w2(32'h3c855612),
	.w3(32'h3aab477d),
	.w4(32'hbc3c8cbb),
	.w5(32'hbc838fb2),
	.w6(32'hb9f69a96),
	.w7(32'hbbcfd98e),
	.w8(32'hbc895e6f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce17266),
	.w1(32'hbbf38d6f),
	.w2(32'h3d1761ed),
	.w3(32'hbcbc169b),
	.w4(32'hbced18ba),
	.w5(32'hbd46092d),
	.w6(32'hbc689887),
	.w7(32'hbccec5bf),
	.w8(32'hbd0d9f7e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db6c3a8),
	.w1(32'h3cdb7502),
	.w2(32'hbc2faebc),
	.w3(32'hbd370267),
	.w4(32'hbb1bec9f),
	.w5(32'h3c2ac405),
	.w6(32'hbd0c13d8),
	.w7(32'hbbf69b42),
	.w8(32'h3bdeed92),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebbd91),
	.w1(32'h3c0ec7fe),
	.w2(32'hba5827fa),
	.w3(32'hbc5dd32f),
	.w4(32'h3ae31bfb),
	.w5(32'h3cc72a39),
	.w6(32'hbc127057),
	.w7(32'h3c8d83d3),
	.w8(32'h3cd4b945),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd701363),
	.w1(32'hbcd33d27),
	.w2(32'hbb82ae42),
	.w3(32'h3c674785),
	.w4(32'h3b37798c),
	.w5(32'hbbc2787f),
	.w6(32'h3c9ebfb4),
	.w7(32'h3c80f928),
	.w8(32'hbc4ab3ae),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d152044),
	.w1(32'h3bc18858),
	.w2(32'hbb4def0d),
	.w3(32'hbc7d25d3),
	.w4(32'hba77dd0c),
	.w5(32'h3b8fa8eb),
	.w6(32'hbcbfaa2a),
	.w7(32'hbb4197f7),
	.w8(32'h3aa3efb6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7922a7),
	.w1(32'h3af0379e),
	.w2(32'h3c980313),
	.w3(32'h3af5ef39),
	.w4(32'hbc13c9eb),
	.w5(32'hbc5e4e15),
	.w6(32'hbacc3721),
	.w7(32'hbc0abb73),
	.w8(32'h3b3ac48d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb50efd),
	.w1(32'hbc118a8f),
	.w2(32'h3c916c89),
	.w3(32'hbc8159aa),
	.w4(32'hbc950e0e),
	.w5(32'hbcdf51b6),
	.w6(32'hbc9ff895),
	.w7(32'hbc8ac0f2),
	.w8(32'hbc8ce380),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d336842),
	.w1(32'h3c8d3be4),
	.w2(32'hbc4a07c8),
	.w3(32'hbcaeffa9),
	.w4(32'hba71011f),
	.w5(32'hbba364c5),
	.w6(32'hbc9366af),
	.w7(32'hbc89616f),
	.w8(32'hbcd2a4b9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9775ba),
	.w1(32'hbb883d23),
	.w2(32'h3c096772),
	.w3(32'hbb62c3c5),
	.w4(32'h3a987524),
	.w5(32'h3c5628ab),
	.w6(32'hbc78ebee),
	.w7(32'h3bc69dfb),
	.w8(32'h3ce84de9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cf15f),
	.w1(32'h3c972d51),
	.w2(32'hbb820dd6),
	.w3(32'hbbd11b17),
	.w4(32'hb9a22e8a),
	.w5(32'h3bede6b9),
	.w6(32'hbb787e77),
	.w7(32'hbbe065bb),
	.w8(32'hba11f37c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33240f),
	.w1(32'h3b865bc3),
	.w2(32'h3c4669ff),
	.w3(32'h3b01d833),
	.w4(32'h3951b040),
	.w5(32'h3ae31c7e),
	.w6(32'hbb877047),
	.w7(32'h3ba24180),
	.w8(32'hbb95ac63),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc16661),
	.w1(32'hba2ad7fb),
	.w2(32'h3cf22b7c),
	.w3(32'hbabc4f4c),
	.w4(32'hbc3a5cbf),
	.w5(32'hbc72e79f),
	.w6(32'hbba06995),
	.w7(32'hba6835b5),
	.w8(32'h3bea6305),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba19114),
	.w1(32'hbc0bfcfa),
	.w2(32'h3c331e10),
	.w3(32'hbb9ffa91),
	.w4(32'hbaae14ed),
	.w5(32'h3a94ad14),
	.w6(32'hbc4bec59),
	.w7(32'h3b84a248),
	.w8(32'h3bd7c725),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd76279),
	.w1(32'h3c119e32),
	.w2(32'h3c2380d4),
	.w3(32'hbb830770),
	.w4(32'h38802f07),
	.w5(32'hbb7ada75),
	.w6(32'h3b8fa42b),
	.w7(32'hbb97307b),
	.w8(32'hbcd28683),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb945f7b),
	.w1(32'h3ae97f28),
	.w2(32'hba801870),
	.w3(32'h3c4212bb),
	.w4(32'hba6de70f),
	.w5(32'h3baa8121),
	.w6(32'h3ba5b05e),
	.w7(32'h3b29934e),
	.w8(32'hbba0d7e7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule