module layer_5 (
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 2048;
	parameter IMG_SIZE = 104;

	wire	valid_out_0,
		valid_out_1,
		valid_out_2,
		valid_out_3,
		valid_out_4,
		valid_out_5,
		valid_out_6,
		valid_out_7,
		valid_out_8,
		valid_out_9,
		valid_out_10,
		valid_out_11,
		valid_out_12,
		valid_out_13,
		valid_out_14,
		valid_out_15,
		valid_out_16,
		valid_out_17,
		valid_out_18,
		valid_out_19,
		valid_out_20,
		valid_out_21,
		valid_out_22,
		valid_out_23,
		valid_out_24,
		valid_out_25,
		valid_out_26,
		valid_out_27,
		valid_out_28,
		valid_out_29,
		valid_out_30,
		valid_out_31,
		valid_out_32,
		valid_out_33,
		valid_out_34,
		valid_out_35,
		valid_out_36,
		valid_out_37,
		valid_out_38,
		valid_out_39,
		valid_out_40,
		valid_out_41,
		valid_out_42,
		valid_out_43,
		valid_out_44,
		valid_out_45,
		valid_out_46,
		valid_out_47,
		valid_out_48,
		valid_out_49,
		valid_out_50,
		valid_out_51,
		valid_out_52,
		valid_out_53,
		valid_out_54,
		valid_out_55,
		valid_out_56,
		valid_out_57,
		valid_out_58,
		valid_out_59,
		valid_out_60,
		valid_out_61,
		valid_out_62,
		valid_out_63;
Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(data_out[31:0]),
	.valid_out(valid_out_0)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(data_out[63:32]),
	.valid_out(valid_out_1)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(data_out[95:64]),
	.valid_out(valid_out_2)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(data_out[127:96]),
	.valid_out(valid_out_3)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(data_out[159:128]),
	.valid_out(valid_out_4)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(data_out[191:160]),
	.valid_out(valid_out_5)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(data_out[223:192]),
	.valid_out(valid_out_6)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(data_out[255:224]),
	.valid_out(valid_out_7)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(data_out[287:256]),
	.valid_out(valid_out_8)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(data_out[319:288]),
	.valid_out(valid_out_9)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(data_out[351:320]),
	.valid_out(valid_out_10)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(data_out[383:352]),
	.valid_out(valid_out_11)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(data_out[415:384]),
	.valid_out(valid_out_12)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(data_out[447:416]),
	.valid_out(valid_out_13)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(data_out[479:448]),
	.valid_out(valid_out_14)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(data_out[511:480]),
	.valid_out(valid_out_15)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(data_out[543:512]),
	.valid_out(valid_out_16)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(data_out[575:544]),
	.valid_out(valid_out_17)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(data_out[607:576]),
	.valid_out(valid_out_18)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(data_out[639:608]),
	.valid_out(valid_out_19)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(data_out[671:640]),
	.valid_out(valid_out_20)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(data_out[703:672]),
	.valid_out(valid_out_21)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(data_out[735:704]),
	.valid_out(valid_out_22)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(data_out[767:736]),
	.valid_out(valid_out_23)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(data_out[799:768]),
	.valid_out(valid_out_24)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(data_out[831:800]),
	.valid_out(valid_out_25)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(data_out[863:832]),
	.valid_out(valid_out_26)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(data_out[895:864]),
	.valid_out(valid_out_27)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(data_out[927:896]),
	.valid_out(valid_out_28)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(data_out[959:928]),
	.valid_out(valid_out_29)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(data_out[991:960]),
	.valid_out(valid_out_30)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(data_out[1023:992]),
	.valid_out(valid_out_31)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(data_out[1055:1024]),
	.valid_out(valid_out_32)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(data_out[1087:1056]),
	.valid_out(valid_out_33)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(data_out[1119:1088]),
	.valid_out(valid_out_34)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(data_out[1151:1120]),
	.valid_out(valid_out_35)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(data_out[1183:1152]),
	.valid_out(valid_out_36)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(data_out[1215:1184]),
	.valid_out(valid_out_37)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(data_out[1247:1216]),
	.valid_out(valid_out_38)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(data_out[1279:1248]),
	.valid_out(valid_out_39)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(data_out[1311:1280]),
	.valid_out(valid_out_40)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(data_out[1343:1312]),
	.valid_out(valid_out_41)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(data_out[1375:1344]),
	.valid_out(valid_out_42)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(data_out[1407:1376]),
	.valid_out(valid_out_43)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(data_out[1439:1408]),
	.valid_out(valid_out_44)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(data_out[1471:1440]),
	.valid_out(valid_out_45)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(data_out[1503:1472]),
	.valid_out(valid_out_46)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(data_out[1535:1504]),
	.valid_out(valid_out_47)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(data_out[1567:1536]),
	.valid_out(valid_out_48)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(data_out[1599:1568]),
	.valid_out(valid_out_49)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(data_out[1631:1600]),
	.valid_out(valid_out_50)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(data_out[1663:1632]),
	.valid_out(valid_out_51)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(data_out[1695:1664]),
	.valid_out(valid_out_52)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(data_out[1727:1696]),
	.valid_out(valid_out_53)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(data_out[1759:1728]),
	.valid_out(valid_out_54)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(data_out[1791:1760]),
	.valid_out(valid_out_55)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(data_out[1823:1792]),
	.valid_out(valid_out_56)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(data_out[1855:1824]),
	.valid_out(valid_out_57)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(data_out[1887:1856]),
	.valid_out(valid_out_58)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(data_out[1919:1888]),
	.valid_out(valid_out_59)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(data_out[1951:1920]),
	.valid_out(valid_out_60)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(data_out[1983:1952]),
	.valid_out(valid_out_61)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(data_out[2015:1984]),
	.valid_out(valid_out_62)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(data_out[2047:2016]),
	.valid_out(valid_out_63)
);

	assign valid_out = valid_out_0 & valid_out_1 & valid_out_2 & valid_out_3 & valid_out_4 & valid_out_5 & valid_out_6 & valid_out_7 & valid_out_8 & valid_out_9 & valid_out_10 & valid_out_11 & valid_out_12 & valid_out_13 & valid_out_14 & valid_out_15 & valid_out_16 & valid_out_17 & valid_out_18 & valid_out_19 & valid_out_20 & valid_out_21 & valid_out_22 & valid_out_23 & valid_out_24 & valid_out_25 & valid_out_26 & valid_out_27 & valid_out_28 & valid_out_29 & valid_out_30 & valid_out_31 & valid_out_32 & valid_out_33 & valid_out_34 & valid_out_35 & valid_out_36 & valid_out_37 & valid_out_38 & valid_out_39 & valid_out_40 & valid_out_41 & valid_out_42 & valid_out_43 & valid_out_44 & valid_out_45 & valid_out_46 & valid_out_47 & valid_out_48 & valid_out_49 & valid_out_50 & valid_out_51 & valid_out_52 & valid_out_53 & valid_out_54 & valid_out_55 & valid_out_56 & valid_out_57 & valid_out_58 & valid_out_59 & valid_out_60 & valid_out_61 & valid_out_62 & valid_out_63;
endmodule