module layer_10_featuremap_131(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d5390),
	.w1(32'hbae9bde2),
	.w2(32'h3b291289),
	.w3(32'hba5e4f1b),
	.w4(32'hbb3ae411),
	.w5(32'h3aa7f9fa),
	.w6(32'hba9a329b),
	.w7(32'h3a919e91),
	.w8(32'h3b106dd7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4c137),
	.w1(32'h3adf0c1c),
	.w2(32'h3a264204),
	.w3(32'h3bc83eb2),
	.w4(32'h3a8840ec),
	.w5(32'hba4b7431),
	.w6(32'h3b1d7faa),
	.w7(32'h3ad735f5),
	.w8(32'hb9fd0f1a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3791c4fb),
	.w1(32'hb8e41a9a),
	.w2(32'h3a169efa),
	.w3(32'hb9b98da1),
	.w4(32'hb97df89f),
	.w5(32'hb8a57cd2),
	.w6(32'hba5b1cd5),
	.w7(32'hb9874809),
	.w8(32'hb9766ab6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f81cf),
	.w1(32'hbb106c91),
	.w2(32'hbb352ee8),
	.w3(32'hba021160),
	.w4(32'hbb722d57),
	.w5(32'hbb20a331),
	.w6(32'hbb10d13c),
	.w7(32'hbb2c228e),
	.w8(32'hbab5a04b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2fbb1),
	.w1(32'hb9951347),
	.w2(32'hba20658b),
	.w3(32'hba9fa728),
	.w4(32'hb9df260a),
	.w5(32'hba8fd0d5),
	.w6(32'hb6a50946),
	.w7(32'hbb0f8b64),
	.w8(32'h39ec850a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81703d),
	.w1(32'h3aca2a87),
	.w2(32'h38aa4e49),
	.w3(32'hbabb55cd),
	.w4(32'h3993aa07),
	.w5(32'hba070089),
	.w6(32'h3a93bea3),
	.w7(32'h38fbb0aa),
	.w8(32'hba8b5434),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853b3b),
	.w1(32'h388bc679),
	.w2(32'h3b8a5d0a),
	.w3(32'hbbba4558),
	.w4(32'h38a0d49e),
	.w5(32'h3b7808e1),
	.w6(32'hbab634b5),
	.w7(32'hb949db70),
	.w8(32'h3ba875f3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a877df2),
	.w1(32'h3a83fb7e),
	.w2(32'h3b8d7f9d),
	.w3(32'h3b626182),
	.w4(32'h3afb1f76),
	.w5(32'h3b321d14),
	.w6(32'hbae6786c),
	.w7(32'h3b4d5e8c),
	.w8(32'h3b4a2b4c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7a715),
	.w1(32'hba9f401c),
	.w2(32'hba08b0e6),
	.w3(32'hba8c2474),
	.w4(32'hba3f42b5),
	.w5(32'hb8872c3b),
	.w6(32'hba751ba9),
	.w7(32'hb8b62c43),
	.w8(32'h3a7a7470),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba44f13),
	.w1(32'h3badc3d6),
	.w2(32'h3bedf737),
	.w3(32'h3a9cd96c),
	.w4(32'hba488614),
	.w5(32'h3a0e51f2),
	.w6(32'h3b1d3792),
	.w7(32'h3b72a772),
	.w8(32'h3b930a60),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e0e13),
	.w1(32'hba9ee1e5),
	.w2(32'hba695ebd),
	.w3(32'hba2fdef2),
	.w4(32'hbb03787f),
	.w5(32'hb9dbbb6e),
	.w6(32'hb9401bc0),
	.w7(32'hb9f6bce9),
	.w8(32'hbac9b804),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78fea8),
	.w1(32'hbb2a67ca),
	.w2(32'h3b7d49f1),
	.w3(32'hbb8ce7b7),
	.w4(32'hbba2f775),
	.w5(32'h3b09dbea),
	.w6(32'hbb6b0251),
	.w7(32'hbb24ab45),
	.w8(32'h3b9e168b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a6003),
	.w1(32'h3b86b588),
	.w2(32'h3bd50db0),
	.w3(32'hba84e6b8),
	.w4(32'h395e4ec2),
	.w5(32'h3afa3e1e),
	.w6(32'h39a30b3f),
	.w7(32'h3b287c4a),
	.w8(32'h3b55f493),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a24e0),
	.w1(32'h3b06670d),
	.w2(32'h3a80d0fd),
	.w3(32'h3a985d0a),
	.w4(32'h3a8a73f7),
	.w5(32'hba468975),
	.w6(32'h3ad62128),
	.w7(32'h3b2e2615),
	.w8(32'h3aef2a79),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e4bc2),
	.w1(32'h3ae8e86f),
	.w2(32'h39ae8437),
	.w3(32'hba6848c8),
	.w4(32'hbb3a4ab8),
	.w5(32'hbb36900b),
	.w6(32'h3b03a45f),
	.w7(32'hba963c80),
	.w8(32'h3aa525f6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ec7d),
	.w1(32'h3bb55377),
	.w2(32'h3bca8a88),
	.w3(32'h39abed82),
	.w4(32'h3af81683),
	.w5(32'h3a94f254),
	.w6(32'h3bb9b315),
	.w7(32'h3baddaca),
	.w8(32'h3b919107),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9188c),
	.w1(32'h3ada47c5),
	.w2(32'h3ae68936),
	.w3(32'h3a2d4923),
	.w4(32'hbb52f89f),
	.w5(32'hbb9c0398),
	.w6(32'hbb4fd6fb),
	.w7(32'hbad8772e),
	.w8(32'hbacd0b9f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8e552),
	.w1(32'h3b7cd2ce),
	.w2(32'h3be06e66),
	.w3(32'hbb22dee1),
	.w4(32'h3ad91eaa),
	.w5(32'h3b8f1a3d),
	.w6(32'h3b598801),
	.w7(32'h3b91cb80),
	.w8(32'h3bfdb3d3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b368944),
	.w1(32'h3aef0935),
	.w2(32'h3b51bd83),
	.w3(32'h3a407d9c),
	.w4(32'hb8490f9a),
	.w5(32'h3aa34958),
	.w6(32'h3a365cdc),
	.w7(32'h3aff5bb6),
	.w8(32'h3b4a5aea),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c243ce),
	.w1(32'hbad6b3b2),
	.w2(32'hbad6846e),
	.w3(32'hb9ebe225),
	.w4(32'hba8a8e8a),
	.w5(32'hbaa22a48),
	.w6(32'hbaacccbe),
	.w7(32'hba9ee8ec),
	.w8(32'h39e71e01),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc6543),
	.w1(32'h3a6c0d8e),
	.w2(32'h39c875ff),
	.w3(32'h3941329f),
	.w4(32'h39f0058a),
	.w5(32'h3a5408bc),
	.w6(32'h399d09d7),
	.w7(32'h38bf10b8),
	.w8(32'h3a579903),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a538dd8),
	.w1(32'hba3c8122),
	.w2(32'hbb3541e6),
	.w3(32'h39d7dc87),
	.w4(32'hbb436308),
	.w5(32'hbb5b13ef),
	.w6(32'hbb124867),
	.w7(32'hbb23455b),
	.w8(32'hbb94d57d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3422ed),
	.w1(32'h3bfae489),
	.w2(32'h3c884704),
	.w3(32'h3b6c74c6),
	.w4(32'hbb7b8445),
	.w5(32'h3b956ea0),
	.w6(32'hbaff01f6),
	.w7(32'h3b9c1ae7),
	.w8(32'h3c1c4e93),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c203718),
	.w1(32'h3b689f34),
	.w2(32'h3b82c630),
	.w3(32'h39555072),
	.w4(32'h381e0ed4),
	.w5(32'h378e9032),
	.w6(32'h3b3f477b),
	.w7(32'h3b3944bf),
	.w8(32'h3af3b51e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95edb5),
	.w1(32'hbb47b08d),
	.w2(32'hbb898165),
	.w3(32'h3b13e05c),
	.w4(32'hbb25513f),
	.w5(32'hbbb85dc2),
	.w6(32'h3b43762b),
	.w7(32'h3975e62d),
	.w8(32'hbb8aa794),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9384d4),
	.w1(32'h38de6962),
	.w2(32'h397d71f3),
	.w3(32'hbac26360),
	.w4(32'hbb2e979c),
	.w5(32'hbb4e1382),
	.w6(32'hbb9529ac),
	.w7(32'hbb66ce59),
	.w8(32'hbb17c0b9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b4d5),
	.w1(32'hba0ecf7a),
	.w2(32'hba6894f4),
	.w3(32'hbb721bd0),
	.w4(32'hb9059d21),
	.w5(32'hba161828),
	.w6(32'hba3e8b7a),
	.w7(32'hba4f4d7c),
	.w8(32'hb94814e3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa8b6f),
	.w1(32'hbb80f29d),
	.w2(32'hba4cefa0),
	.w3(32'h3a81f534),
	.w4(32'hbae08afa),
	.w5(32'hbb20f17a),
	.w6(32'h3abff326),
	.w7(32'h3b1c7d67),
	.w8(32'hba7355ea),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963c960),
	.w1(32'hbaeb7493),
	.w2(32'h3b7c76e9),
	.w3(32'hba4952a8),
	.w4(32'hbbab8189),
	.w5(32'h3a0390d2),
	.w6(32'hbbb0308f),
	.w7(32'h39e96677),
	.w8(32'h39c3447b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc44b78),
	.w1(32'h3b501e58),
	.w2(32'h379c592f),
	.w3(32'hbad01e13),
	.w4(32'hbae629d8),
	.w5(32'hbbd503b8),
	.w6(32'h3b849c99),
	.w7(32'h3b2d0bca),
	.w8(32'hbbb12272),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900f0f),
	.w1(32'h3a2ee17b),
	.w2(32'h3840ea85),
	.w3(32'hbb4b398e),
	.w4(32'h3978a5cb),
	.w5(32'h39a1a248),
	.w6(32'h3a0b9801),
	.w7(32'h38a0542f),
	.w8(32'h39fe7869),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f05e3d),
	.w1(32'h3a5a0e7a),
	.w2(32'h39a483b4),
	.w3(32'h39ff06f7),
	.w4(32'h399263b1),
	.w5(32'h39b2ec22),
	.w6(32'h3933488d),
	.w7(32'hb916a887),
	.w8(32'hba05bd89),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7847d),
	.w1(32'hbae7bcc5),
	.w2(32'hba6e6974),
	.w3(32'h37569ef4),
	.w4(32'hbad93da8),
	.w5(32'hba71ab3e),
	.w6(32'hbb18d2eb),
	.w7(32'hbaa035b7),
	.w8(32'h3a16aa0c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4ea6e),
	.w1(32'hbae12eea),
	.w2(32'h3c220a27),
	.w3(32'h38e92c97),
	.w4(32'hbb12c4a3),
	.w5(32'h3c11678e),
	.w6(32'hbb11c360),
	.w7(32'h3c320e80),
	.w8(32'hbb4d3262),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bfceb),
	.w1(32'h3a85120d),
	.w2(32'h3ad44da0),
	.w3(32'hbbb3e736),
	.w4(32'hba3db40a),
	.w5(32'h3a428b94),
	.w6(32'h3a8e3fc2),
	.w7(32'h3ad27b4c),
	.w8(32'h3aee3cc6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a26d3),
	.w1(32'hbabd4f9f),
	.w2(32'hb91df6dd),
	.w3(32'hbaae0813),
	.w4(32'hba006ac7),
	.w5(32'h3a5618dc),
	.w6(32'hbacfc3b4),
	.w7(32'hba9a3795),
	.w8(32'h3a97089b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83092b),
	.w1(32'hbbcc74da),
	.w2(32'h3bf190c3),
	.w3(32'h3b29a956),
	.w4(32'hbb80e66f),
	.w5(32'h39dff04e),
	.w6(32'h3a4d3de9),
	.w7(32'hbaf9162a),
	.w8(32'h3bb8e54c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211493),
	.w1(32'hbb602044),
	.w2(32'hbb8e10e9),
	.w3(32'hbaa1f40a),
	.w4(32'hbb9aa58a),
	.w5(32'hbc10e7bc),
	.w6(32'h3b05165c),
	.w7(32'hbb758999),
	.w8(32'hbc0035e2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e3bc1),
	.w1(32'h3aac8497),
	.w2(32'hbabac00d),
	.w3(32'hb8ef0ed3),
	.w4(32'hbaa5b4c9),
	.w5(32'hbbae5da1),
	.w6(32'h38c4702d),
	.w7(32'hbb47e735),
	.w8(32'hbbd35d10),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67a74c),
	.w1(32'hbad282f2),
	.w2(32'hbac4f5fa),
	.w3(32'h3965ec5e),
	.w4(32'hbb0a2cde),
	.w5(32'hbb2f0c6d),
	.w6(32'h3a17118d),
	.w7(32'hba871b88),
	.w8(32'hbab8491e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e868d),
	.w1(32'h3c1ff213),
	.w2(32'h3c18485d),
	.w3(32'hba7e79a9),
	.w4(32'h3bacfcea),
	.w5(32'h3b828a86),
	.w6(32'h3bc60192),
	.w7(32'h3bb22763),
	.w8(32'hbade11f8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75ded6),
	.w1(32'hba7898d3),
	.w2(32'hba433d89),
	.w3(32'hbb9dd443),
	.w4(32'hba7792c0),
	.w5(32'hba8de225),
	.w6(32'h3a691078),
	.w7(32'h39e0e3f7),
	.w8(32'hb988d7d5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1214e5),
	.w1(32'h38ea2837),
	.w2(32'h3969be69),
	.w3(32'hbaaa7dcd),
	.w4(32'hba410d43),
	.w5(32'hba0a6f6b),
	.w6(32'hba3de42f),
	.w7(32'hb935141e),
	.w8(32'hb630b9d9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b820993),
	.w1(32'h3bc6058e),
	.w2(32'h3bf2f1ee),
	.w3(32'h3afbfc0c),
	.w4(32'hbae1db0a),
	.w5(32'hba737d9e),
	.w6(32'h3bdda65e),
	.w7(32'h3b90962e),
	.w8(32'h3bea8052),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfc50f),
	.w1(32'h3ac9c619),
	.w2(32'h39dc04a7),
	.w3(32'hb72cb837),
	.w4(32'h39173dd7),
	.w5(32'hba3cae58),
	.w6(32'h3b42bec4),
	.w7(32'h3abf1dba),
	.w8(32'h39fc7819),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00c1d2),
	.w1(32'h3b2a1e18),
	.w2(32'h3b502d6f),
	.w3(32'h3b8c14d8),
	.w4(32'hb93176c3),
	.w5(32'hb994f249),
	.w6(32'h3b20c309),
	.w7(32'h3b200a5f),
	.w8(32'h3ac6cdb4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c9aa),
	.w1(32'h3abeaac9),
	.w2(32'h3af3872a),
	.w3(32'h3b7b14c8),
	.w4(32'hbb291e0d),
	.w5(32'hbb109cfb),
	.w6(32'h3b0e34c8),
	.w7(32'h3a22b136),
	.w8(32'h3b0e8382),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a37c8e),
	.w1(32'h3afe86cb),
	.w2(32'h3c70f980),
	.w3(32'hbbc76d48),
	.w4(32'hbbaea813),
	.w5(32'h3be8e454),
	.w6(32'hbbf60853),
	.w7(32'h3b9fb661),
	.w8(32'h3baebffb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b926158),
	.w1(32'hba20209d),
	.w2(32'hb989d96b),
	.w3(32'hba598ef1),
	.w4(32'hba971aef),
	.w5(32'hba3d4c88),
	.w6(32'hbaa16d3c),
	.w7(32'hba0865a2),
	.w8(32'hba59ab63),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91709c8),
	.w1(32'h3984c01e),
	.w2(32'hb974581d),
	.w3(32'hba2f0d2d),
	.w4(32'hb97e3b99),
	.w5(32'hba9645cf),
	.w6(32'h3a3e177b),
	.w7(32'h368a0d14),
	.w8(32'h39e67e10),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9446e23),
	.w1(32'h38b24e0e),
	.w2(32'h3acb3a8a),
	.w3(32'hba6a6924),
	.w4(32'hba2d81cc),
	.w5(32'h3869be14),
	.w6(32'h3a054e14),
	.w7(32'h3a98f9e7),
	.w8(32'h3ab0cb1a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7f56e),
	.w1(32'hbb2d82a4),
	.w2(32'h3b2673a9),
	.w3(32'h3a9e476a),
	.w4(32'hbac96909),
	.w5(32'h3aa1166b),
	.w6(32'hba8c4829),
	.w7(32'h3a2669b2),
	.w8(32'h3b33f2d9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71a2a7),
	.w1(32'h3b3b1fb0),
	.w2(32'h3a86a1a7),
	.w3(32'h3b0c6fad),
	.w4(32'h3ae16dfb),
	.w5(32'hb8619757),
	.w6(32'h3aa4421c),
	.w7(32'hb813c2b1),
	.w8(32'hba70df91),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f5b86),
	.w1(32'h3befcaf8),
	.w2(32'h3c0e760c),
	.w3(32'hba85802d),
	.w4(32'h3a632b86),
	.w5(32'h3b76a537),
	.w6(32'h3ad409fc),
	.w7(32'h3b4a4628),
	.w8(32'h3c0a3eb5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44de9b),
	.w1(32'hb924087e),
	.w2(32'h3a257672),
	.w3(32'h39cbf284),
	.w4(32'hbb185da8),
	.w5(32'hbafabb64),
	.w6(32'hbb0a797a),
	.w7(32'hbaec3ef3),
	.w8(32'hbae583a5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7eb752),
	.w1(32'h3bc7df36),
	.w2(32'hbb545ff2),
	.w3(32'hbb8b33cb),
	.w4(32'h3b94f7ba),
	.w5(32'hbbb53a62),
	.w6(32'h3bf91cb6),
	.w7(32'hbaba5f69),
	.w8(32'hba9b5b36),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b86531),
	.w1(32'h3b494ada),
	.w2(32'h3b8e0624),
	.w3(32'hbb9f18cc),
	.w4(32'h3a99a521),
	.w5(32'h3ab12e6d),
	.w6(32'h3aa0080f),
	.w7(32'h3adee1e9),
	.w8(32'hbaaf2599),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b036bf4),
	.w1(32'hb825d77a),
	.w2(32'h3b0b22f8),
	.w3(32'hbac71e8f),
	.w4(32'hb94faee8),
	.w5(32'hba176cb1),
	.w6(32'h3ad3dfa5),
	.w7(32'hb9b80f29),
	.w8(32'h3b1b8af4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a964f52),
	.w1(32'hbaf43433),
	.w2(32'hbab77dd0),
	.w3(32'hb874dff5),
	.w4(32'hbb2ab7d0),
	.w5(32'hbb12e0eb),
	.w6(32'hba6fbd3d),
	.w7(32'hb9c0cb49),
	.w8(32'h39b51538),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a91ca8),
	.w1(32'hb9e1ca8f),
	.w2(32'hb794b9d2),
	.w3(32'hba4b50cf),
	.w4(32'hba71dee9),
	.w5(32'hb9e63364),
	.w6(32'hb9778b96),
	.w7(32'h3924a094),
	.w8(32'h3a2f8d5d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd1c2b),
	.w1(32'h39801a58),
	.w2(32'h3b0456a7),
	.w3(32'hba1b8245),
	.w4(32'hbafbce17),
	.w5(32'hb85a1864),
	.w6(32'hba11770f),
	.w7(32'h38f027ff),
	.w8(32'h3afa6b99),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b047d35),
	.w1(32'h3ada979d),
	.w2(32'h3b6faeb9),
	.w3(32'h3a69ee7d),
	.w4(32'h3a426b09),
	.w5(32'h3b0a7630),
	.w6(32'h3b798413),
	.w7(32'h3b461341),
	.w8(32'h3b7e43f1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53bc81),
	.w1(32'hbb817c78),
	.w2(32'h3a0a2eac),
	.w3(32'h3721694b),
	.w4(32'hbb0767cb),
	.w5(32'h3b220f9e),
	.w6(32'hbb654af4),
	.w7(32'h3ad973e2),
	.w8(32'h3a0e0a97),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae12f6c),
	.w1(32'h3992ffd4),
	.w2(32'hb9b68a1a),
	.w3(32'h3a888e28),
	.w4(32'hba9c0702),
	.w5(32'hbb0b77a1),
	.w6(32'h3a911a98),
	.w7(32'h3a509286),
	.w8(32'h3aab0f89),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989c234),
	.w1(32'hba8c3c84),
	.w2(32'hba8b5df1),
	.w3(32'hbaaa09e3),
	.w4(32'hba6f7ddd),
	.w5(32'hba49fc5e),
	.w6(32'hba533589),
	.w7(32'hb9dcbf38),
	.w8(32'hbaa174f1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2be78),
	.w1(32'hbab19d9c),
	.w2(32'h3b0efbb4),
	.w3(32'hba40f0b3),
	.w4(32'hbaed0f78),
	.w5(32'hb934a0b3),
	.w6(32'hba75ff79),
	.w7(32'h3a0c8e63),
	.w8(32'h39d39003),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aa028),
	.w1(32'h3c808aed),
	.w2(32'h3c8abf31),
	.w3(32'hbad104ee),
	.w4(32'h3bcef511),
	.w5(32'h3bc93546),
	.w6(32'h3bc72361),
	.w7(32'h3c0ab296),
	.w8(32'h3bb6ca1b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f2285),
	.w1(32'h3c33e990),
	.w2(32'h3cb952cd),
	.w3(32'hbb86c714),
	.w4(32'h3b549f22),
	.w5(32'h3c7d9d21),
	.w6(32'h39e53d35),
	.w7(32'h3c3a32f9),
	.w8(32'h3b345fe3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29c1ea),
	.w1(32'h3bc7a026),
	.w2(32'h3bc51628),
	.w3(32'hbb3af462),
	.w4(32'h3b7dbce6),
	.w5(32'h3b8d6456),
	.w6(32'h3b470a93),
	.w7(32'h3b4c142f),
	.w8(32'h3bbb3b62),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9d114),
	.w1(32'hbaaef1f0),
	.w2(32'hbac9ea41),
	.w3(32'h3b49a32e),
	.w4(32'hbb029895),
	.w5(32'hbbbd31ad),
	.w6(32'h3bfd4ea0),
	.w7(32'h3b189cb7),
	.w8(32'hbacc4f87),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b28d6),
	.w1(32'hb9568363),
	.w2(32'hb636a9e2),
	.w3(32'h39cb2e03),
	.w4(32'hb9995894),
	.w5(32'hb9f991a3),
	.w6(32'h3a18970e),
	.w7(32'h3a21894f),
	.w8(32'h3a7dd096),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58eba3),
	.w1(32'h3a53bb8a),
	.w2(32'h39c6e1c3),
	.w3(32'hb8dd2105),
	.w4(32'h39f2ab7c),
	.w5(32'hb99a1a70),
	.w6(32'h3a60eaa1),
	.w7(32'h397ff035),
	.w8(32'h3a05087f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfde9a),
	.w1(32'hb9bf373d),
	.w2(32'hb9a4bf0e),
	.w3(32'hb981113b),
	.w4(32'hba15fe8c),
	.w5(32'hba095ac5),
	.w6(32'hb8ed9e9e),
	.w7(32'hb91a4a49),
	.w8(32'h399233ce),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370b2bb5),
	.w1(32'h3a9470a7),
	.w2(32'h3aafd6a9),
	.w3(32'hb9f6bf9f),
	.w4(32'hb9af3331),
	.w5(32'h3a4db040),
	.w6(32'hba2b270a),
	.w7(32'hba210d76),
	.w8(32'h39e8d625),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97054c0),
	.w1(32'hbb0dee22),
	.w2(32'hbb02206b),
	.w3(32'hb9a379cf),
	.w4(32'hbadfa1c6),
	.w5(32'hbaebee9b),
	.w6(32'hbaa8f019),
	.w7(32'hba72a805),
	.w8(32'hba3dd802),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba977581),
	.w1(32'h3a33fe4d),
	.w2(32'h3b076e8e),
	.w3(32'hbb123ec7),
	.w4(32'hbadf4230),
	.w5(32'hba9bfb63),
	.w6(32'hbb1d4c58),
	.w7(32'hbb168a57),
	.w8(32'h3a88592c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4fe4f),
	.w1(32'hb9531e88),
	.w2(32'h3ba1eadf),
	.w3(32'hbb7064b5),
	.w4(32'hbb2ef6bb),
	.w5(32'h3ae8e72d),
	.w6(32'h39e22f6e),
	.w7(32'h38e69548),
	.w8(32'h3b9888cc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b821aee),
	.w1(32'hba2d7ab3),
	.w2(32'hbad84915),
	.w3(32'hb7eeb70c),
	.w4(32'hbacbee8c),
	.w5(32'hbb52565a),
	.w6(32'h3acf2c71),
	.w7(32'h39a367a1),
	.w8(32'hbad8607a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a951ab1),
	.w1(32'h3ac143f4),
	.w2(32'h3b8b0457),
	.w3(32'hb9dca39b),
	.w4(32'hbb664e88),
	.w5(32'hbb1198ae),
	.w6(32'hbb6c4376),
	.w7(32'hbab0d635),
	.w8(32'h39a00451),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba318b3b),
	.w1(32'h3ad68e6f),
	.w2(32'h3b6f0615),
	.w3(32'hbb82919c),
	.w4(32'hba704bc9),
	.w5(32'h3aa5acad),
	.w6(32'h392336e2),
	.w7(32'h3ad08635),
	.w8(32'h3b70f1fd),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d581e),
	.w1(32'h3bf4dba9),
	.w2(32'h3c4924ad),
	.w3(32'h3aac6f42),
	.w4(32'h3b8d7b79),
	.w5(32'h3c1bfd0d),
	.w6(32'h3b457c91),
	.w7(32'h3c02bf26),
	.w8(32'hbb8326a4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f09279),
	.w1(32'hba5f6b8f),
	.w2(32'h3a9a13a1),
	.w3(32'hbbb05277),
	.w4(32'hbb0a69be),
	.w5(32'hba36db6d),
	.w6(32'hbae80bb5),
	.w7(32'hb99963db),
	.w8(32'hb9418895),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4ca61),
	.w1(32'hba067063),
	.w2(32'hba8e299b),
	.w3(32'hbaf489c5),
	.w4(32'hba092a2e),
	.w5(32'hbaeb1e6d),
	.w6(32'hba0eaf40),
	.w7(32'hba3d7652),
	.w8(32'hb94b7582),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a639ee3),
	.w1(32'hba8fbe58),
	.w2(32'hba81240e),
	.w3(32'hba7075e7),
	.w4(32'hba9fe19b),
	.w5(32'hba9b9d0a),
	.w6(32'hba28aebd),
	.w7(32'hb9bc8bfb),
	.w8(32'hba26fc4c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48cd15),
	.w1(32'hba259321),
	.w2(32'h3c7f0e62),
	.w3(32'hba1cfcb9),
	.w4(32'hbb329698),
	.w5(32'h3c572568),
	.w6(32'hbb119045),
	.w7(32'h3c51e0da),
	.w8(32'hbb713f55),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53aa2a),
	.w1(32'h39978102),
	.w2(32'hb9e79fba),
	.w3(32'hbaf2b799),
	.w4(32'h3a162a0e),
	.w5(32'hbacf01f5),
	.w6(32'h3a441bfd),
	.w7(32'hba6132db),
	.w8(32'hbb25d19b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eb1e3),
	.w1(32'hba391c91),
	.w2(32'h37436a2c),
	.w3(32'h3a1ca452),
	.w4(32'hba408687),
	.w5(32'hbabf711b),
	.w6(32'h3b07e401),
	.w7(32'h390830b5),
	.w8(32'h3a2844f3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77073d),
	.w1(32'h39a6a2de),
	.w2(32'h379c55b4),
	.w3(32'hb8253b91),
	.w4(32'hb93e2d67),
	.w5(32'h38e7b4e9),
	.w6(32'h39f6187a),
	.w7(32'hb961b8ab),
	.w8(32'h3a15cccc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98494a),
	.w1(32'h3ac47305),
	.w2(32'h3a5cfb10),
	.w3(32'h3b7d13e3),
	.w4(32'hb9e91197),
	.w5(32'hbb13befd),
	.w6(32'h3b3856e9),
	.w7(32'h3ae41009),
	.w8(32'hbaa7aa4e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24549d),
	.w1(32'h3b6d95b8),
	.w2(32'h3baf74ba),
	.w3(32'hbbba6f85),
	.w4(32'h391d9850),
	.w5(32'h3b19c640),
	.w6(32'h39653fe4),
	.w7(32'h3aa7611f),
	.w8(32'h3b6541a0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2992db),
	.w1(32'h39d621a7),
	.w2(32'hbaf95f5e),
	.w3(32'h3a65f0f3),
	.w4(32'hba9a3291),
	.w5(32'hbb669c7d),
	.w6(32'hb9443712),
	.w7(32'hbb33fdfd),
	.w8(32'hbba6359a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3625a9),
	.w1(32'h3b656c54),
	.w2(32'h3c2af274),
	.w3(32'hbb41cdef),
	.w4(32'hbaf81769),
	.w5(32'h3adb44a4),
	.w6(32'hb96d1b5b),
	.w7(32'hb9b626e9),
	.w8(32'h3b9e030b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fcb2f),
	.w1(32'hba97e711),
	.w2(32'hbb6747b1),
	.w3(32'h3a902474),
	.w4(32'hbb0f8a2f),
	.w5(32'hbb9f449b),
	.w6(32'h3ac03d34),
	.w7(32'hbb51891f),
	.w8(32'hbbb0f204),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9068d0),
	.w1(32'h3c2481c3),
	.w2(32'h3c6be88b),
	.w3(32'hbab81903),
	.w4(32'h3b9d4fe2),
	.w5(32'h3beade74),
	.w6(32'h3b847f2a),
	.w7(32'h3c2c8453),
	.w8(32'h3b9c0dd0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7c967),
	.w1(32'h3b6effc0),
	.w2(32'h3b5989bc),
	.w3(32'h39f29a60),
	.w4(32'h3b0bb02c),
	.w5(32'h3a54df5c),
	.w6(32'h3b75be6b),
	.w7(32'h3b76a7ab),
	.w8(32'h3b2131ce),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82275c),
	.w1(32'h398a706d),
	.w2(32'hbb7d5027),
	.w3(32'h3a7c3f9c),
	.w4(32'hbad99292),
	.w5(32'hbbb04b4a),
	.w6(32'h3b768df7),
	.w7(32'h39091282),
	.w8(32'hbb8219fa),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf36ebf),
	.w1(32'hb98f2d07),
	.w2(32'h3bb61177),
	.w3(32'hba45f779),
	.w4(32'hbb0111bf),
	.w5(32'h3b7e3a42),
	.w6(32'hbb825c91),
	.w7(32'h3b6575d4),
	.w8(32'h39f26e0d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf100c5),
	.w1(32'h39c2d7da),
	.w2(32'h3c213d3b),
	.w3(32'hbab6b046),
	.w4(32'hbb0ea6d3),
	.w5(32'h3bbed7af),
	.w6(32'hba423117),
	.w7(32'h3bf1305c),
	.w8(32'h3bf0b4ce),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d4ba4),
	.w1(32'h3ae3a20e),
	.w2(32'h3bc6f9ca),
	.w3(32'h39a64e6f),
	.w4(32'hba9c63a0),
	.w5(32'h390ea1a6),
	.w6(32'hbb962954),
	.w7(32'h3a9b9172),
	.w8(32'h3b3a2d5c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c26ab),
	.w1(32'hbb96e5d6),
	.w2(32'h3ab8252d),
	.w3(32'h3a0c0952),
	.w4(32'hbb747440),
	.w5(32'h3b14f31d),
	.w6(32'h3b2f7321),
	.w7(32'hbb4ca4bd),
	.w8(32'h3b56d9c8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3564cc),
	.w1(32'hba8faa1c),
	.w2(32'hba8498a6),
	.w3(32'hbb116348),
	.w4(32'hbba40e8f),
	.w5(32'hbc104604),
	.w6(32'h3b582452),
	.w7(32'hbb45445b),
	.w8(32'hbb840723),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd779b9),
	.w1(32'h39ae6af5),
	.w2(32'hbb84a2ee),
	.w3(32'h3b0eeed4),
	.w4(32'hb91bb4ef),
	.w5(32'hbbae907b),
	.w6(32'h3b9afa8c),
	.w7(32'hba369fb0),
	.w8(32'hba8bc914),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39566083),
	.w1(32'h3b2a9cba),
	.w2(32'h3c12f525),
	.w3(32'hba25db7b),
	.w4(32'hbac852cc),
	.w5(32'h398b0536),
	.w6(32'h3a800e4d),
	.w7(32'h3b3841e0),
	.w8(32'h3bed25ec),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9df71c),
	.w1(32'h39af4afb),
	.w2(32'hb983da81),
	.w3(32'hbb61f581),
	.w4(32'hb85d4911),
	.w5(32'hba6d1969),
	.w6(32'h399c7b93),
	.w7(32'hba1d8b2e),
	.w8(32'hb9febb8d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af344d4),
	.w1(32'h3948b6c3),
	.w2(32'h3b859907),
	.w3(32'h3ba455e1),
	.w4(32'h3a8b4438),
	.w5(32'h3aa5a707),
	.w6(32'h3b9e3e1d),
	.w7(32'h3ba3f5c5),
	.w8(32'h3bae2c4f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cb309),
	.w1(32'hbb820388),
	.w2(32'hb915d45d),
	.w3(32'hbb731513),
	.w4(32'hbb774ab1),
	.w5(32'hba3d48ef),
	.w6(32'hbb9beea0),
	.w7(32'hbb7f22b7),
	.w8(32'h3a84b96e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a458b0d),
	.w1(32'hb9db8900),
	.w2(32'hba0872ae),
	.w3(32'h39ba6552),
	.w4(32'hba56ee40),
	.w5(32'hba5333ec),
	.w6(32'hb9c53e72),
	.w7(32'hb90756fb),
	.w8(32'hba8c46e8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b4e6d),
	.w1(32'h3aa5312b),
	.w2(32'h3a3df603),
	.w3(32'hba2dd2e3),
	.w4(32'hb8a815cf),
	.w5(32'h39e3830f),
	.w6(32'h3a9c284a),
	.w7(32'h3a7fc1ac),
	.w8(32'h3a6898a3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fcbb0),
	.w1(32'h3b13ffd3),
	.w2(32'h3b8418c9),
	.w3(32'hb99a1bb6),
	.w4(32'hbae5c028),
	.w5(32'hba1ac1df),
	.w6(32'h3a94a3ad),
	.w7(32'h3af026eb),
	.w8(32'h3b254409),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dbbe9),
	.w1(32'hb9d6b160),
	.w2(32'hbb1073af),
	.w3(32'hb9ae7cf3),
	.w4(32'hba3ae688),
	.w5(32'hbb1a2b6c),
	.w6(32'h3b1a4e76),
	.w7(32'hb9ed811e),
	.w8(32'hba5fa724),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ceac0),
	.w1(32'h3a038cd2),
	.w2(32'hba7d2860),
	.w3(32'h3b55853f),
	.w4(32'hb98eea59),
	.w5(32'hbb47bf8f),
	.w6(32'hb92cd9e5),
	.w7(32'hbad286dc),
	.w8(32'hbb72dd5e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b630c42),
	.w1(32'hbaf898ef),
	.w2(32'hb8af6cbc),
	.w3(32'h3b04464f),
	.w4(32'hbaa4f1ad),
	.w5(32'h38d43c2e),
	.w6(32'hbabd3fff),
	.w7(32'hb8ca3bd2),
	.w8(32'h3aa92d0b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6057d),
	.w1(32'hbb9ad5c9),
	.w2(32'hbb33cafb),
	.w3(32'hbaa4106e),
	.w4(32'hbb60ad93),
	.w5(32'hba6a6acd),
	.w6(32'hb93c7909),
	.w7(32'hbabffadd),
	.w8(32'hb92d21cc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b516127),
	.w1(32'h3bd31032),
	.w2(32'h3bc29ee8),
	.w3(32'h3b1aed90),
	.w4(32'h3b1684f8),
	.w5(32'h3b1086eb),
	.w6(32'h3b93cbdc),
	.w7(32'h3ba60ea9),
	.w8(32'h3bcc6726),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68b98d),
	.w1(32'h3b44b2cb),
	.w2(32'h3b3dce60),
	.w3(32'h3aa4f7b3),
	.w4(32'h3a8de26e),
	.w5(32'h3a6a8fb9),
	.w6(32'h3b329cfc),
	.w7(32'h3b10d186),
	.w8(32'h38a60699),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae592d4),
	.w1(32'h397e329b),
	.w2(32'h39518f1a),
	.w3(32'h3a819959),
	.w4(32'hbaa39b77),
	.w5(32'hbacec93a),
	.w6(32'h3a4a4230),
	.w7(32'h3a4c6834),
	.w8(32'h39f6801d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93748ee),
	.w1(32'h3a3b507e),
	.w2(32'h3a3fb445),
	.w3(32'hbb097bf6),
	.w4(32'h391e9444),
	.w5(32'hb981bc47),
	.w6(32'h3a80caf8),
	.w7(32'h3a7d7e08),
	.w8(32'h39eba8f3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc6760),
	.w1(32'h39768088),
	.w2(32'hb9ec97e7),
	.w3(32'hba844d13),
	.w4(32'hb9abe475),
	.w5(32'hba72ac73),
	.w6(32'h3a08c0d1),
	.w7(32'hb7a1684b),
	.w8(32'hb8ac86a1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16a29a),
	.w1(32'h3a4ac4e7),
	.w2(32'hba361b53),
	.w3(32'hba9ed0be),
	.w4(32'h392f6e73),
	.w5(32'h3a181fd9),
	.w6(32'hb9c890a5),
	.w7(32'h399cfce6),
	.w8(32'h39c64bfa),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b363c3e),
	.w1(32'hb9834a4c),
	.w2(32'h3b676db8),
	.w3(32'h3aecea40),
	.w4(32'hbac9551b),
	.w5(32'h39c04e0c),
	.w6(32'h399306cc),
	.w7(32'h3b1d3829),
	.w8(32'h3abfe373),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03f615),
	.w1(32'h3a06f20b),
	.w2(32'hba6a32b2),
	.w3(32'h3a0c2ab3),
	.w4(32'h3916e45a),
	.w5(32'hb89171c1),
	.w6(32'hb9f713cf),
	.w7(32'hbab4ff76),
	.w8(32'hba8bde11),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7851cee),
	.w1(32'hb8b179cf),
	.w2(32'h3a9323da),
	.w3(32'hba68cced),
	.w4(32'hb9a41491),
	.w5(32'h38b9d920),
	.w6(32'hba7f41dd),
	.w7(32'hba8d41a8),
	.w8(32'h3b08173b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5be85a),
	.w1(32'h3a9cbee5),
	.w2(32'hbac2fdfa),
	.w3(32'h3b0343af),
	.w4(32'h3982981c),
	.w5(32'hbb4d04be),
	.w6(32'h3b2a68a1),
	.w7(32'h3ac4c6a1),
	.w8(32'hbb1e77ee),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7103b13),
	.w1(32'h3ae00d35),
	.w2(32'h393824f3),
	.w3(32'hba0bcd42),
	.w4(32'h3a70ad42),
	.w5(32'h3ac52e9b),
	.w6(32'h3a376fad),
	.w7(32'h3ac0dab4),
	.w8(32'h3b0c74da),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8483b4),
	.w1(32'h3b40147b),
	.w2(32'h3a239ace),
	.w3(32'h3b1b276f),
	.w4(32'h3ac2fcdc),
	.w5(32'h38a45480),
	.w6(32'h3ad5bce5),
	.w7(32'h39d2fd76),
	.w8(32'hbb06c2a7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf1e21),
	.w1(32'h3986e958),
	.w2(32'hb909ddfb),
	.w3(32'hbb0e954c),
	.w4(32'h38a79428),
	.w5(32'h392df59e),
	.w6(32'hb7cc8cbd),
	.w7(32'hb9922e22),
	.w8(32'h3a3011d1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61bc50),
	.w1(32'h3c0b2d65),
	.w2(32'h3b33fdd7),
	.w3(32'h3a522476),
	.w4(32'h3c693305),
	.w5(32'h396a525f),
	.w6(32'h3c0bf4dc),
	.w7(32'hb95507bf),
	.w8(32'h3b72fe75),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14ad99),
	.w1(32'hbbcba0de),
	.w2(32'h3ade48ca),
	.w3(32'hbb0cfb03),
	.w4(32'hbb555272),
	.w5(32'hbc0ea27a),
	.w6(32'h3a00cdf2),
	.w7(32'hbadfea2d),
	.w8(32'h3ad4239c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdea308),
	.w1(32'h3c2f546c),
	.w2(32'h3c212966),
	.w3(32'hbc9cec82),
	.w4(32'hbbe478d4),
	.w5(32'hbbd86261),
	.w6(32'h3b3d54dd),
	.w7(32'hbbb04c0a),
	.w8(32'h3a940600),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3e130),
	.w1(32'h3b6a2b62),
	.w2(32'h3bf89144),
	.w3(32'h3b848554),
	.w4(32'h3a7e5e84),
	.w5(32'h3c52650b),
	.w6(32'hba25344c),
	.w7(32'hbadd7656),
	.w8(32'h3a2262ff),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befe03c),
	.w1(32'hbbc6250b),
	.w2(32'hb9cf1cef),
	.w3(32'h3b6fa96f),
	.w4(32'hbabf3a5a),
	.w5(32'h3c0ff9c1),
	.w6(32'hbbe138bf),
	.w7(32'hbb6853a1),
	.w8(32'h3aed52d6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3669c4),
	.w1(32'h3b34850f),
	.w2(32'h3b1abc04),
	.w3(32'h3b14dbf5),
	.w4(32'hbbc42a1a),
	.w5(32'hbcab4309),
	.w6(32'h3b8f78eb),
	.w7(32'hba286414),
	.w8(32'hbbd9b9a1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed5c1c),
	.w1(32'hbb18d1a0),
	.w2(32'h3c330239),
	.w3(32'hbcb8403e),
	.w4(32'h3b3703eb),
	.w5(32'h3c07946c),
	.w6(32'h3ba6ccd9),
	.w7(32'h3be774fb),
	.w8(32'h3ae861bd),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27e0f9),
	.w1(32'hbc028ef8),
	.w2(32'hbc1d0456),
	.w3(32'hbc46d1a7),
	.w4(32'hbc409303),
	.w5(32'hbce822db),
	.w6(32'hb99ff13e),
	.w7(32'hbbcca5ec),
	.w8(32'hbc1ac63f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90869c),
	.w1(32'h3c0069e8),
	.w2(32'h3c224e62),
	.w3(32'hbd186938),
	.w4(32'h3b13345e),
	.w5(32'h3c60aa87),
	.w6(32'hbbaa1b39),
	.w7(32'hbb46e3dc),
	.w8(32'h391d6e79),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff0b15),
	.w1(32'hbaa4b47d),
	.w2(32'h3b6a07e7),
	.w3(32'h3b3978d1),
	.w4(32'h3b8e1160),
	.w5(32'hbbabe73e),
	.w6(32'h3c00f8a9),
	.w7(32'h3b81da48),
	.w8(32'h3b4f1825),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b206e50),
	.w1(32'hb8c2c7e6),
	.w2(32'h3b09b351),
	.w3(32'hbadbbc18),
	.w4(32'hbb56e8e5),
	.w5(32'hbbac3048),
	.w6(32'h3a3e9348),
	.w7(32'hba91bdd5),
	.w8(32'h39ae02fb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95d8cb),
	.w1(32'hbb1f1782),
	.w2(32'hbb9c6a75),
	.w3(32'hbbec14c3),
	.w4(32'hbb1307d7),
	.w5(32'h3c881796),
	.w6(32'hbc15bf73),
	.w7(32'hbbbb88bd),
	.w8(32'hba24def0),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd1197),
	.w1(32'hbb6629c5),
	.w2(32'hb9dba247),
	.w3(32'h3c793069),
	.w4(32'hba032bb4),
	.w5(32'h3aed597b),
	.w6(32'h3ba6208c),
	.w7(32'h3b4ac166),
	.w8(32'h397c38cd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920cfb),
	.w1(32'hbbf5a8ff),
	.w2(32'hbac0fcd0),
	.w3(32'h3b7f7f0c),
	.w4(32'hbb0a0820),
	.w5(32'hbb04ffc3),
	.w6(32'hb9b5e548),
	.w7(32'hbc1fbb47),
	.w8(32'hbb9a6e3f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc124f1a),
	.w1(32'h3c230ec3),
	.w2(32'h3c585d74),
	.w3(32'hbb2d88a3),
	.w4(32'h3c2c8264),
	.w5(32'h3bc9a3b5),
	.w6(32'h3bccf197),
	.w7(32'h3b9b8951),
	.w8(32'h3b9fb8e9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c412c14),
	.w1(32'hbc919e26),
	.w2(32'hbbfa0742),
	.w3(32'h3c0abfe6),
	.w4(32'hba1d7424),
	.w5(32'h3905af9f),
	.w6(32'hbbda38bf),
	.w7(32'hbbaf8312),
	.w8(32'hbb09df6d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32549a),
	.w1(32'hbbe0963f),
	.w2(32'h3be46338),
	.w3(32'h3cc16204),
	.w4(32'hbc1cb345),
	.w5(32'h3c558602),
	.w6(32'h3ba144bd),
	.w7(32'hbbc97860),
	.w8(32'hbc1520c9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa4fe1),
	.w1(32'hbc0953fe),
	.w2(32'hbbbd9162),
	.w3(32'h3b4d5a7b),
	.w4(32'hbc0bc119),
	.w5(32'hbc43f3ad),
	.w6(32'hbc13e513),
	.w7(32'hbc0b87e8),
	.w8(32'hbbed2e3b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc066424),
	.w1(32'h3b7a2d1e),
	.w2(32'h3b939c1f),
	.w3(32'hbc2fb23c),
	.w4(32'h3ba86cc3),
	.w5(32'h3ba7d94f),
	.w6(32'h3c08bc24),
	.w7(32'h3bc21404),
	.w8(32'h3bc0f58c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b2f32),
	.w1(32'h3b2b5b36),
	.w2(32'hba837077),
	.w3(32'hbbddb6d0),
	.w4(32'h3aeee055),
	.w5(32'h3c6b9e94),
	.w6(32'hbc025ca9),
	.w7(32'hbbd0fdb6),
	.w8(32'hbb4b8b27),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa018d),
	.w1(32'h3aa1a5ce),
	.w2(32'h3bb73b29),
	.w3(32'h3c3187bc),
	.w4(32'h3b5cc1a2),
	.w5(32'h3c71a5a0),
	.w6(32'hbaccae62),
	.w7(32'hbb3e61f4),
	.w8(32'hbb9239f6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb29759),
	.w1(32'hbb0f2b91),
	.w2(32'hb9d15a11),
	.w3(32'h3c0f15cc),
	.w4(32'hbbc7894a),
	.w5(32'hbbf46ff6),
	.w6(32'hbb2acf51),
	.w7(32'hbb7d9d70),
	.w8(32'hbb278be2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7cc6),
	.w1(32'hb9c5a3d6),
	.w2(32'hbad222e9),
	.w3(32'hbb98d9bf),
	.w4(32'h3b59f716),
	.w5(32'hbb1f33c6),
	.w6(32'h3ba1bd92),
	.w7(32'h3a98af8a),
	.w8(32'h3b665a31),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5813ac),
	.w1(32'hbc914d90),
	.w2(32'hbacaf043),
	.w3(32'h3af303c5),
	.w4(32'hbc3428ec),
	.w5(32'h3badd284),
	.w6(32'hbae4eda3),
	.w7(32'h3b8d9d47),
	.w8(32'h3c0c0df2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be36074),
	.w1(32'hba0d44b6),
	.w2(32'h3b06ffea),
	.w3(32'h3caccbb1),
	.w4(32'h39c0973e),
	.w5(32'hbb38ca3b),
	.w6(32'h3b266784),
	.w7(32'h3bbee61b),
	.w8(32'h3bde5f5a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a043f99),
	.w1(32'h3acd5e55),
	.w2(32'h3c2ba8a1),
	.w3(32'hba766e67),
	.w4(32'h3b0fa4fd),
	.w5(32'hbb76e26c),
	.w6(32'h3b994bd2),
	.w7(32'h3ac7a49e),
	.w8(32'h3bba08fa),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13db7b),
	.w1(32'h3bec09f1),
	.w2(32'h3c0792f0),
	.w3(32'hbb9e8473),
	.w4(32'hba87e59f),
	.w5(32'h3a16a59d),
	.w6(32'h3bca6893),
	.w7(32'h3b241795),
	.w8(32'hbb0c4896),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b517460),
	.w1(32'hbb58c0a5),
	.w2(32'h3bf24b10),
	.w3(32'hbb37aab1),
	.w4(32'hbbaa9073),
	.w5(32'hbc00d860),
	.w6(32'h3b86005f),
	.w7(32'h3b8af943),
	.w8(32'h3aca8642),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b33d),
	.w1(32'hbb8c5ec8),
	.w2(32'hbb1cbbde),
	.w3(32'hbbf0a8b4),
	.w4(32'hbb24175d),
	.w5(32'hbbb21a26),
	.w6(32'hbb3c3f74),
	.w7(32'hbb6977f8),
	.w8(32'hbb0287b2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0a46f),
	.w1(32'h3b71957e),
	.w2(32'h3b2e82ea),
	.w3(32'hbb6f4564),
	.w4(32'hba463373),
	.w5(32'hbb92a0cf),
	.w6(32'h3b9b81ea),
	.w7(32'h3a983c29),
	.w8(32'hbae8bba1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942273),
	.w1(32'hbb802cc7),
	.w2(32'hbc2d9890),
	.w3(32'hbc3b67b8),
	.w4(32'h3ae42db3),
	.w5(32'hbbaa7f6e),
	.w6(32'h37ea321d),
	.w7(32'hbbf79c4c),
	.w8(32'hbb19e322),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45239c),
	.w1(32'hbbb630f9),
	.w2(32'hbb85a0a8),
	.w3(32'h3b84b343),
	.w4(32'hbb30c327),
	.w5(32'hba83a0f2),
	.w6(32'h3adfa073),
	.w7(32'hb87d1cc7),
	.w8(32'h3a5e80c2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe7747),
	.w1(32'hbaac85e7),
	.w2(32'h3aa067f1),
	.w3(32'h3b2f9fc5),
	.w4(32'h3938a32d),
	.w5(32'hbb0c6438),
	.w6(32'h39a97bf8),
	.w7(32'hba2af073),
	.w8(32'h3b0c1552),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a048319),
	.w1(32'h3a036d21),
	.w2(32'h392e75a7),
	.w3(32'hbaeb7d61),
	.w4(32'h3ad3658e),
	.w5(32'hbba75b24),
	.w6(32'h3af38b2b),
	.w7(32'hb855163b),
	.w8(32'hb9dfc3e6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8831b),
	.w1(32'h3a91eccc),
	.w2(32'h3bb40672),
	.w3(32'hbbce67b5),
	.w4(32'h3b19a98d),
	.w5(32'h3c16d659),
	.w6(32'hbaba5b99),
	.w7(32'hbb89b304),
	.w8(32'hbb306f71),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb021ce3),
	.w1(32'hbbb33ef9),
	.w2(32'hbb5a194e),
	.w3(32'h3bc24a92),
	.w4(32'hbb62063b),
	.w5(32'h3ac50957),
	.w6(32'h3a9101b5),
	.w7(32'hbc16a3b1),
	.w8(32'hbbff7261),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae31f1f),
	.w1(32'hbb0bca75),
	.w2(32'hbafbf614),
	.w3(32'hbbd3b149),
	.w4(32'hbb83ca17),
	.w5(32'h3be3b659),
	.w6(32'hbb9cf99b),
	.w7(32'hbba89526),
	.w8(32'hbbf6face),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa84b),
	.w1(32'hbb440db4),
	.w2(32'hbaaa254e),
	.w3(32'hba8696b3),
	.w4(32'hbaf99af9),
	.w5(32'hbba17af2),
	.w6(32'hbaeb09dd),
	.w7(32'hbb413643),
	.w8(32'hbb07cd4e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b9bd),
	.w1(32'h3b13bcea),
	.w2(32'h3bd8e85d),
	.w3(32'hbc10d19f),
	.w4(32'hbabdae39),
	.w5(32'h3c5f1359),
	.w6(32'hbadc80f5),
	.w7(32'hbbabf962),
	.w8(32'hbb6ed357),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eddaf),
	.w1(32'h3ac563c7),
	.w2(32'h3b8d75d5),
	.w3(32'h3b9113a8),
	.w4(32'h3aa469c6),
	.w5(32'h3c50437e),
	.w6(32'hbb55b592),
	.w7(32'hbb3290dd),
	.w8(32'h3a1fec5c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba83d25),
	.w1(32'hb9c5535d),
	.w2(32'h3b32d4bc),
	.w3(32'h3b87af3d),
	.w4(32'hba247de3),
	.w5(32'hbc253181),
	.w6(32'h3b7f6c33),
	.w7(32'h3a8ab72a),
	.w8(32'h39e4812d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95ccf2),
	.w1(32'h3b1682ac),
	.w2(32'h3ba8b6ab),
	.w3(32'hbc3a7267),
	.w4(32'h3a84a23a),
	.w5(32'h3c5b7374),
	.w6(32'hbaa8bab8),
	.w7(32'hbadb0015),
	.w8(32'hbb1df37a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb787b5),
	.w1(32'hba298d15),
	.w2(32'h3ab52cd4),
	.w3(32'h3c1df718),
	.w4(32'h3af00f30),
	.w5(32'h3b12f414),
	.w6(32'h3b6b72e3),
	.w7(32'h3b12f563),
	.w8(32'h3bbfb8d5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f9541),
	.w1(32'hbba75162),
	.w2(32'h3b1fcae9),
	.w3(32'h3ae7203e),
	.w4(32'hbc0923da),
	.w5(32'h3b90da30),
	.w6(32'hbc2cfdc6),
	.w7(32'hbc57401d),
	.w8(32'hbc35287b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80fb96),
	.w1(32'h3ba3ca04),
	.w2(32'h3bce4399),
	.w3(32'h3afef01c),
	.w4(32'h3b9d95e2),
	.w5(32'hbad0a7f8),
	.w6(32'h3c0a7f6f),
	.w7(32'h3bb28a38),
	.w8(32'h3b5cb1d0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc12395),
	.w1(32'h3b618e00),
	.w2(32'hbb8c0a93),
	.w3(32'h3a6d62d0),
	.w4(32'h3c6272e1),
	.w5(32'h3cf1439f),
	.w6(32'h3b4ac714),
	.w7(32'h3b35e898),
	.w8(32'h3c20153a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d38dc),
	.w1(32'hbb5b1623),
	.w2(32'h3b39470b),
	.w3(32'h3d0163e4),
	.w4(32'h3c24425e),
	.w5(32'h3d02c844),
	.w6(32'hbcabe1fa),
	.w7(32'hbc7238fc),
	.w8(32'h3b64b22e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4373a),
	.w1(32'h3ae9584a),
	.w2(32'h3c15341c),
	.w3(32'h3d3f4223),
	.w4(32'h3bf1dc00),
	.w5(32'h3ca14893),
	.w6(32'hbca25172),
	.w7(32'hbc18d213),
	.w8(32'hbb63881e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27b716),
	.w1(32'hbad689ea),
	.w2(32'h39076d7d),
	.w3(32'h3cb327fb),
	.w4(32'h3a968a62),
	.w5(32'h3b78b32b),
	.w6(32'hbb2cf687),
	.w7(32'hbbe8b96e),
	.w8(32'h3b1b8763),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4155b),
	.w1(32'hbb857166),
	.w2(32'hbbbde13d),
	.w3(32'h3a812954),
	.w4(32'hbb237587),
	.w5(32'h3aa8428c),
	.w6(32'hb89f2303),
	.w7(32'hbb655afd),
	.w8(32'hb827f052),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c9f67),
	.w1(32'h3b500a65),
	.w2(32'h3bbba309),
	.w3(32'h3bffc690),
	.w4(32'h3b380264),
	.w5(32'hba9e77a0),
	.w6(32'h3b934731),
	.w7(32'h3b829b1d),
	.w8(32'h3b56cd97),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c8a30),
	.w1(32'hbac83d4c),
	.w2(32'h3baed259),
	.w3(32'hbb4043a7),
	.w4(32'h3b95dcf5),
	.w5(32'h3b009638),
	.w6(32'h3aba6ccc),
	.w7(32'h39c48cb7),
	.w8(32'h3b216e1e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86e657),
	.w1(32'hbc79833b),
	.w2(32'hbbe0f7ed),
	.w3(32'h3bac5eef),
	.w4(32'h3b81e85a),
	.w5(32'h3ce313d6),
	.w6(32'hbd0b0279),
	.w7(32'hbcd61d41),
	.w8(32'hbc24667c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd625dc),
	.w1(32'h3ba065c2),
	.w2(32'hbb820643),
	.w3(32'h3d148177),
	.w4(32'hbb5daedc),
	.w5(32'hbc143e1a),
	.w6(32'h3abbf1dc),
	.w7(32'h3a89f797),
	.w8(32'hbc02c237),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48d804),
	.w1(32'hbc92778b),
	.w2(32'hbc48787b),
	.w3(32'hbc54e9bb),
	.w4(32'hbc99bf4a),
	.w5(32'hbcb6276b),
	.w6(32'hbcb9d285),
	.w7(32'hbcbce381),
	.w8(32'hbcabf189),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9eb8d2),
	.w1(32'hbaec3c7f),
	.w2(32'h3ba2e44b),
	.w3(32'hbcdc04af),
	.w4(32'hbab47097),
	.w5(32'hba337f5f),
	.w6(32'h3af4ada9),
	.w7(32'h390c5d7b),
	.w8(32'hbaa1f108),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942200),
	.w1(32'h3be93f08),
	.w2(32'h3c1f71e0),
	.w3(32'hbbf37d45),
	.w4(32'h3b0c47de),
	.w5(32'h3bf591ba),
	.w6(32'h3c19c97c),
	.w7(32'h3c1eb512),
	.w8(32'h3b8d0222),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babff8a),
	.w1(32'hbbcb238f),
	.w2(32'hbbac4488),
	.w3(32'h3b0206d2),
	.w4(32'hbac98799),
	.w5(32'hbb098927),
	.w6(32'h3a71a84f),
	.w7(32'h392b371f),
	.w8(32'h3b0de4c6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33546f),
	.w1(32'hbc2ae65a),
	.w2(32'h3bbe3556),
	.w3(32'hb8ef0214),
	.w4(32'h3ab18d61),
	.w5(32'h3d007837),
	.w6(32'hbcc703c1),
	.w7(32'hbc5e0add),
	.w8(32'h3b97b25f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3548d),
	.w1(32'hbbdf7bf9),
	.w2(32'hb97310ae),
	.w3(32'h3d1937e5),
	.w4(32'h3c5089ca),
	.w5(32'h3c86e05a),
	.w6(32'hbb3d593f),
	.w7(32'hbb82e565),
	.w8(32'hbc435ea4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc900c0b),
	.w1(32'hbac07119),
	.w2(32'h3a58abd0),
	.w3(32'hbb5db088),
	.w4(32'hbb5428d2),
	.w5(32'h3c024cb0),
	.w6(32'hbb96c135),
	.w7(32'hbbb19738),
	.w8(32'hbb85fa8b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9c36a),
	.w1(32'h3b96d6bb),
	.w2(32'h3c3675b6),
	.w3(32'hbb40e0db),
	.w4(32'hb9afb7ff),
	.w5(32'hbb9c6ac9),
	.w6(32'h3bc79eb2),
	.w7(32'h3b7df58b),
	.w8(32'h3c148758),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51f421),
	.w1(32'h3ad05889),
	.w2(32'h3bed4f2b),
	.w3(32'hbbe08f46),
	.w4(32'h3abea937),
	.w5(32'h3c775301),
	.w6(32'hbae94401),
	.w7(32'hbb45ac8b),
	.w8(32'hbb8ae5b3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1820b),
	.w1(32'hbb280210),
	.w2(32'h3ba6b310),
	.w3(32'h3c127b2d),
	.w4(32'hbb2819a1),
	.w5(32'hb905f876),
	.w6(32'hb98f152d),
	.w7(32'hbaad732b),
	.w8(32'h3ba5ee83),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0486a),
	.w1(32'hbc536528),
	.w2(32'hbb4b63db),
	.w3(32'h3b665572),
	.w4(32'hbace5bb2),
	.w5(32'h3c8bbd7d),
	.w6(32'hbc1fd4ba),
	.w7(32'hbc5e6cb9),
	.w8(32'hbcb4fc88),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2a7bb),
	.w1(32'h3ad2580b),
	.w2(32'hbba06273),
	.w3(32'h3cac467e),
	.w4(32'h3be729b6),
	.w5(32'h3c8fd04d),
	.w6(32'h3a1caad6),
	.w7(32'hb9b7e48f),
	.w8(32'h3b4a57ec),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97fb6b),
	.w1(32'h39320945),
	.w2(32'h3aee43ca),
	.w3(32'h3c74d3d7),
	.w4(32'hbab20f80),
	.w5(32'h3c06501a),
	.w6(32'hbb421d4a),
	.w7(32'hbbc85610),
	.w8(32'hbba9f8e2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371b76),
	.w1(32'hbb25d0d2),
	.w2(32'h3c29fbb8),
	.w3(32'h3b4e895a),
	.w4(32'h3c4beab8),
	.w5(32'h3c53be22),
	.w6(32'hbb4293fd),
	.w7(32'h3aa39799),
	.w8(32'h3a7a49a2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf9e91),
	.w1(32'h3b929076),
	.w2(32'hba840fc8),
	.w3(32'hbb080785),
	.w4(32'h3b9a015e),
	.w5(32'hb9e41d88),
	.w6(32'h3bed375a),
	.w7(32'h3b6d5091),
	.w8(32'h3bd4f702),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3499bc),
	.w1(32'h3a19391b),
	.w2(32'hbbb74e9a),
	.w3(32'h3b450732),
	.w4(32'h3b45d96c),
	.w5(32'hbbb6a144),
	.w6(32'h3bc0e40b),
	.w7(32'hb9234022),
	.w8(32'hbb42f0cb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb340621),
	.w1(32'hbc18fa4c),
	.w2(32'hbbd459de),
	.w3(32'h3a097885),
	.w4(32'hbbd9369a),
	.w5(32'hbc3e699b),
	.w6(32'hbc1d0108),
	.w7(32'hbc2c44cc),
	.w8(32'hbc15c85d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb3677),
	.w1(32'hbb09b423),
	.w2(32'h3c1bcac0),
	.w3(32'hbc45f314),
	.w4(32'h3c9ac3a4),
	.w5(32'h3d14e82c),
	.w6(32'hbcbe9363),
	.w7(32'hbc491676),
	.w8(32'hbb72a244),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02d796),
	.w1(32'hba8adacc),
	.w2(32'h398c2514),
	.w3(32'h3d19e4e4),
	.w4(32'hbb08a837),
	.w5(32'h3c22876a),
	.w6(32'hbbd56d6f),
	.w7(32'hbbc27184),
	.w8(32'hbb16abe9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77b9be),
	.w1(32'hba5f5f14),
	.w2(32'h3ba0c88f),
	.w3(32'h3b4fc0a8),
	.w4(32'h3b9de312),
	.w5(32'hbb1b1a49),
	.w6(32'h3a3341a4),
	.w7(32'hbabae155),
	.w8(32'hbaaecece),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0437f),
	.w1(32'hb964a0f9),
	.w2(32'h3b007ee6),
	.w3(32'hbbfdfb7e),
	.w4(32'hba052798),
	.w5(32'hbc20d96e),
	.w6(32'h3b7138d3),
	.w7(32'h3a35342f),
	.w8(32'h39209e28),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba69119),
	.w1(32'hbb3f6685),
	.w2(32'hbb251bd0),
	.w3(32'hbc3dd98d),
	.w4(32'hb9827a5f),
	.w5(32'hbbdd8196),
	.w6(32'hba98f2b6),
	.w7(32'hbb3f4cc2),
	.w8(32'hbb48d1f1),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb075350),
	.w1(32'h3b8d4408),
	.w2(32'h3be9beed),
	.w3(32'hbbccc7e5),
	.w4(32'hba8ff9c1),
	.w5(32'h3c361916),
	.w6(32'hbba1197d),
	.w7(32'hbba7e983),
	.w8(32'hba81fe47),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c181d3a),
	.w1(32'hbbb09913),
	.w2(32'h3b894526),
	.w3(32'h3bd37eeb),
	.w4(32'hbad18f77),
	.w5(32'h3a0f92fd),
	.w6(32'hbc3534ac),
	.w7(32'hbc93a47f),
	.w8(32'hbc3159e1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20b187),
	.w1(32'hb8e2cefe),
	.w2(32'h3b46c62c),
	.w3(32'h3ab7362c),
	.w4(32'h3bdf4dc0),
	.w5(32'hbbc606bf),
	.w6(32'h3c334f15),
	.w7(32'h3be05ef5),
	.w8(32'h3be9c643),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc88f),
	.w1(32'hbc09c4b5),
	.w2(32'hba3d1b9f),
	.w3(32'hba89cf6f),
	.w4(32'hbb75b7a2),
	.w5(32'h3c8f2f5f),
	.w6(32'hbc6a1282),
	.w7(32'hbc396675),
	.w8(32'hbc3638ca),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17b38c),
	.w1(32'h3c0566d2),
	.w2(32'h3c0d544c),
	.w3(32'h3c719a32),
	.w4(32'h3b0deed8),
	.w5(32'hbbbdf378),
	.w6(32'h3c8435f7),
	.w7(32'h3c53842e),
	.w8(32'h3bb9d557),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebbd65),
	.w1(32'h3a469e92),
	.w2(32'hb9e57b08),
	.w3(32'hbc56797f),
	.w4(32'h3b3fa106),
	.w5(32'hbbbac2d7),
	.w6(32'h3b6525bb),
	.w7(32'hba9caaf9),
	.w8(32'h3b32c568),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989a246),
	.w1(32'h3a43d197),
	.w2(32'hbb5c62b6),
	.w3(32'hbb94c574),
	.w4(32'h3b684191),
	.w5(32'hbb1ef64a),
	.w6(32'hbac14f1a),
	.w7(32'hbbb9266e),
	.w8(32'hbafe6666),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18402b),
	.w1(32'hbc120c39),
	.w2(32'hbb0e66f6),
	.w3(32'h3ac0f562),
	.w4(32'hbbdef582),
	.w5(32'h3c373b15),
	.w6(32'hbc8af085),
	.w7(32'hbc819ad7),
	.w8(32'hbc2face3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71c8b3),
	.w1(32'h3a3e9afa),
	.w2(32'h3b8ea6d9),
	.w3(32'h3bf8a5ca),
	.w4(32'hbab0922d),
	.w5(32'h3afc9d37),
	.w6(32'hba113e50),
	.w7(32'hb98631e2),
	.w8(32'hba4fc9c4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c0eb7),
	.w1(32'hbaf53ad8),
	.w2(32'h3b87cd04),
	.w3(32'hbb3b5135),
	.w4(32'hba962827),
	.w5(32'h3c2fb76d),
	.w6(32'hbc05611f),
	.w7(32'hbbb39187),
	.w8(32'h3a42c36f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b0c9b),
	.w1(32'h3c0903e9),
	.w2(32'hbb46e1c1),
	.w3(32'h3bcd923c),
	.w4(32'h3b366520),
	.w5(32'hbb822d6b),
	.w6(32'h3c1d45a7),
	.w7(32'h38d80bdb),
	.w8(32'h3bd88399),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eb886),
	.w1(32'hbb739fbc),
	.w2(32'hbb23eff9),
	.w3(32'h3a6a6887),
	.w4(32'hbb2ccae6),
	.w5(32'h3a9c179e),
	.w6(32'hbab6aa8a),
	.w7(32'hbb6a4b40),
	.w8(32'h3aa91877),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a6189),
	.w1(32'hbc883413),
	.w2(32'h3b44066f),
	.w3(32'hbb4031a8),
	.w4(32'hbb9b888f),
	.w5(32'h3c9242b9),
	.w6(32'hbce07b45),
	.w7(32'hbc575d85),
	.w8(32'hba5142da),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91949d),
	.w1(32'hbb281507),
	.w2(32'hbac63e4c),
	.w3(32'h3d070927),
	.w4(32'hba790102),
	.w5(32'hbb83c121),
	.w6(32'h393c95cb),
	.w7(32'hba92bc2f),
	.w8(32'hb7a07cd5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e8dfa),
	.w1(32'h3c0a65d4),
	.w2(32'h3c44e372),
	.w3(32'hbb1a3b89),
	.w4(32'h3b86f446),
	.w5(32'h3c2676db),
	.w6(32'h3c20919c),
	.w7(32'h3c1ef48c),
	.w8(32'h3bcb33b5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b567fe3),
	.w1(32'hbc299b85),
	.w2(32'h3a419aaa),
	.w3(32'h3b29324f),
	.w4(32'hbb6fa142),
	.w5(32'hbaa6a52a),
	.w6(32'h3adafe33),
	.w7(32'hbbb2e978),
	.w8(32'h3b997b79),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23701b),
	.w1(32'h3954009a),
	.w2(32'h3ba014e5),
	.w3(32'hbbbcabe6),
	.w4(32'hba91a613),
	.w5(32'hbab8dd93),
	.w6(32'h39dbb094),
	.w7(32'h3b32472b),
	.w8(32'h3bb4a588),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7447e),
	.w1(32'hb9b17132),
	.w2(32'h3bc70c15),
	.w3(32'hbb1af267),
	.w4(32'h3c1f606c),
	.w5(32'h3ce43487),
	.w6(32'hbc46b055),
	.w7(32'hbbe6f377),
	.w8(32'h3bc260d0),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c586533),
	.w1(32'hbb68d247),
	.w2(32'hba1f941d),
	.w3(32'h3cceac81),
	.w4(32'hbbcd4c27),
	.w5(32'h39d35343),
	.w6(32'hbaad4160),
	.w7(32'hbb5bb649),
	.w8(32'hbbf8cda8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba35d9f),
	.w1(32'hbbda0cce),
	.w2(32'hbbbd52db),
	.w3(32'hba49d6c9),
	.w4(32'h3a059184),
	.w5(32'hbb48c197),
	.w6(32'hbb08d28c),
	.w7(32'hbb155d68),
	.w8(32'hbb2edf17),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb559873),
	.w1(32'hbb5aed38),
	.w2(32'h3b1d133c),
	.w3(32'h3ad1fa82),
	.w4(32'hbb1aaa26),
	.w5(32'h3b9fdbbe),
	.w6(32'hbb10c38a),
	.w7(32'hba88e578),
	.w8(32'h3a59a90b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2e45),
	.w1(32'hbb28a63f),
	.w2(32'h3b061211),
	.w3(32'h3b8c01d4),
	.w4(32'hbbbb1de1),
	.w5(32'hbc152742),
	.w6(32'hbc3526a0),
	.w7(32'hbc31a7e9),
	.w8(32'hbc88dc64),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc153fc9),
	.w1(32'h3ac42801),
	.w2(32'h3b0009ba),
	.w3(32'hbc79ad83),
	.w4(32'h3b462dcd),
	.w5(32'h3b023c28),
	.w6(32'h3b1f3868),
	.w7(32'h3b2016c0),
	.w8(32'h3b4878d8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f9e58),
	.w1(32'h3b56000d),
	.w2(32'h3b257a73),
	.w3(32'h3b294139),
	.w4(32'h3a3ea315),
	.w5(32'h3b67df8e),
	.w6(32'h3bc2ed5d),
	.w7(32'h3b713833),
	.w8(32'hbb4f342b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cd077),
	.w1(32'hb9d7f3ef),
	.w2(32'h3c307fcf),
	.w3(32'hbc5e88ce),
	.w4(32'h3b56b520),
	.w5(32'h3ce8abdb),
	.w6(32'hbc3cafb3),
	.w7(32'hbbd2d7fa),
	.w8(32'hbb8309c5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5246e3),
	.w1(32'hbbacd3cc),
	.w2(32'h3b84f04a),
	.w3(32'h3cbd24d5),
	.w4(32'hbc1ae973),
	.w5(32'hbb848594),
	.w6(32'hbb19e1d0),
	.w7(32'hbb0d6b2d),
	.w8(32'hbb8bb28c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78e02a),
	.w1(32'hbc1e800d),
	.w2(32'hbbd5a6e4),
	.w3(32'hbc5f3dac),
	.w4(32'h3ba3a56c),
	.w5(32'h3caebac2),
	.w6(32'hbb1845e2),
	.w7(32'hbcba278e),
	.w8(32'hbc4c58f5),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e6aec),
	.w1(32'h3c661b64),
	.w2(32'h3d05af2e),
	.w3(32'h3ca5e92f),
	.w4(32'h3c91fceb),
	.w5(32'h3b009e45),
	.w6(32'h3bf765fc),
	.w7(32'h3c032e24),
	.w8(32'h3b482706),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba22254),
	.w1(32'hbb38bc20),
	.w2(32'h3c1b3cce),
	.w3(32'hbd0d3f1a),
	.w4(32'h3c190f01),
	.w5(32'hbbb18d18),
	.w6(32'h3c489200),
	.w7(32'h3c0caaa2),
	.w8(32'h3c8744b0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2992eb),
	.w1(32'hbb9d150d),
	.w2(32'hba941213),
	.w3(32'hb9c39fbd),
	.w4(32'h39f2b47d),
	.w5(32'hbbd94db0),
	.w6(32'hbb175e11),
	.w7(32'hbbae13a2),
	.w8(32'hbb292db5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c8bee),
	.w1(32'hba92467e),
	.w2(32'h3a6787c6),
	.w3(32'hbc4a851c),
	.w4(32'h3b9760e0),
	.w5(32'hbbaa7379),
	.w6(32'h3be21319),
	.w7(32'h3b839c2c),
	.w8(32'h3b9cd1d1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73b103),
	.w1(32'hbb3973d5),
	.w2(32'h3a857d40),
	.w3(32'hbb647899),
	.w4(32'hbb8db0ce),
	.w5(32'hbb654b3b),
	.w6(32'hbac24e8e),
	.w7(32'hbb0b7a54),
	.w8(32'h3ae19299),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f71b),
	.w1(32'hbc5a4bd1),
	.w2(32'hbbb3a60b),
	.w3(32'hbb0b9b9b),
	.w4(32'hbbe7ad6a),
	.w5(32'h3b505b29),
	.w6(32'hbc619a5b),
	.w7(32'hbc24f879),
	.w8(32'hba6bfadc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0a334),
	.w1(32'hbba7b0cf),
	.w2(32'hbb4f27e3),
	.w3(32'h3ba8b389),
	.w4(32'hbb1e6eb1),
	.w5(32'hbbaf9e94),
	.w6(32'h3ae6b92f),
	.w7(32'h3aa04ad6),
	.w8(32'h3b0f9861),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6d485),
	.w1(32'hbab3c9f5),
	.w2(32'h3af3e68e),
	.w3(32'hbb2f7261),
	.w4(32'h3bc24522),
	.w5(32'hbb6b685c),
	.w6(32'h3bde3ce2),
	.w7(32'h3b959b4d),
	.w8(32'h3bb98bd5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac63282),
	.w1(32'hbc543132),
	.w2(32'hbc7405c3),
	.w3(32'h3931bdf2),
	.w4(32'hbb12c001),
	.w5(32'h3c9d6f24),
	.w6(32'hbcecd565),
	.w7(32'hbce70548),
	.w8(32'hbc0e930b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d53f4),
	.w1(32'hbbdab49e),
	.w2(32'hbc1db16f),
	.w3(32'h3d0af0fd),
	.w4(32'hbc365fef),
	.w5(32'hbca5b1a7),
	.w6(32'hbb76ba22),
	.w7(32'hbbe4d6ce),
	.w8(32'hbc1a6081),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f901a),
	.w1(32'hbb0e364f),
	.w2(32'hbb90cb10),
	.w3(32'hbc804a42),
	.w4(32'hbba30113),
	.w5(32'hba9ec436),
	.w6(32'h370a5f30),
	.w7(32'hbb4b1ce5),
	.w8(32'hbadad10b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc47ffa),
	.w1(32'hbbccaf04),
	.w2(32'hbb6b5aa8),
	.w3(32'h3c91b96d),
	.w4(32'hbc1f34af),
	.w5(32'hbc87ad13),
	.w6(32'hbbeb1f70),
	.w7(32'hbbd127dc),
	.w8(32'hbbb742dd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a0c41),
	.w1(32'hbbd023b2),
	.w2(32'h396d194f),
	.w3(32'hbc9c2298),
	.w4(32'hbc307d77),
	.w5(32'h3b636187),
	.w6(32'hbc7dd371),
	.w7(32'hbc6935b1),
	.w8(32'hbba29234),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e1ddc),
	.w1(32'hbc1b2ccb),
	.w2(32'h3c5084d5),
	.w3(32'h3a1cd7c7),
	.w4(32'hba8cc89b),
	.w5(32'h3ca01472),
	.w6(32'hbc2dc130),
	.w7(32'hbba8d05e),
	.w8(32'h3bb80073),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc12a9d),
	.w1(32'hbab071f4),
	.w2(32'h3b11c94f),
	.w3(32'h3cfdb4bd),
	.w4(32'h3c03029a),
	.w5(32'hbbc51476),
	.w6(32'h3c284d9f),
	.w7(32'h3be0c75c),
	.w8(32'h3c061ba3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb319933),
	.w1(32'hba7bdf8a),
	.w2(32'h3abe5705),
	.w3(32'hba143a3f),
	.w4(32'h3b53b2e8),
	.w5(32'hbbc47c79),
	.w6(32'h3b1e6fdd),
	.w7(32'hbad501a0),
	.w8(32'hba8412ce),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850bae),
	.w1(32'hbb66b24e),
	.w2(32'hbaf01a0d),
	.w3(32'hbc122c0a),
	.w4(32'hb9aa3f39),
	.w5(32'hbc3f9039),
	.w6(32'h3b3fc19a),
	.w7(32'hbae86d24),
	.w8(32'hbb0a16c2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948aaf),
	.w1(32'h3c1a8033),
	.w2(32'h3c70332e),
	.w3(32'hbc3f1d43),
	.w4(32'h3aca82e8),
	.w5(32'h3b94c586),
	.w6(32'h3c773cd0),
	.w7(32'h3c32f3b0),
	.w8(32'h3c9e94b9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e238d),
	.w1(32'h3aae7339),
	.w2(32'h3bc6651d),
	.w3(32'h3c4ba2b1),
	.w4(32'h3c1db25f),
	.w5(32'h3cb95db0),
	.w6(32'hbbcd1909),
	.w7(32'hbc0793d7),
	.w8(32'hbba1a62f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4b097),
	.w1(32'hbc45c4c9),
	.w2(32'hbbeb6e5e),
	.w3(32'h3b928870),
	.w4(32'hbc0930e7),
	.w5(32'hbc1bb4fd),
	.w6(32'hbc64b8d2),
	.w7(32'hbc61aa4e),
	.w8(32'hbc363367),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07438d),
	.w1(32'hbc20f708),
	.w2(32'hbbeb9d40),
	.w3(32'hbc3bcd78),
	.w4(32'hbc157360),
	.w5(32'hbc3754da),
	.w6(32'hbc667ba6),
	.w7(32'hbc5a34f7),
	.w8(32'hbc2ffcb5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ef5e5),
	.w1(32'h3a44c64e),
	.w2(32'h3ba57a3c),
	.w3(32'hbc26c6bc),
	.w4(32'h3b2ae351),
	.w5(32'hbbbd9105),
	.w6(32'h3bc43b99),
	.w7(32'h3ac5d43a),
	.w8(32'h3b1fce65),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6ec3a),
	.w1(32'h3c70d454),
	.w2(32'h3cad2fbf),
	.w3(32'hbc03b3bb),
	.w4(32'h3b1b130d),
	.w5(32'hb9a82bfa),
	.w6(32'h3bfffec2),
	.w7(32'h3b8fadc8),
	.w8(32'h3b506f4e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40cb32),
	.w1(32'hbcb38562),
	.w2(32'hbc91c2d4),
	.w3(32'hbb044a96),
	.w4(32'hbcc01f58),
	.w5(32'hbcdfa2ad),
	.w6(32'hbcb4b5fa),
	.w7(32'hbce34cdf),
	.w8(32'hbcf9bd07),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba165e),
	.w1(32'h3af81941),
	.w2(32'h3bd24b44),
	.w3(32'hbd12844f),
	.w4(32'hbac5eba5),
	.w5(32'hbb91a5be),
	.w6(32'h3b63c5aa),
	.w7(32'h3b07b0db),
	.w8(32'h3b9c3e0e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977f8e),
	.w1(32'h3a2550b4),
	.w2(32'hba06127f),
	.w3(32'hbbe54531),
	.w4(32'h3ac43524),
	.w5(32'h3a8c0345),
	.w6(32'h3aaffdc3),
	.w7(32'h3a1a1dc0),
	.w8(32'h3ab5d966),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0aea3e),
	.w1(32'hbbdfefd9),
	.w2(32'hbba7bddd),
	.w3(32'h3aa78d3d),
	.w4(32'hbba3e025),
	.w5(32'hbba3d587),
	.w6(32'hbb38abaf),
	.w7(32'hbb424c05),
	.w8(32'hbb48733e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule