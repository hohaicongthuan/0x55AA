module layer_6_featuremap_100(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8e2a0),
	.w1(32'h39fdc59f),
	.w2(32'h3b64f1d2),
	.w3(32'h3b5e04fa),
	.w4(32'h3b0d3ead),
	.w5(32'h3b2a8306),
	.w6(32'hb9bf7fc2),
	.w7(32'hba3e798a),
	.w8(32'h3b67b794),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b927da7),
	.w1(32'h38e7557e),
	.w2(32'hba93f19e),
	.w3(32'hbc2a7b7c),
	.w4(32'hbbd51b91),
	.w5(32'hbb4c848f),
	.w6(32'h3bab55f4),
	.w7(32'h3c3296a8),
	.w8(32'h3bb2ec21),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa70131),
	.w1(32'hbb434173),
	.w2(32'h3c7cec51),
	.w3(32'hbbe1b20f),
	.w4(32'hbbbd82c4),
	.w5(32'h3bbcffe4),
	.w6(32'hbc36a59e),
	.w7(32'h3c4ce533),
	.w8(32'h3cca8ce3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97449e),
	.w1(32'h3b0ee480),
	.w2(32'h3b1698d0),
	.w3(32'hb8790960),
	.w4(32'h3b1c8c7d),
	.w5(32'h3b731997),
	.w6(32'h3b38ae48),
	.w7(32'h3b6a75d6),
	.w8(32'h3b29ef15),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c2b9f),
	.w1(32'hbc939ae9),
	.w2(32'hba15f498),
	.w3(32'hbbba59aa),
	.w4(32'hbc39a0da),
	.w5(32'hbcc150b8),
	.w6(32'hbcc925f6),
	.w7(32'hbce58c80),
	.w8(32'hbc3c2596),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f5ee8),
	.w1(32'hbbb899f2),
	.w2(32'h3b68d17e),
	.w3(32'hba324fe5),
	.w4(32'hbc0ac16e),
	.w5(32'hbc2d65b2),
	.w6(32'hbc0caff7),
	.w7(32'hbc38bde0),
	.w8(32'hbae72bd0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c3369),
	.w1(32'hbbe25c3a),
	.w2(32'hbc86967a),
	.w3(32'hbc064c63),
	.w4(32'h3b5b0985),
	.w5(32'hba7beeb2),
	.w6(32'h3b4f62b9),
	.w7(32'h3beb62bb),
	.w8(32'hbc317b6f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc88fa3),
	.w1(32'h3bd404e6),
	.w2(32'h3c9db635),
	.w3(32'h3cb6bee4),
	.w4(32'h3d08d160),
	.w5(32'h3c40fe47),
	.w6(32'h3c165740),
	.w7(32'h3d1257be),
	.w8(32'h3cdf38d7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1572a),
	.w1(32'h3c9527ab),
	.w2(32'h3cc40920),
	.w3(32'hbc9c76a2),
	.w4(32'hbb0e1afe),
	.w5(32'h3b8be994),
	.w6(32'h3c3fa967),
	.w7(32'h3d08df64),
	.w8(32'h3ce7cd2b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fd825),
	.w1(32'hba771cb7),
	.w2(32'h3c6a41cc),
	.w3(32'hbb953533),
	.w4(32'hbc2b9540),
	.w5(32'hbbf0b7f7),
	.w6(32'hbc014a04),
	.w7(32'hba8b4b84),
	.w8(32'h3c1a4813),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1c0ba),
	.w1(32'hbc92658e),
	.w2(32'hbc97c231),
	.w3(32'h3c07352e),
	.w4(32'hbc19d311),
	.w5(32'hbc1b4669),
	.w6(32'hbc674c03),
	.w7(32'hbc8c2753),
	.w8(32'hbc9ed380),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e8d5a),
	.w1(32'hba6c3926),
	.w2(32'h3c85f640),
	.w3(32'hbb7e2680),
	.w4(32'hbc197fa3),
	.w5(32'hbb518f6e),
	.w6(32'hbb964b54),
	.w7(32'hbadb350e),
	.w8(32'h3c24b664),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfd7257),
	.w1(32'hbb8fed17),
	.w2(32'h3bd771bc),
	.w3(32'hba08c6a1),
	.w4(32'h3bb6acf0),
	.w5(32'hbb9a6991),
	.w6(32'h3b4e8047),
	.w7(32'h3c906a29),
	.w8(32'h3aca8945),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0282),
	.w1(32'hbb2b2e51),
	.w2(32'hbc3c258b),
	.w3(32'hbc8645e8),
	.w4(32'hbc9312d7),
	.w5(32'hbb9f7af1),
	.w6(32'hbba6d31a),
	.w7(32'hbc1a5d38),
	.w8(32'hbb8d78a2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b0254),
	.w1(32'hbb7733ab),
	.w2(32'hbb748b9f),
	.w3(32'hbb317139),
	.w4(32'hbb5c25a1),
	.w5(32'hbba21b52),
	.w6(32'hbb2fa526),
	.w7(32'hbbed92f9),
	.w8(32'hbb988baf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b27d1),
	.w1(32'h3b88ea7b),
	.w2(32'h3aa0ee0a),
	.w3(32'h3bbb279e),
	.w4(32'h3bad52ce),
	.w5(32'h3b2a877a),
	.w6(32'h3c37c6e7),
	.w7(32'h3bf3cee5),
	.w8(32'h3b49cf67),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f318a),
	.w1(32'hbb2a80bc),
	.w2(32'h3b00e3ea),
	.w3(32'h3a888c25),
	.w4(32'h3bb01f8d),
	.w5(32'h3cad73a6),
	.w6(32'h3bb13eb5),
	.w7(32'h3bd58b2f),
	.w8(32'h3bda88b5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf0d70),
	.w1(32'h399356a7),
	.w2(32'h3c083809),
	.w3(32'h3a197432),
	.w4(32'hba8c4775),
	.w5(32'h3b3401f9),
	.w6(32'hbb223cb0),
	.w7(32'h3b293eb0),
	.w8(32'h3c2f99d3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c813e27),
	.w1(32'h3925de07),
	.w2(32'hb9c0e4cd),
	.w3(32'hba83f530),
	.w4(32'hbb176f18),
	.w5(32'hbb2c1064),
	.w6(32'hba131d33),
	.w7(32'hbb4d8f97),
	.w8(32'hbb1dbb98),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39f37c),
	.w1(32'h3b48f12c),
	.w2(32'hbbf697bb),
	.w3(32'h3b999deb),
	.w4(32'h3c861670),
	.w5(32'hbc21662c),
	.w6(32'h3c2d924b),
	.w7(32'hbb05035c),
	.w8(32'hbc5a43f7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc142c16),
	.w1(32'h394fe6af),
	.w2(32'hb94e414e),
	.w3(32'h3ad9b6ae),
	.w4(32'h3b93dc7e),
	.w5(32'h3b0d2adb),
	.w6(32'h3b2ff598),
	.w7(32'h3b87b256),
	.w8(32'hb857c05f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977488),
	.w1(32'h3c0d7759),
	.w2(32'h3c694a05),
	.w3(32'h3c560484),
	.w4(32'h3c51e92e),
	.w5(32'h3bec43e4),
	.w6(32'h3c48f45c),
	.w7(32'h3ca1eca0),
	.w8(32'h3c0e5156),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad1739),
	.w1(32'hbac53701),
	.w2(32'h3d22b09d),
	.w3(32'hbd54caee),
	.w4(32'hbd2ce2a7),
	.w5(32'hbcd53f33),
	.w6(32'hbd10862c),
	.w7(32'h3c130d07),
	.w8(32'h3cc6e540),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cea4b84),
	.w1(32'h3c812990),
	.w2(32'h3cd32e55),
	.w3(32'hbc937f1f),
	.w4(32'hb7f037d0),
	.w5(32'h3c9ed430),
	.w6(32'h3bc08eb4),
	.w7(32'h3d3b146f),
	.w8(32'h3c96fdaf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8922fdc),
	.w1(32'hbc9ecaf3),
	.w2(32'hbc1eb68b),
	.w3(32'h3944de2c),
	.w4(32'h3baebd93),
	.w5(32'h3a3150e7),
	.w6(32'hbc845dff),
	.w7(32'h3afd16dd),
	.w8(32'hbbf02d1a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75eda),
	.w1(32'hbb03747f),
	.w2(32'h3af65ea5),
	.w3(32'h3b87aa04),
	.w4(32'hbb192671),
	.w5(32'hbb2948f4),
	.w6(32'h3b085648),
	.w7(32'h3b4b6bc4),
	.w8(32'hbaf03253),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae03da6),
	.w1(32'hba13bd11),
	.w2(32'hbbaed0cc),
	.w3(32'h3b28335e),
	.w4(32'hbb3f36f4),
	.w5(32'hbad92576),
	.w6(32'hbb470e9f),
	.w7(32'hbb8765d2),
	.w8(32'hbb5e0a80),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819963),
	.w1(32'hbaf5ab3c),
	.w2(32'hbc26b6f9),
	.w3(32'hba586ee4),
	.w4(32'h3bfa4e81),
	.w5(32'h3b5cf5e2),
	.w6(32'h3bd14884),
	.w7(32'h3b9215c7),
	.w8(32'hbbed9550),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc659b71),
	.w1(32'h3b2cac6e),
	.w2(32'hbb443e57),
	.w3(32'hbb7e76aa),
	.w4(32'hba0887ad),
	.w5(32'h3acc3560),
	.w6(32'h3a67080f),
	.w7(32'hbac20092),
	.w8(32'hbb3a3c80),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc167fe),
	.w1(32'hb995762b),
	.w2(32'hbba3a636),
	.w3(32'hbc080b9d),
	.w4(32'hbc11368b),
	.w5(32'h3ad593ae),
	.w6(32'hbba049f5),
	.w7(32'hb907dbb5),
	.w8(32'hb8fb744f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c2b1e),
	.w1(32'h3c907325),
	.w2(32'hbc90b7f0),
	.w3(32'h3d2ee6f8),
	.w4(32'h3d85c4fc),
	.w5(32'h3c7f8296),
	.w6(32'h3d999789),
	.w7(32'h3d64a849),
	.w8(32'h3a2b1498),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3cb5cf),
	.w1(32'hbce44656),
	.w2(32'hbc885f41),
	.w3(32'h3ca15bac),
	.w4(32'h394a0e6c),
	.w5(32'hbccc0529),
	.w6(32'hbc0cf45b),
	.w7(32'hbd1b0eb1),
	.w8(32'hbd20f483),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b5f15),
	.w1(32'hbb7bb6ea),
	.w2(32'hbc0118b7),
	.w3(32'h3b773f57),
	.w4(32'h3c10dcd7),
	.w5(32'h3c3e48fe),
	.w6(32'h3c660ffa),
	.w7(32'h3ce1c122),
	.w8(32'hbb438962),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1f49d),
	.w1(32'h3aae1e2f),
	.w2(32'hb99659c3),
	.w3(32'hbc09745e),
	.w4(32'h3c38ff07),
	.w5(32'h3c225913),
	.w6(32'h3b593251),
	.w7(32'h3ca19cf3),
	.w8(32'h3c32792b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1032f9),
	.w1(32'h3aa96b52),
	.w2(32'h3c1427c4),
	.w3(32'h3a985a27),
	.w4(32'hbb8bc496),
	.w5(32'hba806bdc),
	.w6(32'hbbb8a43c),
	.w7(32'hbb90b729),
	.w8(32'h3bddd15d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bfd5e),
	.w1(32'hbbfe1db3),
	.w2(32'hba32107b),
	.w3(32'hbb730ab2),
	.w4(32'hbc0fa8ce),
	.w5(32'hbaa7dc67),
	.w6(32'hbb2a8608),
	.w7(32'hbc305af6),
	.w8(32'h3b9148b8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0779a8),
	.w1(32'hbb9603fd),
	.w2(32'hbb21bb0f),
	.w3(32'h3c19c065),
	.w4(32'h3bd691bb),
	.w5(32'h3b390900),
	.w6(32'hb8500ba4),
	.w7(32'hbbae5403),
	.w8(32'hba45cb7f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9812f8b),
	.w1(32'h3bdda796),
	.w2(32'h3af51031),
	.w3(32'h3b9cb7c1),
	.w4(32'h3b889592),
	.w5(32'h3b96a8c7),
	.w6(32'h3bfd9401),
	.w7(32'h3b950274),
	.w8(32'h3b80cdfa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5a1b0),
	.w1(32'hbc75ff49),
	.w2(32'hbc3870b6),
	.w3(32'h3bdcefa1),
	.w4(32'h3b4b903d),
	.w5(32'hbbbf4335),
	.w6(32'hba8ec144),
	.w7(32'hbb3f9255),
	.w8(32'hbc73b029),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b1d70),
	.w1(32'hbc3f1536),
	.w2(32'hbcb9e833),
	.w3(32'h3ce8ee17),
	.w4(32'h3c1c0b58),
	.w5(32'h3bc89587),
	.w6(32'h3ba9fb06),
	.w7(32'hbb80d952),
	.w8(32'hbcde5c8b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9aefc9),
	.w1(32'h3c248c06),
	.w2(32'h3b8c9db1),
	.w3(32'h3ca9073e),
	.w4(32'h3d0119e8),
	.w5(32'h3cb5977c),
	.w6(32'h3d161553),
	.w7(32'h3d14da52),
	.w8(32'h3cf8f838),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc025a9e),
	.w1(32'h3bb5621d),
	.w2(32'h3b77ae97),
	.w3(32'h3b98f691),
	.w4(32'h3be31f76),
	.w5(32'h3bcffec6),
	.w6(32'h3bcabddd),
	.w7(32'h3bd340e1),
	.w8(32'h3b6df31b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba872b51),
	.w1(32'h3c22ede4),
	.w2(32'h3c76ffd6),
	.w3(32'h3c12f379),
	.w4(32'h3ba0a5cd),
	.w5(32'h3b925839),
	.w6(32'h3c0231cb),
	.w7(32'h3be12d00),
	.w8(32'h3be8ba59),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9af405),
	.w1(32'h3a299547),
	.w2(32'hbbd9cd6e),
	.w3(32'h3c505797),
	.w4(32'h3cd772df),
	.w5(32'h3c2d7b07),
	.w6(32'h3ccd941f),
	.w7(32'h3c83cfdf),
	.w8(32'hbaf21104),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eedce),
	.w1(32'h3ac87bd7),
	.w2(32'h3b99dc80),
	.w3(32'hbc0e19f9),
	.w4(32'hbbffb4af),
	.w5(32'hbb6ce27c),
	.w6(32'hbb263a80),
	.w7(32'h3b5243ae),
	.w8(32'h3b9fa2cd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1299e),
	.w1(32'hbd1efb88),
	.w2(32'hbcc9d20e),
	.w3(32'hbc146c86),
	.w4(32'hbcbe51a4),
	.w5(32'hbcc1c185),
	.w6(32'hbca2009e),
	.w7(32'hbc896b06),
	.w8(32'hbcfe6d46),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb99a48),
	.w1(32'h3c65e9cd),
	.w2(32'h3bcc25f6),
	.w3(32'hbbcf1365),
	.w4(32'hbad9adbd),
	.w5(32'h3cbe191e),
	.w6(32'hbb01f025),
	.w7(32'h3c889860),
	.w8(32'h3ca982a4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f1e5a),
	.w1(32'hbc9ec5ce),
	.w2(32'hbca1f310),
	.w3(32'hbc78e2c2),
	.w4(32'hbb7d76a6),
	.w5(32'hbb933de2),
	.w6(32'hbcb0e0be),
	.w7(32'hbbd79339),
	.w8(32'hbb2ed68b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92b011),
	.w1(32'h399fe500),
	.w2(32'hb99fc4c3),
	.w3(32'hbaa24916),
	.w4(32'hbb9605f3),
	.w5(32'hbb67b9ad),
	.w6(32'hbb065b49),
	.w7(32'hbb374922),
	.w8(32'hba62fa85),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21374d),
	.w1(32'hbcc01289),
	.w2(32'hbd2c8822),
	.w3(32'h3c8c20b4),
	.w4(32'h3c17bb60),
	.w5(32'hbc168cb1),
	.w6(32'hb962e227),
	.w7(32'hbcb7aa16),
	.w8(32'hbcdde093),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc882f6),
	.w1(32'h3b62b27b),
	.w2(32'h3c09fdad),
	.w3(32'hba05b019),
	.w4(32'h3b9daf9a),
	.w5(32'h3b4ab113),
	.w6(32'h3b4e108d),
	.w7(32'h3c632935),
	.w8(32'h3c05ef17),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c0a39),
	.w1(32'h398e2a26),
	.w2(32'h3aac8067),
	.w3(32'hbb818a63),
	.w4(32'h3b1accb0),
	.w5(32'h3b48f2e9),
	.w6(32'h3aeb528f),
	.w7(32'h3c15e375),
	.w8(32'h3c0dea87),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0d4ac),
	.w1(32'h3bca96cd),
	.w2(32'hba3987d5),
	.w3(32'hbbb590e9),
	.w4(32'h3b96a4b3),
	.w5(32'h3c624c06),
	.w6(32'h3bfe9450),
	.w7(32'h3c4a38e9),
	.w8(32'h3c041f34),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28a50d),
	.w1(32'h3acd614e),
	.w2(32'hbbb11ce0),
	.w3(32'hbc9ee154),
	.w4(32'h391d6668),
	.w5(32'h3c370e53),
	.w6(32'h3b3c8a15),
	.w7(32'h3c65f38b),
	.w8(32'h3c2211e5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d8b96),
	.w1(32'hbb029d74),
	.w2(32'h3b5631c4),
	.w3(32'hbc34511c),
	.w4(32'hbb3aeac7),
	.w5(32'hbb0f0469),
	.w6(32'h3b33cf90),
	.w7(32'h3c88d29c),
	.w8(32'h3c6565a5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4c4b6),
	.w1(32'h3a37a2cd),
	.w2(32'h3a51f343),
	.w3(32'h3c167868),
	.w4(32'hbbdde8de),
	.w5(32'hbc09cf9f),
	.w6(32'h3b84cd6f),
	.w7(32'hbb017647),
	.w8(32'hba8240de),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5c127),
	.w1(32'hbc53d8df),
	.w2(32'hbccc9cf4),
	.w3(32'hbc28f93a),
	.w4(32'hbca232c4),
	.w5(32'hbc893b3e),
	.w6(32'hbc8db711),
	.w7(32'hbd0213d1),
	.w8(32'hbcdea685),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca29403),
	.w1(32'h3bb54c9b),
	.w2(32'hba04522a),
	.w3(32'h3a587288),
	.w4(32'h3b495b04),
	.w5(32'hb9c41927),
	.w6(32'h3b86079d),
	.w7(32'h3a14a33d),
	.w8(32'hbb0237e2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970d8eb),
	.w1(32'h3ab19a46),
	.w2(32'h3c0fa45b),
	.w3(32'hbaa0e120),
	.w4(32'h3b7083fb),
	.w5(32'h3bc5158e),
	.w6(32'h3b1872d0),
	.w7(32'h3c130f7d),
	.w8(32'h3c2cdc58),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c222a58),
	.w1(32'hbba5d758),
	.w2(32'h3a0b2d49),
	.w3(32'h3bfb6eb7),
	.w4(32'hbc020d92),
	.w5(32'h3badfdfc),
	.w6(32'hbb986860),
	.w7(32'hbc1d9347),
	.w8(32'h3bd15b3b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6cb210),
	.w1(32'h3b42263f),
	.w2(32'h3bcee7ee),
	.w3(32'hbb39c102),
	.w4(32'hbadda99b),
	.w5(32'h3bba5893),
	.w6(32'h3a927b0c),
	.w7(32'h3bcda9ed),
	.w8(32'h3c8106a4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53616d),
	.w1(32'hbb51c5a3),
	.w2(32'hb919408e),
	.w3(32'hbb7e85a7),
	.w4(32'h3a367b60),
	.w5(32'h39e49ae6),
	.w6(32'h3ab21637),
	.w7(32'h3b9b9b6a),
	.w8(32'h39846d42),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf3fc2),
	.w1(32'hbc420475),
	.w2(32'hbbd68c05),
	.w3(32'h3c16388e),
	.w4(32'h3b25cc99),
	.w5(32'h3c357324),
	.w6(32'hbb8fd0ef),
	.w7(32'hbb9270e2),
	.w8(32'h3a055684),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba30da0),
	.w1(32'hbc9286ee),
	.w2(32'h3d2c383a),
	.w3(32'hbc2b4c50),
	.w4(32'h3d2c0453),
	.w5(32'h3d7ef120),
	.w6(32'hbbaa27b7),
	.w7(32'h3d7f5d8d),
	.w8(32'h3db5f354),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule