module layer_10_featuremap_283(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31dbfa),
	.w1(32'hba87467f),
	.w2(32'hba813df5),
	.w3(32'hb9bbc6c5),
	.w4(32'hb98fd516),
	.w5(32'h37f1797b),
	.w6(32'hbaa984a0),
	.w7(32'hbab99899),
	.w8(32'hb7e39cf0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa23492),
	.w1(32'hba6e0edc),
	.w2(32'hb83ea899),
	.w3(32'hba71f992),
	.w4(32'h3a676e01),
	.w5(32'hb744fc76),
	.w6(32'hba77aa86),
	.w7(32'h3ac050ca),
	.w8(32'h39e5c014),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a6e94),
	.w1(32'hb9c2a709),
	.w2(32'h39c12eff),
	.w3(32'hba62d114),
	.w4(32'hb90bfbcd),
	.w5(32'h39ebf9d4),
	.w6(32'hb764248c),
	.w7(32'h3a26da2f),
	.w8(32'h3a1a56cc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979c116),
	.w1(32'hba32a99f),
	.w2(32'hb9a0b873),
	.w3(32'h3a59e828),
	.w4(32'h3a0d3241),
	.w5(32'hba883bde),
	.w6(32'h3a21c926),
	.w7(32'h39bf2aa3),
	.w8(32'hba33e3a6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18d7ea),
	.w1(32'hba4ce6ff),
	.w2(32'hb9b78e55),
	.w3(32'hb99b9843),
	.w4(32'hb91b06d9),
	.w5(32'h39c51c08),
	.w6(32'h370e606a),
	.w7(32'hb957f19f),
	.w8(32'hb96b87d7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39538e64),
	.w1(32'hb73e9b97),
	.w2(32'hb8ce89c2),
	.w3(32'h3958a30b),
	.w4(32'h3970c79a),
	.w5(32'h3aded9b7),
	.w6(32'hba019882),
	.w7(32'hb9dc3355),
	.w8(32'h3ae50e42),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3ee68),
	.w1(32'h3abf46a4),
	.w2(32'hb90230e1),
	.w3(32'hbb2696d5),
	.w4(32'hbb4a68c2),
	.w5(32'h3a3c7c99),
	.w6(32'hba67034b),
	.w7(32'hbb615ba0),
	.w8(32'hba2a252e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa209c4),
	.w1(32'h3b4646cc),
	.w2(32'h3bb73ed3),
	.w3(32'h3b4c7923),
	.w4(32'h3a4c0806),
	.w5(32'h3bb43584),
	.w6(32'h3bf82ad3),
	.w7(32'hba3049df),
	.w8(32'h39cad139),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d45a1),
	.w1(32'hb9037bd1),
	.w2(32'h389e2dcc),
	.w3(32'h38faedbb),
	.w4(32'hb9807c49),
	.w5(32'hba27321d),
	.w6(32'hbaa8a47d),
	.w7(32'hbaa38136),
	.w8(32'hba7a4882),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd4a74),
	.w1(32'h3b49fa1e),
	.w2(32'h39a9d5cb),
	.w3(32'h3b33de2e),
	.w4(32'h3ae34da6),
	.w5(32'h3a85471e),
	.w6(32'h38bc66a9),
	.w7(32'hbaf9a874),
	.w8(32'h3a6da5ab),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2d8fe),
	.w1(32'h3ab5b6ac),
	.w2(32'h3ac52d10),
	.w3(32'h3a1db2c7),
	.w4(32'h3a95ca51),
	.w5(32'h3a6dad08),
	.w6(32'h381afa93),
	.w7(32'h3a302df3),
	.w8(32'h39094f5b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9229ce0),
	.w1(32'hbb9083b5),
	.w2(32'hbb960b8d),
	.w3(32'hbb906e3e),
	.w4(32'hbc1acf7d),
	.w5(32'hbbc1d399),
	.w6(32'hbaada866),
	.w7(32'hbbd93557),
	.w8(32'hbbb2c5a2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08af17),
	.w1(32'h3b812869),
	.w2(32'hb9bab1ed),
	.w3(32'h3bc6babd),
	.w4(32'h3b32e780),
	.w5(32'h3998e4f1),
	.w6(32'h3b8dd37c),
	.w7(32'h39b544b5),
	.w8(32'h3ae2a84f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6b5db),
	.w1(32'h390ac8e4),
	.w2(32'h3b40140e),
	.w3(32'hbb06a87d),
	.w4(32'hba328958),
	.w5(32'h3afccaea),
	.w6(32'h36bdbc5a),
	.w7(32'hbac1b404),
	.w8(32'h3aaf6508),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13dca4),
	.w1(32'h3b13dfd1),
	.w2(32'h3a0f4912),
	.w3(32'h3a047541),
	.w4(32'hb86adff6),
	.w5(32'hba3efdba),
	.w6(32'hb9e1ffe5),
	.w7(32'hba59cafd),
	.w8(32'hbad624c8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf297b),
	.w1(32'h3ac01f04),
	.w2(32'hbb8aa055),
	.w3(32'h3a161c2f),
	.w4(32'h3b4732e5),
	.w5(32'h3a84e174),
	.w6(32'hbb43d2ab),
	.w7(32'hb9baee92),
	.w8(32'h3b4a85a1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a634f),
	.w1(32'h3a696b1d),
	.w2(32'h3a92a60b),
	.w3(32'h3a3610ad),
	.w4(32'h3a90f93b),
	.w5(32'hb9b6fd15),
	.w6(32'h39da9f00),
	.w7(32'h3a60af7b),
	.w8(32'hba3114cd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82afcc),
	.w1(32'h3bb60fb2),
	.w2(32'h3b2c4ed3),
	.w3(32'hba8a5004),
	.w4(32'hba5f5957),
	.w5(32'h3b597c0b),
	.w6(32'h3b3b69cd),
	.w7(32'hba4129fe),
	.w8(32'h3b161f36),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b828659),
	.w1(32'h3b45cf58),
	.w2(32'h3a9bc1e9),
	.w3(32'h3b1fe08e),
	.w4(32'h3b0634cf),
	.w5(32'h3af0560d),
	.w6(32'h3b46687a),
	.w7(32'h3aaf45c2),
	.w8(32'h3a4a86f6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa529e6),
	.w1(32'hba5d1d9a),
	.w2(32'hba22f946),
	.w3(32'h3932b0cc),
	.w4(32'hb98c160d),
	.w5(32'hb941d125),
	.w6(32'hb9940914),
	.w7(32'hba24ac5b),
	.w8(32'hba0c209b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f493d2),
	.w1(32'h3aca0097),
	.w2(32'h3a122c27),
	.w3(32'h3a9f1a9b),
	.w4(32'hb9813dbe),
	.w5(32'h3ac52e16),
	.w6(32'h3aaf5dd5),
	.w7(32'hba0d2820),
	.w8(32'h3aa7c8f4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8891fb),
	.w1(32'hba4a1f47),
	.w2(32'hb9a9c0f1),
	.w3(32'hb9ba465e),
	.w4(32'h3a364cd8),
	.w5(32'h39225a9c),
	.w6(32'hb902bd16),
	.w7(32'h3abbb3f3),
	.w8(32'h3a163f55),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f196a),
	.w1(32'h3b35eb4b),
	.w2(32'hbb6fdda6),
	.w3(32'h3ba8c4d2),
	.w4(32'hbb9429a5),
	.w5(32'hbbfc84ba),
	.w6(32'hbb3cbcf7),
	.w7(32'hbba97cd7),
	.w8(32'h3a784174),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d2ba9),
	.w1(32'h3b037557),
	.w2(32'hbab222bc),
	.w3(32'h3b2aec4e),
	.w4(32'hba42c0c5),
	.w5(32'hbb2230c2),
	.w6(32'h3a5a162a),
	.w7(32'hbb5a419d),
	.w8(32'hbb1f38ac),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0636ef),
	.w1(32'hbb600ea9),
	.w2(32'hbb4b6784),
	.w3(32'h35bf6061),
	.w4(32'h3a88f71d),
	.w5(32'h3adf3234),
	.w6(32'h39816ff0),
	.w7(32'h3b6c73ed),
	.w8(32'h3b15b536),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33ef2b),
	.w1(32'h39f83b9b),
	.w2(32'h3a16b179),
	.w3(32'h39d6d24c),
	.w4(32'h39b3dd35),
	.w5(32'hba7c19e9),
	.w6(32'h39b5f34b),
	.w7(32'h3a12ce3c),
	.w8(32'hbabfdb08),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba557c89),
	.w1(32'hba623b1c),
	.w2(32'hba08735e),
	.w3(32'hba395a36),
	.w4(32'hba0b3514),
	.w5(32'h3994a516),
	.w6(32'hba889e84),
	.w7(32'hba0826b2),
	.w8(32'hba1096e2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd9506),
	.w1(32'h3aec325c),
	.w2(32'hbb8263ca),
	.w3(32'hbb5179ea),
	.w4(32'h3bdbe346),
	.w5(32'h3b112300),
	.w6(32'hbb98c1ad),
	.w7(32'h3ac53ba2),
	.w8(32'h3a0367c2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9917e6),
	.w1(32'hbb45901f),
	.w2(32'hbb2148c9),
	.w3(32'hbabf6774),
	.w4(32'hbb042a6a),
	.w5(32'h38fb6324),
	.w6(32'hba78ae54),
	.w7(32'hbb0c3846),
	.w8(32'h3a055afd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23201b),
	.w1(32'hb9fd25b6),
	.w2(32'h392f99b4),
	.w3(32'hba8eea70),
	.w4(32'h3bc70b4b),
	.w5(32'h3b60c7ed),
	.w6(32'hbb9d963d),
	.w7(32'h3b18d14c),
	.w8(32'h3acc9ac7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973d9b1),
	.w1(32'h3a39b3d6),
	.w2(32'h38362a95),
	.w3(32'h3a8dfae0),
	.w4(32'h3a9e2e76),
	.w5(32'h38f7bb6b),
	.w6(32'h39e2c15c),
	.w7(32'h39c740c3),
	.w8(32'hb9306bcb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941a031),
	.w1(32'h390dea74),
	.w2(32'hb3f84aae),
	.w3(32'h39862bff),
	.w4(32'h385fdaec),
	.w5(32'hb9bd52ee),
	.w6(32'h39d1e533),
	.w7(32'hb9385331),
	.w8(32'hb9e35536),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0806fe),
	.w1(32'h39b81b9b),
	.w2(32'hb9e892da),
	.w3(32'hba4d1fe2),
	.w4(32'hb95ab495),
	.w5(32'hba5dc536),
	.w6(32'hba4eaf59),
	.w7(32'hbac7ccaa),
	.w8(32'hbadcc63b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c98ae),
	.w1(32'hb9f74396),
	.w2(32'h3a10155a),
	.w3(32'hba9c77a9),
	.w4(32'hb9b9d172),
	.w5(32'h3ab0ac9e),
	.w6(32'hba523585),
	.w7(32'h39f7f77e),
	.w8(32'h3a9b5f1d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bd922),
	.w1(32'h39bff083),
	.w2(32'hba8cb4b1),
	.w3(32'hba5a788d),
	.w4(32'hbaf76e32),
	.w5(32'hbacd18ad),
	.w6(32'hba0bb6b7),
	.w7(32'hbab83cc0),
	.w8(32'hba85d989),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e5321),
	.w1(32'h3af18900),
	.w2(32'h3ab433ea),
	.w3(32'h3ae3b032),
	.w4(32'hbb3e41e4),
	.w5(32'hbb02310f),
	.w6(32'h3b5e487e),
	.w7(32'hb99de193),
	.w8(32'hba0a97f8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06c47c),
	.w1(32'h3be4178c),
	.w2(32'hbb7dbb84),
	.w3(32'h3c0fa5ea),
	.w4(32'hbb86ab07),
	.w5(32'hbc688fce),
	.w6(32'h3ba4d66a),
	.w7(32'hbc113159),
	.w8(32'hbc84b705),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99dd17),
	.w1(32'h39d0bc12),
	.w2(32'hbafb4708),
	.w3(32'hba8c22ca),
	.w4(32'h3b921873),
	.w5(32'hbabb031c),
	.w6(32'h3a7c8305),
	.w7(32'h3bdfdf4c),
	.w8(32'hbacdd1c0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb863c6f),
	.w1(32'hbb49726a),
	.w2(32'hbaab6005),
	.w3(32'hbb8c81fa),
	.w4(32'h3b587efa),
	.w5(32'h3ba9ae88),
	.w6(32'hbb851080),
	.w7(32'h3b883280),
	.w8(32'h3be937bf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc3f13),
	.w1(32'h3a950902),
	.w2(32'hb98ca182),
	.w3(32'h3afff61a),
	.w4(32'h3ae1c4cf),
	.w5(32'h3a8e7b6a),
	.w6(32'h3ae54fd0),
	.w7(32'h3ad31be6),
	.w8(32'h3ac6cb7e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ca339),
	.w1(32'hb92ba230),
	.w2(32'hba64c3fb),
	.w3(32'h3887f29a),
	.w4(32'h3667f65b),
	.w5(32'h39a5df84),
	.w6(32'h398e8daf),
	.w7(32'hba341af4),
	.w8(32'h399fafa4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395dfcb1),
	.w1(32'h390fdef5),
	.w2(32'h3a2b530f),
	.w3(32'h39517b8b),
	.w4(32'h3a5e3638),
	.w5(32'hba45110a),
	.w6(32'h38da5be5),
	.w7(32'h3a90912f),
	.w8(32'hba810f18),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7d8bb),
	.w1(32'h39541312),
	.w2(32'hba1f7b5b),
	.w3(32'hb912b87c),
	.w4(32'hb90357c4),
	.w5(32'hb999b057),
	.w6(32'h3699b21e),
	.w7(32'hb8f46f29),
	.w8(32'hba2dbc5c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fb5b8),
	.w1(32'h3b78dbde),
	.w2(32'hbb15f600),
	.w3(32'h3b160f94),
	.w4(32'h393ed48a),
	.w5(32'h39eef61b),
	.w6(32'h3abac17e),
	.w7(32'hbaf996ae),
	.w8(32'h3b51b401),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49895a),
	.w1(32'h3a8a8d9c),
	.w2(32'hba1e71d6),
	.w3(32'h3b27d397),
	.w4(32'h3ad36af3),
	.w5(32'hbaaf2e2e),
	.w6(32'hba2a8518),
	.w7(32'h38f87777),
	.w8(32'hbb451d9e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add370e),
	.w1(32'h3a10d06d),
	.w2(32'hb9d14500),
	.w3(32'h3b6db9e8),
	.w4(32'hb9f40e26),
	.w5(32'hbb3cf28e),
	.w6(32'h3a804550),
	.w7(32'hba0d6ec7),
	.w8(32'hbb8481f0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398751f1),
	.w1(32'hb928182a),
	.w2(32'hba9e6e1c),
	.w3(32'hba04f046),
	.w4(32'h3a0a072a),
	.w5(32'hba36ceac),
	.w6(32'hbb52ad25),
	.w7(32'hbac4ea17),
	.w8(32'hb9c3cf73),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc620aa),
	.w1(32'h3b935eb8),
	.w2(32'hba95eec6),
	.w3(32'h3bb88ef8),
	.w4(32'h39bb3766),
	.w5(32'h3a50f47c),
	.w6(32'h3c1212ae),
	.w7(32'h3995c5ec),
	.w8(32'h3a37bf12),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365441fa),
	.w1(32'h3981ad65),
	.w2(32'hb9232264),
	.w3(32'hba16d20d),
	.w4(32'hba179bea),
	.w5(32'h3ae71a5f),
	.w6(32'hba0d4a86),
	.w7(32'hba73507c),
	.w8(32'h3ad81bc2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215f1e),
	.w1(32'h3ae223fb),
	.w2(32'h3ab30fc2),
	.w3(32'h3b183c8e),
	.w4(32'h3af0e817),
	.w5(32'hbabaf2b4),
	.w6(32'h3a97b232),
	.w7(32'h3a94a8b3),
	.w8(32'hbaaca6e9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45a163),
	.w1(32'hb982a44a),
	.w2(32'hba2b3f26),
	.w3(32'hba0c35f8),
	.w4(32'hba119326),
	.w5(32'hb9de2656),
	.w6(32'hba5e88c2),
	.w7(32'hba8b2c1c),
	.w8(32'hba855e08),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4f48d),
	.w1(32'h3a6e3b58),
	.w2(32'h39cc9a78),
	.w3(32'h3a11dd54),
	.w4(32'h39e5da7e),
	.w5(32'hba88d3a0),
	.w6(32'hba187fcc),
	.w7(32'h3a943f18),
	.w8(32'h3a1656d2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca656c),
	.w1(32'hba83493d),
	.w2(32'hba8126f6),
	.w3(32'hbaa6cfaa),
	.w4(32'hba06039b),
	.w5(32'h3b00974f),
	.w6(32'hba734621),
	.w7(32'hbaeb471d),
	.w8(32'h3a96c93f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e3768),
	.w1(32'h3b128cd4),
	.w2(32'h3a5791a0),
	.w3(32'h3a4c0a27),
	.w4(32'hb9dc8db8),
	.w5(32'hba314051),
	.w6(32'h3a3b3581),
	.w7(32'hbbac563e),
	.w8(32'hbb7df730),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45ffe2),
	.w1(32'h3943ceb4),
	.w2(32'hbaa5a837),
	.w3(32'hbadf426e),
	.w4(32'hba5806f1),
	.w5(32'h3a188b38),
	.w6(32'hba849941),
	.w7(32'hb9de27cf),
	.w8(32'h3a4d3e0c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86d870),
	.w1(32'h3a28bfd8),
	.w2(32'h37f62a80),
	.w3(32'hb9caf5eb),
	.w4(32'hba6e1b98),
	.w5(32'h39e9324c),
	.w6(32'h39818e2f),
	.w7(32'hba495619),
	.w8(32'h39f78761),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c36759),
	.w1(32'h37e9efe5),
	.w2(32'hb87186ee),
	.w3(32'h386ad1e7),
	.w4(32'hb8ac92ea),
	.w5(32'h3981f4e0),
	.w6(32'h392c769d),
	.w7(32'hb994b60b),
	.w8(32'h3a842265),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38241dfa),
	.w1(32'h39f802a1),
	.w2(32'hb99aaa9e),
	.w3(32'h398fa277),
	.w4(32'h3a2030a2),
	.w5(32'h3af759e1),
	.w6(32'h39bee0b8),
	.w7(32'hb8aaea0a),
	.w8(32'h3affbd53),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd7031),
	.w1(32'h3a937967),
	.w2(32'h3aa9f5f5),
	.w3(32'h3ab6dc18),
	.w4(32'h3ab83f40),
	.w5(32'hb9921e97),
	.w6(32'h3aa74647),
	.w7(32'h3acbec01),
	.w8(32'hba26b5d3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d1b92),
	.w1(32'hb96fdfd1),
	.w2(32'h3a96a925),
	.w3(32'hb9a74585),
	.w4(32'h3a6cb0bf),
	.w5(32'hb6152994),
	.w6(32'hba7ebc99),
	.w7(32'h3aaee864),
	.w8(32'hb901867f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56d637),
	.w1(32'hb8943660),
	.w2(32'hba9cca70),
	.w3(32'h3a1d3fcc),
	.w4(32'hb89de7c8),
	.w5(32'h39bac60d),
	.w6(32'hba5467f7),
	.w7(32'hbb037549),
	.w8(32'h3a8f90d4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafe69d),
	.w1(32'h3b941556),
	.w2(32'hba8ac2b2),
	.w3(32'hbaf3656c),
	.w4(32'h3b86c4e8),
	.w5(32'hba641186),
	.w6(32'hbb56a462),
	.w7(32'h3b28bb1a),
	.w8(32'h3a215b6c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba114708),
	.w1(32'hba9bc924),
	.w2(32'hbaaa5cd3),
	.w3(32'hba8580a4),
	.w4(32'hbab7a1f3),
	.w5(32'h3a407eb0),
	.w6(32'hba120991),
	.w7(32'hba88467e),
	.w8(32'h3a4de7c9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88a803),
	.w1(32'hba391497),
	.w2(32'hba91f2ad),
	.w3(32'hba23a598),
	.w4(32'hba8ab6a1),
	.w5(32'h3ac42eda),
	.w6(32'hba372e01),
	.w7(32'hbad826c0),
	.w8(32'h3a8f8f86),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a400d66),
	.w1(32'h38beb8a3),
	.w2(32'hba0a82ab),
	.w3(32'h39ebde89),
	.w4(32'h39832714),
	.w5(32'hb9ca5622),
	.w6(32'h39c9cb20),
	.w7(32'hb89f4f02),
	.w8(32'hba50e04f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11a79d),
	.w1(32'hbad0396c),
	.w2(32'hbad37f1c),
	.w3(32'h3751172f),
	.w4(32'h39110c47),
	.w5(32'h3a3933a3),
	.w6(32'hba4a71df),
	.w7(32'hba6f62c8),
	.w8(32'h3a0159ae),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfa689),
	.w1(32'h3c0875d8),
	.w2(32'h3abfc56a),
	.w3(32'hbc047d62),
	.w4(32'h3ab26ed3),
	.w5(32'hbae9c7f9),
	.w6(32'hbb925f8b),
	.w7(32'hbba04e4d),
	.w8(32'hba50cec2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd71fe1),
	.w1(32'hbb95aade),
	.w2(32'hbadcdea5),
	.w3(32'hbb897e4c),
	.w4(32'hbbd1e1c2),
	.w5(32'hba293a40),
	.w6(32'hbb200db4),
	.w7(32'hbab0348e),
	.w8(32'h3a67af44),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a9ef5),
	.w1(32'h3a1429bb),
	.w2(32'hbafbf4ba),
	.w3(32'hbb90b8e1),
	.w4(32'hbb94a861),
	.w5(32'h3a415fbf),
	.w6(32'hbb8391b5),
	.w7(32'hbb2575a7),
	.w8(32'h3aa8a8bf),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7d0c0),
	.w1(32'h3a39ec45),
	.w2(32'h3aceada8),
	.w3(32'h3b897a9b),
	.w4(32'h3bacfc6c),
	.w5(32'hbb038a3f),
	.w6(32'h3b4d3070),
	.w7(32'h3bd57263),
	.w8(32'hbaf149c5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf3310),
	.w1(32'h39847f4f),
	.w2(32'hb9afac42),
	.w3(32'h383067d7),
	.w4(32'hb9b2483f),
	.w5(32'hbaa8a906),
	.w6(32'h37556417),
	.w7(32'hb91acf16),
	.w8(32'hbab27524),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba499f39),
	.w1(32'h3a2c2035),
	.w2(32'hba915366),
	.w3(32'h37d63569),
	.w4(32'hb8d5134c),
	.w5(32'hba83abcd),
	.w6(32'h3a827166),
	.w7(32'hba3d7da8),
	.w8(32'h39464c7e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f00369),
	.w1(32'hba9a74fa),
	.w2(32'hbaa33b75),
	.w3(32'hbaa0b0db),
	.w4(32'hba859a92),
	.w5(32'hba7ab14d),
	.w6(32'h3a5f7fc8),
	.w7(32'h3a435ef3),
	.w8(32'hba74391a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6858c5),
	.w1(32'hb9f2eb0a),
	.w2(32'hbab023b4),
	.w3(32'hba83e261),
	.w4(32'hbaa4530e),
	.w5(32'h3a266fc1),
	.w6(32'hb8d9f7ee),
	.w7(32'hb9a4ff66),
	.w8(32'h3a1d13ca),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f37607),
	.w1(32'hb9aafbd8),
	.w2(32'h39a54517),
	.w3(32'hb9310c82),
	.w4(32'h39498568),
	.w5(32'hbaca1784),
	.w6(32'hba71644a),
	.w7(32'hba19e488),
	.w8(32'hbae2cbe5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e4bfa),
	.w1(32'h3b4a1696),
	.w2(32'h3a84bafb),
	.w3(32'hba564ee3),
	.w4(32'hbb14273f),
	.w5(32'h37faa45e),
	.w6(32'hb8ee32a8),
	.w7(32'hbb5b3eea),
	.w8(32'hb9b2bc9f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8190fb),
	.w1(32'h3b567e44),
	.w2(32'hb9e8c10b),
	.w3(32'h3a99886b),
	.w4(32'hbb3c9944),
	.w5(32'hbabe85f9),
	.w6(32'h3b4d371b),
	.w7(32'hbb654ce8),
	.w8(32'hbb2e799f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696583),
	.w1(32'h3ae1bc89),
	.w2(32'hba3eb55f),
	.w3(32'h3bb66bbe),
	.w4(32'h3bae5f42),
	.w5(32'h39ed54c0),
	.w6(32'h3b92057c),
	.w7(32'h3ba8e40d),
	.w8(32'h3a8b1405),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27325d),
	.w1(32'h3ad6b83c),
	.w2(32'h3b041254),
	.w3(32'hbb3e48f8),
	.w4(32'hba03ee6f),
	.w5(32'h3b0e2d21),
	.w6(32'hbadfd87f),
	.w7(32'hba00e471),
	.w8(32'h3a89306e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8f78e),
	.w1(32'h3b92c810),
	.w2(32'h39e52bb3),
	.w3(32'hbb3bc6d2),
	.w4(32'hbaa183f1),
	.w5(32'hba64637a),
	.w6(32'hbb3fae51),
	.w7(32'hbb691ffd),
	.w8(32'hbb0a8145),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab22a0b),
	.w1(32'h3a123a3b),
	.w2(32'hbb113710),
	.w3(32'hb8f61a2d),
	.w4(32'hb89afbf5),
	.w5(32'hbb10627c),
	.w6(32'hbaedef6f),
	.w7(32'hbb0ae5bd),
	.w8(32'hbb173d68),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918082d),
	.w1(32'h3ad13dae),
	.w2(32'h3a500e47),
	.w3(32'h3a052bd2),
	.w4(32'h39ee3d1e),
	.w5(32'h3aaf24d4),
	.w6(32'h3b0fc453),
	.w7(32'h3a7ca930),
	.w8(32'h3b039cb1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39febeb4),
	.w1(32'h39a60663),
	.w2(32'hb9e405b9),
	.w3(32'h3a81bd23),
	.w4(32'h3a211383),
	.w5(32'h3a1e7c5c),
	.w6(32'h3a9d640f),
	.w7(32'h39cf41d5),
	.w8(32'h3a60c9a4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ac672),
	.w1(32'hb98d2070),
	.w2(32'hba2e2e5a),
	.w3(32'hba0b3d79),
	.w4(32'hb930fd9c),
	.w5(32'hb94f6acb),
	.w6(32'hba0f21bb),
	.w7(32'hba5874fe),
	.w8(32'h394a7619),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba143c0c),
	.w1(32'hba016278),
	.w2(32'hba3d5610),
	.w3(32'hb884cbb1),
	.w4(32'hb90ebcf7),
	.w5(32'h3a4520ce),
	.w6(32'hb78f451c),
	.w7(32'hb8fcbbac),
	.w8(32'h39d80e5b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ebecc),
	.w1(32'h398509a4),
	.w2(32'h3a5a6f8f),
	.w3(32'h3a4bba29),
	.w4(32'h3a90187a),
	.w5(32'h3a81c2f9),
	.w6(32'hb9aadfd2),
	.w7(32'h3a15f186),
	.w8(32'h3a7adafe),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59816f),
	.w1(32'h39561be4),
	.w2(32'hb8604c8b),
	.w3(32'h3a3c761d),
	.w4(32'h39dd4c04),
	.w5(32'hbab39027),
	.w6(32'h3a09eb08),
	.w7(32'h3a759a4e),
	.w8(32'hbb0a1087),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bffcdc),
	.w1(32'hba71961c),
	.w2(32'hbab50457),
	.w3(32'h3a8018ac),
	.w4(32'h39e59e3e),
	.w5(32'h391285ca),
	.w6(32'hb8e54f23),
	.w7(32'hb7e57c68),
	.w8(32'hb9395494),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a615bea),
	.w1(32'h3acfe290),
	.w2(32'h3b04fa34),
	.w3(32'h3b97726f),
	.w4(32'h3af07056),
	.w5(32'h3ac3f8c7),
	.w6(32'h3ae7476c),
	.w7(32'h3ad28743),
	.w8(32'h3a616102),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1579b7),
	.w1(32'h3b49e1a2),
	.w2(32'h3b2c169c),
	.w3(32'h3ae5f18a),
	.w4(32'h3af1d096),
	.w5(32'h3aa4dfcf),
	.w6(32'h3b82bb24),
	.w7(32'h3b1158aa),
	.w8(32'h3b12255d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2bed5),
	.w1(32'hb98aa2f9),
	.w2(32'hbadf0a98),
	.w3(32'hbaa0a812),
	.w4(32'h3a0f2010),
	.w5(32'hba737143),
	.w6(32'hbab866ff),
	.w7(32'hb9c6531d),
	.w8(32'hb99eaf19),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12d36f),
	.w1(32'hb9973352),
	.w2(32'hbac8ab61),
	.w3(32'h3add3199),
	.w4(32'hbba31663),
	.w5(32'hbbc7f627),
	.w6(32'hbb5c1c4d),
	.w7(32'hbc109c28),
	.w8(32'hbbcc5404),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacaa86),
	.w1(32'h39d6e9ad),
	.w2(32'hb80a2d96),
	.w3(32'hba99a8f7),
	.w4(32'h3a855d9e),
	.w5(32'hb9a7f021),
	.w6(32'h3a28ff0a),
	.w7(32'h3aa0156a),
	.w8(32'hba5a6cb4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a581d),
	.w1(32'h3ae6d69a),
	.w2(32'h3b0f69f5),
	.w3(32'hbb459762),
	.w4(32'hb91d0bab),
	.w5(32'h3b7bb141),
	.w6(32'hbb887097),
	.w7(32'hbb83b777),
	.w8(32'h3a25ae3c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b054dd9),
	.w1(32'h3a010fb7),
	.w2(32'hba782846),
	.w3(32'hba880d30),
	.w4(32'h3793cfca),
	.w5(32'hba3093f9),
	.w6(32'hbb778c2d),
	.w7(32'hbb388e77),
	.w8(32'hb982c863),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3ebea),
	.w1(32'h3ab54810),
	.w2(32'h39ffbfdf),
	.w3(32'h38b4e0b7),
	.w4(32'h3b88870f),
	.w5(32'h3b049354),
	.w6(32'hba3c29a5),
	.w7(32'h3b76378b),
	.w8(32'h3a6d4c87),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397bc89b),
	.w1(32'h39aae40a),
	.w2(32'h39f36282),
	.w3(32'h3a226fe2),
	.w4(32'h39f73245),
	.w5(32'h3a63bbce),
	.w6(32'hb9152de6),
	.w7(32'h3a19db70),
	.w8(32'h3a0728e5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58b4b8),
	.w1(32'h3b79944f),
	.w2(32'h39689d4b),
	.w3(32'h3a88f5a0),
	.w4(32'hb9d10f11),
	.w5(32'hb8380a75),
	.w6(32'h3ab58954),
	.w7(32'hbb3a238f),
	.w8(32'hb9600826),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf961c9),
	.w1(32'h3bb3fbe6),
	.w2(32'hbb34af16),
	.w3(32'hbb57f4cd),
	.w4(32'hbbaff74c),
	.w5(32'hbc07e410),
	.w6(32'hbb8eedea),
	.w7(32'hbc148204),
	.w8(32'hbbe1d2c4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4450b),
	.w1(32'hba19aaf6),
	.w2(32'hba4dd7be),
	.w3(32'h3c384885),
	.w4(32'hbba665f9),
	.w5(32'hbc530bf7),
	.w6(32'h3c3a1757),
	.w7(32'h3b52b10d),
	.w8(32'hbb6bb149),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c812e),
	.w1(32'h3a9fa40c),
	.w2(32'hbb56b9cd),
	.w3(32'h3b3199ff),
	.w4(32'hbb2670e7),
	.w5(32'hbae6c4a8),
	.w6(32'h3c0d1375),
	.w7(32'h3be9a975),
	.w8(32'hb99eb8cb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf442d6),
	.w1(32'h3b7f9618),
	.w2(32'h3b07317d),
	.w3(32'h3b5681fd),
	.w4(32'h3b099d5f),
	.w5(32'hba74b88f),
	.w6(32'h3be41256),
	.w7(32'h3bd0059f),
	.w8(32'hba46f00d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94c187),
	.w1(32'h3bce262d),
	.w2(32'h3b042b1f),
	.w3(32'hba048e0c),
	.w4(32'hbc1553d5),
	.w5(32'hbb9fe250),
	.w6(32'hb6819966),
	.w7(32'hbc1279e5),
	.w8(32'hbb331c9e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b256da1),
	.w1(32'h3b547668),
	.w2(32'h3ab9a2a6),
	.w3(32'h3aa87886),
	.w4(32'hba84a519),
	.w5(32'h3b8785c9),
	.w6(32'h3b87b45c),
	.w7(32'hba0b1750),
	.w8(32'h3bc50a36),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1341d3),
	.w1(32'h3b688c19),
	.w2(32'h3abf173f),
	.w3(32'h3c8f08e5),
	.w4(32'h39a5ea00),
	.w5(32'hbc061af9),
	.w6(32'h3c06cc7a),
	.w7(32'hbba5096c),
	.w8(32'hbc44ff2e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eb805),
	.w1(32'h3aec58b4),
	.w2(32'h3b3a1a2e),
	.w3(32'h3b1dadd2),
	.w4(32'hba9f54a2),
	.w5(32'hbb937fc8),
	.w6(32'h3a666e1e),
	.w7(32'hb7d2cb48),
	.w8(32'hbb8c9150),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba776d35),
	.w1(32'h3ad63aeb),
	.w2(32'h3b1d778d),
	.w3(32'hb996ebf3),
	.w4(32'h38c3b4ae),
	.w5(32'h3ac6998d),
	.w6(32'h38b6ed4d),
	.w7(32'h3a4506a5),
	.w8(32'h3b9cb779),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92211c),
	.w1(32'hba7a64b9),
	.w2(32'h3a8d0e20),
	.w3(32'h3a1fe7f1),
	.w4(32'h3aa6c05d),
	.w5(32'hbab5e20d),
	.w6(32'h3bba6713),
	.w7(32'h3bd2e9d0),
	.w8(32'hba1b8b56),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e80fc),
	.w1(32'h3b02b0e9),
	.w2(32'hbb05417d),
	.w3(32'h383108ad),
	.w4(32'hbb824c9d),
	.w5(32'h3b969514),
	.w6(32'h3a8a738a),
	.w7(32'hbb07a734),
	.w8(32'h3bc154fc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2094b5),
	.w1(32'h3bdf97d3),
	.w2(32'h3bad9558),
	.w3(32'h3b92578a),
	.w4(32'h3ba1c5f8),
	.w5(32'hbbaaf181),
	.w6(32'h3b142aa1),
	.w7(32'h3b75b822),
	.w8(32'hb9080da6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6356b4),
	.w1(32'h3b182e82),
	.w2(32'hbabc3033),
	.w3(32'h3998c5e1),
	.w4(32'h3b47dbb2),
	.w5(32'h3b910144),
	.w6(32'h3b0c45e4),
	.w7(32'h3b4a345d),
	.w8(32'h3bfeeb2f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb32e2e),
	.w1(32'h3acaf088),
	.w2(32'h3afd9e20),
	.w3(32'h3b1c3358),
	.w4(32'h3baaff4a),
	.w5(32'h3b95d560),
	.w6(32'h3a22f8c6),
	.w7(32'h3b27fc8a),
	.w8(32'hbac1ef99),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba953e4c),
	.w1(32'hbba3fcb5),
	.w2(32'hbba5ddcc),
	.w3(32'h3bca82f1),
	.w4(32'hba91c292),
	.w5(32'h3b47930c),
	.w6(32'hbbb809f6),
	.w7(32'hbc04e2b6),
	.w8(32'hb9968026),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba389b0),
	.w1(32'h3b2f193f),
	.w2(32'h3b225ca7),
	.w3(32'h3c04d4bf),
	.w4(32'h3c1bf791),
	.w5(32'h39aeb2e5),
	.w6(32'hb98ccb60),
	.w7(32'h3b619d39),
	.w8(32'h3b85abdc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba13eb1),
	.w1(32'h3bb6f4eb),
	.w2(32'hba1071c0),
	.w3(32'h3ab58def),
	.w4(32'hba2eb609),
	.w5(32'hbaa67ac8),
	.w6(32'h3b83e4a0),
	.w7(32'h3a156467),
	.w8(32'h3aee516f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eae42),
	.w1(32'hbabc57be),
	.w2(32'h39d49cef),
	.w3(32'hba7e7841),
	.w4(32'hb93aacba),
	.w5(32'h3b96c8d9),
	.w6(32'h3ad9c851),
	.w7(32'hb98038af),
	.w8(32'h3a5e7398),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7db5fe),
	.w1(32'h3b6c9a5c),
	.w2(32'h3bb0038f),
	.w3(32'h3ad40fd6),
	.w4(32'h3ba4b845),
	.w5(32'h3a11fade),
	.w6(32'h3a902aa3),
	.w7(32'h3be20b1a),
	.w8(32'h3be2b14b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e3b8b),
	.w1(32'hbb242329),
	.w2(32'hbb6d85ad),
	.w3(32'hbb269eef),
	.w4(32'hbb8ca572),
	.w5(32'h3b419ecf),
	.w6(32'h3accfd7c),
	.w7(32'h3b1131c5),
	.w8(32'h3994b46b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14d259),
	.w1(32'hbacab064),
	.w2(32'hbbec1c37),
	.w3(32'h3a84f8e4),
	.w4(32'hbb9978d3),
	.w5(32'h3ab84c34),
	.w6(32'hb966ab9a),
	.w7(32'hbba4c079),
	.w8(32'h3b94c4e8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5636df),
	.w1(32'h3bb039c3),
	.w2(32'hbb855299),
	.w3(32'h3c1717b9),
	.w4(32'hbac4a73f),
	.w5(32'hbb8ca16a),
	.w6(32'h3c208323),
	.w7(32'hbaa08207),
	.w8(32'hbb0da088),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b479873),
	.w1(32'h3b417e1f),
	.w2(32'h3b080b55),
	.w3(32'h38d40c7b),
	.w4(32'h3af26c91),
	.w5(32'hbb765139),
	.w6(32'h3aef3f09),
	.w7(32'h3a86fdc8),
	.w8(32'hbbcfcca3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26d1a4),
	.w1(32'hbac5ee8c),
	.w2(32'hbbee393b),
	.w3(32'hbb0f407f),
	.w4(32'hbb81dcd0),
	.w5(32'h3af3bfbd),
	.w6(32'h3a3f61d1),
	.w7(32'hbbfd16cd),
	.w8(32'hbb27b8f7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b8971),
	.w1(32'h3a9a393a),
	.w2(32'h3ba47ead),
	.w3(32'h3bfdc39d),
	.w4(32'h3bf9b8f1),
	.w5(32'h3a646729),
	.w6(32'hba62aef4),
	.w7(32'h3b8e330b),
	.w8(32'hbadad3dc),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4f093),
	.w1(32'hbb231f6f),
	.w2(32'hbae90978),
	.w3(32'hbaa43246),
	.w4(32'h3b093a2e),
	.w5(32'h3a2c40f5),
	.w6(32'hbb180693),
	.w7(32'hbb47fba8),
	.w8(32'hba93f707),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9956ee),
	.w1(32'h3b0050ce),
	.w2(32'h3b5a70c6),
	.w3(32'hbb01edcb),
	.w4(32'hbb1cab72),
	.w5(32'hbb29ac6e),
	.w6(32'h3b5c33c6),
	.w7(32'h3a802874),
	.w8(32'hba425146),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1e637),
	.w1(32'hba87edf1),
	.w2(32'hb8c7fea9),
	.w3(32'hbb53b1aa),
	.w4(32'hbad3967d),
	.w5(32'hba5ab2f6),
	.w6(32'hbaaec36a),
	.w7(32'h3a2843a0),
	.w8(32'h3c0c73b2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87b1a6),
	.w1(32'h3a98e10d),
	.w2(32'hbadc2879),
	.w3(32'hbb184c9b),
	.w4(32'hbb67868f),
	.w5(32'hbaa14e3e),
	.w6(32'h3c5ca7ae),
	.w7(32'h3bd83f72),
	.w8(32'h3a868f5e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ff989),
	.w1(32'hbbd868da),
	.w2(32'hbb9f4dc1),
	.w3(32'hb984c673),
	.w4(32'hbc1c6d8f),
	.w5(32'h3bd46419),
	.w6(32'hbb066d17),
	.w7(32'hbb32696d),
	.w8(32'h3b9dbc59),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcfeef),
	.w1(32'hb8b303af),
	.w2(32'hb9983af9),
	.w3(32'h3b8c989c),
	.w4(32'h3b142d4f),
	.w5(32'hba0330c7),
	.w6(32'h3a09e401),
	.w7(32'hbb56df15),
	.w8(32'hbb274e8e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05ea45),
	.w1(32'h3990f0dc),
	.w2(32'hb99378e1),
	.w3(32'hba9d7cc8),
	.w4(32'hbb2857c0),
	.w5(32'h3a6a5267),
	.w6(32'h3916aa03),
	.w7(32'hbb9bcc88),
	.w8(32'h3b78176b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46b507),
	.w1(32'h3a3b6343),
	.w2(32'hbb982b41),
	.w3(32'hbb111255),
	.w4(32'hbb792dc7),
	.w5(32'hbb1e4493),
	.w6(32'h3be85912),
	.w7(32'h3a6bd38e),
	.w8(32'hbaf0b282),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72bdc2),
	.w1(32'hbaf7a341),
	.w2(32'hbb8b0dea),
	.w3(32'hbb53c427),
	.w4(32'hbba4022a),
	.w5(32'hbbdf5450),
	.w6(32'hbb1038c8),
	.w7(32'hbb77753c),
	.w8(32'hbaffc23a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b327159),
	.w1(32'h3ad349fe),
	.w2(32'h3a43125d),
	.w3(32'hbb655235),
	.w4(32'hbb3cd09b),
	.w5(32'h3b322936),
	.w6(32'h3a29aa36),
	.w7(32'hbaa7a31e),
	.w8(32'h3b8f7469),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd71748),
	.w1(32'h3bd703ec),
	.w2(32'h3b80e3a4),
	.w3(32'hbaa5dbf4),
	.w4(32'h3b0b2133),
	.w5(32'h3b2a59c2),
	.w6(32'h3aaf1c94),
	.w7(32'h3b63316b),
	.w8(32'h3b4215a1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a559b),
	.w1(32'h3ba1a039),
	.w2(32'h3a9e63e4),
	.w3(32'h3a3ffa85),
	.w4(32'hbb37804e),
	.w5(32'h38fcc327),
	.w6(32'h3c3609e9),
	.w7(32'h3b3745bc),
	.w8(32'hbaea7bce),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973b247),
	.w1(32'h3a23cc90),
	.w2(32'h3b24fd34),
	.w3(32'h3b6a964b),
	.w4(32'h3a1759b9),
	.w5(32'h393cdbd3),
	.w6(32'h3ba65b41),
	.w7(32'h3ba313d1),
	.w8(32'hbb866fab),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ab082),
	.w1(32'h3b421eaf),
	.w2(32'h3b16c183),
	.w3(32'h3a5ce5f1),
	.w4(32'h3aa27103),
	.w5(32'h3aa6160c),
	.w6(32'hbbd53c8f),
	.w7(32'hbb3306bb),
	.w8(32'h3ba7d1fd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c154bf8),
	.w1(32'h3bc5fb18),
	.w2(32'h3b2df063),
	.w3(32'h3b30a631),
	.w4(32'hbbae7312),
	.w5(32'hbb44f913),
	.w6(32'h3b997a53),
	.w7(32'hbb3f8346),
	.w8(32'hba7030a9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b0732),
	.w1(32'hbb193a1c),
	.w2(32'hbb126a9b),
	.w3(32'h3abee589),
	.w4(32'hbb92101d),
	.w5(32'h3b14ad35),
	.w6(32'h3ba8231c),
	.w7(32'h3aa30aae),
	.w8(32'h3ac56362),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafac2b),
	.w1(32'h39ca283e),
	.w2(32'hbb8f324d),
	.w3(32'h3bec4c8d),
	.w4(32'h3bab7547),
	.w5(32'h3aa4f053),
	.w6(32'h3b82c89e),
	.w7(32'hbb264b10),
	.w8(32'hbb7b1f45),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1c150),
	.w1(32'hb893118e),
	.w2(32'hb823231f),
	.w3(32'h3bcae218),
	.w4(32'h3bc8d575),
	.w5(32'hbb2ea396),
	.w6(32'hbacc2cdf),
	.w7(32'hbaf7ea0f),
	.w8(32'hbb7d28dc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc173b0),
	.w1(32'hbaa15443),
	.w2(32'hba014baa),
	.w3(32'hb9ebc32c),
	.w4(32'h3c00a3a5),
	.w5(32'h398ca5ea),
	.w6(32'hbbada163),
	.w7(32'h3af7d2c0),
	.w8(32'h3b90c3d1),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39490d82),
	.w1(32'hbb0a7916),
	.w2(32'hbb82435a),
	.w3(32'hb9d6e516),
	.w4(32'hbb0790a5),
	.w5(32'hbb1eb8be),
	.w6(32'h3b38cad0),
	.w7(32'hbb231654),
	.w8(32'hbb715c6c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b0bfd),
	.w1(32'hba88167d),
	.w2(32'hba887867),
	.w3(32'hba8c776e),
	.w4(32'hbb366919),
	.w5(32'h3bb692d0),
	.w6(32'hbb22ab1f),
	.w7(32'hbb6b0d3a),
	.w8(32'h3b292ede),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d2666),
	.w1(32'hbb9ee96e),
	.w2(32'hbaf0f60c),
	.w3(32'h3b2c9148),
	.w4(32'h3b7a9f68),
	.w5(32'h399ec225),
	.w6(32'hbb538d17),
	.w7(32'hbaaecf78),
	.w8(32'h38cd3d03),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b9620),
	.w1(32'h3b0dff2d),
	.w2(32'h3aa34d18),
	.w3(32'h3a831a5c),
	.w4(32'hba4bab9d),
	.w5(32'h3a9f4836),
	.w6(32'h3b044822),
	.w7(32'hba3712ff),
	.w8(32'h3b128c56),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aeadf),
	.w1(32'h38c82153),
	.w2(32'hba96aa30),
	.w3(32'h3bb361bf),
	.w4(32'h3b6e4013),
	.w5(32'h3a829c6c),
	.w6(32'h3ba1fd46),
	.w7(32'h3ace31bf),
	.w8(32'hbb0800fc),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc8d17),
	.w1(32'h3aa8019c),
	.w2(32'hb92f10e7),
	.w3(32'h3bbe967a),
	.w4(32'h3bbc6eca),
	.w5(32'h3a059382),
	.w6(32'h3bc3783d),
	.w7(32'h3bc39407),
	.w8(32'hb99ec884),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a903bee),
	.w1(32'hbb51eb4e),
	.w2(32'hba9a3d6b),
	.w3(32'hbb590109),
	.w4(32'hbb310de1),
	.w5(32'h3bc80e12),
	.w6(32'hbbb5b3ac),
	.w7(32'hbb088f2b),
	.w8(32'h3bc3ca90),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c9ad5),
	.w1(32'h3bc6ba3b),
	.w2(32'h3aee3d3a),
	.w3(32'h3b2d7f80),
	.w4(32'h3b364c38),
	.w5(32'h3b8be74f),
	.w6(32'h3ac03da0),
	.w7(32'h399f3407),
	.w8(32'h3b0c4a16),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00d818),
	.w1(32'h3b1b0852),
	.w2(32'h3980969c),
	.w3(32'h3bccaf44),
	.w4(32'h3ba272ab),
	.w5(32'hbbb27187),
	.w6(32'h3b405d38),
	.w7(32'h3adaf8f3),
	.w8(32'hbc3162e5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b780dd5),
	.w1(32'h3a8c5d40),
	.w2(32'h3ad3552a),
	.w3(32'hbb7a200e),
	.w4(32'hbb92f9bb),
	.w5(32'hba8a5d70),
	.w6(32'h3aae00ad),
	.w7(32'h388fa04a),
	.w8(32'h3adb48dc),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab90fe4),
	.w1(32'h3b78f79f),
	.w2(32'hbb1280a0),
	.w3(32'hba99a6bd),
	.w4(32'h3bbdf118),
	.w5(32'h3a7eb2b6),
	.w6(32'h39e5f6e8),
	.w7(32'h3b500d1a),
	.w8(32'h3beea1f5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0fa9a),
	.w1(32'hb9103a93),
	.w2(32'hba3deb99),
	.w3(32'h3a85c96a),
	.w4(32'hba68face),
	.w5(32'hbb619a2d),
	.w6(32'h3c0f3015),
	.w7(32'h3bf665b5),
	.w8(32'hbb23462e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb053e8),
	.w1(32'hbb8899f5),
	.w2(32'hbbe25cb4),
	.w3(32'hbb2e0c35),
	.w4(32'hbbdde1ed),
	.w5(32'h399fe4e0),
	.w6(32'hbb960a84),
	.w7(32'hbba4b0db),
	.w8(32'hbb5cd720),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8e41e),
	.w1(32'h3b49bb47),
	.w2(32'h3b986e40),
	.w3(32'h3a5379b3),
	.w4(32'h3b51cdd1),
	.w5(32'hbb6f09c9),
	.w6(32'hbba699f6),
	.w7(32'hb9a12a3a),
	.w8(32'hbb8cce03),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fa3d1),
	.w1(32'h3b3cb286),
	.w2(32'h3a1a9896),
	.w3(32'hb9ee42da),
	.w4(32'h39858214),
	.w5(32'hbb7b6ee1),
	.w6(32'hb92079b6),
	.w7(32'h3a7fb259),
	.w8(32'hbba4a690),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd758e2),
	.w1(32'hbb965a84),
	.w2(32'hbba1891e),
	.w3(32'hbb254438),
	.w4(32'hbac4099a),
	.w5(32'hbad20eff),
	.w6(32'hbaf3eda1),
	.w7(32'hbb804211),
	.w8(32'h3bf9d3ad),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0906f2),
	.w1(32'h3c324f59),
	.w2(32'h3c2efd87),
	.w3(32'hbb068a21),
	.w4(32'h3a693cb0),
	.w5(32'h3c255258),
	.w6(32'h3c6d6d9c),
	.w7(32'h3c244808),
	.w8(32'h3b730318),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c04614),
	.w1(32'h3ab5ba28),
	.w2(32'h392e83db),
	.w3(32'h3c2bca8e),
	.w4(32'h3c2a99f5),
	.w5(32'hb9aaff71),
	.w6(32'h3bd8797f),
	.w7(32'h3bcdd012),
	.w8(32'h3af604c7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ebff6),
	.w1(32'h3aeb55c8),
	.w2(32'hbb857118),
	.w3(32'h3b00e466),
	.w4(32'hbb1cba31),
	.w5(32'hbbb14406),
	.w6(32'h3bceb1c4),
	.w7(32'hbadec297),
	.w8(32'hbbb25a2c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f85ec),
	.w1(32'hb9541b8d),
	.w2(32'hb92ba43d),
	.w3(32'hbb57e18e),
	.w4(32'hbb65735e),
	.w5(32'h3ac3c31e),
	.w6(32'hb9b79446),
	.w7(32'hbb4c2294),
	.w8(32'h3a246adb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf1266),
	.w1(32'h3ae4c56d),
	.w2(32'h3913aebf),
	.w3(32'h3a4ea29c),
	.w4(32'h3aa0cd56),
	.w5(32'hbb06a0ef),
	.w6(32'h3a5cd4e9),
	.w7(32'h3b089936),
	.w8(32'hbb6e7181),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bf76a),
	.w1(32'h3ad3531b),
	.w2(32'h3a0a9a0c),
	.w3(32'hba9c62ca),
	.w4(32'hba570b58),
	.w5(32'h3a01c296),
	.w6(32'h3a851e68),
	.w7(32'h3b52d3af),
	.w8(32'h3bb4214a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8a167),
	.w1(32'h39ae3699),
	.w2(32'h3b2e2300),
	.w3(32'hbb45487f),
	.w4(32'hba374dfe),
	.w5(32'h3b30cb80),
	.w6(32'h3bb27605),
	.w7(32'h3bf0d764),
	.w8(32'h3b9d75a7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b096238),
	.w1(32'h3bb17194),
	.w2(32'hb8148c1e),
	.w3(32'h3b714b90),
	.w4(32'hbb2eed4e),
	.w5(32'hba4c3047),
	.w6(32'h3ae5f57d),
	.w7(32'hbb48b24a),
	.w8(32'h3a71f68d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f52fb),
	.w1(32'hba9ccc8e),
	.w2(32'h3af2d404),
	.w3(32'hbabb77ad),
	.w4(32'h3b2d9eb8),
	.w5(32'h3bc72bf2),
	.w6(32'h3b566676),
	.w7(32'h3b42980b),
	.w8(32'h3c0e250a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb1690),
	.w1(32'h3b9c259d),
	.w2(32'h3b32bcdc),
	.w3(32'h3b6663d0),
	.w4(32'h3b0acd0f),
	.w5(32'h3a6cc26a),
	.w6(32'hb9780114),
	.w7(32'hbb2c7763),
	.w8(32'hba95e066),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c1c6c),
	.w1(32'h3a71535a),
	.w2(32'hba8be8f0),
	.w3(32'h3bf12d7d),
	.w4(32'hbb0699e2),
	.w5(32'hbaeb11bb),
	.w6(32'h3b3d6fc9),
	.w7(32'hbb6c3e1a),
	.w8(32'h3ba622ee),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47c58d),
	.w1(32'hbb243a25),
	.w2(32'hbb855a3f),
	.w3(32'h3aced1ea),
	.w4(32'hbb780662),
	.w5(32'hb9197f7c),
	.w6(32'h3c520bb2),
	.w7(32'h3bb7f832),
	.w8(32'h3aabedb6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a0a1f),
	.w1(32'h3b44c2c0),
	.w2(32'h3a62a1d6),
	.w3(32'h3b8b7a3f),
	.w4(32'h3b62dfa4),
	.w5(32'h3ba4313d),
	.w6(32'h3aa71162),
	.w7(32'h3ba549ce),
	.w8(32'h3b6a2204),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03e29e),
	.w1(32'h3a90e222),
	.w2(32'hbb41fbf9),
	.w3(32'hbaf47f9e),
	.w4(32'hbace7db1),
	.w5(32'hbbe94f84),
	.w6(32'hbb034f6c),
	.w7(32'hb9aacd78),
	.w8(32'hbadd0b08),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a5769),
	.w1(32'h39faab3d),
	.w2(32'hbbe6ec1f),
	.w3(32'hba711932),
	.w4(32'hbbc4d5cd),
	.w5(32'h3a49db14),
	.w6(32'h3b8268ce),
	.w7(32'hbb8f37ab),
	.w8(32'h3c551a2f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc97160),
	.w1(32'h3b92acf3),
	.w2(32'h3b6a3dee),
	.w3(32'hbb5cee0a),
	.w4(32'h39cad35c),
	.w5(32'hbbe028b0),
	.w6(32'h3c5c32dd),
	.w7(32'h3c37f48f),
	.w8(32'hbb912d83),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb149980),
	.w1(32'hba53eeef),
	.w2(32'hbbeb391c),
	.w3(32'hbb741e20),
	.w4(32'hbbd84369),
	.w5(32'h3b86441f),
	.w6(32'hbaef2dad),
	.w7(32'hbc04fc1f),
	.w8(32'hbb35d1f4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07d6bd),
	.w1(32'h3961c13f),
	.w2(32'h3a51742f),
	.w3(32'hb9e1b1bb),
	.w4(32'h3b150fe3),
	.w5(32'hbb5a8e3e),
	.w6(32'hbc0632a2),
	.w7(32'hbb72606a),
	.w8(32'hbbc7528d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cc3b3),
	.w1(32'hbb710ec4),
	.w2(32'hbb29de67),
	.w3(32'hbbbb4a8e),
	.w4(32'hba96fef3),
	.w5(32'h3b3ef046),
	.w6(32'hbbfbaf6f),
	.w7(32'hbbb337a9),
	.w8(32'h3bb3b858),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9cfa6),
	.w1(32'h3b19e13c),
	.w2(32'hba30a356),
	.w3(32'h3b2cd221),
	.w4(32'hbab6aa9b),
	.w5(32'hbbc35042),
	.w6(32'h3bde4b0f),
	.w7(32'h3aea86b1),
	.w8(32'hbb90ecb8),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39127d57),
	.w1(32'h3b57dad4),
	.w2(32'h3bb6f6ce),
	.w3(32'hbad151d4),
	.w4(32'h3ab28a8d),
	.w5(32'h3ac8ed97),
	.w6(32'h3913c1b7),
	.w7(32'h3b87b36b),
	.w8(32'h3b83624e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeab323),
	.w1(32'h39b6096b),
	.w2(32'h37e94f03),
	.w3(32'hba02defa),
	.w4(32'hbb002123),
	.w5(32'hbb83f215),
	.w6(32'h3a99b141),
	.w7(32'h3ab7da70),
	.w8(32'hba05b2bc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b7602),
	.w1(32'h39dfb0fd),
	.w2(32'hbb86f078),
	.w3(32'hbb23e1dd),
	.w4(32'h39e076ec),
	.w5(32'h3b01b5bf),
	.w6(32'hba21bc68),
	.w7(32'h398fe6d7),
	.w8(32'h3bdc5e66),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ecfc8),
	.w1(32'h3b8d2d27),
	.w2(32'h3b400f5a),
	.w3(32'h3b2b050a),
	.w4(32'h3b1583fa),
	.w5(32'h3b7fb650),
	.w6(32'h3c1147c8),
	.w7(32'h3b4d98f7),
	.w8(32'h3b393f8c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02f2ca),
	.w1(32'h3a267492),
	.w2(32'h3aa9d3af),
	.w3(32'h3abc84b8),
	.w4(32'hba796f8c),
	.w5(32'hbb63007a),
	.w6(32'h3b4f3c40),
	.w7(32'h3a94ac16),
	.w8(32'hbb3fc8ba),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e6e77),
	.w1(32'h38cf9f35),
	.w2(32'h3a8c1e3e),
	.w3(32'hbb2e4e2c),
	.w4(32'hbb6a5962),
	.w5(32'h3b276c89),
	.w6(32'h37d3b940),
	.w7(32'h3adba168),
	.w8(32'h3a846fa4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f039f),
	.w1(32'h39057a60),
	.w2(32'h3988ea34),
	.w3(32'hbb6d69d4),
	.w4(32'hbba6592b),
	.w5(32'h3b2020de),
	.w6(32'hbc0003b5),
	.w7(32'hbbaf5537),
	.w8(32'h3bba802e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd47c7),
	.w1(32'h3c0336ae),
	.w2(32'hb9257228),
	.w3(32'h3c102c0e),
	.w4(32'hbb3bd096),
	.w5(32'hbb2a58e1),
	.w6(32'h3ba6fc13),
	.w7(32'hbbb70ab7),
	.w8(32'hbb91a2df),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba211f07),
	.w1(32'h3abb95d6),
	.w2(32'h3a404126),
	.w3(32'h3b799b12),
	.w4(32'h3a003844),
	.w5(32'hbb373aad),
	.w6(32'h3bf469a3),
	.w7(32'h3bac0de6),
	.w8(32'hbbd102bd),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2603f3),
	.w1(32'h3b0aebb9),
	.w2(32'hbb933ddf),
	.w3(32'h3acf7678),
	.w4(32'hbbec0bae),
	.w5(32'h3b170a91),
	.w6(32'hbc2410f9),
	.w7(32'hbc87f6be),
	.w8(32'h3a3081ef),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ef867),
	.w1(32'h3b6ec384),
	.w2(32'hbb1c79e5),
	.w3(32'hbb32b194),
	.w4(32'h3b9e8ad4),
	.w5(32'hbb519b81),
	.w6(32'hbb2dbd87),
	.w7(32'hb9bff0c4),
	.w8(32'h3bc3ec11),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0905),
	.w1(32'h3b11ddb7),
	.w2(32'hb98c8141),
	.w3(32'h3b04ea33),
	.w4(32'hbaacb42e),
	.w5(32'hbb51a476),
	.w6(32'h3c3860e0),
	.w7(32'h3b8324ee),
	.w8(32'h39f5ecf7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d5110),
	.w1(32'hbae5781a),
	.w2(32'hba8ab588),
	.w3(32'hbb5e87f4),
	.w4(32'hbb655ea5),
	.w5(32'hba8d5000),
	.w6(32'h3b08defd),
	.w7(32'h3a09ffda),
	.w8(32'hbad9856b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad88420),
	.w1(32'h3a0cfff6),
	.w2(32'h3a4371b0),
	.w3(32'h396b3db6),
	.w4(32'hba9c1b59),
	.w5(32'hbb858f8f),
	.w6(32'hbaa04b43),
	.w7(32'hba581362),
	.w8(32'hbb8aef81),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb548f4),
	.w1(32'h3b0c226a),
	.w2(32'h3b6e66f0),
	.w3(32'hb88dc4dc),
	.w4(32'hba95a720),
	.w5(32'hbb11bf9e),
	.w6(32'h3b3cfcbc),
	.w7(32'h3b5990d6),
	.w8(32'hba0549f0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9edcfe),
	.w1(32'hba64aa3b),
	.w2(32'hba8b16ff),
	.w3(32'hbb34391e),
	.w4(32'hbbe776c5),
	.w5(32'h3ba1a9c5),
	.w6(32'h3abb2ae3),
	.w7(32'hbb6b0da8),
	.w8(32'h3c19c7d4),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd61169),
	.w1(32'h3b328f52),
	.w2(32'hbac4f72f),
	.w3(32'h3a87063f),
	.w4(32'hbb4e090c),
	.w5(32'hbb76d460),
	.w6(32'h3bc970ac),
	.w7(32'hbb4fdc65),
	.w8(32'hbba8f3e6),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dc95b),
	.w1(32'h3b26c3e0),
	.w2(32'h3ade994c),
	.w3(32'h3a8d08cd),
	.w4(32'h39819430),
	.w5(32'hb9fe7bef),
	.w6(32'hbaa77120),
	.w7(32'h3b2445cd),
	.w8(32'h39a24db4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5da2a2),
	.w1(32'h3b1c0994),
	.w2(32'h3b935ddf),
	.w3(32'h3b99c18b),
	.w4(32'h3b962b7f),
	.w5(32'hbb0bf1ef),
	.w6(32'h3bc88e0a),
	.w7(32'h3b84fbb0),
	.w8(32'h3aff0c1f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81851f),
	.w1(32'h3ac09c91),
	.w2(32'hbaeb9dd0),
	.w3(32'h3b093d7c),
	.w4(32'hbac22879),
	.w5(32'hbb15d344),
	.w6(32'h3b354a12),
	.w7(32'hb9e2f402),
	.w8(32'hbaeb8b80),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11afba),
	.w1(32'hbb01db39),
	.w2(32'hbb89dd1e),
	.w3(32'h3b4b7c5d),
	.w4(32'hbb031577),
	.w5(32'h3b12abfd),
	.w6(32'h3aeb8dac),
	.w7(32'hb9c2e5a4),
	.w8(32'hbb07ff04),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d15868),
	.w1(32'hbbe2e1a0),
	.w2(32'hbaad655f),
	.w3(32'hbb69a7a3),
	.w4(32'hbb2be07a),
	.w5(32'h3c0e2a96),
	.w6(32'hbbe46405),
	.w7(32'hbb345a48),
	.w8(32'hbb8436fe),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedebb2),
	.w1(32'h3ba143df),
	.w2(32'h3b6bc34a),
	.w3(32'h3c37634d),
	.w4(32'h3c25fd25),
	.w5(32'h39e62ea7),
	.w6(32'hbbc0ee97),
	.w7(32'hb993b607),
	.w8(32'h3a18cf4d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab623ef),
	.w1(32'h3b036662),
	.w2(32'h3b297eb8),
	.w3(32'hb9654aef),
	.w4(32'h393dcccd),
	.w5(32'h3c0e05b9),
	.w6(32'h3ab8c7c7),
	.w7(32'h39660ad6),
	.w8(32'h3bba22ea),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ac87),
	.w1(32'h38e71f49),
	.w2(32'hbb84adb1),
	.w3(32'h3bf67fc1),
	.w4(32'h3abeb974),
	.w5(32'h3aefa8e2),
	.w6(32'hb9341abe),
	.w7(32'hbbdb2049),
	.w8(32'hbac5c250),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0dcf),
	.w1(32'h3a5cad50),
	.w2(32'h3acf3a1d),
	.w3(32'h3a1b6f7e),
	.w4(32'h3a9d17e1),
	.w5(32'hbb9d195a),
	.w6(32'hbb1c008c),
	.w7(32'h39e9853f),
	.w8(32'hbae06a47),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e3db8),
	.w1(32'h3a96dbe8),
	.w2(32'hba19e986),
	.w3(32'hbaadabcd),
	.w4(32'hb9e13b2f),
	.w5(32'hbb8d8e80),
	.w6(32'h3a5a201e),
	.w7(32'h3a944cb8),
	.w8(32'hba1b4647),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fe4e8),
	.w1(32'hba4319cd),
	.w2(32'hbb576ab1),
	.w3(32'hbb453ebc),
	.w4(32'hbb9fd7a7),
	.w5(32'hbac798c8),
	.w6(32'h3a4f2a80),
	.w7(32'hbb0f1b22),
	.w8(32'hbb0de26f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0f3ba),
	.w1(32'h3acbad01),
	.w2(32'hb989782a),
	.w3(32'hb9b16e51),
	.w4(32'h3b278a9d),
	.w5(32'h3b486bd8),
	.w6(32'hb9f1a899),
	.w7(32'h3866dfea),
	.w8(32'h3baa8762),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8900),
	.w1(32'h3be44f41),
	.w2(32'h3bbf418a),
	.w3(32'h39e4eee9),
	.w4(32'h3ae9a111),
	.w5(32'hbb4604b5),
	.w6(32'h3b44250e),
	.w7(32'h3a92e4c7),
	.w8(32'hbbbe96f3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21633c),
	.w1(32'hbb8f5d19),
	.w2(32'hbb5fa1f4),
	.w3(32'h3b0f06d4),
	.w4(32'hba8baaea),
	.w5(32'h3b71cb93),
	.w6(32'hbacead8e),
	.w7(32'hba4381d4),
	.w8(32'h3b61384b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2d499),
	.w1(32'h3a3e5e5f),
	.w2(32'h3abe7b21),
	.w3(32'h3aaef190),
	.w4(32'h3aacee43),
	.w5(32'hba30e504),
	.w6(32'h3aeafb8f),
	.w7(32'h3a449061),
	.w8(32'hbac7e3da),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39809a4e),
	.w1(32'h3b17f087),
	.w2(32'h3ac3134c),
	.w3(32'h399932a9),
	.w4(32'hb97a8b7f),
	.w5(32'h3ad2a8f2),
	.w6(32'h3a33d453),
	.w7(32'hba92eaa7),
	.w8(32'hbac217fd),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6514b6),
	.w1(32'hbac93cf7),
	.w2(32'hbba91197),
	.w3(32'h3ad69012),
	.w4(32'hbbbcf33f),
	.w5(32'hbb8d7e1d),
	.w6(32'h3ac8967b),
	.w7(32'hbb9bd8b4),
	.w8(32'hbb9a3a42),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af355f0),
	.w1(32'hb7c2361e),
	.w2(32'hbad754ed),
	.w3(32'hba18eb13),
	.w4(32'hbbaeaabf),
	.w5(32'hbb344adc),
	.w6(32'hbb42f3ca),
	.w7(32'hbbc50778),
	.w8(32'hbac8175a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf0b6f),
	.w1(32'hb99f6e87),
	.w2(32'hba557524),
	.w3(32'h3a52a292),
	.w4(32'hbabbad25),
	.w5(32'hbb65defd),
	.w6(32'h3c1f1a20),
	.w7(32'h3c16586b),
	.w8(32'h3afcd398),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8fb5c),
	.w1(32'h398fd424),
	.w2(32'hbc0659b7),
	.w3(32'hbb90114e),
	.w4(32'hbbf9c03e),
	.w5(32'hbc0b1665),
	.w6(32'h3b3ad50b),
	.w7(32'hbbf235e9),
	.w8(32'hbba8720b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382145dd),
	.w1(32'hbaa3a252),
	.w2(32'hba986ac5),
	.w3(32'hbb9ef28c),
	.w4(32'hbb9340f8),
	.w5(32'h3b76ed60),
	.w6(32'hb8f19183),
	.w7(32'h3a38cf5c),
	.w8(32'h3ba71ddf),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c379f),
	.w1(32'h3b3b9529),
	.w2(32'h3af5b2f0),
	.w3(32'h3ac56e4f),
	.w4(32'h3a38cf55),
	.w5(32'hbb709e28),
	.w6(32'h3b939cdf),
	.w7(32'h3b4cc624),
	.w8(32'hbaf191a2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc4cb0),
	.w1(32'hbbc629df),
	.w2(32'hbb82502b),
	.w3(32'h3b0603e5),
	.w4(32'hbc2fc8d2),
	.w5(32'hbc44f28a),
	.w6(32'h3b7c8711),
	.w7(32'hbbe46d44),
	.w8(32'hbc8cf54d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e81aa),
	.w1(32'h398f73b1),
	.w2(32'hbb0026bb),
	.w3(32'hbb1da784),
	.w4(32'hbaeda81c),
	.w5(32'h39c74c4d),
	.w6(32'hbaf4e918),
	.w7(32'hbb78f729),
	.w8(32'h39f8eba3),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26fc3a),
	.w1(32'h3b221f84),
	.w2(32'h3a8e0872),
	.w3(32'h3b863a33),
	.w4(32'hbb93223c),
	.w5(32'hba73d39a),
	.w6(32'h3ba71be4),
	.w7(32'hbab9eae9),
	.w8(32'hba7499a3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5b849),
	.w1(32'hb8b66dce),
	.w2(32'hbb4283fb),
	.w3(32'h3bda2643),
	.w4(32'h3b2b58c4),
	.w5(32'h3bd66c2f),
	.w6(32'h3c60262b),
	.w7(32'h3bef2bf3),
	.w8(32'h3b9cff8f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14455f),
	.w1(32'h3a69c2fd),
	.w2(32'hbbf58459),
	.w3(32'h3bc088ff),
	.w4(32'hb8faccae),
	.w5(32'h3b94378d),
	.w6(32'hb9adc4a3),
	.w7(32'hbb90a8c5),
	.w8(32'h3b70427b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befd8d4),
	.w1(32'h3b72fc43),
	.w2(32'h3a9804c4),
	.w3(32'h3b9e5dc3),
	.w4(32'hba53ed4e),
	.w5(32'hbb5d7387),
	.w6(32'h3ae5191e),
	.w7(32'hb9d31b0f),
	.w8(32'hbaafffa8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aee94),
	.w1(32'hba0e2464),
	.w2(32'hbab0e784),
	.w3(32'hbaabf3e0),
	.w4(32'hbae8be25),
	.w5(32'hb9912e0e),
	.w6(32'hba8dfd6d),
	.w7(32'hb9d854b8),
	.w8(32'hba751790),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c6a3a),
	.w1(32'h3a4a886e),
	.w2(32'h3b03cc80),
	.w3(32'hbaa08026),
	.w4(32'h3a8a30d2),
	.w5(32'hbaa5c05c),
	.w6(32'hbac5f508),
	.w7(32'hbb08d053),
	.w8(32'h3ae8b561),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca9706),
	.w1(32'hba8289c0),
	.w2(32'h3a15d6f8),
	.w3(32'hbabad458),
	.w4(32'hbb24e02b),
	.w5(32'h395b1f3f),
	.w6(32'h3bb05c45),
	.w7(32'h3b98e667),
	.w8(32'hba0b295e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20d301),
	.w1(32'h3b0dc668),
	.w2(32'h3b0888b6),
	.w3(32'h3a8fd6fb),
	.w4(32'h3998b249),
	.w5(32'h3afe6f22),
	.w6(32'h3b8635c7),
	.w7(32'h3a667632),
	.w8(32'h3aaa8a71),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ed6f7),
	.w1(32'hba6f2102),
	.w2(32'hbad97f11),
	.w3(32'h3895eadd),
	.w4(32'hbadf554f),
	.w5(32'hbb941f59),
	.w6(32'hbac14106),
	.w7(32'hbb3de3fe),
	.w8(32'hbbbc06d5),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1115a),
	.w1(32'h3a43a528),
	.w2(32'hbb30b4d0),
	.w3(32'h3ad2f63a),
	.w4(32'hbb4e2b28),
	.w5(32'hbb2c7a7a),
	.w6(32'hb9e72a39),
	.w7(32'hbb197eef),
	.w8(32'hbba03ab4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb882a6),
	.w1(32'hbba903d3),
	.w2(32'hbacd4f4f),
	.w3(32'hb7fb595b),
	.w4(32'hbb752230),
	.w5(32'h3b1a0831),
	.w6(32'hbb8d970d),
	.w7(32'hbac1cc99),
	.w8(32'h3aa2e406),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0df8cb),
	.w1(32'hba47c331),
	.w2(32'hb97101b9),
	.w3(32'h3ba6ec22),
	.w4(32'hbc09c449),
	.w5(32'hbbb85d32),
	.w6(32'h3b77842c),
	.w7(32'hbbc4fb06),
	.w8(32'hbc2a9d53),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75a74d),
	.w1(32'hbbbc469d),
	.w2(32'hbb840d3e),
	.w3(32'hbb742449),
	.w4(32'hbb283681),
	.w5(32'hb8d2a56a),
	.w6(32'hbb5562ac),
	.w7(32'hbbdfb659),
	.w8(32'h3aa9c3fb),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba882821),
	.w1(32'h3b19944e),
	.w2(32'h3aa4647f),
	.w3(32'h3ace5c65),
	.w4(32'h3b4497c4),
	.w5(32'h3ae9dcf9),
	.w6(32'h3bdd5160),
	.w7(32'h3bff7b2c),
	.w8(32'h3b57c9a6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d808b),
	.w1(32'h3bb28d0a),
	.w2(32'h3b4dbf57),
	.w3(32'h3b8b74d4),
	.w4(32'h3b924132),
	.w5(32'hba6258c3),
	.w6(32'h3bd39723),
	.w7(32'h3b631131),
	.w8(32'hbaf0bd75),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb450f1e),
	.w1(32'h3afac3f9),
	.w2(32'h3ac0ea29),
	.w3(32'h3a78af02),
	.w4(32'h3a863d75),
	.w5(32'h3aaa7b3a),
	.w6(32'hbacfe261),
	.w7(32'h3b9f63fe),
	.w8(32'h3a931bed),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3f8fa),
	.w1(32'h3aa11f8f),
	.w2(32'h3a879057),
	.w3(32'h39399d3d),
	.w4(32'hba623a35),
	.w5(32'hbb16a576),
	.w6(32'h3a9a3641),
	.w7(32'h3958e11e),
	.w8(32'hbb493bdb),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0615c),
	.w1(32'h3b14d306),
	.w2(32'h3a65ea04),
	.w3(32'h3aeec343),
	.w4(32'h3ad29d59),
	.w5(32'hbb4d55f9),
	.w6(32'h3b6a5823),
	.w7(32'h3af0f13e),
	.w8(32'hbb0056d1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb848d78),
	.w1(32'hbad4e952),
	.w2(32'hb9f93a05),
	.w3(32'hbb2084fb),
	.w4(32'hbb0fdfa4),
	.w5(32'h3b6b0701),
	.w6(32'hba560545),
	.w7(32'h3a6f3a01),
	.w8(32'h384396fc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fc9f8),
	.w1(32'h39561224),
	.w2(32'h3b19ec8e),
	.w3(32'h3b576cee),
	.w4(32'h3b01bda6),
	.w5(32'hbac6bb25),
	.w6(32'h3b8342ef),
	.w7(32'h3b5204e1),
	.w8(32'hbba8ca0b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c9b83),
	.w1(32'h3b0664b1),
	.w2(32'h3b855b5c),
	.w3(32'hbb73ebb8),
	.w4(32'h3ba58c94),
	.w5(32'hbb48668f),
	.w6(32'hbc3c2ab1),
	.w7(32'hbae57c66),
	.w8(32'h3a1bd80f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3268f4),
	.w1(32'h3b7d4697),
	.w2(32'h3b62b01d),
	.w3(32'h3a5d0f81),
	.w4(32'hbad52461),
	.w5(32'h3b9bbf90),
	.w6(32'h3b900f31),
	.w7(32'h3a63dcd6),
	.w8(32'hbb554625),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad3d06),
	.w1(32'h3b0bc0ed),
	.w2(32'hba8f93da),
	.w3(32'h3bb6c133),
	.w4(32'h3b0a2ef2),
	.w5(32'hba60b458),
	.w6(32'hba969c1f),
	.w7(32'hbb723236),
	.w8(32'h3b6abc4c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b249ba7),
	.w1(32'h3b26b703),
	.w2(32'hba6ed8b0),
	.w3(32'h3af8de04),
	.w4(32'h3bc71712),
	.w5(32'hbb06de59),
	.w6(32'h3a1493b6),
	.w7(32'h3980f717),
	.w8(32'hbb90a034),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d1419),
	.w1(32'hbb604cc6),
	.w2(32'hbb15e7a0),
	.w3(32'hbb804eae),
	.w4(32'hbb12502f),
	.w5(32'hbab74057),
	.w6(32'hbbf5c80f),
	.w7(32'hbb80897f),
	.w8(32'hba2f4c93),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39145239),
	.w1(32'hba9b3d59),
	.w2(32'hba24a171),
	.w3(32'hbb022bb1),
	.w4(32'hba2e4433),
	.w5(32'h394ead2c),
	.w6(32'hbb1083d2),
	.w7(32'hbade15e9),
	.w8(32'hba165197),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83e4d3),
	.w1(32'h3aafe5d7),
	.w2(32'h3a3f71bc),
	.w3(32'hb95b88b4),
	.w4(32'h3a8b1d76),
	.w5(32'h3b31f93e),
	.w6(32'h3b56631f),
	.w7(32'h3a4ca70d),
	.w8(32'h3b3c1829),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4c8db),
	.w1(32'h3a9c183c),
	.w2(32'h3990ca0a),
	.w3(32'hba723825),
	.w4(32'hb9df6bda),
	.w5(32'h3b1efbd3),
	.w6(32'hba5cb329),
	.w7(32'hbabd2ad3),
	.w8(32'hba1b0b32),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc1b56),
	.w1(32'h3b9ad30d),
	.w2(32'h3b724103),
	.w3(32'h3b4292e9),
	.w4(32'h3b64fc1d),
	.w5(32'h38bfdb5b),
	.w6(32'h3a8fddef),
	.w7(32'h3a65af24),
	.w8(32'hbaa74485),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad14aa),
	.w1(32'h3b89268f),
	.w2(32'h3c2dfa4f),
	.w3(32'hbadf8359),
	.w4(32'h3beb9f22),
	.w5(32'hba73e245),
	.w6(32'hbbd42fe6),
	.w7(32'h3ba29ceb),
	.w8(32'hb8fb5db2),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeeb0ad),
	.w1(32'h3aa7f77b),
	.w2(32'h3bb9a961),
	.w3(32'h3b8e3766),
	.w4(32'h3bab5d5d),
	.w5(32'h3b013d40),
	.w6(32'h3a0740a4),
	.w7(32'h3b74bef1),
	.w8(32'h3a3d10cc),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed6e7e),
	.w1(32'h3b55df82),
	.w2(32'h3b4c6d5c),
	.w3(32'hbb2f02bd),
	.w4(32'hbb80316f),
	.w5(32'hba86cda5),
	.w6(32'hb825525f),
	.w7(32'h3af7a029),
	.w8(32'hbae83276),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36be81d1),
	.w1(32'hb9acb033),
	.w2(32'h3b7f6a9c),
	.w3(32'h39ab6b3d),
	.w4(32'hb900c463),
	.w5(32'hba137364),
	.w6(32'h3acc4ff9),
	.w7(32'h3b7ce862),
	.w8(32'h3af25d51),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3514cc),
	.w1(32'h38ca8f9a),
	.w2(32'h398455b4),
	.w3(32'hb9720010),
	.w4(32'h3aa9221e),
	.w5(32'h3bdd29ad),
	.w6(32'hb921859a),
	.w7(32'h3a8397a5),
	.w8(32'h3a550c4e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf73ef2),
	.w1(32'h3b679020),
	.w2(32'h3c043639),
	.w3(32'h3c116baf),
	.w4(32'h3c675d74),
	.w5(32'hb9e666e3),
	.w6(32'hbb9d9002),
	.w7(32'h3c4e58c7),
	.w8(32'h3b71ed10),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb103af2),
	.w1(32'hba138a7c),
	.w2(32'hba21c479),
	.w3(32'hba6e0b2b),
	.w4(32'hb9a1d8fe),
	.w5(32'hbaf336f1),
	.w6(32'h3a0ea080),
	.w7(32'hba9f30d7),
	.w8(32'hbb169b43),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8878bb),
	.w1(32'hbb4a9888),
	.w2(32'hbb2f41d1),
	.w3(32'h3ac51bb2),
	.w4(32'h3a508d3c),
	.w5(32'hbb8d6556),
	.w6(32'hbb80a075),
	.w7(32'hba1c7ae2),
	.w8(32'hbb81a358),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule