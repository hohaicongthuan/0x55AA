module layer_8_featuremap_92(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afef8cf),
	.w1(32'hbd3bffdd),
	.w2(32'hbc58e785),
	.w3(32'hbcae381e),
	.w4(32'hbc496066),
	.w5(32'h3c97bf13),
	.w6(32'hbcc83590),
	.w7(32'h3b0b6745),
	.w8(32'h3cdcb4dc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76d1f6),
	.w1(32'hbbfddb8f),
	.w2(32'hbd1bb687),
	.w3(32'h3bcc8dcf),
	.w4(32'hbc2ddd68),
	.w5(32'hbc167970),
	.w6(32'hbab50017),
	.w7(32'hbbc9d70e),
	.w8(32'hbbc3e42b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd07a2f),
	.w1(32'h3c8e2605),
	.w2(32'h3c2ea872),
	.w3(32'hbd25ef43),
	.w4(32'hbba3608e),
	.w5(32'h3d1c0f65),
	.w6(32'hbc01671e),
	.w7(32'h3b8d1fb5),
	.w8(32'hbb84df20),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5685cc),
	.w1(32'h3cb5bc88),
	.w2(32'h3ce4c2ab),
	.w3(32'hbcc3b495),
	.w4(32'h3b3ff3ff),
	.w5(32'h3d24acf6),
	.w6(32'hbd2128b9),
	.w7(32'hbd234c4a),
	.w8(32'hbc6eac3c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05449f),
	.w1(32'h3bccbb81),
	.w2(32'hbc03eac8),
	.w3(32'hbb3729a9),
	.w4(32'hbc61f802),
	.w5(32'h3aadd399),
	.w6(32'hbb2bf8aa),
	.w7(32'hbd461fae),
	.w8(32'h3c32f570),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d0fd8),
	.w1(32'hbd1ef9fb),
	.w2(32'h3d06f012),
	.w3(32'hb9d386b1),
	.w4(32'hbba39644),
	.w5(32'h3c2000f3),
	.w6(32'hbbdefea4),
	.w7(32'hb9cc1a66),
	.w8(32'hb8cc5ba6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd37e1c5),
	.w1(32'hbc4fd57a),
	.w2(32'h3c754d0b),
	.w3(32'h3d458e96),
	.w4(32'h3c2c2c47),
	.w5(32'h3c151ae8),
	.w6(32'hbcc866a4),
	.w7(32'h3ca23c0c),
	.w8(32'hbb9c881e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b744d74),
	.w1(32'h3c8ecacb),
	.w2(32'h3ce09b3f),
	.w3(32'hbc291d16),
	.w4(32'hbd6f9f10),
	.w5(32'hbd01c8a3),
	.w6(32'hbd1ea798),
	.w7(32'hbb8f3bef),
	.w8(32'hbcf0a6f8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31ead2),
	.w1(32'h3cf6ca94),
	.w2(32'h3ba11eb8),
	.w3(32'hbc5f2d27),
	.w4(32'hbc260f23),
	.w5(32'hbadb76ca),
	.w6(32'h3bd4a703),
	.w7(32'hbd43c7c7),
	.w8(32'hbc4537e8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c72fd),
	.w1(32'hbb982cac),
	.w2(32'hbbf85356),
	.w3(32'h3c50db11),
	.w4(32'h3bb0c4c1),
	.w5(32'hbd986f61),
	.w6(32'hbbf88fc5),
	.w7(32'hbca76a0a),
	.w8(32'h3b96fd27),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3774b1),
	.w1(32'hbcae6007),
	.w2(32'hbd88344d),
	.w3(32'hbc42792d),
	.w4(32'hba80c1f6),
	.w5(32'h3b1097aa),
	.w6(32'h3cdc42a9),
	.w7(32'hbc01cdb3),
	.w8(32'hbc9e87d3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb544c4),
	.w1(32'hbbf9513a),
	.w2(32'h3c80f0e7),
	.w3(32'hbc73f247),
	.w4(32'hbcbd6eda),
	.w5(32'hbd33f295),
	.w6(32'hbbb0de2a),
	.w7(32'hbc762e19),
	.w8(32'h3b92b2b2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b339b1a),
	.w1(32'h3d2595e7),
	.w2(32'hbd4b715f),
	.w3(32'hbc1e2664),
	.w4(32'h3ba2effc),
	.w5(32'hbc312893),
	.w6(32'hbc1f3b12),
	.w7(32'h3cc03cfd),
	.w8(32'h3bcc2c29),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97ab76),
	.w1(32'h3a000678),
	.w2(32'h3c03e417),
	.w3(32'h3b9c868e),
	.w4(32'h3c042fb1),
	.w5(32'hbd130eea),
	.w6(32'hbd269232),
	.w7(32'hbb4b4c64),
	.w8(32'hbbc68205),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4149d8),
	.w1(32'hbd36cd79),
	.w2(32'h3c5fc153),
	.w3(32'h3b38dd83),
	.w4(32'hbc4fcce6),
	.w5(32'h3b3add36),
	.w6(32'h3bf27585),
	.w7(32'h3c25351b),
	.w8(32'h3b6cba0f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fc1aa),
	.w1(32'h3b092930),
	.w2(32'hbbdec59a),
	.w3(32'h3ac847f6),
	.w4(32'h3bd9ee8f),
	.w5(32'hbb05f0d3),
	.w6(32'h3b8c6c48),
	.w7(32'h3bb5f143),
	.w8(32'h3c83ae2a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa988bf),
	.w1(32'h3b09a86a),
	.w2(32'hbadda4ad),
	.w3(32'hbc2be0a9),
	.w4(32'h3b9111a2),
	.w5(32'h3c6b0552),
	.w6(32'hbc972f18),
	.w7(32'h3c824026),
	.w8(32'h3d0a6088),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f0dd8),
	.w1(32'hbbbb42ea),
	.w2(32'hbcb15ba7),
	.w3(32'hbbafc740),
	.w4(32'h3c1dfd65),
	.w5(32'h3afaa510),
	.w6(32'h3c3300f8),
	.w7(32'hbc525f22),
	.w8(32'h3c239abc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391da2be),
	.w1(32'hbc44da0a),
	.w2(32'h3b96f60c),
	.w3(32'hbb57e1bc),
	.w4(32'hbc6080fa),
	.w5(32'hbc702431),
	.w6(32'h3c7b2223),
	.w7(32'h3d520878),
	.w8(32'hbcade259),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed3d52),
	.w1(32'hbc483330),
	.w2(32'hbbd0ef13),
	.w3(32'hbc39481d),
	.w4(32'hbbebacb8),
	.w5(32'hb8553776),
	.w6(32'hbbb8a126),
	.w7(32'h3bfea53a),
	.w8(32'h3c40a37b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c6133),
	.w1(32'hbb2a4ce9),
	.w2(32'hbb990373),
	.w3(32'h3cb46f2c),
	.w4(32'hbce5cf34),
	.w5(32'hbb484813),
	.w6(32'h3b956d8f),
	.w7(32'h3b81b147),
	.w8(32'hbcf91e0e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8209d),
	.w1(32'h3bdb21e4),
	.w2(32'hbb81aa0a),
	.w3(32'h3b521048),
	.w4(32'h3b4c5cd0),
	.w5(32'h3bdf8193),
	.w6(32'h3b8c38e0),
	.w7(32'h3cda085d),
	.w8(32'h3db51143),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59e445),
	.w1(32'h3caebb2a),
	.w2(32'h3b242870),
	.w3(32'hbc8faa86),
	.w4(32'hbb43240e),
	.w5(32'hbc5e5cc2),
	.w6(32'hbbb15ca6),
	.w7(32'hbc01c586),
	.w8(32'hbc97d8a4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f7d65),
	.w1(32'h3d5f3b5d),
	.w2(32'hbc80bf22),
	.w3(32'hbde2c069),
	.w4(32'h3c77b70e),
	.w5(32'h3d354938),
	.w6(32'hbc385b39),
	.w7(32'h3c512a64),
	.w8(32'hbd6dfdd5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ad794),
	.w1(32'hbc373769),
	.w2(32'h3d06cf70),
	.w3(32'hbb8f6ee7),
	.w4(32'hbc51fc93),
	.w5(32'hbbd127c5),
	.w6(32'h3d1ad5bc),
	.w7(32'hbcaa3cf9),
	.w8(32'hbc1d7972),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb700848a),
	.w1(32'h3c7f4ece),
	.w2(32'h3c92a935),
	.w3(32'h3cc128fe),
	.w4(32'hbc4596b1),
	.w5(32'hbc9d5bac),
	.w6(32'h3969709c),
	.w7(32'h3c8b0aec),
	.w8(32'h3cfb100a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3b81),
	.w1(32'h3c472510),
	.w2(32'h3b04c74a),
	.w3(32'h3c412d60),
	.w4(32'hbc727084),
	.w5(32'h3c064506),
	.w6(32'h3b94047d),
	.w7(32'h3bd12d5f),
	.w8(32'hbc97a45f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe72020),
	.w1(32'hbc3a3f38),
	.w2(32'hbc8d6534),
	.w3(32'hbc0891ca),
	.w4(32'hbc807b6d),
	.w5(32'hbc92b759),
	.w6(32'h3c6db868),
	.w7(32'h3a30639c),
	.w8(32'h3bc3babc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be95f80),
	.w1(32'hbc802db7),
	.w2(32'hbc8db9bb),
	.w3(32'hb6dc45e5),
	.w4(32'h3be082e0),
	.w5(32'hbbf49dcf),
	.w6(32'hbc7520b1),
	.w7(32'hbc29ae3c),
	.w8(32'hbc29a517),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb959745),
	.w1(32'h3bc07345),
	.w2(32'hbc138c84),
	.w3(32'h3cad8966),
	.w4(32'hbcbf5d81),
	.w5(32'hbc0bbecd),
	.w6(32'hbcba4b10),
	.w7(32'h3c87d7ee),
	.w8(32'hbc92e520),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c212ae6),
	.w1(32'hbbbf5a2f),
	.w2(32'hbb6d84a9),
	.w3(32'hbc4c1e25),
	.w4(32'hbd17789d),
	.w5(32'h3bcfccd2),
	.w6(32'h3d042802),
	.w7(32'hbc5c18ef),
	.w8(32'hbad63b32),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b01f),
	.w1(32'hbb374044),
	.w2(32'h3b657979),
	.w3(32'hbc3834ba),
	.w4(32'hbc4f025e),
	.w5(32'h3ce0a686),
	.w6(32'hbc436504),
	.w7(32'hbc8eb4fe),
	.w8(32'hbca51385),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7a888),
	.w1(32'hbc58a8ca),
	.w2(32'hbb3005b8),
	.w3(32'h3bb75142),
	.w4(32'hbbf6c296),
	.w5(32'hbc1e1275),
	.w6(32'h3ceaef65),
	.w7(32'hbc0a1904),
	.w8(32'hbcbc872f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0aab0b),
	.w1(32'hbbb67b5c),
	.w2(32'hbd01c339),
	.w3(32'hbc2a2784),
	.w4(32'hbc79b887),
	.w5(32'h3bdec56f),
	.w6(32'hbb7a72c8),
	.w7(32'hbcbb7386),
	.w8(32'h3c0d77b9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dd4f5),
	.w1(32'hbc825827),
	.w2(32'hbc801e84),
	.w3(32'hbc498535),
	.w4(32'hbc6661c0),
	.w5(32'h3c219722),
	.w6(32'h3d15fd9c),
	.w7(32'h3cb948f0),
	.w8(32'h3cac5e0e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc122a6),
	.w1(32'h3bc7771d),
	.w2(32'hbc189f37),
	.w3(32'h3c70ccaa),
	.w4(32'hbc115f5a),
	.w5(32'hba4a5600),
	.w6(32'hbc94cd2a),
	.w7(32'h3c853775),
	.w8(32'hbcaa27cb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6ea85),
	.w1(32'h3b8a09ad),
	.w2(32'h3c3e2de3),
	.w3(32'h3bd4d68e),
	.w4(32'h3bdd4dd5),
	.w5(32'h3c164bce),
	.w6(32'hbb9bf3bd),
	.w7(32'hbcabe9dd),
	.w8(32'hbb0f5f97),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2e260),
	.w1(32'h3ccb7837),
	.w2(32'hbc411c0f),
	.w3(32'hbb437f4c),
	.w4(32'h3b24aa07),
	.w5(32'hbc8af528),
	.w6(32'hbba3496b),
	.w7(32'h3c3d71fe),
	.w8(32'hbbda7dee),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cba20),
	.w1(32'h3c5a8786),
	.w2(32'h3d45c84a),
	.w3(32'hbc97cfb4),
	.w4(32'hbc207ed4),
	.w5(32'hbc29d839),
	.w6(32'hbaa3593f),
	.w7(32'hbc212b07),
	.w8(32'hbc2da908),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2ddf),
	.w1(32'h3be9bfdb),
	.w2(32'hbbb06963),
	.w3(32'hbb8f5b29),
	.w4(32'hbbc34b88),
	.w5(32'hbb5a2692),
	.w6(32'hbc374043),
	.w7(32'h3ca40087),
	.w8(32'h3b15bb1a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb479c5c),
	.w1(32'hbcb5861a),
	.w2(32'hbc8a118a),
	.w3(32'h3b601949),
	.w4(32'hbb8919be),
	.w5(32'h3bfecc52),
	.w6(32'hbbf44296),
	.w7(32'hbacec66d),
	.w8(32'h3b5a7f19),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b972695),
	.w1(32'hbb9f6724),
	.w2(32'h3c892097),
	.w3(32'hbc36cc1f),
	.w4(32'h3cb5f668),
	.w5(32'hb9caa2d2),
	.w6(32'hbc05820c),
	.w7(32'hbb4452a6),
	.w8(32'hbb9f1228),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca7790),
	.w1(32'hb9729cd4),
	.w2(32'h3b785fcf),
	.w3(32'h3c77f8f8),
	.w4(32'h3d21e43d),
	.w5(32'h3bb7dda6),
	.w6(32'h3d45e20d),
	.w7(32'hbd1ea5d6),
	.w8(32'hbbb1daa4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5c9c0),
	.w1(32'hbcf4d857),
	.w2(32'h3ace3eec),
	.w3(32'h3d91ed4f),
	.w4(32'h3c3ec35c),
	.w5(32'h3c18671b),
	.w6(32'hbb09babf),
	.w7(32'hbd4b9289),
	.w8(32'hbc9c85c8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9ac7e),
	.w1(32'h3d10b8ae),
	.w2(32'hbe34ce11),
	.w3(32'hbd50a628),
	.w4(32'hb834ee80),
	.w5(32'hbca1c53f),
	.w6(32'hbbb957d0),
	.w7(32'h3d76f1b1),
	.w8(32'h3ccd0660),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b7c8d),
	.w1(32'h3ca80aeb),
	.w2(32'hbbf80834),
	.w3(32'h3c21c28b),
	.w4(32'h3ca67cf3),
	.w5(32'hbcd9b48a),
	.w6(32'hbcb4c68a),
	.w7(32'h3c1a6d2e),
	.w8(32'hbd140ee0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cde2f93),
	.w1(32'h3cc217b2),
	.w2(32'h3c1ac391),
	.w3(32'hbb8e075d),
	.w4(32'h3d0cf87d),
	.w5(32'h3ca28d18),
	.w6(32'hbcdac340),
	.w7(32'hbcfde3be),
	.w8(32'h3c2f0715),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae0d9b),
	.w1(32'h3aea424b),
	.w2(32'hbb43b2cd),
	.w3(32'hbd5e28fe),
	.w4(32'h3c6aa171),
	.w5(32'hbc171b95),
	.w6(32'hbd8df07b),
	.w7(32'hbb0d66af),
	.w8(32'h3c553882),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bcea5),
	.w1(32'h3c9f9c03),
	.w2(32'hbd13548a),
	.w3(32'hbbb7b55f),
	.w4(32'hba10648f),
	.w5(32'h3d7cd063),
	.w6(32'h394d13ac),
	.w7(32'hbc6ee39b),
	.w8(32'h3a8a54b0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd8738),
	.w1(32'hbb2157c5),
	.w2(32'hbb142539),
	.w3(32'hb9f2261a),
	.w4(32'h3cfd8585),
	.w5(32'hbce0fa45),
	.w6(32'h3c9479b4),
	.w7(32'h3d166f6d),
	.w8(32'hbd284e1d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5f36ae),
	.w1(32'hbc76a39e),
	.w2(32'h3c54a59b),
	.w3(32'hbd3cfb4b),
	.w4(32'hbd9b27d6),
	.w5(32'h3c7707cd),
	.w6(32'h3d13ea5d),
	.w7(32'hbbe05fca),
	.w8(32'h3a6d4961),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae240de),
	.w1(32'hbbd2c311),
	.w2(32'hbc4e443d),
	.w3(32'hbc195ec2),
	.w4(32'hbc2aada4),
	.w5(32'hbc68987b),
	.w6(32'hbcc1115f),
	.w7(32'hbc2c81af),
	.w8(32'h3c96584d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72c03e),
	.w1(32'hbc8f2e7f),
	.w2(32'hba0ae8d8),
	.w3(32'h3b7c0bd0),
	.w4(32'hbd1ea815),
	.w5(32'hbc08ee50),
	.w6(32'hbd0b0cca),
	.w7(32'h3c4b76f8),
	.w8(32'h3c266234),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80370e),
	.w1(32'hbd330852),
	.w2(32'h3ca6b89e),
	.w3(32'h3cb03614),
	.w4(32'hbba1ff94),
	.w5(32'h3cc31ad5),
	.w6(32'h3b95791f),
	.w7(32'h3b874f7a),
	.w8(32'h3bb96676),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f85e9),
	.w1(32'h3cd6d1d2),
	.w2(32'h38c422b1),
	.w3(32'hbb3e6b11),
	.w4(32'hbd2b734c),
	.w5(32'h3c10626a),
	.w6(32'hbd29f907),
	.w7(32'h3d2e6b39),
	.w8(32'hbc74df7d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fd1e2),
	.w1(32'h3b8600dc),
	.w2(32'hbb2c17e7),
	.w3(32'h3c2c1aba),
	.w4(32'h3baa5fa3),
	.w5(32'h3b88e8c9),
	.w6(32'h3c3bedbe),
	.w7(32'h3c91cef2),
	.w8(32'hbc0e58a0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5628e),
	.w1(32'hbd186024),
	.w2(32'hbdb71c22),
	.w3(32'hbc45635f),
	.w4(32'hbd56485d),
	.w5(32'h3b9e703c),
	.w6(32'hbb900c90),
	.w7(32'hbd0bcdb1),
	.w8(32'h3afcfb8c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c0a2a),
	.w1(32'hbd8fc6c9),
	.w2(32'hbb6e51a0),
	.w3(32'h3b8ad581),
	.w4(32'hbb78a533),
	.w5(32'hbc0b467e),
	.w6(32'h3cc09ab5),
	.w7(32'hbc9ffeca),
	.w8(32'hbbfb9e03),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84bbd8),
	.w1(32'h3d1952a5),
	.w2(32'hbcb5654e),
	.w3(32'hbc5156b5),
	.w4(32'hb9bd2e3e),
	.w5(32'hbd05d58e),
	.w6(32'hbc42beab),
	.w7(32'h3d1ae8e0),
	.w8(32'h3c9cb32a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c960e5a),
	.w1(32'hbcf6b0cc),
	.w2(32'h3c4cd414),
	.w3(32'hbbf915a5),
	.w4(32'h3a68c575),
	.w5(32'hbcaa304a),
	.w6(32'hbbd72fec),
	.w7(32'hbc473c0a),
	.w8(32'hbc88f552),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2a1997),
	.w1(32'hbc329348),
	.w2(32'hbaa0162f),
	.w3(32'h3ba100da),
	.w4(32'h3d627a4e),
	.w5(32'h3c906548),
	.w6(32'hbc437356),
	.w7(32'h3bc3ec23),
	.w8(32'hbca32471),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc21f05),
	.w1(32'hbcb192a9),
	.w2(32'hbc2d337a),
	.w3(32'hbc771988),
	.w4(32'hb9a889de),
	.w5(32'hbc214e77),
	.w6(32'hbc8bce7d),
	.w7(32'hbcf81a76),
	.w8(32'h3bbec391),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09b6a2),
	.w1(32'hbc8e8c75),
	.w2(32'hbcc81d1c),
	.w3(32'h3c252811),
	.w4(32'hbb080480),
	.w5(32'hbb85fe31),
	.w6(32'hbcacba01),
	.w7(32'h3c1bf5f2),
	.w8(32'hbc7057b2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb23bb8),
	.w1(32'h3bb0c7b1),
	.w2(32'hbd08efa6),
	.w3(32'h3bcf938b),
	.w4(32'hbca2766b),
	.w5(32'hba6f0c4f),
	.w6(32'h3c822dd2),
	.w7(32'hbc97a9b8),
	.w8(32'hbc491d7b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28dac6),
	.w1(32'h3b4450ac),
	.w2(32'h3a9fd723),
	.w3(32'hbbc80ce8),
	.w4(32'hbd12207c),
	.w5(32'hbc7b37fc),
	.w6(32'h3d5a4748),
	.w7(32'hbc62b5af),
	.w8(32'h3b17f15a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaeb0dd),
	.w1(32'h3bfb4551),
	.w2(32'h3cb5cc43),
	.w3(32'h39417cb1),
	.w4(32'h3c953f3f),
	.w5(32'h3d5f760f),
	.w6(32'hbca9f8b4),
	.w7(32'hbc8537f4),
	.w8(32'hbc475794),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d037d96),
	.w1(32'hbb3c9f9a),
	.w2(32'h3cd2e617),
	.w3(32'hba8460a1),
	.w4(32'hbcd40c82),
	.w5(32'h39a22959),
	.w6(32'h3b330185),
	.w7(32'hbc4b021f),
	.w8(32'hbcc8f319),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6eaa8),
	.w1(32'h3d01141f),
	.w2(32'h3ca1c9cb),
	.w3(32'hbce22600),
	.w4(32'hbacb4f68),
	.w5(32'h3c8090a5),
	.w6(32'h3c879183),
	.w7(32'h3cc6daae),
	.w8(32'hbc07d14b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05a10c),
	.w1(32'h3bd02a59),
	.w2(32'h3bad20f1),
	.w3(32'hbba874a2),
	.w4(32'h3b441a0c),
	.w5(32'h3c6b79be),
	.w6(32'hbc609c43),
	.w7(32'hbccda7d2),
	.w8(32'hbb86a5c1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b09cc),
	.w1(32'hbbf6259c),
	.w2(32'hbbcc9005),
	.w3(32'hbcec6297),
	.w4(32'hbc311e65),
	.w5(32'hbc5d0630),
	.w6(32'hbc18dbb2),
	.w7(32'h3b140b19),
	.w8(32'h3c0258b3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d11b43),
	.w1(32'hbcb1dd08),
	.w2(32'hbc688734),
	.w3(32'hbd47d9f5),
	.w4(32'hbbc43a6d),
	.w5(32'h3cbb5367),
	.w6(32'hbb9fc191),
	.w7(32'h3bf379d9),
	.w8(32'h3c298334),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc301a6d),
	.w1(32'h3ca4bc8b),
	.w2(32'hbadea0b8),
	.w3(32'h3b8e3974),
	.w4(32'h3c0284b7),
	.w5(32'hba6a2a45),
	.w6(32'hbc48d59d),
	.w7(32'hbc601f5f),
	.w8(32'hbcae0757),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd89220),
	.w1(32'h3b6ed754),
	.w2(32'hbb542701),
	.w3(32'h3c3fc407),
	.w4(32'h3c40e9f6),
	.w5(32'hbb458797),
	.w6(32'hbb776702),
	.w7(32'hbc821013),
	.w8(32'hbb9d6f08),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0161b2),
	.w1(32'hb72e0a20),
	.w2(32'h3c231d6f),
	.w3(32'hbb157f38),
	.w4(32'hbc2c09b7),
	.w5(32'hbce597cd),
	.w6(32'h3b61f11a),
	.w7(32'h3b7a9645),
	.w8(32'h3ca0d81b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0dcc2),
	.w1(32'hbcae35ba),
	.w2(32'h3b3c496c),
	.w3(32'h3c7b2e20),
	.w4(32'h3bfeae4b),
	.w5(32'hbb0d6486),
	.w6(32'hbc43d5f1),
	.w7(32'hbbc00c56),
	.w8(32'hbb04308f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e6413),
	.w1(32'hbb318fdb),
	.w2(32'h3aa78ca9),
	.w3(32'h3ba10bd9),
	.w4(32'h3d0a54ef),
	.w5(32'h3d58f2fd),
	.w6(32'h3b993cf0),
	.w7(32'hbb662504),
	.w8(32'h3c8b0436),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bc494),
	.w1(32'h3c940370),
	.w2(32'h3b68b8b5),
	.w3(32'h3c24d48e),
	.w4(32'h3ba83e98),
	.w5(32'h3c98bb62),
	.w6(32'hbbce72ba),
	.w7(32'hbb47e99a),
	.w8(32'h3c719360),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee19ba),
	.w1(32'h3c5d87cc),
	.w2(32'h3ba3cf79),
	.w3(32'h3ba52497),
	.w4(32'hbb6c26bd),
	.w5(32'hbbcc3a2f),
	.w6(32'h3aab6f51),
	.w7(32'hbb8316b6),
	.w8(32'hbb803ad4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d6301),
	.w1(32'hbc2df03c),
	.w2(32'hbd5c1451),
	.w3(32'h3bc75a2d),
	.w4(32'h3c422e9d),
	.w5(32'h3a086064),
	.w6(32'h3c466ab1),
	.w7(32'hbbbdff3b),
	.w8(32'h3b63c475),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc585a5d),
	.w1(32'h3a98d76d),
	.w2(32'hbb000809),
	.w3(32'hbade2102),
	.w4(32'hb9076402),
	.w5(32'hbb885c10),
	.w6(32'h3bc69ac8),
	.w7(32'hbb593fd6),
	.w8(32'h3b20dea8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7804a3),
	.w1(32'hbc84aea6),
	.w2(32'h3b8dca45),
	.w3(32'h3a8ae0c6),
	.w4(32'h3d25a6a2),
	.w5(32'hbd48bd61),
	.w6(32'h3d34544d),
	.w7(32'h3cdaf6ca),
	.w8(32'hbad00794),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb86c12),
	.w1(32'hbb909eac),
	.w2(32'hbb234761),
	.w3(32'h3d8ef260),
	.w4(32'hbc6c23d3),
	.w5(32'hbad1cb68),
	.w6(32'hbc0bf087),
	.w7(32'h3c8a3367),
	.w8(32'hbc04f439),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86c19e),
	.w1(32'hbb7444e3),
	.w2(32'h3c26bd08),
	.w3(32'h3ca71bb1),
	.w4(32'h383e8674),
	.w5(32'h3c2838b9),
	.w6(32'h3b894d81),
	.w7(32'h3bb5a529),
	.w8(32'h3b798923),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc4654),
	.w1(32'hbb74819b),
	.w2(32'hbf490b9e),
	.w3(32'hbb2572db),
	.w4(32'hbc821bdb),
	.w5(32'hbf6d57e5),
	.w6(32'h3ac41113),
	.w7(32'hbe999cce),
	.w8(32'hbdaee5fd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbefd9a88),
	.w1(32'hbf0156df),
	.w2(32'hbf2af6eb),
	.w3(32'hbf1e9258),
	.w4(32'hbf0886be),
	.w5(32'hbe24af7b),
	.w6(32'hbf2d790a),
	.w7(32'h4002ec61),
	.w8(32'hbecbfef7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf9c0f14),
	.w1(32'hbee81f28),
	.w2(32'hbf1fd238),
	.w3(32'hbecaab95),
	.w4(32'h3f1a6931),
	.w5(32'hbef3c47d),
	.w6(32'hbf3a5f3f),
	.w7(32'hbdb7787e),
	.w8(32'hbf122797),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf4bc0c3),
	.w1(32'hbf6bd0b4),
	.w2(32'hbea4cb0e),
	.w3(32'hbf58a331),
	.w4(32'hbf7ef799),
	.w5(32'hbeeaf5a3),
	.w6(32'hbeb95b4a),
	.w7(32'hbf6bf631),
	.w8(32'hbf38eae3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf06767d),
	.w1(32'hbefb4c1d),
	.w2(32'hbf3f23d5),
	.w3(32'hbec0a993),
	.w4(32'hbf989f30),
	.w5(32'hbc8e31f5),
	.w6(32'hbcd48c70),
	.w7(32'hbf07b078),
	.w8(32'hbf08c15f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeb3352d),
	.w1(32'hbf69a298),
	.w2(32'hbf2fb052),
	.w3(32'hbeb31071),
	.w4(32'hbf0af074),
	.w5(32'hbee15517),
	.w6(32'hbfa23505),
	.w7(32'hbecf2117),
	.w8(32'hbf2792ba),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf83af2d),
	.w1(32'hbf13ec40),
	.w2(32'hbf3cc427),
	.w3(32'hbf46aadc),
	.w4(32'hbe044755),
	.w5(32'hbf1549b5),
	.w6(32'hbf23e590),
	.w7(32'hbee0b1dd),
	.w8(32'hbf3b5cd7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf272dbf),
	.w1(32'hbf6a3ea9),
	.w2(32'hbeea532d),
	.w3(32'hbf4d9cf2),
	.w4(32'h3ebd9a16),
	.w5(32'hbf000dc6),
	.w6(32'hbeb9e100),
	.w7(32'hbc1e3b47),
	.w8(32'hbfb4e900),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeffbd52),
	.w1(32'hbf550e19),
	.w2(32'hbf063c1d),
	.w3(32'hbf855cbc),
	.w4(32'hbf1ecf21),
	.w5(32'hbf17ee47),
	.w6(32'hbf5a83f1),
	.w7(32'hbf64b149),
	.w8(32'hbf316f80),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf4dc859),
	.w1(32'hbf067eda),
	.w2(32'hbf0c1e8d),
	.w3(32'hbf05f073),
	.w4(32'hbf4aedca),
	.w5(32'hbf7775ee),
	.w6(32'hbf251055),
	.w7(32'hbf29cbe0),
	.w8(32'hbf670fb9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbde37768),
	.w1(32'h3d0c691e),
	.w2(32'hbf0dd977),
	.w3(32'hbeaeb2fd),
	.w4(32'hbe39e80a),
	.w5(32'hbf16f0e6),
	.w6(32'h3c3da993),
	.w7(32'hbf44a589),
	.w8(32'hbef4ca81),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec2865c),
	.w1(32'h3c215255),
	.w2(32'hbeb0a761),
	.w3(32'hbeda08bf),
	.w4(32'hbf27b706),
	.w5(32'hbe92deca),
	.w6(32'hbe336afd),
	.w7(32'hbf366323),
	.w8(32'hbc161fdc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf5f3b44),
	.w1(32'hbf49260a),
	.w2(32'hbf8b80ec),
	.w3(32'hbf88704a),
	.w4(32'hbeddcd2d),
	.w5(32'hbdf8004d),
	.w6(32'hbf37e480),
	.w7(32'hbf82c319),
	.w8(32'hbf607d8b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf45360d),
	.w1(32'hbf14e08c),
	.w2(32'hbed074a6),
	.w3(32'h3e238718),
	.w4(32'hbf37faf1),
	.w5(32'hbf96417c),
	.w6(32'hbf9d4b7c),
	.w7(32'hbefae887),
	.w8(32'hbf18b7d1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbefa7c3d),
	.w1(32'hbf06269a),
	.w2(32'hbf47fecd),
	.w3(32'hbf780c39),
	.w4(32'hbf90cdc5),
	.w5(32'h3751463a),
	.w6(32'hbccf4612),
	.w7(32'hbf0ff08b),
	.w8(32'h3f240b15),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fe3b90f),
	.w1(32'h3fac24fa),
	.w2(32'h3805b7be),
	.w3(32'h36ebf425),
	.w4(32'h38ac4861),
	.w5(32'h3f78da31),
	.w6(32'h3fbb7194),
	.w7(32'h3fb48ef2),
	.w8(32'h38331af5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fc506b1),
	.w1(32'h3f82e0f0),
	.w2(32'h3f74308b),
	.w3(32'h3f9794d2),
	.w4(32'h3fd49839),
	.w5(32'h3fcb3a44),
	.w6(32'h3f64832d),
	.w7(32'h3619cdc6),
	.w8(32'h3fd4421f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fd65526),
	.w1(32'h3fcf22d6),
	.w2(32'h3f673027),
	.w3(32'hb7f31bb2),
	.w4(32'h3fc84f74),
	.w5(32'h3fd12776),
	.w6(32'h3fb2a2d8),
	.w7(32'h3fbf5a65),
	.w8(32'h3fbb099f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fbc9ca0),
	.w1(32'h3f1119a6),
	.w2(32'h3f5ad7f8),
	.w3(32'hb7ca4658),
	.w4(32'h3f330a36),
	.w5(32'h3f8523b7),
	.w6(32'h3e9ed84e),
	.w7(32'h3f81f079),
	.w8(32'h3f84ca1e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ee66335),
	.w1(32'h3e8114aa),
	.w2(32'h3f1d3a7f),
	.w3(32'h37d8e73e),
	.w4(32'h3f96844e),
	.w5(32'h3f8909a9),
	.w6(32'h3f550e5c),
	.w7(32'h3f47a742),
	.w8(32'h3f87b18c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc0b58),
	.w1(32'h3fdf067f),
	.w2(32'h3ef0b202),
	.w3(32'h3e991592),
	.w4(32'h3f9c31f5),
	.w5(32'h39311c38),
	.w6(32'h3fd19179),
	.w7(32'h39553046),
	.w8(32'h3fd2005f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fcd3650),
	.w1(32'h3f48c71f),
	.w2(32'h3f3262df),
	.w3(32'h3faf3eb7),
	.w4(32'h38f3db0f),
	.w5(32'h3e542305),
	.w6(32'h3fd8962b),
	.w7(32'h3fcd58a7),
	.w8(32'h3e8cc06a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e9629d2),
	.w1(32'h3fe13378),
	.w2(32'h3fd5de26),
	.w3(32'hba63ff89),
	.w4(32'h3f6ae1e2),
	.w5(32'hba99408b),
	.w6(32'hba4d6215),
	.w7(32'h3fdab7fd),
	.w8(32'h3f990703),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fa790fc),
	.w1(32'h3fb65781),
	.w2(32'h3f49acbf),
	.w3(32'h3f4c1931),
	.w4(32'h3f3513ce),
	.w5(32'h3fa61424),
	.w6(32'h3f5199e9),
	.w7(32'h3f1e665a),
	.w8(32'h3fb7d14d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fceb01e),
	.w1(32'h3faa140a),
	.w2(32'hb7ad7261),
	.w3(32'h3fd470f7),
	.w4(32'h3fa41fe3),
	.w5(32'h3f2f3006),
	.w6(32'h3fa1524a),
	.w7(32'h3ee577ab),
	.w8(32'h3fd20b02),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f851322),
	.w1(32'h3904272e),
	.w2(32'h3fe50b7e),
	.w3(32'h3d4520b7),
	.w4(32'h3fbd5158),
	.w5(32'h3fcae436),
	.w6(32'h3d7ce7fd),
	.w7(32'h3ed0c60c),
	.w8(32'h3f6a6276),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fc33312),
	.w1(32'h3fc6ff8b),
	.w2(32'hb796ca91),
	.w3(32'h3fa458d6),
	.w4(32'h3fd654da),
	.w5(32'h3f611436),
	.w6(32'h3f70e24e),
	.w7(32'h3fcbc0b6),
	.w8(32'h3f7f4e02),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4ffe87),
	.w1(32'h389417e0),
	.w2(32'h3f282c99),
	.w3(32'h38586949),
	.w4(32'h3f3592a3),
	.w5(32'hba17d138),
	.w6(32'h3f9bc487),
	.w7(32'h3fcd588b),
	.w8(32'h3f751517),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f6592f7),
	.w1(32'h3fc5de13),
	.w2(32'h3f7ec055),
	.w3(32'h3fcfbbec),
	.w4(32'h3e85507e),
	.w5(32'h3fcb0cd9),
	.w6(32'h3eece892),
	.w7(32'hba14909a),
	.w8(32'h3fbb5ed6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfc2a1),
	.w1(32'h3a8e835e),
	.w2(32'hb996c89f),
	.w3(32'h3cac7136),
	.w4(32'hbd8a8e2f),
	.w5(32'hbe13fad1),
	.w6(32'hbe066fa2),
	.w7(32'hbe08cace),
	.w8(32'h39119e64),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd4478e),
	.w1(32'hbda9ca10),
	.w2(32'hbdd603d6),
	.w3(32'h3911573d),
	.w4(32'hbded6064),
	.w5(32'h378e722e),
	.w6(32'hbdb50019),
	.w7(32'hbe6cb828),
	.w8(32'h3e27613f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdf36e5d),
	.w1(32'hba8157d9),
	.w2(32'h3d7a126d),
	.w3(32'hbd66c4ba),
	.w4(32'hbe6b34f8),
	.w5(32'hbe33df1f),
	.w6(32'hbd09900e),
	.w7(32'hbe522089),
	.w8(32'hbd24296f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdd6c9b9),
	.w1(32'hb78faf53),
	.w2(32'hbdf94fb9),
	.w3(32'hbd75f42d),
	.w4(32'hbe1b9bc8),
	.w5(32'hbdf10e6c),
	.w6(32'hbdc47abc),
	.w7(32'h3d421edf),
	.w8(32'hbe3b6ea4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda3ef69),
	.w1(32'h394b089b),
	.w2(32'hbe64bc32),
	.w3(32'hbe461b90),
	.w4(32'hbd908193),
	.w5(32'h3a9b736b),
	.w6(32'hbd82809d),
	.w7(32'h3d5646fa),
	.w8(32'hbab0b9f1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe21d18b),
	.w1(32'hbde723e8),
	.w2(32'hbe021ac7),
	.w3(32'hbe0ae13c),
	.w4(32'hbe56148a),
	.w5(32'hba30322e),
	.w6(32'hb982fdec),
	.w7(32'hbe04f1a0),
	.w8(32'hbe3d672c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9d4ee),
	.w1(32'hbe3346fe),
	.w2(32'h36f61d62),
	.w3(32'hbe21dc2a),
	.w4(32'hbe2bca00),
	.w5(32'hbe1c7f7e),
	.w6(32'hbdeb50f4),
	.w7(32'hbd974981),
	.w8(32'h3bb0e144),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe571786),
	.w1(32'hb937713e),
	.w2(32'hbe3ac071),
	.w3(32'h3e84dad2),
	.w4(32'hb8129d06),
	.w5(32'hbe170a40),
	.w6(32'hbcb1b021),
	.w7(32'hbe8e52c1),
	.w8(32'hbd4e731d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f5c5a2),
	.w1(32'h3e7025c4),
	.w2(32'h3d962f1e),
	.w3(32'hbe53ad80),
	.w4(32'h3e003b2f),
	.w5(32'hbde34d4d),
	.w6(32'hbe09ad2e),
	.w7(32'hbe78f6b8),
	.w8(32'h3e077367),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6685a6),
	.w1(32'hbd7fad90),
	.w2(32'hbdabe56b),
	.w3(32'hbbd9eefb),
	.w4(32'hbda77ef1),
	.w5(32'hbe88c0da),
	.w6(32'hbe3750fc),
	.w7(32'hbd6e6461),
	.w8(32'hb94768b6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdd6ff59),
	.w1(32'hbc6a7e30),
	.w2(32'hbe2dd753),
	.w3(32'hbdc20d99),
	.w4(32'hbccee838),
	.w5(32'hbe02ef03),
	.w6(32'hbe73eb71),
	.w7(32'h37445b57),
	.w8(32'hbc5a98cd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbde82281),
	.w1(32'h3dcf13c0),
	.w2(32'hbccb9735),
	.w3(32'hbe486b01),
	.w4(32'hbe6f5a16),
	.w5(32'hbe678d20),
	.w6(32'hbda0633c),
	.w7(32'hbe43fac3),
	.w8(32'h37c49999),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3de7a4f9),
	.w1(32'h39312006),
	.w2(32'h3d2b6afb),
	.w3(32'h3e325ba0),
	.w4(32'hbe507051),
	.w5(32'hbb8dfe41),
	.w6(32'hbc1c71ee),
	.w7(32'hb9beec4e),
	.w8(32'hbcdfce9e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39491d1c),
	.w1(32'h3b0ccf7c),
	.w2(32'hbd8e8754),
	.w3(32'hbe10e5dc),
	.w4(32'h3dea759f),
	.w5(32'hb9d13a2c),
	.w6(32'hbdd4eb62),
	.w7(32'hbe3face6),
	.w8(32'hbd910b37),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd005cf0),
	.w1(32'h3cdb3537),
	.w2(32'h3dd4fe07),
	.w3(32'hbe2a6998),
	.w4(32'h3d6bcc8f),
	.w5(32'h3d545812),
	.w6(32'hb7a8135e),
	.w7(32'h3826529a),
	.w8(32'hb8adea5b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5f7fe6),
	.w1(32'hb97f1c26),
	.w2(32'h3c0e7f42),
	.w3(32'hb9198e18),
	.w4(32'h3d8a1d3c),
	.w5(32'h3d397392),
	.w6(32'h3d84337e),
	.w7(32'h3d2a2a24),
	.w8(32'h3dfbadc7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule