module layer_8_featuremap_29(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac049a7),
	.w1(32'h3b235926),
	.w2(32'hbbd03012),
	.w3(32'hbac5888d),
	.w4(32'h3a5c9aa2),
	.w5(32'hbbc3d07d),
	.w6(32'hbbed0efc),
	.w7(32'hbb96d5f8),
	.w8(32'hbc1434a2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b0212),
	.w1(32'hb9499d7e),
	.w2(32'h39b2f1e2),
	.w3(32'hbab19083),
	.w4(32'h3973414d),
	.w5(32'h3a664131),
	.w6(32'hba1f0618),
	.w7(32'hb923efb3),
	.w8(32'h3a23d8e7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7e2b1),
	.w1(32'h3b21c4b4),
	.w2(32'h3b1571bc),
	.w3(32'hbb31d8bc),
	.w4(32'hbaa2ecb4),
	.w5(32'hba60947b),
	.w6(32'hbb78132a),
	.w7(32'hbb1b077e),
	.w8(32'hbae64f6d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1023),
	.w1(32'h3a917dba),
	.w2(32'hbca99ee3),
	.w3(32'hbbbddb42),
	.w4(32'hbae66b5f),
	.w5(32'hbc1c66b1),
	.w6(32'hbc3497ec),
	.w7(32'hbbb8c279),
	.w8(32'hbca2af32),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc284388),
	.w1(32'hbb927d32),
	.w2(32'hbb887909),
	.w3(32'hbba486cd),
	.w4(32'h3b0ab40e),
	.w5(32'h3b152bf8),
	.w6(32'hbb8741ed),
	.w7(32'h3b3859e4),
	.w8(32'h3b4fa570),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9a565),
	.w1(32'h3c41d6d8),
	.w2(32'h3c847e73),
	.w3(32'hbc6b27f1),
	.w4(32'h3c9c2200),
	.w5(32'h3cb85804),
	.w6(32'hbc7147b6),
	.w7(32'h3c7cbff0),
	.w8(32'h3cd6ebd1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c683e),
	.w1(32'hb812fa0c),
	.w2(32'h38a82bb1),
	.w3(32'h397706fe),
	.w4(32'h39305161),
	.w5(32'h38ad0a51),
	.w6(32'h39e309e0),
	.w7(32'h391cacb8),
	.w8(32'h37bdd832),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d4207),
	.w1(32'h3b4e1047),
	.w2(32'h3b501c7f),
	.w3(32'hbae66af9),
	.w4(32'h3b757962),
	.w5(32'h3aae6874),
	.w6(32'hbaefb08e),
	.w7(32'h39bc86f1),
	.w8(32'hbb67c016),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54c55b),
	.w1(32'hbb6514bd),
	.w2(32'hba75b244),
	.w3(32'hbb4d6c5f),
	.w4(32'hbba10cbc),
	.w5(32'hba65fe0a),
	.w6(32'hbb155ee4),
	.w7(32'hbb60153e),
	.w8(32'h396559fa),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb2e4),
	.w1(32'hba7c3125),
	.w2(32'hbb99ff84),
	.w3(32'h3b2914ee),
	.w4(32'h3be361d6),
	.w5(32'h3a5cca76),
	.w6(32'hbb0b40c7),
	.w7(32'hbb1373ae),
	.w8(32'hbba936ef),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe58a12),
	.w1(32'hbabb69d0),
	.w2(32'hbc0377b8),
	.w3(32'hbbba8167),
	.w4(32'hbb66684b),
	.w5(32'hbbbaa2c7),
	.w6(32'hbc080831),
	.w7(32'hbba6cd01),
	.w8(32'hbc21f4a2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61a005),
	.w1(32'hbb689f48),
	.w2(32'hbba6fc1d),
	.w3(32'hbbacbce8),
	.w4(32'h3b1ff0f8),
	.w5(32'hbb068562),
	.w6(32'hbc483f84),
	.w7(32'hbb1407d2),
	.w8(32'hbbc16914),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0948b4),
	.w1(32'h3b0119f6),
	.w2(32'h3ad44495),
	.w3(32'hbbd71b9f),
	.w4(32'h3b8324a4),
	.w5(32'h3b93f6bc),
	.w6(32'hbc02f553),
	.w7(32'h3ae57f83),
	.w8(32'h3aaf640d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cffa2),
	.w1(32'h39bf68eb),
	.w2(32'h3886360b),
	.w3(32'h39f7e8b2),
	.w4(32'h399336ea),
	.w5(32'hb911cdb4),
	.w6(32'h3a0fe0de),
	.w7(32'hb773e6d9),
	.w8(32'hb9eb5d3e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b4c19),
	.w1(32'h37b78983),
	.w2(32'hb89060c2),
	.w3(32'h38d9e302),
	.w4(32'hb8a8dcf3),
	.w5(32'hb8ed66af),
	.w6(32'h38d4d943),
	.w7(32'hb9070e51),
	.w8(32'hb903bb38),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba444e04),
	.w1(32'hba937d66),
	.w2(32'hb976dd4c),
	.w3(32'hba517baa),
	.w4(32'hbac115f4),
	.w5(32'hba5c1cf2),
	.w6(32'hba08f423),
	.w7(32'hba8eab3b),
	.w8(32'hba0a5020),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b9e1c),
	.w1(32'h3a800a31),
	.w2(32'h3b10c636),
	.w3(32'hb9f4f46e),
	.w4(32'h3a1ce5ac),
	.w5(32'h3ad7a6e8),
	.w6(32'hba9140bb),
	.w7(32'hba8bf8a6),
	.w8(32'h3afcf0bd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43411d),
	.w1(32'hbc0f8e46),
	.w2(32'hbc275c9a),
	.w3(32'hbb237dd2),
	.w4(32'hbb229a81),
	.w5(32'hbbb8a8b3),
	.w6(32'hbc050261),
	.w7(32'hbbd8cd65),
	.w8(32'hbbccc1db),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd11dad2),
	.w1(32'hbbdcc870),
	.w2(32'hbc8a9591),
	.w3(32'hbd2895dc),
	.w4(32'hbc810df2),
	.w5(32'hbccea7bb),
	.w6(32'hbd0ee4b6),
	.w7(32'hbc396087),
	.w8(32'hbc9a21e9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd525a8b),
	.w1(32'hbce379eb),
	.w2(32'hbd06f068),
	.w3(32'hbcefff8b),
	.w4(32'hbbc296c9),
	.w5(32'hbc3aa825),
	.w6(32'hbd0fbf73),
	.w7(32'hbc02fdec),
	.w8(32'hbc792743),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c4a16),
	.w1(32'hbb08f498),
	.w2(32'h3ba863d6),
	.w3(32'hbba63030),
	.w4(32'h3c112829),
	.w5(32'h3c346f00),
	.w6(32'hbc2fa103),
	.w7(32'h3bff27a8),
	.w8(32'h3c455d12),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a9c7),
	.w1(32'h3bb567aa),
	.w2(32'h3a5dc592),
	.w3(32'hbbc65682),
	.w4(32'h3b9e0329),
	.w5(32'h3b5d589a),
	.w6(32'h39804836),
	.w7(32'h3bd73b64),
	.w8(32'h3b67ce00),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c614976),
	.w1(32'h3b6ee1fd),
	.w2(32'h3bab61e8),
	.w3(32'h3c983825),
	.w4(32'hba8d45ef),
	.w5(32'hba86cf8f),
	.w6(32'h3b9ab464),
	.w7(32'hbbdb45d3),
	.w8(32'hbc6cbc7f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc048a19),
	.w1(32'hbb72afe9),
	.w2(32'hb84e95f0),
	.w3(32'hbbcc9bca),
	.w4(32'hbab88c17),
	.w5(32'h3b8d6865),
	.w6(32'hbc14e280),
	.w7(32'hbb9f6f16),
	.w8(32'h3adf22dc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a382ce3),
	.w1(32'hba17d485),
	.w2(32'h3a7ce6d2),
	.w3(32'h3af498a9),
	.w4(32'hbabbdd31),
	.w5(32'hba128323),
	.w6(32'h3b43ac5d),
	.w7(32'hbabe2593),
	.w8(32'hba26ad2f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b90db),
	.w1(32'h3a285011),
	.w2(32'hba7efe7c),
	.w3(32'hbb324d82),
	.w4(32'h3c1c5ab1),
	.w5(32'h3bb9611f),
	.w6(32'hbbac72c9),
	.w7(32'h3bde81d7),
	.w8(32'h3a510d4e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad91557),
	.w1(32'h3ae96772),
	.w2(32'h3af0329f),
	.w3(32'h3a9dc9f1),
	.w4(32'h3aacddc0),
	.w5(32'h3adb8dc0),
	.w6(32'h3aa7597b),
	.w7(32'h3abd0fc8),
	.w8(32'h3ab317ad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd822418),
	.w1(32'h3c9ec5f9),
	.w2(32'h3cd70504),
	.w3(32'hbb81fd52),
	.w4(32'h3da3f954),
	.w5(32'h3cd77aab),
	.w6(32'hbd857ed8),
	.w7(32'h3cd9d485),
	.w8(32'hbcef2822),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c4775),
	.w1(32'hbb1b5e08),
	.w2(32'hbb8cf295),
	.w3(32'hbb9f8ab5),
	.w4(32'h3b0d1208),
	.w5(32'h38c60f1b),
	.w6(32'hbc1f5007),
	.w7(32'hba00115b),
	.w8(32'hbb71d588),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94fa5f),
	.w1(32'hba7bc79f),
	.w2(32'hbb0d6f7d),
	.w3(32'hbb192b6f),
	.w4(32'h3a8f6c37),
	.w5(32'hb8626377),
	.w6(32'hbb1227c3),
	.w7(32'h3a5adebc),
	.w8(32'hb9b3e6eb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835713),
	.w1(32'h3bc0d430),
	.w2(32'h3b7b0579),
	.w3(32'h3b715429),
	.w4(32'h3bafa781),
	.w5(32'h3b55f33a),
	.w6(32'h3b3b7e25),
	.w7(32'h3b4657de),
	.w8(32'h39a56e32),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba2c18),
	.w1(32'h3b7388d2),
	.w2(32'h3bbad03b),
	.w3(32'hbb835f77),
	.w4(32'h3bbd1b1d),
	.w5(32'h3c17d902),
	.w6(32'h3868e7a7),
	.w7(32'h3c3aec48),
	.w8(32'h3c5d58ab),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c8edd),
	.w1(32'h38c9e1d5),
	.w2(32'h381b2307),
	.w3(32'h3a0ee292),
	.w4(32'h384d9c5e),
	.w5(32'hb88fdc2b),
	.w6(32'h39d52713),
	.w7(32'hb9094a4b),
	.w8(32'hb98945f9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ba22b),
	.w1(32'h39055255),
	.w2(32'h388cd0c7),
	.w3(32'h39d86761),
	.w4(32'h37aa0e1b),
	.w5(32'hb8adad92),
	.w6(32'h39d75d60),
	.w7(32'h378db807),
	.w8(32'hb840f7aa),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61f4a4),
	.w1(32'hbb1b04f7),
	.w2(32'hbbc2a1a3),
	.w3(32'hbc53f410),
	.w4(32'h3af1573a),
	.w5(32'h39129a9e),
	.w6(32'hbc5d0220),
	.w7(32'hb9c4cfb1),
	.w8(32'hbaa6b41a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf63db),
	.w1(32'hbab6d960),
	.w2(32'h39f5b744),
	.w3(32'hbbc89d45),
	.w4(32'hbaaa97f3),
	.w5(32'h39be9f79),
	.w6(32'hbba5ca9b),
	.w7(32'h3aa02faa),
	.w8(32'hb9d942b2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39958aa1),
	.w1(32'hb98b3798),
	.w2(32'h39b0b81c),
	.w3(32'hb8a4fc09),
	.w4(32'hba1182df),
	.w5(32'h39753a67),
	.w6(32'hb899845e),
	.w7(32'hb9b3d717),
	.w8(32'h391f01fb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae58341),
	.w1(32'h3ac4694c),
	.w2(32'h397adc73),
	.w3(32'h3b333a1a),
	.w4(32'h3b2ad345),
	.w5(32'h3ac27a53),
	.w6(32'h3b856cf8),
	.w7(32'h3b53bfa3),
	.w8(32'h3b4c3603),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61bd4b),
	.w1(32'h38498fb7),
	.w2(32'h397840cd),
	.w3(32'h39f380cb),
	.w4(32'hb9e8b12b),
	.w5(32'hb91a573c),
	.w6(32'h39d5e994),
	.w7(32'hb9f2ddfe),
	.w8(32'hb9a69f99),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a5a8f),
	.w1(32'h3a48a628),
	.w2(32'h3a543994),
	.w3(32'h3a30c69e),
	.w4(32'h39597e2b),
	.w5(32'h397f5c1f),
	.w6(32'h3a769e92),
	.w7(32'hb9f789e2),
	.w8(32'hba84c6e0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd745ced),
	.w1(32'h3c858f75),
	.w2(32'hbb3adb06),
	.w3(32'hbcf45691),
	.w4(32'h3d031ad5),
	.w5(32'h3c96be48),
	.w6(32'hbd519a48),
	.w7(32'h3c26daa8),
	.w8(32'hba20993e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9269a0),
	.w1(32'h3aba8732),
	.w2(32'h3b8be5d8),
	.w3(32'hbb82d8d4),
	.w4(32'h3b2c7b16),
	.w5(32'h3b49e9ec),
	.w6(32'hbb9c3423),
	.w7(32'h3b805c5c),
	.w8(32'hbae8cd17),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc252048),
	.w1(32'h3b1725e0),
	.w2(32'h3bdd8869),
	.w3(32'hbc053671),
	.w4(32'h3a6267d6),
	.w5(32'h3b8a2bbe),
	.w6(32'hb9383807),
	.w7(32'h3bca0ec4),
	.w8(32'h39febbf4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e6535),
	.w1(32'hbb52e9b5),
	.w2(32'hbb6fd484),
	.w3(32'hbbf7ce61),
	.w4(32'h3af67e99),
	.w5(32'h3aa95cc6),
	.w6(32'hbc509b8b),
	.w7(32'hbb230350),
	.w8(32'hbba7e309),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72ef16),
	.w1(32'hba953ae7),
	.w2(32'hbc01e5a6),
	.w3(32'hbbd76df2),
	.w4(32'h3af8d733),
	.w5(32'hbbaa6d91),
	.w6(32'hbc1a7eb8),
	.w7(32'hbbdd2383),
	.w8(32'hbcb45d65),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4904e8),
	.w1(32'h3a82f3b7),
	.w2(32'hbbb4e527),
	.w3(32'hbbda26b9),
	.w4(32'h3b962f9c),
	.w5(32'h3b893384),
	.w6(32'hbbfe0eac),
	.w7(32'h3a5ff17e),
	.w8(32'hbc22dd7e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1dd5e),
	.w1(32'hb8ff9fd2),
	.w2(32'h3b61b7ae),
	.w3(32'h3ae4a075),
	.w4(32'h3b39a7d8),
	.w5(32'h3bb363ff),
	.w6(32'hbb56a627),
	.w7(32'h3ae51bed),
	.w8(32'hbb4b4408),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc430ec9),
	.w1(32'hbbdf3919),
	.w2(32'hbb57be2f),
	.w3(32'hbc5cb1b8),
	.w4(32'hbc2f4d39),
	.w5(32'hbc08c323),
	.w6(32'hbbef6c70),
	.w7(32'hbb961265),
	.w8(32'h3af73c1a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeed6d0),
	.w1(32'hba30f220),
	.w2(32'h3b213022),
	.w3(32'hbafca7b7),
	.w4(32'h3b8b3a63),
	.w5(32'h3bc1ced1),
	.w6(32'hbb6eee9d),
	.w7(32'h3bf5e6f5),
	.w8(32'hbab7ca93),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc191b14),
	.w1(32'h3b4256bc),
	.w2(32'hbc2b79ea),
	.w3(32'hbbfa8dce),
	.w4(32'h3b1fa795),
	.w5(32'hbb2df486),
	.w6(32'hbc276a9c),
	.w7(32'hbac92d29),
	.w8(32'hbc367dbc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20a452),
	.w1(32'h3c945d1f),
	.w2(32'h3c9835a3),
	.w3(32'h3a975f77),
	.w4(32'h3cb10b64),
	.w5(32'h3cbd43b4),
	.w6(32'h3b36dc88),
	.w7(32'h3ca9a715),
	.w8(32'h3cb99f50),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd588141),
	.w1(32'hbbc62ac5),
	.w2(32'hbc254310),
	.w3(32'hbd09d372),
	.w4(32'h3c2fa376),
	.w5(32'h3c6be7d0),
	.w6(32'hbd02bde5),
	.w7(32'hbbef9565),
	.w8(32'hbc1a6942),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc878b7e),
	.w1(32'hbbdcefa8),
	.w2(32'hbbb66d1c),
	.w3(32'hbc5f217c),
	.w4(32'hbaef7434),
	.w5(32'h3acb1a37),
	.w6(32'hbc04207e),
	.w7(32'hbba73d0e),
	.w8(32'h3b224362),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1df3ff),
	.w1(32'hbbcaafa0),
	.w2(32'hbc990e21),
	.w3(32'h3b4527fa),
	.w4(32'h3c0f287e),
	.w5(32'hbabb21aa),
	.w6(32'hbc1d4dff),
	.w7(32'hbc2abe32),
	.w8(32'hbc8ce273),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4268d4),
	.w1(32'hb9fbe9e2),
	.w2(32'h3b5a2c09),
	.w3(32'h3a8128b0),
	.w4(32'hbadee033),
	.w5(32'h3b28c096),
	.w6(32'hba58240c),
	.w7(32'h3b7d47b1),
	.w8(32'h3b666d24),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b25b0),
	.w1(32'hbbee42bd),
	.w2(32'hbc35ef6b),
	.w3(32'hbbc67d09),
	.w4(32'h3c18272d),
	.w5(32'hba0122a2),
	.w6(32'hbc1fb503),
	.w7(32'h3b40de24),
	.w8(32'hba2b4700),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b197599),
	.w1(32'h3aa2ad0b),
	.w2(32'h3b06c533),
	.w3(32'h3bbe0238),
	.w4(32'h3b8f7202),
	.w5(32'h3ba99c24),
	.w6(32'hba5a9cf5),
	.w7(32'h3a03816f),
	.w8(32'h396cfc3a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86fc71),
	.w1(32'hbb202122),
	.w2(32'h3b8a78f3),
	.w3(32'hbc668be5),
	.w4(32'hbaae4e48),
	.w5(32'h3c1c9e50),
	.w6(32'hbbcedd1d),
	.w7(32'h3ba2e991),
	.w8(32'hb9a1dfff),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba390a),
	.w1(32'hbb329879),
	.w2(32'hba213011),
	.w3(32'hba8e42a8),
	.w4(32'h39974d20),
	.w5(32'h3acda445),
	.w6(32'hbb923c44),
	.w7(32'hbb0639bc),
	.w8(32'hbbdc2283),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95bb06),
	.w1(32'hbc547e3b),
	.w2(32'hbba697e8),
	.w3(32'hbc4438a7),
	.w4(32'hbb868a3a),
	.w5(32'hbbb43014),
	.w6(32'hbc7ec533),
	.w7(32'hbbcc8205),
	.w8(32'hbb9a8782),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cb796),
	.w1(32'h38ac1f05),
	.w2(32'h3b6e50ae),
	.w3(32'hbb32da1a),
	.w4(32'hbb5c55d5),
	.w5(32'h3b1e2c1f),
	.w6(32'hbb2f7115),
	.w7(32'hbb4a7ea7),
	.w8(32'h3a1ea13b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba938a70),
	.w1(32'h377552c2),
	.w2(32'hbb1278ba),
	.w3(32'hbac8d096),
	.w4(32'hba9946ab),
	.w5(32'hbb0eb0bf),
	.w6(32'h3a2657a5),
	.w7(32'hbb042cc4),
	.w8(32'hbbc04e35),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd26614c),
	.w1(32'hbaa6f758),
	.w2(32'hbbf3bfb4),
	.w3(32'hbcc0f82f),
	.w4(32'h3c7a762d),
	.w5(32'h3c3fbe92),
	.w6(32'hbcd27525),
	.w7(32'h3c2cadfe),
	.w8(32'h3c1d90ee),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb484172),
	.w1(32'hba131efd),
	.w2(32'hbb283fd2),
	.w3(32'hbbddc3e7),
	.w4(32'hbbe1a9fb),
	.w5(32'hbba7ecb8),
	.w6(32'hbb8068b3),
	.w7(32'hbbab4973),
	.w8(32'hbb94bc3f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4db2f5),
	.w1(32'h38181924),
	.w2(32'h3a23ab97),
	.w3(32'hb9dcaaad),
	.w4(32'hba9def8d),
	.w5(32'hb9cf02cd),
	.w6(32'hba65f3e5),
	.w7(32'hbab4d9c4),
	.w8(32'hbac54b7e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860ad1),
	.w1(32'hbaa21dde),
	.w2(32'h3b629902),
	.w3(32'hbb97b04e),
	.w4(32'hbb18d3f5),
	.w5(32'h393be5f3),
	.w6(32'hbbb90e78),
	.w7(32'hbb0b1d7b),
	.w8(32'hbae89d6c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91aa2a),
	.w1(32'hbb8fdd38),
	.w2(32'hbb087e0d),
	.w3(32'hbc21e58c),
	.w4(32'h3b1704ca),
	.w5(32'h3b07f376),
	.w6(32'hbc4f63b3),
	.w7(32'h39c0ead2),
	.w8(32'h3bc3f712),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c0752),
	.w1(32'h3ba43e12),
	.w2(32'h3b826fbc),
	.w3(32'hbbd26146),
	.w4(32'h3c6092f0),
	.w5(32'h3c3b199c),
	.w6(32'hbbea77d4),
	.w7(32'h3c2dfa11),
	.w8(32'h3c29f728),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8221bc),
	.w1(32'hba833ddb),
	.w2(32'hb90606cc),
	.w3(32'hbad14b3f),
	.w4(32'hbaad0b01),
	.w5(32'h385b2609),
	.w6(32'hbae3ed2e),
	.w7(32'hbad984ce),
	.w8(32'hbb914ae2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1141e9),
	.w1(32'hbc439e27),
	.w2(32'hbca377e3),
	.w3(32'hbcd3c4c3),
	.w4(32'hbc1e70b6),
	.w5(32'hbc3ec507),
	.w6(32'hbd04da59),
	.w7(32'hbc8c71ed),
	.w8(32'hbc9c5e8c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab23dd7),
	.w1(32'hbae54e22),
	.w2(32'hba3c6c5d),
	.w3(32'hba9285e5),
	.w4(32'hba90967f),
	.w5(32'hba5ec110),
	.w6(32'hbafd67ea),
	.w7(32'hb9b37b0b),
	.w8(32'hb9ab497b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98d55c),
	.w1(32'hbc081bd5),
	.w2(32'hbc159bb3),
	.w3(32'hbc35ce78),
	.w4(32'hbb412ebd),
	.w5(32'hbb78b7dd),
	.w6(32'hbc365d0c),
	.w7(32'hbb420da7),
	.w8(32'hbc056b79),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba61692),
	.w1(32'hbbc182c3),
	.w2(32'hbb0fb640),
	.w3(32'hbb94add5),
	.w4(32'hbb89419d),
	.w5(32'hbaea3a5f),
	.w6(32'hbbbcfd84),
	.w7(32'hbb4b1423),
	.w8(32'h3b364630),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964d5c7),
	.w1(32'hbb9b568f),
	.w2(32'hbc646a87),
	.w3(32'h3ab8a3f6),
	.w4(32'h3b525e4c),
	.w5(32'hbc041746),
	.w6(32'hbc34b0c1),
	.w7(32'hbc4a4db1),
	.w8(32'hbc4bc90e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e3f5e),
	.w1(32'hbb2147bb),
	.w2(32'hbaf12f4e),
	.w3(32'hbb3b17e9),
	.w4(32'hbabb102d),
	.w5(32'hbab24268),
	.w6(32'hbb51a62f),
	.w7(32'hbb19f7b4),
	.w8(32'hbb216fd9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc300343),
	.w1(32'hbb6ee955),
	.w2(32'hbad9da00),
	.w3(32'hbb7b2d2f),
	.w4(32'h3b2e69bb),
	.w5(32'h3b035a08),
	.w6(32'hbb876158),
	.w7(32'h3a2eeb7b),
	.w8(32'hba7a089a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a3ff1),
	.w1(32'hbb4318eb),
	.w2(32'hbad4be8c),
	.w3(32'hbb352c30),
	.w4(32'hbb167f35),
	.w5(32'hbab033b4),
	.w6(32'hbb678116),
	.w7(32'hbb0c0bf8),
	.w8(32'hbbabad8b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa1f71),
	.w1(32'hbb20642e),
	.w2(32'hbb9cbd15),
	.w3(32'hbcbc919d),
	.w4(32'hbbb784c5),
	.w5(32'hbbf04f4c),
	.w6(32'hbcb9d9fb),
	.w7(32'hbb391b83),
	.w8(32'h3aecd331),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc063cba),
	.w1(32'hbb17e08e),
	.w2(32'hbb70665e),
	.w3(32'hbba91056),
	.w4(32'h3b236cb1),
	.w5(32'hba9e074a),
	.w6(32'hbbb11dbe),
	.w7(32'hbb61f1e9),
	.w8(32'hbb90f791),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990c887),
	.w1(32'hba4ae75d),
	.w2(32'hba9f60b3),
	.w3(32'hb8a7c823),
	.w4(32'hba2bf828),
	.w5(32'hba2937ec),
	.w6(32'hbade337e),
	.w7(32'hbaedf995),
	.w8(32'hbb95197b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15537b),
	.w1(32'h3a8f0518),
	.w2(32'h3b29c907),
	.w3(32'hbb0ec7a4),
	.w4(32'hbb9f8de2),
	.w5(32'hbbb6fc38),
	.w6(32'hbbe6dedc),
	.w7(32'hbbb4a18b),
	.w8(32'hbb0e57a7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca84120),
	.w1(32'hbc14beea),
	.w2(32'hbbde767e),
	.w3(32'hbc133b03),
	.w4(32'h3aee4a59),
	.w5(32'h3aaf4e37),
	.w6(32'hbc6fc08b),
	.w7(32'hbbc11cc7),
	.w8(32'hbb913ef7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6b456),
	.w1(32'hbb1be0a5),
	.w2(32'hbb818bea),
	.w3(32'hbc9f898b),
	.w4(32'h3b5dea88),
	.w5(32'h3b4ecdb8),
	.w6(32'hbcc7fe25),
	.w7(32'h3a9d804c),
	.w8(32'h3b149bd8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd64c073),
	.w1(32'h3c2b2522),
	.w2(32'h3b624607),
	.w3(32'hbd29b574),
	.w4(32'h3cee9a5d),
	.w5(32'h3cb69b99),
	.w6(32'hbd580c86),
	.w7(32'h3c91d445),
	.w8(32'h3c2ba1b4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd313404),
	.w1(32'hbb6e0b7b),
	.w2(32'hbc0ebb32),
	.w3(32'hbc9bbda0),
	.w4(32'h3c4d3e20),
	.w5(32'h3c0db2c4),
	.w6(32'hbcfae4aa),
	.w7(32'h3b4af7b9),
	.w8(32'hbc390d13),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca662ec),
	.w1(32'hbc88805c),
	.w2(32'hbc7ad3b1),
	.w3(32'hbc36eb12),
	.w4(32'hbbd57e9e),
	.w5(32'hbb5deef4),
	.w6(32'hbc70a067),
	.w7(32'hbc855484),
	.w8(32'hbb379538),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c371fe8),
	.w1(32'h3bd26b7c),
	.w2(32'h3c06591c),
	.w3(32'h3c4b26af),
	.w4(32'h3bf890e5),
	.w5(32'h3c036c76),
	.w6(32'h3c209616),
	.w7(32'h3c3c7a54),
	.w8(32'hbb20afe1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca1989),
	.w1(32'hba075810),
	.w2(32'hb976e66e),
	.w3(32'hb8c50a87),
	.w4(32'hb851221d),
	.w5(32'hb98ead85),
	.w6(32'hbb0576c9),
	.w7(32'hbad0a134),
	.w8(32'hbb6a390b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb661c6e),
	.w1(32'hbb39566a),
	.w2(32'hbb1822a0),
	.w3(32'hba03bff4),
	.w4(32'hbb08a184),
	.w5(32'hbab4b56c),
	.w6(32'hbabb84ad),
	.w7(32'hba82be52),
	.w8(32'h3c42a183),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bd16e),
	.w1(32'h3b9113bd),
	.w2(32'h3bdea249),
	.w3(32'h3c4991f7),
	.w4(32'h3b911186),
	.w5(32'h3bccdd89),
	.w6(32'h3c29580f),
	.w7(32'h3c143602),
	.w8(32'h3c157663),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc564ad5),
	.w1(32'hbb284072),
	.w2(32'h3913b0d9),
	.w3(32'hbadbf2e1),
	.w4(32'h3bdb821f),
	.w5(32'h3c4ce1d7),
	.w6(32'hbb96c1b5),
	.w7(32'h3c048a98),
	.w8(32'h3b0a0fb5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97de2e),
	.w1(32'hba2c2c08),
	.w2(32'h3b2662ec),
	.w3(32'h3b543e41),
	.w4(32'h3b1bfaba),
	.w5(32'h3b590833),
	.w6(32'h3af950dc),
	.w7(32'h3b982eb2),
	.w8(32'h3bc627eb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc365f64),
	.w1(32'hbaea046d),
	.w2(32'hbb967532),
	.w3(32'hbb6c2ea4),
	.w4(32'h3c0d6eb3),
	.w5(32'h3bc5aafb),
	.w6(32'hbc4ae6b2),
	.w7(32'h3b55982c),
	.w8(32'h3aa49002),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc869bbb),
	.w1(32'hbbb0f9b6),
	.w2(32'hbbcfd765),
	.w3(32'hbc21a8c7),
	.w4(32'hbaa2fa64),
	.w5(32'hbb2d1b6e),
	.w6(32'hbc486d1f),
	.w7(32'hbb7c83d0),
	.w8(32'hba34aa77),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4446f7),
	.w1(32'h3bcaac0f),
	.w2(32'h3b50c7f4),
	.w3(32'h3b4520fa),
	.w4(32'h3b9d9655),
	.w5(32'h3bbd4d1a),
	.w6(32'h3b95a606),
	.w7(32'h3bade8ba),
	.w8(32'hbbe503d1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88f16c),
	.w1(32'hbb7be22b),
	.w2(32'hba88190a),
	.w3(32'hbc7abddc),
	.w4(32'hbb3e63f4),
	.w5(32'hbb9165e0),
	.w6(32'hbcad9624),
	.w7(32'hbbe0e835),
	.w8(32'hbae7db08),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf453f5),
	.w1(32'hbbfc5c07),
	.w2(32'hbb9febc7),
	.w3(32'hbc86b80a),
	.w4(32'h3ac26aa1),
	.w5(32'h3b9ed895),
	.w6(32'hbc45ffcc),
	.w7(32'h3948b263),
	.w8(32'h3b6bf824),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05349b),
	.w1(32'hbaca4537),
	.w2(32'hba2c0032),
	.w3(32'h3b8add68),
	.w4(32'h3a47e3fe),
	.w5(32'h39e41dbe),
	.w6(32'hbaf8f338),
	.w7(32'hbb160941),
	.w8(32'hbb97fe03),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0de05),
	.w1(32'hbbce5db0),
	.w2(32'hbbd2ec13),
	.w3(32'hbba4b9c5),
	.w4(32'hbbd94528),
	.w5(32'hbbcc5682),
	.w6(32'hbb9e00e2),
	.w7(32'hbbd54490),
	.w8(32'hbb3b0e38),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aa406),
	.w1(32'hbb057457),
	.w2(32'hba2ac2b8),
	.w3(32'hba5ed03c),
	.w4(32'hbae27365),
	.w5(32'hba7229e4),
	.w6(32'hbb3ef841),
	.w7(32'hbb16b22c),
	.w8(32'hbaaebef6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba234d25),
	.w1(32'hb9eeebd2),
	.w2(32'hba386e44),
	.w3(32'h39b04702),
	.w4(32'hb83e2b75),
	.w5(32'hb9df4319),
	.w6(32'hba0ed667),
	.w7(32'hba82ba37),
	.w8(32'hbb3be168),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf65b6e),
	.w1(32'hbb4e5b81),
	.w2(32'hbb9aa045),
	.w3(32'hbb393f20),
	.w4(32'hbb3307b1),
	.w5(32'hbb7631ac),
	.w6(32'hbb4cbbce),
	.w7(32'hbb3bca35),
	.w8(32'hbc4a96ab),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2029d2),
	.w1(32'hbbbae42f),
	.w2(32'hbb8f3778),
	.w3(32'hbc4c7a54),
	.w4(32'hbc19b823),
	.w5(32'hbb97cd96),
	.w6(32'hbbd92d66),
	.w7(32'hbbee8ae7),
	.w8(32'h3b63b2b3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb97c10),
	.w1(32'hbc7b7563),
	.w2(32'hbc1ba569),
	.w3(32'hbc4684a1),
	.w4(32'hba32560f),
	.w5(32'hba9f9942),
	.w6(32'hbc9797c9),
	.w7(32'hbb981edc),
	.w8(32'hba962294),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d71f8),
	.w1(32'hb9adf6ee),
	.w2(32'hbb413236),
	.w3(32'hbaee8e56),
	.w4(32'h3ac63508),
	.w5(32'hba52cd32),
	.w6(32'hbb1a5e6f),
	.w7(32'h3b3fcb5a),
	.w8(32'hbba080ed),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88acdc),
	.w1(32'hbbb3b866),
	.w2(32'hba97d5d6),
	.w3(32'hbc68b242),
	.w4(32'hbb69218f),
	.w5(32'h3b35f1ca),
	.w6(32'hbc813f64),
	.w7(32'hbc05f8ee),
	.w8(32'hbc070612),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05d055),
	.w1(32'hbb88bcb8),
	.w2(32'hbbce2636),
	.w3(32'h3b058af1),
	.w4(32'hbbc03118),
	.w5(32'hbbe104e2),
	.w6(32'hbb30e345),
	.w7(32'hbc231b7c),
	.w8(32'hbb5a0bee),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc813e6c),
	.w1(32'hbb648359),
	.w2(32'hbc15bec0),
	.w3(32'hbc4219b5),
	.w4(32'h3a7985bc),
	.w5(32'hbb5d66f2),
	.w6(32'hbc2025ab),
	.w7(32'h3a0dc48c),
	.w8(32'hbb3d8697),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ac975),
	.w1(32'h3a69f0e1),
	.w2(32'hbb55cbbf),
	.w3(32'hbb0ee616),
	.w4(32'h3b10354d),
	.w5(32'hbaa2253f),
	.w6(32'hba799621),
	.w7(32'h3ad1915e),
	.w8(32'hbb4c108c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb013288),
	.w1(32'hbb762a03),
	.w2(32'hbb48e8c6),
	.w3(32'h3a33403b),
	.w4(32'hbba253cb),
	.w5(32'hba682f2e),
	.w6(32'h3a2800fc),
	.w7(32'hbbb011de),
	.w8(32'hbb860695),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca62143),
	.w1(32'h3b593c48),
	.w2(32'h3adb2d29),
	.w3(32'hbb99e9d1),
	.w4(32'h3c3f7eaa),
	.w5(32'h3bdb59b3),
	.w6(32'hbc91e386),
	.w7(32'h3c0fdad7),
	.w8(32'h3c08d74d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcefc759),
	.w1(32'hbbb70236),
	.w2(32'hbbefb893),
	.w3(32'hbcbd9800),
	.w4(32'h38fd98ca),
	.w5(32'h3aa6ecdc),
	.w6(32'hbc8d2c3e),
	.w7(32'h3bb27248),
	.w8(32'h3ac7b5d0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe386ef),
	.w1(32'hbb178d88),
	.w2(32'hbc0bbce9),
	.w3(32'hbb8bfe86),
	.w4(32'h3affd175),
	.w5(32'hbb81e999),
	.w6(32'hbb96d3e1),
	.w7(32'h3a734f92),
	.w8(32'hbc053c82),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5056d),
	.w1(32'h3a289a78),
	.w2(32'h399c7ce2),
	.w3(32'h3a9c8782),
	.w4(32'hba78fcb9),
	.w5(32'hba640f95),
	.w6(32'h3b01d613),
	.w7(32'hb91ab08b),
	.w8(32'hbab2a3db),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b6ae5),
	.w1(32'h3a221416),
	.w2(32'hbae2eeb9),
	.w3(32'hb90ecf5d),
	.w4(32'hba0ad99a),
	.w5(32'hbabe4b3d),
	.w6(32'hb8891532),
	.w7(32'hb7341a22),
	.w8(32'hbb9a020f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4abb32),
	.w1(32'h3a1321ab),
	.w2(32'hb8d28e72),
	.w3(32'hba29d7f5),
	.w4(32'hb9cd645a),
	.w5(32'hba89efb2),
	.w6(32'h3aee1678),
	.w7(32'h389cab75),
	.w8(32'h3afcf5b8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a48f2),
	.w1(32'hbb058755),
	.w2(32'hbb9502cc),
	.w3(32'hbc15dc3c),
	.w4(32'h3b1beb22),
	.w5(32'h3b62e4ff),
	.w6(32'hbc0d2838),
	.w7(32'hb935a0a4),
	.w8(32'hba987dda),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa57ac),
	.w1(32'h3b25a6a2),
	.w2(32'h3a93b6fd),
	.w3(32'hbc3fc93f),
	.w4(32'h3bb87fa7),
	.w5(32'h3b7bafe8),
	.w6(32'hbc452ec7),
	.w7(32'h3bdc24c6),
	.w8(32'hba865504),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ff429),
	.w1(32'h3ae447a2),
	.w2(32'h3ba49f30),
	.w3(32'hbac53209),
	.w4(32'h3b24e7a7),
	.w5(32'h3b12a5d1),
	.w6(32'hba8fb7fc),
	.w7(32'h3a85c2a6),
	.w8(32'h3a8cc235),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb276f27),
	.w1(32'h3b5cf723),
	.w2(32'h3ba85796),
	.w3(32'h3b2960a2),
	.w4(32'h3bb29520),
	.w5(32'h3b74a57b),
	.w6(32'h3b8e50c6),
	.w7(32'h3bbf4b53),
	.w8(32'hbab0f66d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ff846),
	.w1(32'hbc3fb078),
	.w2(32'hbc002e2c),
	.w3(32'hbae653ad),
	.w4(32'h3c0d8a98),
	.w5(32'h3b60bbd8),
	.w6(32'hbc8c3507),
	.w7(32'hbbf519a5),
	.w8(32'hbbc53524),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32391c),
	.w1(32'hba117b43),
	.w2(32'h3a1128bd),
	.w3(32'hbb903270),
	.w4(32'hbba789c5),
	.w5(32'h3a9c87bd),
	.w6(32'hbabd4976),
	.w7(32'hbc29bd1f),
	.w8(32'hbbdc3211),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd625d),
	.w1(32'hb926b7d9),
	.w2(32'hba591dcf),
	.w3(32'h3aa1311d),
	.w4(32'h3a8bbb2d),
	.w5(32'h399ea681),
	.w6(32'h3a0b7b43),
	.w7(32'hba954a0b),
	.w8(32'h3a0f74d9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f5d6f),
	.w1(32'h3bb922ad),
	.w2(32'h3a3abb89),
	.w3(32'h3b47bcc9),
	.w4(32'h3b748e28),
	.w5(32'hba1226c0),
	.w6(32'h3ab43213),
	.w7(32'h3ae454aa),
	.w8(32'h3b5aa240),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a2362),
	.w1(32'hbb23b54d),
	.w2(32'h3b4e09e0),
	.w3(32'h3a5ab9ea),
	.w4(32'h3b95d115),
	.w5(32'hbb55a073),
	.w6(32'hbbb5021a),
	.w7(32'h3b06dc63),
	.w8(32'hbaa1e77f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9baabf),
	.w1(32'h3a8c00d7),
	.w2(32'hbb668c69),
	.w3(32'hbba52349),
	.w4(32'h39f3c823),
	.w5(32'hbaa101e9),
	.w6(32'hbb41bf29),
	.w7(32'h3b474e6a),
	.w8(32'h3afb9ec0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb541a76),
	.w1(32'h3a4646e0),
	.w2(32'hb8b8eac8),
	.w3(32'hb8af0713),
	.w4(32'h3afb8032),
	.w5(32'hbab370c8),
	.w6(32'hbaa74fbd),
	.w7(32'h3a7d7f39),
	.w8(32'h3a9c2b71),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93c60b),
	.w1(32'h3b391ab7),
	.w2(32'h3ba4d073),
	.w3(32'hbba99cbe),
	.w4(32'hbb631325),
	.w5(32'h3b84e179),
	.w6(32'h3b18569d),
	.w7(32'hbb118720),
	.w8(32'hb8afe01f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule