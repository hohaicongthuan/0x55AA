module layer_8_featuremap_3(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba829dc),
	.w1(32'h39a52aef),
	.w2(32'h3b5e5b42),
	.w3(32'h3c3c2d3e),
	.w4(32'hbb3056c3),
	.w5(32'h39761e43),
	.w6(32'h3b665913),
	.w7(32'hbb9c194b),
	.w8(32'h3ad7b614),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e968e2),
	.w1(32'hbbd0f4b7),
	.w2(32'hba687bbf),
	.w3(32'h3ba076e9),
	.w4(32'hbbdca72f),
	.w5(32'hba1a8816),
	.w6(32'h3a9257c6),
	.w7(32'hbba8cfd8),
	.w8(32'hba8feb0f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7edb5),
	.w1(32'h3a7d31bf),
	.w2(32'h3ae34bba),
	.w3(32'h3bf739ea),
	.w4(32'hbb2fc061),
	.w5(32'hbb2b4257),
	.w6(32'h3b928df2),
	.w7(32'hbb387129),
	.w8(32'hbb09a351),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b136),
	.w1(32'hbbe3eb23),
	.w2(32'hbbd2a73f),
	.w3(32'h3b4fc495),
	.w4(32'hbc091d9a),
	.w5(32'hbbc5e7c7),
	.w6(32'h3b178ccd),
	.w7(32'hbbc26037),
	.w8(32'hbaac8a83),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabca437),
	.w1(32'h3aaef7f3),
	.w2(32'h3b45e220),
	.w3(32'h368b4bd5),
	.w4(32'hbb226e4a),
	.w5(32'h38104648),
	.w6(32'h3b8e5320),
	.w7(32'hbb0fdd6b),
	.w8(32'h3aa71f2e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab63314),
	.w1(32'h3bb12947),
	.w2(32'hba00151f),
	.w3(32'hb90ba244),
	.w4(32'h3bd4d8f6),
	.w5(32'h3b25b571),
	.w6(32'h3aff3bf6),
	.w7(32'h3bfc812f),
	.w8(32'h3c0789f4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898c360),
	.w1(32'hbd53778c),
	.w2(32'hbd8b0e72),
	.w3(32'hbb3b8a60),
	.w4(32'hbd9a1910),
	.w5(32'hbdbe09a3),
	.w6(32'h3abb4605),
	.w7(32'hbd82a257),
	.w8(32'hbd9d9470),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd626617),
	.w1(32'hbab0aafa),
	.w2(32'h3c06ecdd),
	.w3(32'hbd97f3de),
	.w4(32'h3c05bed9),
	.w5(32'h3c5f6c27),
	.w6(32'hbd83ae2c),
	.w7(32'h3bb2bed3),
	.w8(32'h3c06ef14),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89c131),
	.w1(32'h3b8f3ddf),
	.w2(32'h3b2a7cbc),
	.w3(32'h3bd33039),
	.w4(32'h3b8ca295),
	.w5(32'h3b939d8e),
	.w6(32'h3b7a7db8),
	.w7(32'h3bcae9b3),
	.w8(32'h3bdfa369),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c50b1),
	.w1(32'h3b9560cf),
	.w2(32'h3b1d9a4a),
	.w3(32'h3bbad653),
	.w4(32'h3b4a6f1b),
	.w5(32'h3b95185f),
	.w6(32'h3c1b1e1f),
	.w7(32'h3bd51744),
	.w8(32'h3ba31ab1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dde31),
	.w1(32'h3cc89915),
	.w2(32'h3d05bebf),
	.w3(32'h3c3ced2d),
	.w4(32'h3cf4897d),
	.w5(32'h3d1b0cd8),
	.w6(32'h3ba44649),
	.w7(32'h3cc82d5b),
	.w8(32'h3d075798),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd44ab),
	.w1(32'hbb0d72bf),
	.w2(32'h3ac5ed88),
	.w3(32'h3d02b040),
	.w4(32'h3b10f761),
	.w5(32'hbaef83f6),
	.w6(32'h3cce79d3),
	.w7(32'h3ab26a01),
	.w8(32'hbad1732c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54f33c),
	.w1(32'hbc0316c3),
	.w2(32'h3bce3fab),
	.w3(32'hbbbec254),
	.w4(32'hbc13495f),
	.w5(32'h3b04a8e8),
	.w6(32'hba83a8a2),
	.w7(32'h3c0f4395),
	.w8(32'h3c0fe756),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d4482),
	.w1(32'hbd56f8a1),
	.w2(32'hbd9098ad),
	.w3(32'h3abc21d8),
	.w4(32'hbda0a2f0),
	.w5(32'hbddd906f),
	.w6(32'hbadfd886),
	.w7(32'hbd877665),
	.w8(32'hbdaf4438),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3b94db),
	.w1(32'h3c1b3cb6),
	.w2(32'h3ca76132),
	.w3(32'hbd9c756a),
	.w4(32'h3c9eb3c7),
	.w5(32'h3d0009c6),
	.w6(32'hbd61f7d3),
	.w7(32'h3c6f3b3c),
	.w8(32'h3ce12d69),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c375585),
	.w1(32'hba403e3b),
	.w2(32'hb9ee46ab),
	.w3(32'h3cba1712),
	.w4(32'h3c215374),
	.w5(32'h3bf976de),
	.w6(32'h3c9e461f),
	.w7(32'hbaab798a),
	.w8(32'hba287ccf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaecd7),
	.w1(32'h3b11ac2b),
	.w2(32'h3b2e897c),
	.w3(32'h3c41738f),
	.w4(32'h3bea9f5a),
	.w5(32'h3b3367fb),
	.w6(32'h38d654aa),
	.w7(32'h3a834406),
	.w8(32'h3b16e0f0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9fa5d),
	.w1(32'hbbda4b44),
	.w2(32'hbc12688d),
	.w3(32'hbbcadf6a),
	.w4(32'hbc08efae),
	.w5(32'hbc805e70),
	.w6(32'h3aed61d6),
	.w7(32'hbc0ab26f),
	.w8(32'hbc36bd98),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb384c22),
	.w1(32'hbc64b430),
	.w2(32'hbc02f5b4),
	.w3(32'hbbc4d59f),
	.w4(32'hbc1c81c3),
	.w5(32'h3927e5c6),
	.w6(32'hbbdb7d51),
	.w7(32'hbc5cefca),
	.w8(32'h39269c2a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0669a7),
	.w1(32'hbbf27f9f),
	.w2(32'hbc2131af),
	.w3(32'h3c42119c),
	.w4(32'hbc7890f0),
	.w5(32'hbc7e7739),
	.w6(32'hba01e98c),
	.w7(32'hbc2c9a6d),
	.w8(32'hbbe5d209),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff2c47),
	.w1(32'h3c61b967),
	.w2(32'h3cf4ea45),
	.w3(32'hbab900c2),
	.w4(32'h3cce485e),
	.w5(32'h3d21a121),
	.w6(32'h3bc5282e),
	.w7(32'h3c9f2ef1),
	.w8(32'h3d0d1aa4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb887b6),
	.w1(32'hbb0afa12),
	.w2(32'h3baf8f39),
	.w3(32'h3cf55cde),
	.w4(32'h3b91e641),
	.w5(32'h3c310f8d),
	.w6(32'h3cde921d),
	.w7(32'hbc29c888),
	.w8(32'h3b77b36d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb342000),
	.w1(32'hbc1ce644),
	.w2(32'h3b66bc01),
	.w3(32'h3b45836e),
	.w4(32'hba3f8868),
	.w5(32'h3ca24b85),
	.w6(32'hba5a66a6),
	.w7(32'hba1b53c1),
	.w8(32'h3c0ac980),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0e9ce),
	.w1(32'hbcf8eb1a),
	.w2(32'hbd061369),
	.w3(32'h3c34f33b),
	.w4(32'hbd3c75b1),
	.w5(32'hbd4fca33),
	.w6(32'h3c2e8116),
	.w7(32'hbd1bfd19),
	.w8(32'hbd2be6dd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda55e7),
	.w1(32'h3b1dc73a),
	.w2(32'h3befa420),
	.w3(32'hbd2ae1dc),
	.w4(32'h3b8ce90a),
	.w5(32'h3c0d4a76),
	.w6(32'hbd0fd9a4),
	.w7(32'hbbc260d1),
	.w8(32'h3adaea6b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36deb3),
	.w1(32'hb8c8393c),
	.w2(32'hbba6d4d8),
	.w3(32'h3c0dd2fd),
	.w4(32'hb893efa5),
	.w5(32'hbbb8eea3),
	.w6(32'h3c0d5698),
	.w7(32'h3b8a6141),
	.w8(32'h39302c33),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0967dc),
	.w1(32'hbc312de1),
	.w2(32'h3d9222df),
	.w3(32'hbb56e5eb),
	.w4(32'h3cd28977),
	.w5(32'h3e04cf91),
	.w6(32'h3ae3cd18),
	.w7(32'hbbc7eedd),
	.w8(32'h3db24737),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ee441),
	.w1(32'h3b1abd19),
	.w2(32'hbcb30e01),
	.w3(32'h3d36b44a),
	.w4(32'h3c68a193),
	.w5(32'hba99b22c),
	.w6(32'h3bde6a96),
	.w7(32'hbb3ed2ec),
	.w8(32'hbc14c9e9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee607),
	.w1(32'hba9e59d8),
	.w2(32'hbbcb5db8),
	.w3(32'h3a104f00),
	.w4(32'hbb35fa8d),
	.w5(32'hbbe2695e),
	.w6(32'hbba01310),
	.w7(32'h3aa15e12),
	.w8(32'hbbb86193),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba38bdf),
	.w1(32'hbc0b98dc),
	.w2(32'hbc2c006c),
	.w3(32'hbbe2c5ff),
	.w4(32'hbc435d8e),
	.w5(32'hbc636591),
	.w6(32'hbbb04d61),
	.w7(32'hbbd62e6d),
	.w8(32'hbbc9d94c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d5453),
	.w1(32'hbb86475a),
	.w2(32'h38eb95b8),
	.w3(32'hbbb8cae1),
	.w4(32'hb88afc57),
	.w5(32'h3a6bb37c),
	.w6(32'hb76d8c4d),
	.w7(32'hbb02860a),
	.w8(32'h3aa3fa13),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04fca9),
	.w1(32'hbc8f6668),
	.w2(32'hbc84e28e),
	.w3(32'h3b9fd65c),
	.w4(32'hbcac0694),
	.w5(32'hbc95473f),
	.w6(32'h3b8e2fce),
	.w7(32'hbc45864e),
	.w8(32'hbc1c8401),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39aa38),
	.w1(32'hbd0266d5),
	.w2(32'hbd513711),
	.w3(32'hbc52ee35),
	.w4(32'hbd6561f4),
	.w5(32'hbda85be2),
	.w6(32'hbb642a8b),
	.w7(32'hbd43530f),
	.w8(32'hbd87bfad),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ad7d8),
	.w1(32'h3b6e171e),
	.w2(32'h3be1bc17),
	.w3(32'hbd6ddd99),
	.w4(32'h3b631518),
	.w5(32'h3c09f28e),
	.w6(32'hbd35fac9),
	.w7(32'h3a33391b),
	.w8(32'h3be347a5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eb596),
	.w1(32'h3b7bf1ea),
	.w2(32'h3c4c01d2),
	.w3(32'h3b79c7be),
	.w4(32'h3c1ef3b1),
	.w5(32'h3c5b22e4),
	.w6(32'hbb60eb6d),
	.w7(32'h3c036e03),
	.w8(32'h3c8436dd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8c843),
	.w1(32'h3b1b2188),
	.w2(32'h3aea8ef2),
	.w3(32'h3c5667c2),
	.w4(32'h3afa178a),
	.w5(32'h3bbead75),
	.w6(32'h3c2499cd),
	.w7(32'h3b44e874),
	.w8(32'h3be214ae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb675b6),
	.w1(32'hbc4fba95),
	.w2(32'h3bd1962e),
	.w3(32'h3c1202ed),
	.w4(32'hbb5d7c48),
	.w5(32'h3c7f2eaf),
	.w6(32'h3c16adfc),
	.w7(32'hbbdd081f),
	.w8(32'h3c6b8ec1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6bde3),
	.w1(32'h3b045bfc),
	.w2(32'h3b3ef095),
	.w3(32'h3bf96b8a),
	.w4(32'h3b1f480c),
	.w5(32'h3b5bbd91),
	.w6(32'hbaee933a),
	.w7(32'h3bc46900),
	.w8(32'hbb3a2fec),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4ab2d),
	.w1(32'h3bc79fe5),
	.w2(32'h3b752359),
	.w3(32'h3b2344f6),
	.w4(32'h3bb773ba),
	.w5(32'hba0d63b8),
	.w6(32'hbb667548),
	.w7(32'h3c0395c1),
	.w8(32'h3bd96a5d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b596f31),
	.w1(32'h3abb12f8),
	.w2(32'h3b3f7833),
	.w3(32'h3be72eb9),
	.w4(32'h3b8a45c2),
	.w5(32'h3b93bdcf),
	.w6(32'h3b4eee72),
	.w7(32'h3bbc9ed9),
	.w8(32'h3b045d8a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3a7bc),
	.w1(32'hbafcbed7),
	.w2(32'h3b46242f),
	.w3(32'h3aa3ce5b),
	.w4(32'h3adb816d),
	.w5(32'h3a96ae76),
	.w6(32'hba8915d7),
	.w7(32'hbbe702d6),
	.w8(32'h3b6ebc1f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c0295f),
	.w1(32'hbc72d853),
	.w2(32'hbc692333),
	.w3(32'h399e8a08),
	.w4(32'hbcb976bd),
	.w5(32'hbcd24e36),
	.w6(32'h3aa32027),
	.w7(32'hbc9a4cb5),
	.w8(32'hbc903063),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02cfdc),
	.w1(32'hbbcbe1ec),
	.w2(32'hbc07cdb8),
	.w3(32'hbc7c6654),
	.w4(32'hbb8fdcaf),
	.w5(32'hbbe3f2a5),
	.w6(32'hbbf72171),
	.w7(32'hbb8c6cb6),
	.w8(32'hbbb98b0a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7d14e),
	.w1(32'h3b61bdd8),
	.w2(32'h3c05046a),
	.w3(32'hbb4ec52c),
	.w4(32'h3c3523e0),
	.w5(32'h3c0e9624),
	.w6(32'hbb3dfe08),
	.w7(32'h3b541199),
	.w8(32'h3c0de412),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c345133),
	.w1(32'hbb69770a),
	.w2(32'hba3b8c68),
	.w3(32'h3c329b50),
	.w4(32'hbbb989cc),
	.w5(32'h37555506),
	.w6(32'h3c269215),
	.w7(32'hbca6eec7),
	.w8(32'hbc1de31a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5fab2),
	.w1(32'hb96a65cc),
	.w2(32'h3bf74308),
	.w3(32'h3b6c4077),
	.w4(32'h3b559e95),
	.w5(32'h3c3ec09a),
	.w6(32'h3aee771d),
	.w7(32'hbbce898a),
	.w8(32'h3b70f0d5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade9679),
	.w1(32'hbbac020b),
	.w2(32'h3aa3f370),
	.w3(32'h3bd06c6b),
	.w4(32'hbb68e248),
	.w5(32'h3b0f57fc),
	.w6(32'hba5c86ef),
	.w7(32'hbc278dbd),
	.w8(32'hba2b0b7e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b068642),
	.w1(32'hba00154b),
	.w2(32'h3b92c671),
	.w3(32'hbb0651dc),
	.w4(32'h39b9c1c9),
	.w5(32'h3c1498dc),
	.w6(32'hbb2e57c2),
	.w7(32'hbb1835c5),
	.w8(32'h3c2bafbc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9854cc),
	.w1(32'hbcb7da1d),
	.w2(32'hbcf01f03),
	.w3(32'h3b6083ca),
	.w4(32'hbcfc2f4c),
	.w5(32'hbd21c4cf),
	.w6(32'h3b24e2a0),
	.w7(32'hbd030925),
	.w8(32'hbd2323f0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce43d22),
	.w1(32'hbc800d13),
	.w2(32'hbb4c37b0),
	.w3(32'hbd13263e),
	.w4(32'hbc82cfd5),
	.w5(32'h3baabe3c),
	.w6(32'hbd14b9ca),
	.w7(32'hbb624e71),
	.w8(32'h3b6ae615),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a482d),
	.w1(32'hbc5767c2),
	.w2(32'hbc4019f4),
	.w3(32'h3c166221),
	.w4(32'hbc518281),
	.w5(32'hbc6cd569),
	.w6(32'hba5ff067),
	.w7(32'hbc4c5c52),
	.w8(32'hbc55080f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6caea5),
	.w1(32'hbc373138),
	.w2(32'hbc8b4738),
	.w3(32'hbc4803f1),
	.w4(32'hbc0e8e92),
	.w5(32'hbc78e174),
	.w6(32'hbc8424bf),
	.w7(32'hbc45fe90),
	.w8(32'hbc93802f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34e092),
	.w1(32'h3a9a76e2),
	.w2(32'h3abb8fef),
	.w3(32'hbc763947),
	.w4(32'hbaa84aa7),
	.w5(32'h3c1b5a5a),
	.w6(32'hbc4f1aa7),
	.w7(32'hbaf28b2a),
	.w8(32'h3c019111),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5994bd),
	.w1(32'hbc03d120),
	.w2(32'hbb5d9174),
	.w3(32'h3b3757f5),
	.w4(32'hbb8011ac),
	.w5(32'h3bab7b73),
	.w6(32'h3c14ef98),
	.w7(32'hbbd017aa),
	.w8(32'h3c15635c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60ae87),
	.w1(32'h3b4b1236),
	.w2(32'hbbb2d3e8),
	.w3(32'h3b870af4),
	.w4(32'h3b3b7ae3),
	.w5(32'hbbab3d77),
	.w6(32'h3c830372),
	.w7(32'h3a92afe1),
	.w8(32'h39bbed65),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae95c57),
	.w1(32'hbbe064a6),
	.w2(32'hbc13b62d),
	.w3(32'h3ba4000c),
	.w4(32'hbc15fd2d),
	.w5(32'hbc6b210a),
	.w6(32'h3c6be10a),
	.w7(32'hbc1e4ccc),
	.w8(32'hbc370da8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc1e60),
	.w1(32'hbbc3ea71),
	.w2(32'hbbce9bf9),
	.w3(32'hbbd7eeb6),
	.w4(32'hbb49b055),
	.w5(32'hbc1440cb),
	.w6(32'hbb746eeb),
	.w7(32'hbbc9355b),
	.w8(32'hbc12aa53),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3b597),
	.w1(32'h3ba0efd8),
	.w2(32'h3b4d6a34),
	.w3(32'hbb85e377),
	.w4(32'h3bee33e9),
	.w5(32'h3bfff594),
	.w6(32'hbbbf353b),
	.w7(32'hba776b61),
	.w8(32'h3b3a165f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed7e01),
	.w1(32'hbac68c58),
	.w2(32'hba7f4c28),
	.w3(32'h3c053586),
	.w4(32'h3afa1400),
	.w5(32'h3a8fcc2a),
	.w6(32'h38d35ed3),
	.w7(32'h3a4b1ef2),
	.w8(32'h3abf1487),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1e770),
	.w1(32'hbc284237),
	.w2(32'hbbd90739),
	.w3(32'h3b25bb90),
	.w4(32'hbbb3d339),
	.w5(32'h3b949925),
	.w6(32'h3aec1140),
	.w7(32'hbb4e3ae7),
	.w8(32'hbbacf317),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc331b52),
	.w1(32'h39880fe9),
	.w2(32'h3c2e391b),
	.w3(32'h396617a1),
	.w4(32'h3c2b4753),
	.w5(32'h3ca1a7d1),
	.w6(32'h3ac95b77),
	.w7(32'hbb414b7b),
	.w8(32'h3c410a63),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b893ec8),
	.w1(32'hbb45a475),
	.w2(32'h3b8b8cce),
	.w3(32'h3ca4c8f5),
	.w4(32'h3a9a934b),
	.w5(32'h3beac6fd),
	.w6(32'h3c2d3ec1),
	.w7(32'h3a0d8d87),
	.w8(32'h3b38cd64),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb827b8c),
	.w1(32'hbc176471),
	.w2(32'hbc97964f),
	.w3(32'h3b095afc),
	.w4(32'hbc4fe02f),
	.w5(32'hbc94a5c4),
	.w6(32'hba7a1c19),
	.w7(32'hbc6cef33),
	.w8(32'hbc8e2f55),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc466e37),
	.w1(32'hbbe76ee0),
	.w2(32'h3b80c099),
	.w3(32'hbc37e183),
	.w4(32'hbabcdc1c),
	.w5(32'h3c16f700),
	.w6(32'hbc11e864),
	.w7(32'hbbab8c9c),
	.w8(32'h3c6ed745),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2adb7c),
	.w1(32'hbb169e9f),
	.w2(32'h3c04167b),
	.w3(32'h3c668c64),
	.w4(32'h3b67d325),
	.w5(32'h3c263c4f),
	.w6(32'h3bb20266),
	.w7(32'h3a473d67),
	.w8(32'h3c27fc70),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c5555),
	.w1(32'hbb559bff),
	.w2(32'h3b1aeede),
	.w3(32'h3bbd18de),
	.w4(32'hba7a6666),
	.w5(32'h3b811eac),
	.w6(32'h3b5dd1b4),
	.w7(32'h3b0f6422),
	.w8(32'h3bdde9a0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2513),
	.w1(32'hbc3e4d8c),
	.w2(32'hbc98c4d6),
	.w3(32'h3b519a98),
	.w4(32'hbca04d5b),
	.w5(32'hbce3b43b),
	.w6(32'h3c03c793),
	.w7(32'hbc7c4afb),
	.w8(32'hbc85eac1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b9aa1),
	.w1(32'hbae66537),
	.w2(32'h3c06f14f),
	.w3(32'hbc6d9cb6),
	.w4(32'h3c123303),
	.w5(32'h3cfc1371),
	.w6(32'hbb504da1),
	.w7(32'hbb222a86),
	.w8(32'h3c830684),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80405d),
	.w1(32'h3a9626af),
	.w2(32'h3c02528f),
	.w3(32'h3cbdd90b),
	.w4(32'h3c1aa671),
	.w5(32'h3c6dce61),
	.w6(32'h3c73d59f),
	.w7(32'h3bbd6557),
	.w8(32'h3c2c4268),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5575b),
	.w1(32'hbae76c21),
	.w2(32'h395c0b9b),
	.w3(32'h3c8b9230),
	.w4(32'h3b4dcdd0),
	.w5(32'h3bdfe5d2),
	.w6(32'h3bc13aa6),
	.w7(32'hbc1446cc),
	.w8(32'hbc05bcc6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd5d98),
	.w1(32'hbc0d0a01),
	.w2(32'hbc4b5c83),
	.w3(32'h3b07d292),
	.w4(32'hbb9bd299),
	.w5(32'hbc06036a),
	.w6(32'hbb1bc28c),
	.w7(32'h3795c5d2),
	.w8(32'hba8f7829),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc273f03),
	.w1(32'h3b8ec406),
	.w2(32'h3b4323de),
	.w3(32'hbbb257d4),
	.w4(32'h3ac61777),
	.w5(32'h3bab9f85),
	.w6(32'hba459daf),
	.w7(32'hbb75a9e8),
	.w8(32'h3b8af7cf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb239179),
	.w1(32'hbafc76ff),
	.w2(32'hbb262f10),
	.w3(32'h3a430fe7),
	.w4(32'hbb80e187),
	.w5(32'hbb98d0ad),
	.w6(32'hbae4cbca),
	.w7(32'hbbd65873),
	.w8(32'hbbe28c97),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb141d1a),
	.w1(32'hbc0e9729),
	.w2(32'hbc45d222),
	.w3(32'hbbaf6003),
	.w4(32'hbb9a0702),
	.w5(32'hbc2c221c),
	.w6(32'hbc0f7e85),
	.w7(32'h3a6b88b1),
	.w8(32'hba26341f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5d415),
	.w1(32'h3a9b4189),
	.w2(32'h3a296a22),
	.w3(32'hbbc417c1),
	.w4(32'hbae3493d),
	.w5(32'hbace87eb),
	.w6(32'hb9561b1e),
	.w7(32'hbad55c58),
	.w8(32'hbb4c15d9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e36eb),
	.w1(32'hba9b9618),
	.w2(32'hbbff6a7c),
	.w3(32'hbb4f0be9),
	.w4(32'h3a8c7187),
	.w5(32'hbbc3cfd6),
	.w6(32'hbb6c72cf),
	.w7(32'h3c1d1c73),
	.w8(32'h3bcfb804),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e9919),
	.w1(32'h3a5576df),
	.w2(32'h3bcb3bae),
	.w3(32'hbc151563),
	.w4(32'h3ba36dfa),
	.w5(32'h3c004c1d),
	.w6(32'h3bec917a),
	.w7(32'h3bb830b3),
	.w8(32'h3b9a254b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8958b8),
	.w1(32'hbafd15ec),
	.w2(32'h3bd222da),
	.w3(32'h3c28a1c6),
	.w4(32'h3c145cc2),
	.w5(32'h3c882180),
	.w6(32'h3a93b90b),
	.w7(32'h3b960a38),
	.w8(32'h3bd3a882),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3b4a6),
	.w1(32'h3b09b85a),
	.w2(32'h39cbd465),
	.w3(32'h3c8f7531),
	.w4(32'h3989b7c1),
	.w5(32'hba042902),
	.w6(32'h3c0b230d),
	.w7(32'hbb26a1e5),
	.w8(32'hbb1c4cb0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3782b8),
	.w1(32'h3aff5d3c),
	.w2(32'h39b0f44a),
	.w3(32'hbaa2ffaf),
	.w4(32'h3c138510),
	.w5(32'h3c0e6f10),
	.w6(32'hbb6ddad4),
	.w7(32'hbc04def8),
	.w8(32'hbbfb82f2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d425d),
	.w1(32'h3b92fb59),
	.w2(32'h3b93e725),
	.w3(32'h3c0b77c3),
	.w4(32'h3b73faca),
	.w5(32'h3c856fb6),
	.w6(32'hbbe88246),
	.w7(32'h3c17b443),
	.w8(32'h3c03dd47),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6898ee),
	.w1(32'h3946cc3a),
	.w2(32'h3b7371f9),
	.w3(32'h3b02d4a2),
	.w4(32'h3baddcbd),
	.w5(32'h3c06521d),
	.w6(32'hbbbd620c),
	.w7(32'h3b4065a0),
	.w8(32'h3b8e86be),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56b52b),
	.w1(32'h3c041757),
	.w2(32'hb9082d2d),
	.w3(32'h3bf2064d),
	.w4(32'h3bec1110),
	.w5(32'h3b829c58),
	.w6(32'h3ae2a137),
	.w7(32'hbaf67e81),
	.w8(32'h3bc75cf9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0be5d),
	.w1(32'hbad30b19),
	.w2(32'hbc132e4d),
	.w3(32'hbb9c0b34),
	.w4(32'hbbc949ce),
	.w5(32'hbc3f85c6),
	.w6(32'hbbee1460),
	.w7(32'hbb8166ab),
	.w8(32'hbbbe7c6a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb100e7),
	.w1(32'hbb5cd739),
	.w2(32'h3b4aed48),
	.w3(32'hbbaff7e8),
	.w4(32'h3b9f79cd),
	.w5(32'h3c4b9f67),
	.w6(32'hbbbe9810),
	.w7(32'hbbcdf3c1),
	.w8(32'hbafa8391),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b597f44),
	.w1(32'hbc82e94a),
	.w2(32'hbc9285b5),
	.w3(32'h3c4674f9),
	.w4(32'hbb8b92c6),
	.w5(32'h3ad73299),
	.w6(32'h3ac96ebe),
	.w7(32'hbc1b0414),
	.w8(32'h3b833541),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b0f7),
	.w1(32'h3bc984ea),
	.w2(32'h3b8db684),
	.w3(32'h3a197510),
	.w4(32'h3b493363),
	.w5(32'h3c5ac326),
	.w6(32'h3be2a7de),
	.w7(32'hbc0172a3),
	.w8(32'hbb928537),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f9e7),
	.w1(32'hbc16dff1),
	.w2(32'hbc3fd27c),
	.w3(32'h3b0bd2c6),
	.w4(32'hbba8c0ab),
	.w5(32'hbbb79d72),
	.w6(32'h3aec67a8),
	.w7(32'hba4ac8bb),
	.w8(32'h3abcb733),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26c7a2),
	.w1(32'h3a9cbf7f),
	.w2(32'hbb173464),
	.w3(32'hbb710a97),
	.w4(32'h3bc5e8fe),
	.w5(32'h3add21de),
	.w6(32'h3b3bbecb),
	.w7(32'h3c294acb),
	.w8(32'h3c17aa36),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29b216),
	.w1(32'hba83555f),
	.w2(32'h39cea35b),
	.w3(32'h3b0f3f38),
	.w4(32'hbb851039),
	.w5(32'hb96fbdc8),
	.w6(32'h3c0fe838),
	.w7(32'hbc2e0296),
	.w8(32'hbbc54013),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb667d9d),
	.w1(32'h3b754932),
	.w2(32'h3bcb0319),
	.w3(32'hbb5f00d6),
	.w4(32'h3a2d1e87),
	.w5(32'h3b8fc802),
	.w6(32'hbba102e2),
	.w7(32'h3aee1502),
	.w8(32'h3b87e1d6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ec049),
	.w1(32'h3ba42823),
	.w2(32'h3c2b70f0),
	.w3(32'h3ae630cf),
	.w4(32'h3b832654),
	.w5(32'hba7cc186),
	.w6(32'h3b4db1e3),
	.w7(32'hbb23a680),
	.w8(32'hbaf7a7fd),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ee940),
	.w1(32'h3c004822),
	.w2(32'h3bfb6fd6),
	.w3(32'h3b28ea1e),
	.w4(32'h3c3120c9),
	.w5(32'h3c5f1a49),
	.w6(32'hbaf4cade),
	.w7(32'h3ac02e43),
	.w8(32'h3b9a629a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3d20a),
	.w1(32'hbb12cbfa),
	.w2(32'hbb874f27),
	.w3(32'h3c023180),
	.w4(32'hb89fca9d),
	.w5(32'hbb06506d),
	.w6(32'hbab055ce),
	.w7(32'hb9dc8dd2),
	.w8(32'hbad76808),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f500c),
	.w1(32'hbb312d9e),
	.w2(32'hbc027b09),
	.w3(32'hba86f734),
	.w4(32'hbb2afbac),
	.w5(32'hbc016907),
	.w6(32'hbaec4f3c),
	.w7(32'h3b0bc3fc),
	.w8(32'hbacc3631),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefe02d),
	.w1(32'hbb2abdf2),
	.w2(32'hbb8b81fa),
	.w3(32'hbbf0fa1b),
	.w4(32'hba6f56c9),
	.w5(32'hbab69917),
	.w6(32'hba7af959),
	.w7(32'hbb61d97a),
	.w8(32'hbb434d07),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb765411),
	.w1(32'hb8e9ec04),
	.w2(32'hbb070c32),
	.w3(32'h3996634b),
	.w4(32'h3b0c66b8),
	.w5(32'hba303e41),
	.w6(32'hba9e65ad),
	.w7(32'h3b51c060),
	.w8(32'h3aa4647b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87aa9a),
	.w1(32'h3b3bc87a),
	.w2(32'h3af1c829),
	.w3(32'h3a916a5e),
	.w4(32'h3b7ae6df),
	.w5(32'hba5c5d25),
	.w6(32'h3adc6135),
	.w7(32'hba6007d4),
	.w8(32'h3af7abc1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf89c7b),
	.w1(32'h3b99e2b4),
	.w2(32'h3bd3b16c),
	.w3(32'hbbab5510),
	.w4(32'h3b97c8c0),
	.w5(32'h3bfedd85),
	.w6(32'h3a675326),
	.w7(32'hb9244886),
	.w8(32'h3af0a881),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babd4a3),
	.w1(32'h3b5d8418),
	.w2(32'h3bfc1602),
	.w3(32'h3bcb124f),
	.w4(32'h3c5aad33),
	.w5(32'h3c68f662),
	.w6(32'h39f5dc7a),
	.w7(32'h3c60a9c4),
	.w8(32'h3c7d3f89),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cbf2f),
	.w1(32'hbb5d4da4),
	.w2(32'h3b4fc311),
	.w3(32'h3c3e799f),
	.w4(32'h399c5026),
	.w5(32'h3b8bf5f1),
	.w6(32'h3c16db75),
	.w7(32'hbb3d837f),
	.w8(32'h3b9ab492),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bd494),
	.w1(32'hbb7879cc),
	.w2(32'hbb507202),
	.w3(32'h3c865225),
	.w4(32'h3b5d9347),
	.w5(32'h3c3fc72f),
	.w6(32'h3c1bd50a),
	.w7(32'hba1b57f5),
	.w8(32'h3b6ecaf1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf47ff),
	.w1(32'h3ae4c54d),
	.w2(32'h3abd4647),
	.w3(32'h3bd56693),
	.w4(32'hbb3224c5),
	.w5(32'hb87d675d),
	.w6(32'hbb87dd3a),
	.w7(32'h3a5ea319),
	.w8(32'hbaed65a9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccb467),
	.w1(32'hbb29fb6a),
	.w2(32'hbb4bbdd8),
	.w3(32'hba654277),
	.w4(32'hba3fbbbc),
	.w5(32'hbada288b),
	.w6(32'hba614696),
	.w7(32'h3913127d),
	.w8(32'hbaca090d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995a0da),
	.w1(32'hbb21fe29),
	.w2(32'hbb0b80ee),
	.w3(32'hbb0dacdd),
	.w4(32'h3c2e28a3),
	.w5(32'h3c28ccf3),
	.w6(32'hba9a30d4),
	.w7(32'h3abb31f0),
	.w8(32'hb9fa43bc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb835e440),
	.w1(32'hbb0bd9ec),
	.w2(32'h38b64bed),
	.w3(32'h3c76553a),
	.w4(32'h3b5b745f),
	.w5(32'h3b9d4294),
	.w6(32'hbb81a7e2),
	.w7(32'hbaed1e73),
	.w8(32'hbad685a0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fef92),
	.w1(32'hbb4097be),
	.w2(32'hbacc6f8d),
	.w3(32'h3b273cd9),
	.w4(32'hbaec7750),
	.w5(32'hb743f667),
	.w6(32'h380586db),
	.w7(32'hbb018454),
	.w8(32'hbae01266),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67e560),
	.w1(32'hba42361a),
	.w2(32'hbb55e14d),
	.w3(32'h3a0a1db4),
	.w4(32'h3b614dc1),
	.w5(32'h3ac08b27),
	.w6(32'hbaf94509),
	.w7(32'hb9881a9e),
	.w8(32'hbb744358),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea585f),
	.w1(32'hbb3f9f10),
	.w2(32'hbb6fa5bd),
	.w3(32'hb97b0408),
	.w4(32'h3a8dd796),
	.w5(32'hbb882430),
	.w6(32'h3aac26b5),
	.w7(32'hbb2efecb),
	.w8(32'hbcb62818),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b68c),
	.w1(32'hbc29f97e),
	.w2(32'hbbaaa3eb),
	.w3(32'hbb745829),
	.w4(32'hbc414ae5),
	.w5(32'hbc5736a6),
	.w6(32'hbcc95fec),
	.w7(32'hbc23c125),
	.w8(32'hbc04efad),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7191b5),
	.w1(32'hbc0d074a),
	.w2(32'hbb927765),
	.w3(32'hbc944d40),
	.w4(32'h3a74e7a4),
	.w5(32'h3bb40761),
	.w6(32'hbc10471d),
	.w7(32'h3a1cfc12),
	.w8(32'hbb9f1b3b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b7a19),
	.w1(32'hbbccd388),
	.w2(32'hbbbe36e0),
	.w3(32'hbc9887a6),
	.w4(32'hba596215),
	.w5(32'hbc255fb8),
	.w6(32'hbc2f92a9),
	.w7(32'h3adec8ea),
	.w8(32'hbb4945cc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc032926),
	.w1(32'hba6c6bc5),
	.w2(32'hbb1735ae),
	.w3(32'hbc1a97e4),
	.w4(32'hb997c2be),
	.w5(32'hbaae7274),
	.w6(32'hbb2048ef),
	.w7(32'hb936e2af),
	.w8(32'hbaf3e96b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb570b98),
	.w1(32'hba0e96b0),
	.w2(32'h3c065557),
	.w3(32'hbb806b2a),
	.w4(32'hbbc0eda9),
	.w5(32'hbbd7f9b3),
	.w6(32'hbb7f9524),
	.w7(32'hbb834342),
	.w8(32'h3bd8ecc6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2289a5),
	.w1(32'h3b99e08d),
	.w2(32'h3b36ba8b),
	.w3(32'h3b353dee),
	.w4(32'h3b0cc394),
	.w5(32'h3a68d71f),
	.w6(32'h3bb811ad),
	.w7(32'h3a635017),
	.w8(32'h3a4e89c9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76433d),
	.w1(32'h3ad60c8e),
	.w2(32'h3a8451d9),
	.w3(32'h3a3de914),
	.w4(32'h3b83afe4),
	.w5(32'h3b3542e7),
	.w6(32'hba1659dc),
	.w7(32'h3b6bea84),
	.w8(32'h3b0432c0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbe311),
	.w1(32'h3b6b9600),
	.w2(32'h3be63e27),
	.w3(32'h3b3da2dd),
	.w4(32'h3bc17566),
	.w5(32'h3bf73cec),
	.w6(32'h3ad6a37f),
	.w7(32'h3c5d5ed3),
	.w8(32'h3c4223f3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75b921),
	.w1(32'h3a50f4f0),
	.w2(32'h3b86c544),
	.w3(32'h3b513ac2),
	.w4(32'h39f0f0e7),
	.w5(32'h3aa58a8c),
	.w6(32'h3c4419be),
	.w7(32'h3b4840a8),
	.w8(32'h3bbf0cc6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29adef),
	.w1(32'hbbd4e1b6),
	.w2(32'hbbcbb322),
	.w3(32'hbb82cefb),
	.w4(32'hbc6b0900),
	.w5(32'hbc82e204),
	.w6(32'h3b4287e4),
	.w7(32'hbbaf9071),
	.w8(32'hbbd7e2bb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b576d6b),
	.w1(32'h3b5340e0),
	.w2(32'h3bb135fb),
	.w3(32'hbbcf6f52),
	.w4(32'h3ba95a00),
	.w5(32'h3bfeeba2),
	.w6(32'hb9265299),
	.w7(32'h3b1826d9),
	.w8(32'h3b1bd731),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a45cf),
	.w1(32'h3af0d84d),
	.w2(32'hb850f8df),
	.w3(32'h3bdaa283),
	.w4(32'h3aa1f149),
	.w5(32'hb9575133),
	.w6(32'h3b020a60),
	.w7(32'hb9bba2f9),
	.w8(32'hbb2684d8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b202800),
	.w1(32'h3bd39d6c),
	.w2(32'h3bfc0314),
	.w3(32'h3a8e0200),
	.w4(32'h3be24e3c),
	.w5(32'hbaf6f159),
	.w6(32'h3a64ef1c),
	.w7(32'hb8b71eb9),
	.w8(32'hbba7fb4f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8683ca),
	.w1(32'hba1959d8),
	.w2(32'h3a036aec),
	.w3(32'hbb3cabf4),
	.w4(32'hbb0597b9),
	.w5(32'hba8f8c45),
	.w6(32'hbb9b41f6),
	.w7(32'hbb376416),
	.w8(32'hba85023c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b38d7),
	.w1(32'h3b5f6612),
	.w2(32'h3b349f07),
	.w3(32'hba49cc8e),
	.w4(32'h3bbc614d),
	.w5(32'h3c14d6b0),
	.w6(32'h3a203211),
	.w7(32'h3c04c1cd),
	.w8(32'h3bfe0ce5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5a840),
	.w1(32'h3af1b91f),
	.w2(32'h3b2250ef),
	.w3(32'h3b1c07fc),
	.w4(32'hbb260e1b),
	.w5(32'h3aff6d4c),
	.w6(32'hb9002015),
	.w7(32'hbc209dc2),
	.w8(32'hbc5483f4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53f389),
	.w1(32'h3b9959b7),
	.w2(32'hbc5bc1bb),
	.w3(32'hba788776),
	.w4(32'h390224a7),
	.w5(32'hbc8a72f9),
	.w6(32'hbc6c1401),
	.w7(32'h3a9b8a05),
	.w8(32'h3ab358e3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85bb23),
	.w1(32'h3a09d160),
	.w2(32'hbae77908),
	.w3(32'hbc938e74),
	.w4(32'hba45768f),
	.w5(32'hbb3d3355),
	.w6(32'hbbf1e5a5),
	.w7(32'hbb5c3249),
	.w8(32'hbb8f2f31),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cec53),
	.w1(32'hbc521475),
	.w2(32'hbc10cae7),
	.w3(32'hbb555cba),
	.w4(32'hba62321d),
	.w5(32'hbc751abd),
	.w6(32'hbba31280),
	.w7(32'h394fa527),
	.w8(32'hbba8353a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule