module layer_10_featuremap_37(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4ac7f),
	.w1(32'hbc29e0df),
	.w2(32'h3bd1f5c4),
	.w3(32'h3aa0b855),
	.w4(32'hbc44d596),
	.w5(32'h3c7a47c8),
	.w6(32'h3be299d6),
	.w7(32'hbc1099a0),
	.w8(32'h3c6d5219),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1cde2),
	.w1(32'hbb9bf63f),
	.w2(32'hbbdb7c10),
	.w3(32'h3c9058c7),
	.w4(32'h3af5b829),
	.w5(32'h3a00ddf5),
	.w6(32'h3c9ee77b),
	.w7(32'h3bc5ec11),
	.w8(32'h3a58c7ee),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb343f25),
	.w1(32'hbc043730),
	.w2(32'h3b83d4f1),
	.w3(32'hbafdf85b),
	.w4(32'hbba56a95),
	.w5(32'h3ba9169e),
	.w6(32'hb8eb6667),
	.w7(32'hbbc5983c),
	.w8(32'hbb11d9a4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd13ea2),
	.w1(32'h3a4c4072),
	.w2(32'h3bd9d029),
	.w3(32'h3bfb20e7),
	.w4(32'h3bf94297),
	.w5(32'h3b1b2726),
	.w6(32'h3bb3aef6),
	.w7(32'h3c21b4eb),
	.w8(32'h3c10f173),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6b321),
	.w1(32'hbb17c7bc),
	.w2(32'h3bd47095),
	.w3(32'h3b07bbef),
	.w4(32'hbba2266f),
	.w5(32'h3c33a0d7),
	.w6(32'h3af00e56),
	.w7(32'hbb153346),
	.w8(32'h3c545f62),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc374),
	.w1(32'hbc0c3682),
	.w2(32'hba47fb6f),
	.w3(32'h3af4be46),
	.w4(32'hbc1a001d),
	.w5(32'hba943049),
	.w6(32'h3c282fbe),
	.w7(32'hbca1564c),
	.w8(32'hbb6d77ae),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe11bf),
	.w1(32'h3b06cdb4),
	.w2(32'h3c20f532),
	.w3(32'h3bf5e287),
	.w4(32'hbab6d440),
	.w5(32'h3c1cb03d),
	.w6(32'h3b86fd2d),
	.w7(32'hbb88ed9f),
	.w8(32'h3ae198e2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49361f),
	.w1(32'hbb3b007e),
	.w2(32'h3be40bdb),
	.w3(32'h3acf3f09),
	.w4(32'hbc0ca181),
	.w5(32'h3c6b2845),
	.w6(32'hbadf062f),
	.w7(32'hbb22eb99),
	.w8(32'h3c1dd740),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cc40d),
	.w1(32'hbbac8c50),
	.w2(32'hbc292c96),
	.w3(32'hba8fc5a1),
	.w4(32'hbc28e963),
	.w5(32'hbc90d019),
	.w6(32'h3b12f335),
	.w7(32'hbb37b4b9),
	.w8(32'hbc57538a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8346fa),
	.w1(32'h3af1c78b),
	.w2(32'hbaba622f),
	.w3(32'hbbef5393),
	.w4(32'h3b7f43ea),
	.w5(32'hbb98f7b8),
	.w6(32'hbbcc433f),
	.w7(32'h3b71c5d0),
	.w8(32'hbab7d70d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f91e3a),
	.w1(32'h3b013585),
	.w2(32'h3b12a5e0),
	.w3(32'h37c8b16b),
	.w4(32'h3b2f7d43),
	.w5(32'h39f322ed),
	.w6(32'h3b1abe55),
	.w7(32'h3b8a9632),
	.w8(32'h3af47465),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15f8f0),
	.w1(32'hba7f0cd3),
	.w2(32'h3ba911a4),
	.w3(32'h3bf53391),
	.w4(32'h3a91eaf1),
	.w5(32'h3c0b6662),
	.w6(32'h3bca7517),
	.w7(32'h3bf32d4c),
	.w8(32'h3be855b1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5fc9d),
	.w1(32'h3b4dfb8c),
	.w2(32'h3babc0fa),
	.w3(32'h3c14d084),
	.w4(32'h3b9946bf),
	.w5(32'h3c45a075),
	.w6(32'h3bf919ff),
	.w7(32'h3b184468),
	.w8(32'h3c17fb26),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb292b6),
	.w1(32'h3c3dc3dd),
	.w2(32'h3b9a0597),
	.w3(32'h3c49a3bb),
	.w4(32'h39b51f94),
	.w5(32'h3c30953b),
	.w6(32'h3b858f2b),
	.w7(32'h3b092da2),
	.w8(32'h3c0645d1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab66164),
	.w1(32'hbafd802d),
	.w2(32'hbb2516cc),
	.w3(32'h3c0d595c),
	.w4(32'hbc023510),
	.w5(32'hba9e72d4),
	.w6(32'h3c24722e),
	.w7(32'hbb6e06cb),
	.w8(32'hbb85248e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42e54a),
	.w1(32'hbb244138),
	.w2(32'hbb212828),
	.w3(32'h39cccc85),
	.w4(32'hbb784b40),
	.w5(32'hbb5de22f),
	.w6(32'hba9ea822),
	.w7(32'hbba919dd),
	.w8(32'hba86d2ca),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ef08f),
	.w1(32'hb99e5842),
	.w2(32'hbb41e952),
	.w3(32'h3957a176),
	.w4(32'hb99b7995),
	.w5(32'hbaa0c2c8),
	.w6(32'h3b041a57),
	.w7(32'h3a00de49),
	.w8(32'h3aa56a27),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f2b94),
	.w1(32'hbbe7a2bd),
	.w2(32'h3c209a48),
	.w3(32'h3b227cf3),
	.w4(32'hbc0962e6),
	.w5(32'h3c0325fb),
	.w6(32'h3b849446),
	.w7(32'hbba0e6b0),
	.w8(32'h3c1d7206),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87cccc),
	.w1(32'h3b03975f),
	.w2(32'hba007572),
	.w3(32'h3ab7483d),
	.w4(32'h3b63c9da),
	.w5(32'h3bfe71d2),
	.w6(32'h3badc7a2),
	.w7(32'h3bc38f94),
	.w8(32'h3c0905e0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba664953),
	.w1(32'hbb488ee9),
	.w2(32'h3bc5c8ce),
	.w3(32'h3be26254),
	.w4(32'hbba1fe2d),
	.w5(32'h3bea3e75),
	.w6(32'h3c647084),
	.w7(32'hbafaa219),
	.w8(32'h3b94a1aa),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86b0b6),
	.w1(32'hbb0a92f2),
	.w2(32'hba0d0b78),
	.w3(32'h3b697915),
	.w4(32'hbb820014),
	.w5(32'h3b0cbd4b),
	.w6(32'h3baf9c9f),
	.w7(32'hbbcd24cb),
	.w8(32'h3bf062ec),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca3a62),
	.w1(32'h3bc04f35),
	.w2(32'h39df3363),
	.w3(32'h3c1628a3),
	.w4(32'h3c128e2a),
	.w5(32'h3b6b6452),
	.w6(32'h3c24e226),
	.w7(32'h3b9f7040),
	.w8(32'h3b8e8bb8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80044a),
	.w1(32'h3b318385),
	.w2(32'h3ac101d5),
	.w3(32'h3b2573a2),
	.w4(32'hbb4c7629),
	.w5(32'h3b10bb42),
	.w6(32'h3b0f7955),
	.w7(32'hbb4188f8),
	.w8(32'h3b741b3c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9089cc),
	.w1(32'hbb668c9e),
	.w2(32'h3c469e25),
	.w3(32'h3ab2b3cf),
	.w4(32'hbb779b33),
	.w5(32'h3b318e90),
	.w6(32'h3b303648),
	.w7(32'hbb44dde7),
	.w8(32'h3b084935),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9514fb4),
	.w1(32'h3aea3765),
	.w2(32'hbbd6216d),
	.w3(32'h3ba6b1ad),
	.w4(32'h3b24dd17),
	.w5(32'h3bfe325c),
	.w6(32'h3b8b45f8),
	.w7(32'h3af1dec1),
	.w8(32'h3c6e3e51),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf661bb),
	.w1(32'h3b86144f),
	.w2(32'h3bba75e4),
	.w3(32'h3bb55574),
	.w4(32'h3ac914e9),
	.w5(32'hb9cc97c7),
	.w6(32'h3c322303),
	.w7(32'h3aad081a),
	.w8(32'hb9181718),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb90497),
	.w1(32'h3b2c56a7),
	.w2(32'hbb2f37b3),
	.w3(32'h3bbcbd96),
	.w4(32'h3b27db5a),
	.w5(32'hbb28779b),
	.w6(32'h3a45c700),
	.w7(32'h3baac905),
	.w8(32'hbb14049b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b865f69),
	.w1(32'hb9cef9c4),
	.w2(32'hb96648ee),
	.w3(32'h3abb278d),
	.w4(32'hbaf1e7ea),
	.w5(32'h3c93bdfb),
	.w6(32'h3b91d583),
	.w7(32'hbb10c652),
	.w8(32'h3c3b7442),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38547f0a),
	.w1(32'hbc064960),
	.w2(32'h3b8e6089),
	.w3(32'h3c9b9314),
	.w4(32'h3c07b50e),
	.w5(32'h3bd8df54),
	.w6(32'h3c1cf684),
	.w7(32'hba2d2519),
	.w8(32'h3b56978c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402abf),
	.w1(32'hbb8d7970),
	.w2(32'h3d5b2036),
	.w3(32'h3ae55f4f),
	.w4(32'hbaa94b84),
	.w5(32'h3debdbe3),
	.w6(32'h3ae176ea),
	.w7(32'h3b63a170),
	.w8(32'h3d662fde),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3824d),
	.w1(32'hbd458c16),
	.w2(32'h3bd24c35),
	.w3(32'h3ae63cfe),
	.w4(32'hbddff406),
	.w5(32'hbaddb171),
	.w6(32'hbc9ce6a5),
	.w7(32'hbda48b42),
	.w8(32'h3b9606f4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b288759),
	.w1(32'h3b2af35c),
	.w2(32'h3c06d15f),
	.w3(32'h3b588213),
	.w4(32'h398d8ccd),
	.w5(32'hb9846386),
	.w6(32'h3bc2ec15),
	.w7(32'h3bb79bbd),
	.w8(32'h3b336518),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819017),
	.w1(32'h3ba2b180),
	.w2(32'h3dbf72f1),
	.w3(32'h3b66b91d),
	.w4(32'h398a6e5f),
	.w5(32'h3e1b21f2),
	.w6(32'h3acc1fea),
	.w7(32'hb96fe66c),
	.w8(32'h3d9d9414),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94cdc5),
	.w1(32'hbd8eb76b),
	.w2(32'hbbc1f0eb),
	.w3(32'hbc626199),
	.w4(32'hbe2c25f2),
	.w5(32'hba0c6688),
	.w6(32'hbd2d1e42),
	.w7(32'hbe056abb),
	.w8(32'h3c2d03e9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39385dbe),
	.w1(32'h3c73dae1),
	.w2(32'hbd0cc635),
	.w3(32'h3c1dc4f6),
	.w4(32'h3bea7636),
	.w5(32'hbd6ef6be),
	.w6(32'h3c363677),
	.w7(32'h3a97165d),
	.w8(32'hbd143cf0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23425c),
	.w1(32'h3c5ab614),
	.w2(32'h3b62c078),
	.w3(32'hb95556c0),
	.w4(32'h3d541a1a),
	.w5(32'h38cd718e),
	.w6(32'h3c087571),
	.w7(32'h3d20d4ba),
	.w8(32'h3ab43a24),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf11b3),
	.w1(32'hb91691e4),
	.w2(32'h3dd09366),
	.w3(32'hbb2bcdc4),
	.w4(32'hbb8b9358),
	.w5(32'h3e28d76c),
	.w6(32'hba135470),
	.w7(32'h3b945ab5),
	.w8(32'h3dc6c1f6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce06e60),
	.w1(32'hbd5edbb3),
	.w2(32'hbb9d5dce),
	.w3(32'h3c19d37a),
	.w4(32'hbdf9dc34),
	.w5(32'h3c3d7fc5),
	.w6(32'hbc7d46ec),
	.w7(32'hbdb00de7),
	.w8(32'h3c987ba6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacce5e5),
	.w1(32'hba21c8ba),
	.w2(32'hbb989789),
	.w3(32'h3b150d89),
	.w4(32'hbbf16ba8),
	.w5(32'h3acc7e98),
	.w6(32'h3bde98df),
	.w7(32'hbb6eb958),
	.w8(32'h3b8bd6bb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d4c4d),
	.w1(32'hbb16f05d),
	.w2(32'hbab911f3),
	.w3(32'hbc1336f9),
	.w4(32'hbb6b9669),
	.w5(32'hbb175910),
	.w6(32'hbbbf2b07),
	.w7(32'h3a657cf3),
	.w8(32'hbb88046d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814dff),
	.w1(32'h3c1883f8),
	.w2(32'h3aff7142),
	.w3(32'h3bb700e6),
	.w4(32'h3c559002),
	.w5(32'h3c71f913),
	.w6(32'h3ab7715f),
	.w7(32'h3bbb4786),
	.w8(32'h3b4e330a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02f4f4),
	.w1(32'h3aa4fa86),
	.w2(32'hb98413bb),
	.w3(32'h3b7c32ae),
	.w4(32'hbbe274de),
	.w5(32'h3939f3b0),
	.w6(32'hbb332042),
	.w7(32'h39c443de),
	.w8(32'h39b65371),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b913bed),
	.w1(32'hbab4adfa),
	.w2(32'hbd8810b3),
	.w3(32'hbb7938ed),
	.w4(32'h3b85fcd2),
	.w5(32'hbddc98fe),
	.w6(32'h3b5fa07f),
	.w7(32'h3ab6b6a9),
	.w8(32'hbd4454e0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9849f9),
	.w1(32'h3d0ce132),
	.w2(32'hbbf6ec08),
	.w3(32'h3c11614b),
	.w4(32'h3ddd31d9),
	.w5(32'hbc27e33a),
	.w6(32'h3cd23e9f),
	.w7(32'h3d9b591a),
	.w8(32'hbc0c50d9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397eada9),
	.w1(32'h3b573f49),
	.w2(32'hbb9c2395),
	.w3(32'hbb00bf5e),
	.w4(32'hba58ed8d),
	.w5(32'h3b2e534e),
	.w6(32'hba8ff6fa),
	.w7(32'h3996d8e7),
	.w8(32'hbb93f42a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab34c33),
	.w1(32'h3b0626fe),
	.w2(32'h3b61f1cf),
	.w3(32'h3bc59331),
	.w4(32'h3b2b9315),
	.w5(32'h3bc17631),
	.w6(32'hbb18f790),
	.w7(32'hbb9d81d1),
	.w8(32'h3b910d31),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983862c),
	.w1(32'h3abb7b6e),
	.w2(32'hbb9fb288),
	.w3(32'hbad9cd61),
	.w4(32'hba088412),
	.w5(32'h3b1ff99b),
	.w6(32'h3b7d5e80),
	.w7(32'hba26a589),
	.w8(32'h3c17a9e4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b026691),
	.w1(32'h3b6f1a4d),
	.w2(32'hbda4f682),
	.w3(32'hbc1726f1),
	.w4(32'hbbc9b1c7),
	.w5(32'hbe042d50),
	.w6(32'hbb6d1177),
	.w7(32'h3a8bd085),
	.w8(32'hbd89ceab),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb8ece),
	.w1(32'h3d1f56f7),
	.w2(32'h3a951777),
	.w3(32'hbac72278),
	.w4(32'h3df539ad),
	.w5(32'hba8185bb),
	.w6(32'h3cb254d9),
	.w7(32'h3dad3d75),
	.w8(32'h3aafbe0c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fefec),
	.w1(32'h3c160128),
	.w2(32'h3ae3c41b),
	.w3(32'h3c281828),
	.w4(32'h3b8a0dc0),
	.w5(32'h3b2866ab),
	.w6(32'h3c2017a9),
	.w7(32'h3c07ff8c),
	.w8(32'h39ecb3cf),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b645fd3),
	.w1(32'h3b1a4eaa),
	.w2(32'hbb777905),
	.w3(32'hba131708),
	.w4(32'h3bfc7805),
	.w5(32'hbbc703ef),
	.w6(32'hbaebe31c),
	.w7(32'h3b93b657),
	.w8(32'h3a50d034),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3725ab),
	.w1(32'hbc13b3cf),
	.w2(32'h3b1f20b7),
	.w3(32'hbc950381),
	.w4(32'hbb4e367e),
	.w5(32'h3a363ef4),
	.w6(32'hbbbc1dcb),
	.w7(32'h3c670686),
	.w8(32'h3ab3e463),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15906f),
	.w1(32'h39a9753d),
	.w2(32'h3aaed6fb),
	.w3(32'hbc2c6e4d),
	.w4(32'hbb906590),
	.w5(32'hbbf4ce56),
	.w6(32'hbb5e3c6f),
	.w7(32'hbacbd797),
	.w8(32'hbbfffd72),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b9a01),
	.w1(32'h3b816604),
	.w2(32'hbac92419),
	.w3(32'hbbe3f0b1),
	.w4(32'h3afd70b3),
	.w5(32'hbc43670e),
	.w6(32'h3b7e31ad),
	.w7(32'h3be17c09),
	.w8(32'hbb505857),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84a92e9),
	.w1(32'h3aba74dc),
	.w2(32'h3a7245be),
	.w3(32'h3a3340ff),
	.w4(32'hbb14937e),
	.w5(32'hba88daf9),
	.w6(32'h36e1b794),
	.w7(32'h3b97f469),
	.w8(32'hbb385eb6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dfd77),
	.w1(32'h3b962649),
	.w2(32'hbbc8c48d),
	.w3(32'h3a79a137),
	.w4(32'h3b211469),
	.w5(32'h39acf6b5),
	.w6(32'h3b41fbff),
	.w7(32'h3bc85dbc),
	.w8(32'h3baa1440),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb0043),
	.w1(32'h3b5bce95),
	.w2(32'hba99114c),
	.w3(32'h3c11a2bc),
	.w4(32'h3b3d095a),
	.w5(32'h3c3c7df4),
	.w6(32'h3bc3e46d),
	.w7(32'h3bc98a1d),
	.w8(32'h3c272eca),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed14a2),
	.w1(32'h3b5ae75f),
	.w2(32'h3b7a7cff),
	.w3(32'h3c6efcd4),
	.w4(32'h3b904dc0),
	.w5(32'h3c289a46),
	.w6(32'h3c63c6eb),
	.w7(32'h3b614799),
	.w8(32'hbbeef192),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee0990),
	.w1(32'h3c8f4b87),
	.w2(32'hbbff6647),
	.w3(32'hb9ce6c27),
	.w4(32'h3c5d7b57),
	.w5(32'h3b9c0809),
	.w6(32'hbc3e3e2f),
	.w7(32'h3c0cb3a2),
	.w8(32'h3c1dbe50),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6df6b5),
	.w1(32'h3bbb7e9e),
	.w2(32'hbaea9caf),
	.w3(32'h3be8164f),
	.w4(32'h3b5f5526),
	.w5(32'h3c75b0b3),
	.w6(32'h3bd9fe5d),
	.w7(32'hbb179a23),
	.w8(32'h3be6e53f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c004182),
	.w1(32'hba9673ae),
	.w2(32'hb92ae7e4),
	.w3(32'h3bab10e3),
	.w4(32'h3a8bcba4),
	.w5(32'hbbb5462e),
	.w6(32'hbac11e70),
	.w7(32'h3ba59422),
	.w8(32'h3ae8e88b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443ece),
	.w1(32'h3b304a5b),
	.w2(32'hba1a5a89),
	.w3(32'hbc1e787b),
	.w4(32'h3a7c5e76),
	.w5(32'hb86f6578),
	.w6(32'hbb50c684),
	.w7(32'hba97e8d0),
	.w8(32'hbb45b2be),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae2c53),
	.w1(32'hbb8970eb),
	.w2(32'h3a8f5b6d),
	.w3(32'h3c153100),
	.w4(32'h3b0e3e6e),
	.w5(32'h3c3d9f5c),
	.w6(32'h3bb8c22b),
	.w7(32'hbb8177b3),
	.w8(32'h3abe7904),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaa407),
	.w1(32'h3b846704),
	.w2(32'h3a16c63f),
	.w3(32'hbbc08388),
	.w4(32'hbc7f8b56),
	.w5(32'h3a0a6f6b),
	.w6(32'hba853e1c),
	.w7(32'h3a74640a),
	.w8(32'h3b820ded),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4ee14),
	.w1(32'hba5107ee),
	.w2(32'h3bbf7d76),
	.w3(32'h3af1539b),
	.w4(32'hba4b500e),
	.w5(32'h3c1a4c97),
	.w6(32'h39be7d88),
	.w7(32'h3b915f74),
	.w8(32'h3bb54799),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b787),
	.w1(32'h3bc10a23),
	.w2(32'h3c0e8a2a),
	.w3(32'h3c3387da),
	.w4(32'h3c0b7b87),
	.w5(32'h3c840fc6),
	.w6(32'h3c293d14),
	.w7(32'h3c2c688f),
	.w8(32'h3c8f7117),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1ccec),
	.w1(32'hbc8bc657),
	.w2(32'hbacd2720),
	.w3(32'hbbba8e56),
	.w4(32'hbcda2bdc),
	.w5(32'hbb1ff68b),
	.w6(32'hbb1c827e),
	.w7(32'hbc7680c1),
	.w8(32'h3b2689c8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb7bfb),
	.w1(32'h3aa5ba4c),
	.w2(32'hb997f3a0),
	.w3(32'hbaa9c084),
	.w4(32'h38308e47),
	.w5(32'h3ae2a1a7),
	.w6(32'hbc18b714),
	.w7(32'hbba72660),
	.w8(32'h3ab0fd5a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18618d),
	.w1(32'h398caf42),
	.w2(32'hbb9839c2),
	.w3(32'hbaca132e),
	.w4(32'hbbedd20f),
	.w5(32'hbb84fe12),
	.w6(32'hba21b135),
	.w7(32'hbbde29ef),
	.w8(32'hbc44abf7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8be512),
	.w1(32'h3b62d4ae),
	.w2(32'hbc27658d),
	.w3(32'h3bd37993),
	.w4(32'h3bf7a60b),
	.w5(32'hbc776dfb),
	.w6(32'hb8b21c86),
	.w7(32'hbaa58ffb),
	.w8(32'hbb951a1d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4ee1f),
	.w1(32'hb7a2673e),
	.w2(32'h3b75a145),
	.w3(32'hbd185589),
	.w4(32'h37a7141d),
	.w5(32'h3b9101a8),
	.w6(32'hbcac28eb),
	.w7(32'h3b93985e),
	.w8(32'h381e9162),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99022f),
	.w1(32'hbb51111d),
	.w2(32'h3a13ec21),
	.w3(32'h3b622bcd),
	.w4(32'h3b832f47),
	.w5(32'h3ae8283a),
	.w6(32'hbb9eff10),
	.w7(32'h3b480fb3),
	.w8(32'h3aa06bda),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b882b),
	.w1(32'hbb8716b8),
	.w2(32'h3b8ee749),
	.w3(32'hbc1bedee),
	.w4(32'h3b88290e),
	.w5(32'h3c368cbc),
	.w6(32'hbbc14b20),
	.w7(32'hbb8c6a2e),
	.w8(32'h3c145b67),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4afb0a),
	.w1(32'h3bcc249e),
	.w2(32'hbda0f2f8),
	.w3(32'h388aafa7),
	.w4(32'h3bd1f0a7),
	.w5(32'hbdbb909a),
	.w6(32'h3bc7d784),
	.w7(32'h3bf213ee),
	.w8(32'hbd792324),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb657fd),
	.w1(32'h3cfd619e),
	.w2(32'h3bd5bca7),
	.w3(32'h3c9616f2),
	.w4(32'h3dded550),
	.w5(32'h3c1e966f),
	.w6(32'h3cc08a45),
	.w7(32'h3d9e04d5),
	.w8(32'h3ba32036),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf1b9c),
	.w1(32'hba42359a),
	.w2(32'hbc043701),
	.w3(32'h3b550099),
	.w4(32'hbb6b24ec),
	.w5(32'hbb5f3a51),
	.w6(32'h3b9b367a),
	.w7(32'hba0ffff5),
	.w8(32'hbba0eee3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc321bfd),
	.w1(32'hbbb3eff8),
	.w2(32'hbb839471),
	.w3(32'hbc1a89f7),
	.w4(32'hbc06fa1d),
	.w5(32'hbc0f2add),
	.w6(32'hbba075c0),
	.w7(32'hba4be708),
	.w8(32'h3ad80327),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d49de),
	.w1(32'h3aed8137),
	.w2(32'h3bb250a2),
	.w3(32'hbc0c4cce),
	.w4(32'hbbb48883),
	.w5(32'h3b5b80fd),
	.w6(32'hbbc23484),
	.w7(32'hbb6f2422),
	.w8(32'h3a95f5fa),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c215b),
	.w1(32'hbb35cca3),
	.w2(32'hbb4b3973),
	.w3(32'h3b55ef2d),
	.w4(32'h3bb6b0bb),
	.w5(32'h3bfe6fb6),
	.w6(32'h3aac626d),
	.w7(32'h3b555079),
	.w8(32'hbb5392bc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad19493),
	.w1(32'hbb40be0b),
	.w2(32'h3b01f70e),
	.w3(32'h3c73719c),
	.w4(32'h3c8c9c21),
	.w5(32'hbba8c5f3),
	.w6(32'h3b9f27e9),
	.w7(32'hbb880403),
	.w8(32'h3b377f45),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6484b6),
	.w1(32'h3afff09b),
	.w2(32'h3d0780cd),
	.w3(32'hbc9ddf00),
	.w4(32'hbb81da54),
	.w5(32'h3d9b6d33),
	.w6(32'hbb1846ea),
	.w7(32'h3b629409),
	.w8(32'h3d0babae),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bc5c8),
	.w1(32'hbc9d580d),
	.w2(32'hbbf6b8bd),
	.w3(32'h3c3170a6),
	.w4(32'hbd6542e0),
	.w5(32'hbc0b1fb9),
	.w6(32'hbbf5b57e),
	.w7(32'hbd2237f3),
	.w8(32'hbc1d9c89),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ae2a),
	.w1(32'hbb890e6a),
	.w2(32'hbba03ff6),
	.w3(32'hbb143e7b),
	.w4(32'hb8a6639e),
	.w5(32'hbc051274),
	.w6(32'hbb19b3f8),
	.w7(32'hbab76b51),
	.w8(32'hbb20533b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf243d3),
	.w1(32'hbb41c6f9),
	.w2(32'h3b768e93),
	.w3(32'hbc8dc650),
	.w4(32'hbbc2665f),
	.w5(32'h3bc5cbce),
	.w6(32'hbc0b5c45),
	.w7(32'h3b170a98),
	.w8(32'h3a040ee8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb874a3c2),
	.w1(32'hbb43750e),
	.w2(32'hbc5d926e),
	.w3(32'h3b40c749),
	.w4(32'h3b60c90d),
	.w5(32'hbc86eb1f),
	.w6(32'hbb9ddb2b),
	.w7(32'h3b6aca30),
	.w8(32'hbb33f746),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4caec1),
	.w1(32'hba998ddc),
	.w2(32'h3bc9cfbe),
	.w3(32'hbbb22340),
	.w4(32'hbb7a5ab1),
	.w5(32'h3c609f80),
	.w6(32'hbbc07fff),
	.w7(32'hba97d4f1),
	.w8(32'h3c10fbc2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7b037),
	.w1(32'h3c029751),
	.w2(32'hbbb40424),
	.w3(32'h3c64a77d),
	.w4(32'h3c63a5e3),
	.w5(32'hbbc4f753),
	.w6(32'h3bf02eba),
	.w7(32'h3c5289de),
	.w8(32'hbb5bb9c8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e227),
	.w1(32'h3b024817),
	.w2(32'hbb85bfb1),
	.w3(32'h3b651035),
	.w4(32'h3c48299c),
	.w5(32'h3b95d0b2),
	.w6(32'h3c2c1bd9),
	.w7(32'h3c903afe),
	.w8(32'h3bb2cd89),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9174f),
	.w1(32'hbb968f86),
	.w2(32'hbb36cea8),
	.w3(32'hbb3cfe2e),
	.w4(32'hb96a4db2),
	.w5(32'h39f80ba3),
	.w6(32'h38878f95),
	.w7(32'hbadf50df),
	.w8(32'h3c41ce6e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea2cef),
	.w1(32'hb907909f),
	.w2(32'h3c2746d0),
	.w3(32'hb8891701),
	.w4(32'hbb9d674b),
	.w5(32'h3c2cf0f2),
	.w6(32'h3ae61ab6),
	.w7(32'hbb1359d8),
	.w8(32'hbab61122),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c552),
	.w1(32'hbc2f1b38),
	.w2(32'hbbcb9705),
	.w3(32'hbac517ca),
	.w4(32'hba390907),
	.w5(32'hbbd9f2d5),
	.w6(32'h3b5519af),
	.w7(32'h3c4afbaa),
	.w8(32'hbb9709fe),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad038bf),
	.w1(32'h3ae58771),
	.w2(32'hbc0dcb9d),
	.w3(32'h3b39f39b),
	.w4(32'h3c7da144),
	.w5(32'hbb456a54),
	.w6(32'h3a085dc8),
	.w7(32'h3c21175d),
	.w8(32'hbc22ee32),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2110b3),
	.w1(32'hb7b85e87),
	.w2(32'hbd107579),
	.w3(32'h39ab0bf2),
	.w4(32'h398bd069),
	.w5(32'hbd2e4615),
	.w6(32'hbbdc9279),
	.w7(32'hbb06ee3c),
	.w8(32'hbcafe2ea),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf61b09),
	.w1(32'h3c956b05),
	.w2(32'hbba6aa69),
	.w3(32'h3c1ac132),
	.w4(32'h3d408424),
	.w5(32'h3badfaf3),
	.w6(32'h3c707b5c),
	.w7(32'h3d1a1a22),
	.w8(32'hbb998957),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98420b3),
	.w1(32'h39d452db),
	.w2(32'h3a93bbe7),
	.w3(32'hbbb22975),
	.w4(32'h3b870a80),
	.w5(32'h3bbb4db0),
	.w6(32'h39646db0),
	.w7(32'hba09bf49),
	.w8(32'h3b969189),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b910ebf),
	.w1(32'hbb46ef72),
	.w2(32'hbb342f62),
	.w3(32'hb92f779e),
	.w4(32'hbb9bec95),
	.w5(32'h3a870a51),
	.w6(32'h3bb32c8c),
	.w7(32'hbc2d501e),
	.w8(32'hbc120dbe),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44f5a0),
	.w1(32'hbaa5ba0e),
	.w2(32'hbb1fc946),
	.w3(32'hbb53f179),
	.w4(32'hbbc6ab04),
	.w5(32'hb9277e20),
	.w6(32'hbc1fedd5),
	.w7(32'h3b356f9b),
	.w8(32'hbac9fa39),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80c0f6),
	.w1(32'hbb178367),
	.w2(32'h39096e66),
	.w3(32'hbb4a86fa),
	.w4(32'hbbb96196),
	.w5(32'hbb7017dd),
	.w6(32'hbab3ceda),
	.w7(32'hbbba5f23),
	.w8(32'h3b5ea1a6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37a73),
	.w1(32'h3c06876f),
	.w2(32'hbc24dcf3),
	.w3(32'h3acf7e13),
	.w4(32'h3b4e2eef),
	.w5(32'hbc940f5d),
	.w6(32'h3b6affa0),
	.w7(32'hbb143439),
	.w8(32'hbc3b2be7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce18d23),
	.w1(32'hbba15847),
	.w2(32'hbb419d31),
	.w3(32'hbd1ba49b),
	.w4(32'hbba0db6e),
	.w5(32'hbb802944),
	.w6(32'hbcfda00b),
	.w7(32'hbba7908e),
	.w8(32'hb8bfc269),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7412e),
	.w1(32'h3c0d8e7a),
	.w2(32'h3b6b1e4a),
	.w3(32'h3a9789f4),
	.w4(32'hb95045b8),
	.w5(32'hbba2db65),
	.w6(32'hbb8874c8),
	.w7(32'h3aeb4f0c),
	.w8(32'h3b0eacbb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44faf3),
	.w1(32'hbaa89996),
	.w2(32'hbb244c8b),
	.w3(32'h3c161964),
	.w4(32'h3b09a516),
	.w5(32'hbba12615),
	.w6(32'hbb6c1038),
	.w7(32'h3bb5fc03),
	.w8(32'hbb19e1cc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2308d1),
	.w1(32'h3ab73f4f),
	.w2(32'hbbbe47ec),
	.w3(32'hbc1f958d),
	.w4(32'h3b319773),
	.w5(32'hbca27ddc),
	.w6(32'hbba97450),
	.w7(32'hbad9c406),
	.w8(32'hbc9cc186),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc229fe),
	.w1(32'hbbcb5b76),
	.w2(32'hbbebe031),
	.w3(32'hbd1a4915),
	.w4(32'hbb0f8e6f),
	.w5(32'hbbc7f9b9),
	.w6(32'hbcbfc681),
	.w7(32'h3b340bc5),
	.w8(32'hbba7b0d7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895138),
	.w1(32'hbbcda416),
	.w2(32'hbb7785bf),
	.w3(32'hbb648414),
	.w4(32'hbbbe86c6),
	.w5(32'hbbc00e88),
	.w6(32'hbbb2be51),
	.w7(32'hbc194b7c),
	.w8(32'hbbdfddeb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2406b),
	.w1(32'h3ac02180),
	.w2(32'hbba0b69d),
	.w3(32'hbbc9ec8a),
	.w4(32'h3b2be368),
	.w5(32'h3a20a8f5),
	.w6(32'hbbb44a54),
	.w7(32'h3aaab4a6),
	.w8(32'h3a21da66),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93979c),
	.w1(32'h3a59590d),
	.w2(32'hba3b16d2),
	.w3(32'h39c9cb42),
	.w4(32'h3bb0471d),
	.w5(32'hbc424acd),
	.w6(32'hba37af0f),
	.w7(32'h3ba412a0),
	.w8(32'h39b91715),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00229a),
	.w1(32'h3b1b2260),
	.w2(32'hbb427fe8),
	.w3(32'hbc30881d),
	.w4(32'hbb4ff1f5),
	.w5(32'hb98b88fb),
	.w6(32'hbc5d822f),
	.w7(32'hbbf3c220),
	.w8(32'hbb6a365a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2932a6),
	.w1(32'h3a93c45a),
	.w2(32'hba902663),
	.w3(32'h39c36a36),
	.w4(32'h381a2644),
	.w5(32'hbb8f4c19),
	.w6(32'hbc0b8e5f),
	.w7(32'hb9ae6b12),
	.w8(32'h3ba06e19),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a811cac),
	.w1(32'h3b066afc),
	.w2(32'hbbe9aa4e),
	.w3(32'h3b791834),
	.w4(32'h3b04a7c8),
	.w5(32'hbba0c954),
	.w6(32'hbb7eba21),
	.w7(32'hba9cf06b),
	.w8(32'hbb5642a4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e45232),
	.w1(32'hbb98db2c),
	.w2(32'hb91a3f46),
	.w3(32'hbaac0ca0),
	.w4(32'h396146e4),
	.w5(32'h3bbaf570),
	.w6(32'hbb837ab3),
	.w7(32'h3b258210),
	.w8(32'h3c14980f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0d6b1),
	.w1(32'h3ba35529),
	.w2(32'h3b11dcd6),
	.w3(32'h3b3398ac),
	.w4(32'h3c0dd08a),
	.w5(32'hbb1b6a78),
	.w6(32'h3b8eac06),
	.w7(32'h3b4dc8c7),
	.w8(32'hbc1d5a85),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48aace),
	.w1(32'hbbd835a2),
	.w2(32'hbb26981a),
	.w3(32'hbc1ec601),
	.w4(32'hbc144883),
	.w5(32'h3b2ad277),
	.w6(32'hbc1a543b),
	.w7(32'hbbb7639c),
	.w8(32'h3ad67172),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeeaa24),
	.w1(32'h3c350f37),
	.w2(32'hbc0b0c20),
	.w3(32'h3ba238f8),
	.w4(32'h3bad99dc),
	.w5(32'hbb22a78e),
	.w6(32'hb922115f),
	.w7(32'h3b433af9),
	.w8(32'h3b66eca7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba45bdc),
	.w1(32'h3a93844e),
	.w2(32'hbbe81da8),
	.w3(32'h3b849ee7),
	.w4(32'hbb0cbdfe),
	.w5(32'h3a3bd382),
	.w6(32'h3a1911fb),
	.w7(32'hbb3858a5),
	.w8(32'hba21d5e2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b343a),
	.w1(32'h399afb2c),
	.w2(32'h3ac19dbb),
	.w3(32'hb9149070),
	.w4(32'hba0c64e7),
	.w5(32'hb9bb1ae4),
	.w6(32'hbbb27274),
	.w7(32'hbbb9c31f),
	.w8(32'hbc158b02),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe27544),
	.w1(32'hbb7b1c54),
	.w2(32'h3b35f61c),
	.w3(32'hbb2fed0e),
	.w4(32'h3b3dbd3d),
	.w5(32'h3bc84c61),
	.w6(32'h3a1e2725),
	.w7(32'h3c0dde3f),
	.w8(32'hbb7c3a00),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0cb86),
	.w1(32'h3bd1b1f8),
	.w2(32'h3ba12403),
	.w3(32'h3ba58438),
	.w4(32'h382ae577),
	.w5(32'h3b64a0c4),
	.w6(32'h39f178d3),
	.w7(32'hbb1894b6),
	.w8(32'h3be9b5c0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c09b04),
	.w1(32'h3bcbb759),
	.w2(32'h3a8f5a88),
	.w3(32'h3ae11276),
	.w4(32'h3bbd506f),
	.w5(32'hbb8cbe1e),
	.w6(32'h3b997cc9),
	.w7(32'h3bd39cc2),
	.w8(32'h3b26ee96),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ebdb),
	.w1(32'h3b8fa103),
	.w2(32'hbb7b8c6c),
	.w3(32'hbbf924d3),
	.w4(32'h3b5b6ab1),
	.w5(32'h3b568c2d),
	.w6(32'hbbb61ff4),
	.w7(32'h3a781683),
	.w8(32'hbad64d38),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53355d),
	.w1(32'h3b17acdb),
	.w2(32'h3c000560),
	.w3(32'hbb06ea92),
	.w4(32'h3b99f4d9),
	.w5(32'h3cb79927),
	.w6(32'hb98f5c91),
	.w7(32'h3bc520f9),
	.w8(32'h3c32a721),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b389a53),
	.w1(32'hbb7a4292),
	.w2(32'h3c65cc02),
	.w3(32'hba771fc6),
	.w4(32'hbc76c9ae),
	.w5(32'h3d2c03a0),
	.w6(32'hbac7fa52),
	.w7(32'hbc237301),
	.w8(32'h3c67b879),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a169c6b),
	.w1(32'hbca33dc3),
	.w2(32'hbc3ed375),
	.w3(32'hbaf4b850),
	.w4(32'hbd40e2f6),
	.w5(32'hba426763),
	.w6(32'hbc1a9fd2),
	.w7(32'hbd023b39),
	.w8(32'hbbd3a4eb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a4758),
	.w1(32'hbc9e0602),
	.w2(32'h3bc6b0b9),
	.w3(32'hbcbb34cb),
	.w4(32'hbc7d8dc5),
	.w5(32'h3c9c0f1a),
	.w6(32'hbc3016b7),
	.w7(32'hbc088924),
	.w8(32'h3c176ef6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c0bea),
	.w1(32'h3bec46a9),
	.w2(32'hbc2e1fe7),
	.w3(32'h3caa5604),
	.w4(32'h3c7eef08),
	.w5(32'hbc2a1033),
	.w6(32'h3c53a441),
	.w7(32'h3bc9733c),
	.w8(32'hbba38594),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9f3f),
	.w1(32'h3ac68481),
	.w2(32'hbbb7d201),
	.w3(32'hbbcfef6f),
	.w4(32'h3b90637f),
	.w5(32'hbab2c9d9),
	.w6(32'hbb803224),
	.w7(32'h3c13ccc5),
	.w8(32'hba9d343c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b148959),
	.w1(32'h3a3d76e3),
	.w2(32'hbb75a66e),
	.w3(32'hbbd3e4d0),
	.w4(32'hbc049ef8),
	.w5(32'h3a9ff0c1),
	.w6(32'hbc209e2b),
	.w7(32'hbb86bf1d),
	.w8(32'h3a9bba67),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00df61),
	.w1(32'hbba3a30c),
	.w2(32'h3a420a2c),
	.w3(32'hbc047f75),
	.w4(32'hbbebae67),
	.w5(32'h3be6a288),
	.w6(32'hbc17a32c),
	.w7(32'h3b04a921),
	.w8(32'h3b945d54),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04587b),
	.w1(32'h3c1479e9),
	.w2(32'hbbfdacd2),
	.w3(32'h3a9df035),
	.w4(32'hba1f58ef),
	.w5(32'hbbf79db5),
	.w6(32'hbb1e9c5d),
	.w7(32'hbc2ff568),
	.w8(32'hbb920811),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dad2e),
	.w1(32'hbb7bf05a),
	.w2(32'h3bbe5366),
	.w3(32'hbbe7f8bc),
	.w4(32'hba455938),
	.w5(32'h3c2b5bb5),
	.w6(32'hbc21c99d),
	.w7(32'h3b99d35a),
	.w8(32'h3bd84e6c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badc404),
	.w1(32'h3b16ef9e),
	.w2(32'hbba0e4ec),
	.w3(32'h3be2d9a3),
	.w4(32'h3bc2eeca),
	.w5(32'hbb882c22),
	.w6(32'h3bf26282),
	.w7(32'h3bd7722a),
	.w8(32'h3a075fb5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2095e6),
	.w1(32'hbad1a2a2),
	.w2(32'hbc13d0db),
	.w3(32'hbbbd33a9),
	.w4(32'h3b9e63f2),
	.w5(32'hbb8184ad),
	.w6(32'hba39d93c),
	.w7(32'hbbc51354),
	.w8(32'h3b8d4eaa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1d672),
	.w1(32'hba894469),
	.w2(32'hbbb58ba6),
	.w3(32'h3b48fabd),
	.w4(32'h3b5db581),
	.w5(32'hbc9b4876),
	.w6(32'hbba4dc40),
	.w7(32'hba799e09),
	.w8(32'hbc0d380b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc205a4e),
	.w1(32'hb78499fe),
	.w2(32'hbd8c6cae),
	.w3(32'hbc6b3d36),
	.w4(32'h39cbdd2b),
	.w5(32'hbdbc0aa9),
	.w6(32'hbc0d73fc),
	.w7(32'hba3e1e4e),
	.w8(32'hbd436a9a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72364a),
	.w1(32'h3d183b9a),
	.w2(32'hbbadb081),
	.w3(32'h3cbc3910),
	.w4(32'h3de678cc),
	.w5(32'h3a342ed7),
	.w6(32'h3cdb942e),
	.w7(32'h3d9d2058),
	.w8(32'hba7d42ae),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38ee73),
	.w1(32'h3b76973c),
	.w2(32'hbb8641ff),
	.w3(32'h3b6506f1),
	.w4(32'h3acb15b3),
	.w5(32'h3a511c6c),
	.w6(32'h3bc3e4f6),
	.w7(32'hbbe5b673),
	.w8(32'hbb34e1d3),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab420c7),
	.w1(32'h3b6fd624),
	.w2(32'h3bb4f21a),
	.w3(32'h3bbe4cb0),
	.w4(32'hbb2a750c),
	.w5(32'h3c26ec19),
	.w6(32'hbbae41e0),
	.w7(32'hbb0ac560),
	.w8(32'h3c260c61),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e78718),
	.w1(32'h3a3a7b01),
	.w2(32'h3d0b98cc),
	.w3(32'h3bdcdd21),
	.w4(32'hb9ff1716),
	.w5(32'h3d82f6a5),
	.w6(32'hb9db2567),
	.w7(32'h399c9b7b),
	.w8(32'h3d072998),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0edde2),
	.w1(32'hbce5f69f),
	.w2(32'hb9ae26c8),
	.w3(32'hbb12ece5),
	.w4(32'hbd819bf6),
	.w5(32'h3b3f9c02),
	.w6(32'hbc34883d),
	.w7(32'hbd297b3b),
	.w8(32'h39972aad),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb748e80),
	.w1(32'hba98166d),
	.w2(32'hbcc2a8cb),
	.w3(32'hbb98dd93),
	.w4(32'h3b888bfd),
	.w5(32'hbccf7833),
	.w6(32'hba6b052a),
	.w7(32'h3beacc73),
	.w8(32'hbc81aac0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4b82f),
	.w1(32'h3ccdafc2),
	.w2(32'hb8266cb0),
	.w3(32'h3c8e1525),
	.w4(32'h3d5cbd21),
	.w5(32'hb885dded),
	.w6(32'h3c94f2f5),
	.w7(32'h3d2d23f7),
	.w8(32'hbab59650),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ff21),
	.w1(32'hbb05554e),
	.w2(32'hbbcc8242),
	.w3(32'hbbc3e478),
	.w4(32'h3b95ecb9),
	.w5(32'hbbb18605),
	.w6(32'h39ae5d6f),
	.w7(32'h3afb2aa3),
	.w8(32'h3b7fb28d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49e15c),
	.w1(32'h3b6b798d),
	.w2(32'h3b287f95),
	.w3(32'hbc11101f),
	.w4(32'hbb24b923),
	.w5(32'hbac8d2ef),
	.w6(32'h3c08cbe0),
	.w7(32'h3bd9244a),
	.w8(32'h3959e2dd),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ea738c),
	.w1(32'h3c0d640c),
	.w2(32'h3c875298),
	.w3(32'hbc103ede),
	.w4(32'hbb6cbd0f),
	.w5(32'h3d102a6e),
	.w6(32'hbc5d6d5a),
	.w7(32'hbbd08815),
	.w8(32'h3ca6d439),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39356382),
	.w1(32'hbc5d2283),
	.w2(32'hbab87d7d),
	.w3(32'h3ac44247),
	.w4(32'hbd07834e),
	.w5(32'h3a92a154),
	.w6(32'hbb065f54),
	.w7(32'hbca6d73b),
	.w8(32'h3c01c4c2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b031fea),
	.w1(32'h3c89526d),
	.w2(32'hba3cc416),
	.w3(32'hbb66879e),
	.w4(32'h3c151cc3),
	.w5(32'hba709d9a),
	.w6(32'hbba2f067),
	.w7(32'h3a9ed460),
	.w8(32'hbb8fd857),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9b8f5),
	.w1(32'hb7c8172e),
	.w2(32'h3bc52fe4),
	.w3(32'hbb9981d8),
	.w4(32'h3b970b6f),
	.w5(32'h3ba1fb40),
	.w6(32'hba4716dd),
	.w7(32'hbabe05a5),
	.w8(32'h3bfce827),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0526d7),
	.w1(32'hbbf02f7b),
	.w2(32'hb992b0fa),
	.w3(32'hbb184779),
	.w4(32'hbbb8bd3d),
	.w5(32'hbc1734fc),
	.w6(32'h3bc96ad7),
	.w7(32'h3a14ce17),
	.w8(32'hbc262458),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdacd83),
	.w1(32'hba5e93bf),
	.w2(32'hba68b2e4),
	.w3(32'hbc9e7003),
	.w4(32'hba4ab8f2),
	.w5(32'h3b885bf6),
	.w6(32'hbc7105ac),
	.w7(32'hbb308c89),
	.w8(32'h3b8cb50a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ae55f),
	.w1(32'hbab925ce),
	.w2(32'h3a29cf03),
	.w3(32'h397ca1db),
	.w4(32'h3ad2c9c5),
	.w5(32'h3c0910bc),
	.w6(32'h3b4f8747),
	.w7(32'hbb134d2c),
	.w8(32'h3c45d170),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b420561),
	.w1(32'hbb827a2c),
	.w2(32'h3ca0a556),
	.w3(32'h3981b93b),
	.w4(32'hbbeaa041),
	.w5(32'h3d7dded4),
	.w6(32'hbb115149),
	.w7(32'hbb9aa187),
	.w8(32'h3caf3660),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1d564),
	.w1(32'hbca0176a),
	.w2(32'hbab5cb23),
	.w3(32'h3b2922a4),
	.w4(32'hbd595565),
	.w5(32'h3ae6e869),
	.w6(32'hbc2a8918),
	.w7(32'hbd1d814b),
	.w8(32'hbb268f20),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05940b),
	.w1(32'hbb7c8dc4),
	.w2(32'hbb4be21e),
	.w3(32'hbbdcb8e1),
	.w4(32'h3a8afcf9),
	.w5(32'h3b9e766c),
	.w6(32'hba85a9cd),
	.w7(32'hbaa12668),
	.w8(32'h3b169f28),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadeea3c),
	.w1(32'hbb6dca56),
	.w2(32'h3b9bfa71),
	.w3(32'hbb868fc2),
	.w4(32'hbc11080f),
	.w5(32'hbb8ddfe3),
	.w6(32'h3b085547),
	.w7(32'hba0d4f90),
	.w8(32'h3bcc2728),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16274c),
	.w1(32'hbc25619c),
	.w2(32'h3b475dc3),
	.w3(32'hbbd13b43),
	.w4(32'hbbfd04a0),
	.w5(32'h3b8b077b),
	.w6(32'hbb6bcda6),
	.w7(32'hbb6ad2b2),
	.w8(32'hbb19d408),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3e9fa),
	.w1(32'h39c2b19c),
	.w2(32'hbac98be8),
	.w3(32'hbbf08b6b),
	.w4(32'hba7ce686),
	.w5(32'h3bd2da33),
	.w6(32'hbb7379ca),
	.w7(32'hbb99727a),
	.w8(32'hba1b956d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cdd2c),
	.w1(32'h398905ff),
	.w2(32'h3949b147),
	.w3(32'hbb84fda6),
	.w4(32'hbb9ca1a4),
	.w5(32'h3c0494cc),
	.w6(32'hbc751282),
	.w7(32'hbc1ca064),
	.w8(32'h3a81533e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9027c1b),
	.w1(32'hbbad27f7),
	.w2(32'h3c6c9bc4),
	.w3(32'h3b74ba5f),
	.w4(32'hbb241785),
	.w5(32'h3c9f11b4),
	.w6(32'h3bcc49e1),
	.w7(32'h3ba04899),
	.w8(32'h3c5042b2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca35100),
	.w1(32'h3c86ac3a),
	.w2(32'hbbc2459f),
	.w3(32'h3c9190d7),
	.w4(32'h3c83c568),
	.w5(32'hbb252070),
	.w6(32'h3c3382f7),
	.w7(32'h3c0e4d6a),
	.w8(32'h3bfa0994),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc42a9f),
	.w1(32'h3bbb032a),
	.w2(32'hbbdeb6f1),
	.w3(32'h3a4849e5),
	.w4(32'hba5aa0f0),
	.w5(32'hbb5f6adf),
	.w6(32'hbabfc094),
	.w7(32'h3bb1c8af),
	.w8(32'h3c5b9cd9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f6e70),
	.w1(32'hbb1559e5),
	.w2(32'hbc03b8e5),
	.w3(32'hbac788db),
	.w4(32'h3b1ee9ae),
	.w5(32'hbbe8ae74),
	.w6(32'h3c360f05),
	.w7(32'hba0a9259),
	.w8(32'hbbd28f4a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e5276),
	.w1(32'hbb12ed66),
	.w2(32'h395aacbd),
	.w3(32'hbb9d96ec),
	.w4(32'hba18bc90),
	.w5(32'h3bce86d1),
	.w6(32'hbc12e4b4),
	.w7(32'hbb8f5764),
	.w8(32'h3b75e505),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4c135),
	.w1(32'hbbdf3ccb),
	.w2(32'hbb7e68f9),
	.w3(32'h3b629cdd),
	.w4(32'hba2c67fb),
	.w5(32'h3ba341a1),
	.w6(32'h3bba9ab9),
	.w7(32'hbc23800e),
	.w8(32'h3bf16c75),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d692),
	.w1(32'hbb0ac500),
	.w2(32'hbb1826d5),
	.w3(32'h3c988be9),
	.w4(32'h3bf33a5c),
	.w5(32'hbb88d831),
	.w6(32'h3ca55d1a),
	.w7(32'h3c40f2e9),
	.w8(32'hb9a6bb15),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac962),
	.w1(32'hb9bbe4ae),
	.w2(32'hbcd984d2),
	.w3(32'hbbf20057),
	.w4(32'h3b81f3d6),
	.w5(32'hbb97e2e1),
	.w6(32'h3bdb9b6c),
	.w7(32'h3c3c1538),
	.w8(32'hbc1ccafc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c6a86),
	.w1(32'hbc10a64e),
	.w2(32'hbbdebf4e),
	.w3(32'h3c00fb94),
	.w4(32'h3bba6236),
	.w5(32'hbb44bb1e),
	.w6(32'hb8d76225),
	.w7(32'hba626896),
	.w8(32'h3ae39159),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc014c7d),
	.w1(32'hbab29844),
	.w2(32'hbc247786),
	.w3(32'hbb3ce10d),
	.w4(32'hbbcd391a),
	.w5(32'hb9bdbcd4),
	.w6(32'hbb96920e),
	.w7(32'hbbe39a70),
	.w8(32'hbba4d028),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5af01a),
	.w1(32'h3ba976da),
	.w2(32'h38b4daca),
	.w3(32'h3b94a0fd),
	.w4(32'h3bd4998a),
	.w5(32'h3aaf9dc5),
	.w6(32'h3b755dba),
	.w7(32'h3bf2e808),
	.w8(32'h3c0c8281),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28920a),
	.w1(32'hbb0f3d9f),
	.w2(32'hbc6a928b),
	.w3(32'h3b8d40ed),
	.w4(32'hbbb4cd40),
	.w5(32'hbb8f8eae),
	.w6(32'h3bacfc09),
	.w7(32'hbb3a30ef),
	.w8(32'h3aca5553),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e9a8b),
	.w1(32'hbbe0ba5e),
	.w2(32'hbaf59dd3),
	.w3(32'hbb2bbc4f),
	.w4(32'hbb3214cd),
	.w5(32'h3bcb15ec),
	.w6(32'h3babc910),
	.w7(32'hba61e58e),
	.w8(32'h398fb05e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9376d4a),
	.w1(32'h3a3b8af0),
	.w2(32'hbc8d4571),
	.w3(32'h3c38d72e),
	.w4(32'h3bb94dba),
	.w5(32'hbcdcade5),
	.w6(32'h3b4aeb7a),
	.w7(32'h3bd54598),
	.w8(32'hbca6d25c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5ef34),
	.w1(32'hbca184d1),
	.w2(32'h38ab7216),
	.w3(32'hbd40e87c),
	.w4(32'hbd15a03a),
	.w5(32'h3bc2eec2),
	.w6(32'hbd15bfd6),
	.w7(32'hbcd2d2ae),
	.w8(32'h3c172493),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5e031),
	.w1(32'hbad6c867),
	.w2(32'h3b6bebf3),
	.w3(32'h3bdd3f0d),
	.w4(32'hba55df2f),
	.w5(32'h3b075759),
	.w6(32'h3b9faed5),
	.w7(32'h3b611a63),
	.w8(32'h3bcf1771),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3698a3),
	.w1(32'hbb23a2a2),
	.w2(32'h3b1df058),
	.w3(32'hbc410a90),
	.w4(32'hbc37434d),
	.w5(32'h3be0645b),
	.w6(32'hbc1d3bad),
	.w7(32'hbb176811),
	.w8(32'h3be9a9b4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e6dd7),
	.w1(32'h3b498972),
	.w2(32'hb99d7d35),
	.w3(32'h3be23208),
	.w4(32'h3b71e071),
	.w5(32'h3be0fa4c),
	.w6(32'h3c0740c5),
	.w7(32'h3b8d6655),
	.w8(32'h3bce3e39),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eb0f4),
	.w1(32'hbbda7a3f),
	.w2(32'hbca21dad),
	.w3(32'h3bc38872),
	.w4(32'h3ba6cc14),
	.w5(32'hbb799c3a),
	.w6(32'h3be6b2c4),
	.w7(32'hbbf15015),
	.w8(32'hbb83333b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b7896),
	.w1(32'hbc99c124),
	.w2(32'h3c2947f4),
	.w3(32'h3c423cb1),
	.w4(32'h3a14a882),
	.w5(32'h3bb7fd2e),
	.w6(32'h3c3d678a),
	.w7(32'h3afc4b05),
	.w8(32'h3c0692ab),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b540e0f),
	.w1(32'h3b7da82d),
	.w2(32'hbbf18527),
	.w3(32'hbb63117a),
	.w4(32'h3c008241),
	.w5(32'hb93cfb18),
	.w6(32'hba84bf48),
	.w7(32'hbb6c4842),
	.w8(32'hbb642349),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3b68),
	.w1(32'h3bd8afde),
	.w2(32'hbbcf358b),
	.w3(32'h3b87d1c2),
	.w4(32'hbb713d54),
	.w5(32'h39d9f4e8),
	.w6(32'h3b4f52a0),
	.w7(32'hbabf8f9f),
	.w8(32'hbae2c813),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b159fad),
	.w1(32'hbb893116),
	.w2(32'hb9a4d993),
	.w3(32'h3bb1b329),
	.w4(32'h3c35c483),
	.w5(32'h3a4ebe5f),
	.w6(32'h3bc81f7f),
	.w7(32'h3bc0b2b9),
	.w8(32'h3c1f2108),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803324),
	.w1(32'hbb1f333a),
	.w2(32'h39be5f43),
	.w3(32'h3b682913),
	.w4(32'h3b9cfcb7),
	.w5(32'hb51ea2e7),
	.w6(32'h3be3e1e0),
	.w7(32'hbaf840c5),
	.w8(32'hbb9302cd),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f7c0c),
	.w1(32'h3b22fd77),
	.w2(32'h3bebe343),
	.w3(32'hbabd9b85),
	.w4(32'hba39017a),
	.w5(32'h3c246105),
	.w6(32'h38440951),
	.w7(32'hbb3d89aa),
	.w8(32'h3a0a2ca0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b548968),
	.w1(32'h3a68bfbe),
	.w2(32'hbb9968fc),
	.w3(32'h3b08e0df),
	.w4(32'h39c88035),
	.w5(32'h3b792edd),
	.w6(32'h3bfdd98a),
	.w7(32'h3b568b9d),
	.w8(32'h3b3c2fe7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35aac7),
	.w1(32'hb9cbabe5),
	.w2(32'h3b933f60),
	.w3(32'h3c0bf7b1),
	.w4(32'h3b345008),
	.w5(32'h3c02d3db),
	.w6(32'h3c05cb8d),
	.w7(32'h3ba8b890),
	.w8(32'h3c48aa6f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9913ba),
	.w1(32'h39d2d295),
	.w2(32'hbc26f094),
	.w3(32'hbb37265c),
	.w4(32'hb91bcf80),
	.w5(32'hbb003888),
	.w6(32'h3b41999f),
	.w7(32'hbb9d02a6),
	.w8(32'h3ad79a46),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a1806),
	.w1(32'hbbb2669c),
	.w2(32'h3b24c4b8),
	.w3(32'h3c033836),
	.w4(32'hbb25582d),
	.w5(32'h3af72f2d),
	.w6(32'h3c062f5c),
	.w7(32'hbb882039),
	.w8(32'h3c147d6c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb68a7),
	.w1(32'h3b2c7138),
	.w2(32'hbc15f285),
	.w3(32'hbbf4eb21),
	.w4(32'hbbfbad5a),
	.w5(32'hbab1dc2b),
	.w6(32'hba923429),
	.w7(32'hbbf79b67),
	.w8(32'h3b04ec0a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8766c9),
	.w1(32'hbba8d0c3),
	.w2(32'hb9e82cf0),
	.w3(32'h3b8eea5f),
	.w4(32'h3a6ed030),
	.w5(32'h3be29c25),
	.w6(32'h3b2021d2),
	.w7(32'hbb04041a),
	.w8(32'h3c3b6038),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8c9e5),
	.w1(32'h3b9505b0),
	.w2(32'h3a984ffe),
	.w3(32'h3c08a499),
	.w4(32'h3bed555f),
	.w5(32'hb9ca3ac0),
	.w6(32'h3c2fd23d),
	.w7(32'h3bcc0d38),
	.w8(32'h3a8220c3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba600d4e),
	.w1(32'hba02becd),
	.w2(32'hbaf48351),
	.w3(32'h3b0c23cc),
	.w4(32'h3b05e632),
	.w5(32'hbbc1a146),
	.w6(32'h3aaea6e2),
	.w7(32'hbb1d17ae),
	.w8(32'hbbffd759),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2e4dd),
	.w1(32'hbb633115),
	.w2(32'hbaa42ba5),
	.w3(32'hbbae9e36),
	.w4(32'hbba46b3a),
	.w5(32'hbb47d11c),
	.w6(32'hbc06b236),
	.w7(32'hbbba804a),
	.w8(32'h3b0f9ae7),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b538b),
	.w1(32'hba9728d3),
	.w2(32'hbb07b54a),
	.w3(32'hbb4fa678),
	.w4(32'hbbce3eea),
	.w5(32'h3b6f5682),
	.w6(32'h3baa8739),
	.w7(32'h3b32b711),
	.w8(32'h3b91a4bb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc85a8f),
	.w1(32'hbb5df109),
	.w2(32'h3b29c57b),
	.w3(32'h3ba427c4),
	.w4(32'h3c089e04),
	.w5(32'h3bfc9a68),
	.w6(32'h3b43b069),
	.w7(32'hbabfab8f),
	.w8(32'h3c86e89b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9feef),
	.w1(32'hbbffb957),
	.w2(32'hbcdcc2c7),
	.w3(32'h3b4e3dab),
	.w4(32'hbb846945),
	.w5(32'hbd635593),
	.w6(32'h3c38cb97),
	.w7(32'h3b4305f9),
	.w8(32'hbd399a44),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd492a26),
	.w1(32'hbcc94cb5),
	.w2(32'hbb61c247),
	.w3(32'hbdd0a4d5),
	.w4(32'hbd818821),
	.w5(32'hbb8a2259),
	.w6(32'hbdb1e547),
	.w7(32'hbd58bba2),
	.w8(32'h3813d835),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09e49f),
	.w1(32'h3c114831),
	.w2(32'h3ba19c37),
	.w3(32'h3be75b6e),
	.w4(32'hbb0a92b2),
	.w5(32'h3b804e4c),
	.w6(32'h3b82701b),
	.w7(32'h3c194552),
	.w8(32'hbacc0c14),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6aebe),
	.w1(32'hba600d70),
	.w2(32'h3bc2e4f8),
	.w3(32'h38fa59af),
	.w4(32'h3a88c868),
	.w5(32'h3ba4b551),
	.w6(32'hbb4123a2),
	.w7(32'hbb6d9109),
	.w8(32'h3bddeae7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd94419),
	.w1(32'h3b9bf21d),
	.w2(32'hbbfea6c9),
	.w3(32'h3b027767),
	.w4(32'h3b0042e0),
	.w5(32'hbaea8e7c),
	.w6(32'h3b539788),
	.w7(32'h3b999e17),
	.w8(32'h3a5b8e23),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa36e3c),
	.w1(32'hbb0463c1),
	.w2(32'hbba29757),
	.w3(32'h3987dc24),
	.w4(32'h3b8042a5),
	.w5(32'hbbcfac29),
	.w6(32'h3bbd71a2),
	.w7(32'h3baaa58e),
	.w8(32'hbc0cfee0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53a741),
	.w1(32'hbaa7236d),
	.w2(32'hbb6c25da),
	.w3(32'hbba1525a),
	.w4(32'hbbd9a8ff),
	.w5(32'hbb0a41a0),
	.w6(32'hbba2738f),
	.w7(32'hbbd5a0ad),
	.w8(32'h3b8a3147),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74d2d1),
	.w1(32'hbb7e065c),
	.w2(32'hb7a7a565),
	.w3(32'hba7936c8),
	.w4(32'hbb35b779),
	.w5(32'h3b08e040),
	.w6(32'hbad51e1e),
	.w7(32'h3b803667),
	.w8(32'h3b1df311),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc43b3c),
	.w1(32'h387de088),
	.w2(32'hbbfc1b30),
	.w3(32'h3c5f5815),
	.w4(32'h3c14591a),
	.w5(32'h3c91bdd1),
	.w6(32'h3b95e299),
	.w7(32'hbb3d190e),
	.w8(32'h3bf2b78d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd76327),
	.w1(32'hbafe8447),
	.w2(32'hbb5db19e),
	.w3(32'h3d66582b),
	.w4(32'h3cd66e9d),
	.w5(32'hbb73259e),
	.w6(32'h3d389578),
	.w7(32'h3c9aa8db),
	.w8(32'hbbf13f46),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2d1e1),
	.w1(32'hbb709caa),
	.w2(32'hbb47397a),
	.w3(32'hbaa911eb),
	.w4(32'hbbac8dd3),
	.w5(32'h3bbf924b),
	.w6(32'hbbc10cb7),
	.w7(32'hbc0f11b1),
	.w8(32'h3b864d07),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c815a),
	.w1(32'hba107fda),
	.w2(32'hbb76adf6),
	.w3(32'h3c08ad87),
	.w4(32'h3c1ba4c4),
	.w5(32'h3a88965e),
	.w6(32'h3b998ba6),
	.w7(32'hbb76c45a),
	.w8(32'hbb6b35b1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1366fc),
	.w1(32'hbaf4f73e),
	.w2(32'h3b212e0c),
	.w3(32'hb832c0a8),
	.w4(32'h3a94d399),
	.w5(32'h3b41cace),
	.w6(32'h3b367aad),
	.w7(32'hbb9754d1),
	.w8(32'h3c1aad93),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde68c4),
	.w1(32'h39eeee9c),
	.w2(32'h3b3c2b03),
	.w3(32'h3b992d40),
	.w4(32'hbb2ebafd),
	.w5(32'h3c0091e0),
	.w6(32'h3b8d4b31),
	.w7(32'h3a62b3f8),
	.w8(32'hbbe7de41),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0dae1),
	.w1(32'hbac4e1a2),
	.w2(32'h3b55cc8e),
	.w3(32'hbc39ceae),
	.w4(32'hbb015c31),
	.w5(32'h3a7f9414),
	.w6(32'hbc449f46),
	.w7(32'hbc2ea8ec),
	.w8(32'h3989f46d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcde1cf),
	.w1(32'h3bb77163),
	.w2(32'h3b90a150),
	.w3(32'h3b7fb25b),
	.w4(32'h3c03222e),
	.w5(32'hbbbc5f23),
	.w6(32'h3b9e348c),
	.w7(32'h3c1eb7ba),
	.w8(32'hbc97a717),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9afbcf),
	.w1(32'h39af8b59),
	.w2(32'hbb640f1e),
	.w3(32'hbd07281c),
	.w4(32'hbcca5a38),
	.w5(32'hbbea72a7),
	.w6(32'hbd28def7),
	.w7(32'hbd00313d),
	.w8(32'hbbacd62b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcda9b3),
	.w1(32'hb9c41504),
	.w2(32'hbb84fd8a),
	.w3(32'hbc02bea2),
	.w4(32'hbb96ff68),
	.w5(32'hbb1cbe2a),
	.w6(32'hbb922b57),
	.w7(32'h3a3f5590),
	.w8(32'hbb429b13),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea31db),
	.w1(32'h3c1cd41f),
	.w2(32'h3b0e048e),
	.w3(32'h3b0579b7),
	.w4(32'h3bf16ed2),
	.w5(32'hb9650e7c),
	.w6(32'h3b0e188e),
	.w7(32'h3becdcaa),
	.w8(32'h3a4e021e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93b610),
	.w1(32'h3b7d7b7c),
	.w2(32'hbadab2f3),
	.w3(32'h3b90f699),
	.w4(32'h3b558fe9),
	.w5(32'h3bc8564e),
	.w6(32'h3bd048a0),
	.w7(32'h3c04f9c1),
	.w8(32'h3bb0455d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16e4b3),
	.w1(32'hbc2ba86c),
	.w2(32'h3bdc944b),
	.w3(32'hbc0153e0),
	.w4(32'hbc6c7d59),
	.w5(32'h3c085178),
	.w6(32'h39a7ea13),
	.w7(32'hbb6e699f),
	.w8(32'h3c1c242e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89f809),
	.w1(32'hbab2b462),
	.w2(32'hbbc913fe),
	.w3(32'hbb0ba1fd),
	.w4(32'hbb9b5c1b),
	.w5(32'hbc3d9e8f),
	.w6(32'hbb59f77c),
	.w7(32'hbbd94e6c),
	.w8(32'hbc2e7e61),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc233f1a),
	.w1(32'hbbe1e634),
	.w2(32'hbada5cb6),
	.w3(32'hbc869cfa),
	.w4(32'hbc6660bc),
	.w5(32'h3bed920e),
	.w6(32'hbc819987),
	.w7(32'hbc648273),
	.w8(32'hbab39147),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b8fa),
	.w1(32'h3a8110b0),
	.w2(32'h3a59bfd1),
	.w3(32'h3b9db1cb),
	.w4(32'h3b0b1c78),
	.w5(32'h3bb6c375),
	.w6(32'h3bfa2609),
	.w7(32'hba216637),
	.w8(32'h3aa5fe01),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09811b),
	.w1(32'h3b5f826e),
	.w2(32'hbc64e87f),
	.w3(32'h3b3555bf),
	.w4(32'hbb57d972),
	.w5(32'hbc0549a6),
	.w6(32'h38d845d1),
	.w7(32'hbbed06ed),
	.w8(32'h3b92b984),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86ec5a),
	.w1(32'hbc96b016),
	.w2(32'hbac4b2d7),
	.w3(32'hbc170161),
	.w4(32'hbc1be26f),
	.w5(32'h3b94180d),
	.w6(32'h3c0b4919),
	.w7(32'h3b58012f),
	.w8(32'h3c10c5b1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70072d),
	.w1(32'h39993630),
	.w2(32'hbb140662),
	.w3(32'h3b6120b7),
	.w4(32'hbb11d484),
	.w5(32'hbb84afc0),
	.w6(32'h3bf097b8),
	.w7(32'hb941fa5a),
	.w8(32'hbb4a5615),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc078e82),
	.w1(32'hbbf752e6),
	.w2(32'hbba1d5bd),
	.w3(32'hbc514386),
	.w4(32'hbc37879c),
	.w5(32'hbc5f819a),
	.w6(32'hbc14ce61),
	.w7(32'hbc184074),
	.w8(32'hbc1e5326),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0625d5),
	.w1(32'hbb1392ef),
	.w2(32'hbb5c2498),
	.w3(32'hbd04fa83),
	.w4(32'hbc989993),
	.w5(32'h3b133902),
	.w6(32'hbcd3d1fd),
	.w7(32'hbc70f02b),
	.w8(32'h39d2428a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b612ba5),
	.w1(32'h3b239d39),
	.w2(32'hba6086f2),
	.w3(32'hb9370ac6),
	.w4(32'h3b0b934b),
	.w5(32'hba39f820),
	.w6(32'h3abd0b14),
	.w7(32'hbacd6154),
	.w8(32'h39a5d580),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86684c),
	.w1(32'hbb3a0923),
	.w2(32'h3bd041c8),
	.w3(32'h3c45b904),
	.w4(32'hbb28854a),
	.w5(32'h3bfa6874),
	.w6(32'h3b865247),
	.w7(32'hbb37b657),
	.w8(32'hbb7fc224),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffdc1a),
	.w1(32'hbaa3eb34),
	.w2(32'h3b95074c),
	.w3(32'h3be26ae7),
	.w4(32'h3b060821),
	.w5(32'h3b067dba),
	.w6(32'hbae2f473),
	.w7(32'hbb3712bd),
	.w8(32'hba50a4cf),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb1bad),
	.w1(32'h3b4c3449),
	.w2(32'hbb87d799),
	.w3(32'h3c08f06b),
	.w4(32'h3bdc5b95),
	.w5(32'hbb16969a),
	.w6(32'hb70a941b),
	.w7(32'hbac986fc),
	.w8(32'hbb02ed39),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93c89c),
	.w1(32'h3b5769fb),
	.w2(32'hbc947f73),
	.w3(32'h3bd5c797),
	.w4(32'h3b709efb),
	.w5(32'hbc9ae423),
	.w6(32'h3b97a779),
	.w7(32'h398b1801),
	.w8(32'hbcc4fcf6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07c17e),
	.w1(32'h3c01be80),
	.w2(32'hbba6b122),
	.w3(32'hbb3073f9),
	.w4(32'h3c23c9e5),
	.w5(32'h3b6b4d06),
	.w6(32'hbbedd069),
	.w7(32'h3bb386de),
	.w8(32'hba89fa24),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55b7e1),
	.w1(32'hbb1e5cd1),
	.w2(32'hbc22bb5f),
	.w3(32'h3c0208ae),
	.w4(32'h3bce049e),
	.w5(32'hbbee4f20),
	.w6(32'h3a921d71),
	.w7(32'h3b27eaff),
	.w8(32'hba014a51),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf88072),
	.w1(32'hbbe41f74),
	.w2(32'hbb06d14c),
	.w3(32'hb980d4e2),
	.w4(32'h3b307ac5),
	.w5(32'h3b9df89c),
	.w6(32'h3b230e8c),
	.w7(32'h3b5ca369),
	.w8(32'h3b085114),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a692c36),
	.w1(32'h3c041967),
	.w2(32'h39a5fddf),
	.w3(32'h3be5a31d),
	.w4(32'h3c4cb2a5),
	.w5(32'h3b265f5e),
	.w6(32'h3b608c43),
	.w7(32'h3c1b85ac),
	.w8(32'h3be08912),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfd881),
	.w1(32'h3bd816c7),
	.w2(32'hbb90e09a),
	.w3(32'h3c3bc69f),
	.w4(32'h3c40d450),
	.w5(32'h3a60c441),
	.w6(32'h3c71940c),
	.w7(32'h3c8ee9c2),
	.w8(32'h37ebbe1a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91719d),
	.w1(32'hbb9dadcc),
	.w2(32'hb992d391),
	.w3(32'h3b99875b),
	.w4(32'hba99dccc),
	.w5(32'h3b211c1b),
	.w6(32'h3a847041),
	.w7(32'h3bb9a6e4),
	.w8(32'h3b3d9a61),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71e94e),
	.w1(32'h3b991398),
	.w2(32'h3b51784c),
	.w3(32'h3c179aef),
	.w4(32'h3c019484),
	.w5(32'h3baaa2ef),
	.w6(32'h3c576e46),
	.w7(32'h3c1e143b),
	.w8(32'h3bfea86d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1187ed),
	.w1(32'hbba888a4),
	.w2(32'hbb72935a),
	.w3(32'h3ac52d84),
	.w4(32'hbbe6eafd),
	.w5(32'h3b9c3e9e),
	.w6(32'h3a9b6b88),
	.w7(32'hbba9ed61),
	.w8(32'hba0ee93f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d6de),
	.w1(32'h3c06e619),
	.w2(32'h3b8323ab),
	.w3(32'h3c06ab03),
	.w4(32'h3c2b7f65),
	.w5(32'hbb26033f),
	.w6(32'h3b937fc4),
	.w7(32'h3aaaa8d5),
	.w8(32'hbb31cfb3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be639c2),
	.w1(32'h3b3886dd),
	.w2(32'hba3ffc3c),
	.w3(32'h3bab6669),
	.w4(32'h3bb93127),
	.w5(32'h3a5a58fa),
	.w6(32'h3c0d93a8),
	.w7(32'h3b823de6),
	.w8(32'hbbb9454d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54f1d2),
	.w1(32'hbb33d5e6),
	.w2(32'hbae3be02),
	.w3(32'hba2d8500),
	.w4(32'h3bd4ace8),
	.w5(32'hbb469250),
	.w6(32'hbace15bd),
	.w7(32'h3bbb6c9b),
	.w8(32'hbb80b9cf),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb464807),
	.w1(32'h3bbf7546),
	.w2(32'hbb7e6207),
	.w3(32'h3bda80c5),
	.w4(32'h3a12ee97),
	.w5(32'h3baebfb6),
	.w6(32'h3b1e64d3),
	.w7(32'h3b9cc2ea),
	.w8(32'hbb746b9c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1419c2),
	.w1(32'hbb64e6eb),
	.w2(32'h3b200b69),
	.w3(32'h3c3c1632),
	.w4(32'h3bb951b6),
	.w5(32'hb90b30ed),
	.w6(32'h3b27d89d),
	.w7(32'hba8beae6),
	.w8(32'h3afa782c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab89602),
	.w1(32'h38fcd089),
	.w2(32'hbbaa7019),
	.w3(32'h3b762d46),
	.w4(32'h3bc26500),
	.w5(32'h3b16011c),
	.w6(32'hba5c84c7),
	.w7(32'h3b43624a),
	.w8(32'hbad73d6a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2f591),
	.w1(32'h3bd4c02e),
	.w2(32'h3ad5164c),
	.w3(32'h3be11fb4),
	.w4(32'h3b644ced),
	.w5(32'h3ad040f5),
	.w6(32'h3a97e297),
	.w7(32'h3b99c1be),
	.w8(32'h3b99e85c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b856dd4),
	.w1(32'h3b89e682),
	.w2(32'h3c1a1d42),
	.w3(32'h3bae03fb),
	.w4(32'h39fc08ca),
	.w5(32'h3c01efd9),
	.w6(32'h3b4be2a4),
	.w7(32'hbaded2a0),
	.w8(32'hbbd75421),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8367fd),
	.w1(32'h3c8636c4),
	.w2(32'hbc54cc09),
	.w3(32'h3c20fe4c),
	.w4(32'h3c0b7dfc),
	.w5(32'hbbc4e5d8),
	.w6(32'hbbd20547),
	.w7(32'hbbc822a3),
	.w8(32'h3addfcaf),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe23919),
	.w1(32'hbbfb2b8d),
	.w2(32'h3bd8ed32),
	.w3(32'hbaa68b94),
	.w4(32'hbb25896c),
	.w5(32'h3b6533fd),
	.w6(32'h3bde5c7d),
	.w7(32'h3b833962),
	.w8(32'h3b9ea661),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3002a4),
	.w1(32'h3c1927e4),
	.w2(32'hb9903c32),
	.w3(32'h3b00138d),
	.w4(32'hbab3c099),
	.w5(32'h3bd9bbf5),
	.w6(32'h3a67b84b),
	.w7(32'hbb36f988),
	.w8(32'h3aa9b4d5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c467),
	.w1(32'h3a16075f),
	.w2(32'hba438039),
	.w3(32'h3c2a9dad),
	.w4(32'h3ad77c82),
	.w5(32'h3af29798),
	.w6(32'h3b9564e8),
	.w7(32'h3b62d989),
	.w8(32'h3a641d9d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba937425),
	.w1(32'hbad285a0),
	.w2(32'hbac7209c),
	.w3(32'hbb0823f9),
	.w4(32'hbb274616),
	.w5(32'hba837d9f),
	.w6(32'h3bab757f),
	.w7(32'h3b88541f),
	.w8(32'h3ab34312),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7daaf8),
	.w1(32'h3a9e4d58),
	.w2(32'h3b0b5d32),
	.w3(32'hbb4b59cc),
	.w4(32'hbb2cfd4a),
	.w5(32'h3c5e655e),
	.w6(32'hbb8a0698),
	.w7(32'h3b4dbe20),
	.w8(32'h3c6f07dc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35012e),
	.w1(32'h3c51ca20),
	.w2(32'h38bc2cb3),
	.w3(32'h3d0a321a),
	.w4(32'h3cf69310),
	.w5(32'h3bc49cd6),
	.w6(32'h3d0c76bf),
	.w7(32'h3cf417ea),
	.w8(32'h3b7aaeff),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd3a18),
	.w1(32'h3b9ddc9b),
	.w2(32'h3ade9714),
	.w3(32'h3c5d31c5),
	.w4(32'h3c1f1143),
	.w5(32'h3beb727a),
	.w6(32'h3c269c86),
	.w7(32'h3be208a9),
	.w8(32'h3bc5967c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad31cb2),
	.w1(32'h39b495ea),
	.w2(32'h3c56ea0f),
	.w3(32'h3a182a2c),
	.w4(32'hbc08f987),
	.w5(32'h3c72c241),
	.w6(32'h3b913046),
	.w7(32'h393b7b7e),
	.w8(32'h3bb8ca69),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2162ef),
	.w1(32'h39f99093),
	.w2(32'h3be478b3),
	.w3(32'h3c10128e),
	.w4(32'hbae0cac6),
	.w5(32'h38b0d7a0),
	.w6(32'hba868770),
	.w7(32'hbc167b5c),
	.w8(32'h3bae0eda),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82316b),
	.w1(32'h3b08b9a7),
	.w2(32'hba80f941),
	.w3(32'hbb9ad2ef),
	.w4(32'hbb4842ce),
	.w5(32'h38c7c626),
	.w6(32'h3b3a6534),
	.w7(32'h3b01a79f),
	.w8(32'hbb0415c3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c2a19),
	.w1(32'hbb7a6335),
	.w2(32'hbbed1ea8),
	.w3(32'h3ba2146b),
	.w4(32'hb98b4a94),
	.w5(32'hbb1fe706),
	.w6(32'h3b285b3d),
	.w7(32'hb7b1144c),
	.w8(32'h399123e4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4f3e7),
	.w1(32'hbbbc2d0b),
	.w2(32'hbc26fadc),
	.w3(32'h3b6a2167),
	.w4(32'hbb580d16),
	.w5(32'h3a96461c),
	.w6(32'h3be0f249),
	.w7(32'hbb5b22fb),
	.w8(32'hbbd25497),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule