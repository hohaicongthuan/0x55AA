module layer_8_featuremap_191(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84d89a),
	.w1(32'h3bd4f08b),
	.w2(32'hbae301fc),
	.w3(32'hb9e83f09),
	.w4(32'h3c663bbf),
	.w5(32'h3b14aceb),
	.w6(32'h3b492316),
	.w7(32'hbcb6a81c),
	.w8(32'hbc226c8f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc881be3),
	.w1(32'hb823208b),
	.w2(32'h3ba9af9e),
	.w3(32'h3ba9eedb),
	.w4(32'hba81cfef),
	.w5(32'h3bc81d32),
	.w6(32'hbba6ba24),
	.w7(32'h3a0e0380),
	.w8(32'hbb417733),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac58f8c),
	.w1(32'hbbf12f5c),
	.w2(32'h3c58b28d),
	.w3(32'h3adb6212),
	.w4(32'hbc121411),
	.w5(32'h3bbde088),
	.w6(32'hbb85652b),
	.w7(32'h3c350ec6),
	.w8(32'h3bc7ed66),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0494c5),
	.w1(32'h3b4cd5d3),
	.w2(32'h3c38678c),
	.w3(32'h3b9b241a),
	.w4(32'h3b6ed435),
	.w5(32'h3cb72a10),
	.w6(32'h3a12bd7b),
	.w7(32'hbb750fa7),
	.w8(32'hbc6b649e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab48e6),
	.w1(32'hbbaaaf24),
	.w2(32'hbb5703a4),
	.w3(32'h3ba599bb),
	.w4(32'hbbe2084f),
	.w5(32'h399afdbe),
	.w6(32'hbb98341d),
	.w7(32'hbb7c5e80),
	.w8(32'hbbf89694),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb953d48),
	.w1(32'h3c22b08c),
	.w2(32'h3ccc15d7),
	.w3(32'hbb527a0c),
	.w4(32'h3bff55f4),
	.w5(32'h3ba64fef),
	.w6(32'hbbf5c392),
	.w7(32'h3cbb62ea),
	.w8(32'hbc6a7b3d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6a132),
	.w1(32'hbb467eba),
	.w2(32'hbb922703),
	.w3(32'hbc73c11d),
	.w4(32'hbb3c8422),
	.w5(32'hbba7dfef),
	.w6(32'h3a2ba8c6),
	.w7(32'hbaefcd11),
	.w8(32'hbaca0f18),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb430807),
	.w1(32'h3ca6c4f6),
	.w2(32'h3cf971a7),
	.w3(32'hbb79e7a8),
	.w4(32'h3a613bb5),
	.w5(32'h3cc75d46),
	.w6(32'h3cd3e243),
	.w7(32'h3c73301c),
	.w8(32'hbc8d62b4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d9a5f),
	.w1(32'hbc0d17d2),
	.w2(32'h3bbb2e14),
	.w3(32'hb68f0235),
	.w4(32'hbc367ec7),
	.w5(32'h3b9d3a0a),
	.w6(32'hbc4c1500),
	.w7(32'h3aa28fd0),
	.w8(32'hbb01e32a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc3fcf),
	.w1(32'hbc3a8767),
	.w2(32'hbc2438c0),
	.w3(32'hbac057ac),
	.w4(32'h3a49139f),
	.w5(32'hbb4d5124),
	.w6(32'hbbb623e5),
	.w7(32'h3a84c7d9),
	.w8(32'h3b7c3e21),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d44c1),
	.w1(32'h3b18e489),
	.w2(32'hbc47b237),
	.w3(32'hb9f5f3d7),
	.w4(32'h3b802949),
	.w5(32'hbb94c4fc),
	.w6(32'hbc5286db),
	.w7(32'hbc79a5c1),
	.w8(32'hbc0c8954),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3981e9),
	.w1(32'hba49caf6),
	.w2(32'h3c17ccad),
	.w3(32'hbc3fe120),
	.w4(32'h3a711e6b),
	.w5(32'h3c093aae),
	.w6(32'h3a408f00),
	.w7(32'h3c351c03),
	.w8(32'hbb4e8e92),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe662b6),
	.w1(32'h3995d628),
	.w2(32'hbc22053e),
	.w3(32'hbbb14e16),
	.w4(32'h3c03fe20),
	.w5(32'hbb8759d3),
	.w6(32'hb9f4941d),
	.w7(32'hbbaa9807),
	.w8(32'hbaa12ec4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c867bd),
	.w1(32'hbc20a5ab),
	.w2(32'h3cb5af2e),
	.w3(32'h3a4c6302),
	.w4(32'hbc1293a7),
	.w5(32'h3bc568dc),
	.w6(32'h392e4e73),
	.w7(32'h3c34fa82),
	.w8(32'hbb74c907),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c892531),
	.w1(32'hbc23e4db),
	.w2(32'h3a4290ea),
	.w3(32'h3c830674),
	.w4(32'hbb865498),
	.w5(32'h399b6d6d),
	.w6(32'hbbb3bafa),
	.w7(32'h3a21ae80),
	.w8(32'h3ae625f3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b4bd0),
	.w1(32'hbbb626f0),
	.w2(32'hbd08f0c5),
	.w3(32'h3b36c335),
	.w4(32'hbb3dc6f2),
	.w5(32'hbcb9a13d),
	.w6(32'hbc3173c5),
	.w7(32'hbc20240a),
	.w8(32'h3c681658),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fe11d),
	.w1(32'hbc39270f),
	.w2(32'hbaeabf40),
	.w3(32'hbbe4adec),
	.w4(32'hbb7aebf2),
	.w5(32'h3b1d74b4),
	.w6(32'hbc7b1dd7),
	.w7(32'h3bce3b2e),
	.w8(32'h3c1da1ad),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb250f54),
	.w1(32'h3bf38087),
	.w2(32'h3bf9925e),
	.w3(32'hbc88bba3),
	.w4(32'h3b7b8079),
	.w5(32'h3b41aa08),
	.w6(32'hbad76dae),
	.w7(32'hbba6e562),
	.w8(32'h3b9c38af),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb67d4c),
	.w1(32'hbc241646),
	.w2(32'h3c66ff71),
	.w3(32'hbbf7aa94),
	.w4(32'hbc348b5f),
	.w5(32'h39d95e77),
	.w6(32'hbbb42946),
	.w7(32'h3c98a840),
	.w8(32'h3c2143b5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3463d9),
	.w1(32'hbb4f02f8),
	.w2(32'hbad88dd4),
	.w3(32'hbc175f0b),
	.w4(32'h3a55ecee),
	.w5(32'hbb35d528),
	.w6(32'hbb453731),
	.w7(32'h3a49d501),
	.w8(32'h3b85bcc7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb13d3a),
	.w1(32'hbc424d74),
	.w2(32'h3c286574),
	.w3(32'h3b201c84),
	.w4(32'hbc0cb878),
	.w5(32'hbb92bbee),
	.w6(32'hbb9f39ca),
	.w7(32'h3b578807),
	.w8(32'h3b9ffafa),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a932aa8),
	.w1(32'hbc32b7b5),
	.w2(32'hbceaf656),
	.w3(32'h3abf00b5),
	.w4(32'h3aa5c8d9),
	.w5(32'hbc89c378),
	.w6(32'hbc8f5952),
	.w7(32'hbc9f0479),
	.w8(32'hbba2b4bb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18b2cb),
	.w1(32'hbc64439a),
	.w2(32'hbc37a7e2),
	.w3(32'h3ac1bae5),
	.w4(32'hbc63f9e8),
	.w5(32'hbc79d4b3),
	.w6(32'hbc114e25),
	.w7(32'hbc57648e),
	.w8(32'h3b636538),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacbee6),
	.w1(32'hbb82d059),
	.w2(32'hbd0678f5),
	.w3(32'hba95a213),
	.w4(32'h3abf18d8),
	.w5(32'hbcb26afc),
	.w6(32'hbc6fcc0e),
	.w7(32'hbc2c4471),
	.w8(32'h3bcfd10b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f26e63),
	.w1(32'hbb3ae7b5),
	.w2(32'h3bcc494b),
	.w3(32'h3c2ec7ce),
	.w4(32'h3b115e04),
	.w5(32'h3b0364c3),
	.w6(32'hbb92f81f),
	.w7(32'h3b7eb0f2),
	.w8(32'h3b039f67),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b906b61),
	.w1(32'h3b441afb),
	.w2(32'hbb2e9608),
	.w3(32'hbb5d9fad),
	.w4(32'h3bd96537),
	.w5(32'hbc0d2563),
	.w6(32'h3b8f4566),
	.w7(32'hbc962cbb),
	.w8(32'hbc82d786),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf72d60),
	.w1(32'hbb70a4ea),
	.w2(32'h3b2cb977),
	.w3(32'hbbc9e87b),
	.w4(32'hbc3432fb),
	.w5(32'hbbfdefec),
	.w6(32'h3b8eba1e),
	.w7(32'hb907f70f),
	.w8(32'hbbe28b1f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fe17b),
	.w1(32'h3bffd693),
	.w2(32'hbc9c2f61),
	.w3(32'h3c00a8b5),
	.w4(32'h3bbd0e86),
	.w5(32'hbc8090a5),
	.w6(32'hbbd675b2),
	.w7(32'hbc98d593),
	.w8(32'hbb528c0b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdca40),
	.w1(32'h38f28a33),
	.w2(32'hb9a1436a),
	.w3(32'hbc53ca17),
	.w4(32'hba9c1457),
	.w5(32'hbb0a4166),
	.w6(32'hbbceb3e1),
	.w7(32'hbb1eb54b),
	.w8(32'hbb7d4706),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e226a),
	.w1(32'hba9103e4),
	.w2(32'hbb5604e0),
	.w3(32'hbaa8bddd),
	.w4(32'hbb857386),
	.w5(32'h3b9b234d),
	.w6(32'hbaf14389),
	.w7(32'hbab7a275),
	.w8(32'hba5a3631),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e956fb),
	.w1(32'hbbc7e61d),
	.w2(32'h3bc57f1f),
	.w3(32'h3b8f64e9),
	.w4(32'hbb9acedc),
	.w5(32'h3b56eda3),
	.w6(32'hbb9f520c),
	.w7(32'hba809b60),
	.w8(32'hbaf4a484),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba36504),
	.w1(32'hbb2462c8),
	.w2(32'h3c20083d),
	.w3(32'h3b50a7ef),
	.w4(32'hbb2ad560),
	.w5(32'h3b97434a),
	.w6(32'hbb7636f7),
	.w7(32'h3c1dd465),
	.w8(32'h3b341bfe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8e36d),
	.w1(32'hbba6e075),
	.w2(32'h39961620),
	.w3(32'h3b915a7f),
	.w4(32'h39cdf30f),
	.w5(32'hbb8f7701),
	.w6(32'hbc2f3902),
	.w7(32'hbab362d9),
	.w8(32'h3b96eb93),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98df60),
	.w1(32'h3c5529c4),
	.w2(32'h3c9db05a),
	.w3(32'hbba48d25),
	.w4(32'hbbc7a675),
	.w5(32'h3a7c8875),
	.w6(32'h3b93888c),
	.w7(32'h3a1ee917),
	.w8(32'hbbf47ed3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb284409),
	.w1(32'h3b24a308),
	.w2(32'hbbee8e7a),
	.w3(32'hba9e9845),
	.w4(32'h3b9c9330),
	.w5(32'hbbc2d396),
	.w6(32'h3b04def0),
	.w7(32'hbc151232),
	.w8(32'h3ba92646),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30dac4),
	.w1(32'hbc8b857d),
	.w2(32'h3b97165c),
	.w3(32'h3af293f7),
	.w4(32'hbca3a13f),
	.w5(32'hbc87157c),
	.w6(32'hbbd22ac9),
	.w7(32'h3be382e8),
	.w8(32'h3c1b0275),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbbd91),
	.w1(32'hbba6842c),
	.w2(32'hbbcc8044),
	.w3(32'h3bf3ffbb),
	.w4(32'hbb33b8fc),
	.w5(32'hbbf89e24),
	.w6(32'hbbb4451a),
	.w7(32'hbb8dec2b),
	.w8(32'hbad25c34),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9645e40),
	.w1(32'hbb86dff2),
	.w2(32'h3b661765),
	.w3(32'hbb2af27d),
	.w4(32'h3b0a87ed),
	.w5(32'h3c00c8d9),
	.w6(32'hbbcc0fbd),
	.w7(32'hbb3491e2),
	.w8(32'h3ad7867c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52804),
	.w1(32'h3b6b9a3b),
	.w2(32'hba8a6f41),
	.w3(32'h3c19e619),
	.w4(32'h3c5d5870),
	.w5(32'hbab14300),
	.w6(32'hbaaafda2),
	.w7(32'hb80dec5e),
	.w8(32'hbc72e0c0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92c7c9),
	.w1(32'hbb88e496),
	.w2(32'hbc38146b),
	.w3(32'hbb7ff26b),
	.w4(32'h3b190e78),
	.w5(32'hbb91ad72),
	.w6(32'hbbaf4bd3),
	.w7(32'h3a3324e9),
	.w8(32'h3c07b3cd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e01b6),
	.w1(32'h3b1d102c),
	.w2(32'hbbdd9fcb),
	.w3(32'h3c0f941a),
	.w4(32'h3bd3fd7a),
	.w5(32'hbb28eff3),
	.w6(32'h3af4983b),
	.w7(32'hbbf05e5b),
	.w8(32'h3ab78d73),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d84a78),
	.w1(32'hba9e3eac),
	.w2(32'hbbe0150a),
	.w3(32'h3aa85faa),
	.w4(32'h3a8bd418),
	.w5(32'hbbef5ddc),
	.w6(32'hbb25edf4),
	.w7(32'hbc676d4a),
	.w8(32'hb9bb5f74),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fd898),
	.w1(32'h3bd2b481),
	.w2(32'h3c1927d7),
	.w3(32'h3ba87774),
	.w4(32'h3bccab23),
	.w5(32'h3b98cb9a),
	.w6(32'h3ba7da7f),
	.w7(32'h3baf0a2e),
	.w8(32'h3bc0486f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba7d0f),
	.w1(32'h3bc9b3fa),
	.w2(32'h3b93b5b7),
	.w3(32'h3b9b9b28),
	.w4(32'hba8ecd77),
	.w5(32'h3bd69b9c),
	.w6(32'h3c0dbd7e),
	.w7(32'h3c4ae9e2),
	.w8(32'hbc400f45),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c874c),
	.w1(32'hbd295510),
	.w2(32'hbb21f423),
	.w3(32'hbc554d93),
	.w4(32'hbd0661b5),
	.w5(32'hbc988250),
	.w6(32'hbd01b5cf),
	.w7(32'h3ae4adb3),
	.w8(32'h3cfd4923),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d253776),
	.w1(32'hbb95d03e),
	.w2(32'hbb60f335),
	.w3(32'h3cb50279),
	.w4(32'h3a014d95),
	.w5(32'hbabfc82f),
	.w6(32'hbb1116c9),
	.w7(32'h38bbc539),
	.w8(32'h3bdd49fc),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb18dc7),
	.w1(32'h3b46345b),
	.w2(32'hbb24fc09),
	.w3(32'h3b459d52),
	.w4(32'h3840c9ca),
	.w5(32'hba25cc12),
	.w6(32'h3bed73e6),
	.w7(32'h3b0fa4cc),
	.w8(32'hbc3ad2d8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6ee08),
	.w1(32'hbc52a329),
	.w2(32'hbcb08065),
	.w3(32'hbbc2019a),
	.w4(32'hbc10ba11),
	.w5(32'hbc43f939),
	.w6(32'hbc7344d6),
	.w7(32'hbb64030f),
	.w8(32'h3c678784),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bc58a),
	.w1(32'hbcbd241d),
	.w2(32'hbc86a2ed),
	.w3(32'h3ba51abc),
	.w4(32'hbc5d684a),
	.w5(32'hbc41f73d),
	.w6(32'hbbfe09b7),
	.w7(32'hbb9f84e8),
	.w8(32'h3c263783),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd397f),
	.w1(32'hb9959077),
	.w2(32'h3c02cbe6),
	.w3(32'h398b759a),
	.w4(32'hba9551db),
	.w5(32'h3ba7f59d),
	.w6(32'hbb4a7d35),
	.w7(32'h3ba70982),
	.w8(32'hbbf65d87),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92c473),
	.w1(32'h3aced99e),
	.w2(32'hbbc2f2ed),
	.w3(32'hbbc9bfba),
	.w4(32'h3b154d12),
	.w5(32'hbc084113),
	.w6(32'h3ada8c50),
	.w7(32'hbbfdf626),
	.w8(32'h3b0b5294),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9978d1c),
	.w1(32'hbbc3d2e6),
	.w2(32'h3b0d2bc8),
	.w3(32'h3ae7ee40),
	.w4(32'h3b2c6316),
	.w5(32'h3bd132a5),
	.w6(32'hbba50951),
	.w7(32'hb97b85f8),
	.w8(32'h3c07f2a2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdbbfd),
	.w1(32'hbb1e29ff),
	.w2(32'h3b252ce8),
	.w3(32'h3c0fee74),
	.w4(32'h38d9f298),
	.w5(32'h3bd4ba34),
	.w6(32'hbb77d352),
	.w7(32'hb9908e34),
	.w8(32'hba9eaf96),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb879a),
	.w1(32'h3ca1379f),
	.w2(32'h3ce04334),
	.w3(32'h3bb7ef71),
	.w4(32'h3c7bcfa1),
	.w5(32'h3cae8775),
	.w6(32'h3d0061ed),
	.w7(32'h3ce73a3f),
	.w8(32'hbb2f497c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba563f8),
	.w1(32'h3b83c358),
	.w2(32'h3c482ff0),
	.w3(32'hbb73e0a0),
	.w4(32'hbc1cc3df),
	.w5(32'h3bb07532),
	.w6(32'h3b23c75b),
	.w7(32'h3c8248da),
	.w8(32'h3babca10),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62d59f),
	.w1(32'h3c803ab0),
	.w2(32'hbb216605),
	.w3(32'hbaeba5d0),
	.w4(32'h3b27593d),
	.w5(32'h39e2bb77),
	.w6(32'h3c01c0d2),
	.w7(32'hbb81cc3d),
	.w8(32'hbba75377),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb009d8),
	.w1(32'hbbf361b0),
	.w2(32'hbca7860b),
	.w3(32'hbc896fce),
	.w4(32'h3b69900c),
	.w5(32'hbc27af78),
	.w6(32'hbba8d298),
	.w7(32'hbc10fabd),
	.w8(32'h3c311ef3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be22f0b),
	.w1(32'hbb8db3ee),
	.w2(32'hbb35e1d4),
	.w3(32'h3a4788fd),
	.w4(32'hba9cee37),
	.w5(32'hbc16c8ac),
	.w6(32'hbb9b2878),
	.w7(32'h3b136c98),
	.w8(32'hb9f03f12),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39276d2c),
	.w1(32'hbb49cc26),
	.w2(32'hbc03f961),
	.w3(32'hba88584b),
	.w4(32'hbb3a285c),
	.w5(32'hbb271031),
	.w6(32'hbb0e8ef6),
	.w7(32'hbb85e4c5),
	.w8(32'hbaa5b2ba),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4c233),
	.w1(32'hbc3f894b),
	.w2(32'hbcefa594),
	.w3(32'hba5d51af),
	.w4(32'h3b3c3ae3),
	.w5(32'hbcaa2da6),
	.w6(32'hbc127373),
	.w7(32'hbc3fda28),
	.w8(32'h374f60d5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba429c50),
	.w1(32'h3c010e08),
	.w2(32'h3a690cef),
	.w3(32'hbb6f4475),
	.w4(32'h3c849813),
	.w5(32'h3b981d51),
	.w6(32'h3c2bee63),
	.w7(32'hba919be5),
	.w8(32'hbc32c395),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3683be),
	.w1(32'hba67d762),
	.w2(32'h3aa3d0a0),
	.w3(32'hbb95ebfd),
	.w4(32'h39b7a9b5),
	.w5(32'hbbc06099),
	.w6(32'hba584356),
	.w7(32'hbb1d3058),
	.w8(32'hbba2ca56),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51149f),
	.w1(32'h3b9bdda6),
	.w2(32'h3c6e26c3),
	.w3(32'hbbc61c5a),
	.w4(32'h3a3017f3),
	.w5(32'h3c1e0853),
	.w6(32'hba241f12),
	.w7(32'h3c089cdc),
	.w8(32'h3c2f417b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47cf4b),
	.w1(32'h3bba91ca),
	.w2(32'hbbaf560d),
	.w3(32'h3c1cc0d5),
	.w4(32'h3b95949b),
	.w5(32'hbbe53852),
	.w6(32'h3c13da53),
	.w7(32'hbb297fc0),
	.w8(32'h3b1ed8b3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb31013),
	.w1(32'hba8f19c6),
	.w2(32'h3a865ffd),
	.w3(32'hbb9e98ab),
	.w4(32'hb9680104),
	.w5(32'h3ab75b3d),
	.w6(32'hbada2bfa),
	.w7(32'h3aa9f02b),
	.w8(32'h3b298351),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbe87a),
	.w1(32'hbb12f567),
	.w2(32'hbc864a5a),
	.w3(32'hba193805),
	.w4(32'hbb29e41c),
	.w5(32'hbc8e77a5),
	.w6(32'hbb1a9848),
	.w7(32'hbb0e9069),
	.w8(32'h3b539ed9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb136ddd),
	.w1(32'hbc0778b7),
	.w2(32'hbb458229),
	.w3(32'h3bcd2f96),
	.w4(32'h3bc1eea5),
	.w5(32'h39a5ec05),
	.w6(32'hbbcf9a2b),
	.w7(32'hba5dec85),
	.w8(32'h3bd5c587),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2b75e),
	.w1(32'h3bc9be5a),
	.w2(32'hbbaf2ce7),
	.w3(32'hbbb15f21),
	.w4(32'h3bce710f),
	.w5(32'hbbabae3b),
	.w6(32'h3bdf0fcb),
	.w7(32'hbbb74618),
	.w8(32'hbc16566c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b22d1),
	.w1(32'h3caa797c),
	.w2(32'h3cc2985e),
	.w3(32'hbc0df0ed),
	.w4(32'h3b77c516),
	.w5(32'h3c975c27),
	.w6(32'h3bdbfcad),
	.w7(32'h3c38d289),
	.w8(32'hbc52b9df),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe828d8),
	.w1(32'hbc107202),
	.w2(32'hbc906693),
	.w3(32'hba8d8bc7),
	.w4(32'hbc8ad316),
	.w5(32'hbc6f6507),
	.w6(32'hbc625e56),
	.w7(32'h3b12e763),
	.w8(32'h3bfb5d5c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c124f),
	.w1(32'hbb2f1289),
	.w2(32'h3a974bb2),
	.w3(32'hbbac9d56),
	.w4(32'h3a0f36c6),
	.w5(32'h3b8e3915),
	.w6(32'hbac9d3af),
	.w7(32'h39939a2d),
	.w8(32'h3c104e77),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80b45f),
	.w1(32'hbd02a539),
	.w2(32'h3bfd9e9f),
	.w3(32'h3c1032f4),
	.w4(32'hbcae0f93),
	.w5(32'hbbbc6598),
	.w6(32'hbc209c71),
	.w7(32'h3c2e5d48),
	.w8(32'h3b82cdcc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a351f),
	.w1(32'hbd00cda1),
	.w2(32'hbbf09d92),
	.w3(32'h3b2daeab),
	.w4(32'hbc8ba4cb),
	.w5(32'hbc21f73c),
	.w6(32'hbc8aac27),
	.w7(32'h3c52affb),
	.w8(32'h3c8bd8d6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e8b09),
	.w1(32'hbbf20168),
	.w2(32'hbb64b0e3),
	.w3(32'hb922909e),
	.w4(32'hbb202dae),
	.w5(32'hba2ff617),
	.w6(32'hbb2283fd),
	.w7(32'hbb2c1732),
	.w8(32'hbb0e9716),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ebfda6),
	.w1(32'hbae68202),
	.w2(32'h3ae081f7),
	.w3(32'h39302503),
	.w4(32'hba79a302),
	.w5(32'hba37cb70),
	.w6(32'h3b2ae046),
	.w7(32'h3b7eaceb),
	.w8(32'h3af76d6c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29bcde),
	.w1(32'h3bc14d6c),
	.w2(32'hbbbf54d6),
	.w3(32'hbb987b7e),
	.w4(32'h3b2d7ad6),
	.w5(32'hbb9a2972),
	.w6(32'hba74598c),
	.w7(32'hbb612c0b),
	.w8(32'h39b3350b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1ce6b),
	.w1(32'h3bafe3d9),
	.w2(32'h3ba42d08),
	.w3(32'hbc106e21),
	.w4(32'h3b52253e),
	.w5(32'h3a7dff53),
	.w6(32'h3beedf0f),
	.w7(32'h3bc845f5),
	.w8(32'h3be3c19f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92f61d),
	.w1(32'h3afa284e),
	.w2(32'hbbf0937e),
	.w3(32'h3aafdfeb),
	.w4(32'h3a123817),
	.w5(32'hbc402cba),
	.w6(32'h3b36848d),
	.w7(32'hbbc7b633),
	.w8(32'h38f3edf5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87b99b),
	.w1(32'h3b32fa98),
	.w2(32'hbbd370f8),
	.w3(32'hbb940900),
	.w4(32'h3bfeed8c),
	.w5(32'hbb19ecd0),
	.w6(32'hbb6f90c0),
	.w7(32'hbb6b8cca),
	.w8(32'hbaab097e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc531),
	.w1(32'h3c8f27f7),
	.w2(32'hbc9c4279),
	.w3(32'h3b72eef8),
	.w4(32'h3b48f1cf),
	.w5(32'hbc9a0341),
	.w6(32'h3c098f8c),
	.w7(32'hbc9a2ba8),
	.w8(32'hbb90e543),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d4d8e),
	.w1(32'hbc82fe62),
	.w2(32'h3c1fa366),
	.w3(32'hbcc2f9b0),
	.w4(32'h38d57538),
	.w5(32'h3bd08384),
	.w6(32'hbbd6cd1b),
	.w7(32'h3c3fb80b),
	.w8(32'h3a906808),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87038c),
	.w1(32'h3bb0fcce),
	.w2(32'h3c91aba5),
	.w3(32'h3a5d41bf),
	.w4(32'h39898188),
	.w5(32'h3c44c832),
	.w6(32'hbb7b8694),
	.w7(32'h3c2ceaed),
	.w8(32'hbb498458),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab64ee8),
	.w1(32'h3b0dd75d),
	.w2(32'hbbbb4474),
	.w3(32'h3bd29db7),
	.w4(32'h3b87070b),
	.w5(32'hbbeb6302),
	.w6(32'h3b41c74d),
	.w7(32'hbc2e81f9),
	.w8(32'h3bc72656),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939bee3),
	.w1(32'h3c980145),
	.w2(32'h3cd6071e),
	.w3(32'h3b1d9848),
	.w4(32'h3c2d0843),
	.w5(32'h3c14a205),
	.w6(32'h3c8ee5a4),
	.w7(32'h3cadb9c6),
	.w8(32'h3ba81cc7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb467ca),
	.w1(32'hbaee56b0),
	.w2(32'h3cf1a22a),
	.w3(32'hba92055e),
	.w4(32'h3ba31e06),
	.w5(32'h3c958ce1),
	.w6(32'h3aa74c03),
	.w7(32'h3c9935d3),
	.w8(32'h3b89ec4a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cf7e5),
	.w1(32'hba17b081),
	.w2(32'hbc46ead3),
	.w3(32'h3bdda7e8),
	.w4(32'hbbdae63c),
	.w5(32'hbc8037a5),
	.w6(32'h3bed1881),
	.w7(32'h3afa41f4),
	.w8(32'hba2b9134),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b26ed),
	.w1(32'hbb196baa),
	.w2(32'hbb7b1b8d),
	.w3(32'h3bc06d32),
	.w4(32'h3a2da7b4),
	.w5(32'hbaff6e2c),
	.w6(32'hbbbd4ff5),
	.w7(32'hbb2a10ca),
	.w8(32'h3aad8336),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea929a),
	.w1(32'h3b28bbea),
	.w2(32'h3a2205cc),
	.w3(32'hba34e000),
	.w4(32'h3b89a24d),
	.w5(32'h3abd1569),
	.w6(32'h3a69e378),
	.w7(32'h3a3123a4),
	.w8(32'hba9f12a2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48d86a),
	.w1(32'hbba3864e),
	.w2(32'h3a0c1564),
	.w3(32'hbb40bfc3),
	.w4(32'h3a9d2225),
	.w5(32'h3b2bc181),
	.w6(32'hbb902c05),
	.w7(32'hb9ad89eb),
	.w8(32'h3afd9dc3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78f185),
	.w1(32'hbcbc6c82),
	.w2(32'hbc20c1c5),
	.w3(32'h3a35dfdd),
	.w4(32'hbabc3264),
	.w5(32'hbbd203ad),
	.w6(32'h3a30f1fd),
	.w7(32'h3bc79f89),
	.w8(32'h3b4d99d6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dc581),
	.w1(32'hbd0563ab),
	.w2(32'h3bbaa201),
	.w3(32'h3c06c35a),
	.w4(32'hbcf3820e),
	.w5(32'hbbf98748),
	.w6(32'hba67a12f),
	.w7(32'h3bf73f75),
	.w8(32'h3c27e1c2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2e0f8),
	.w1(32'h3b901ade),
	.w2(32'h3c62a83b),
	.w3(32'h3c2caa1e),
	.w4(32'hbbb1d6c3),
	.w5(32'h3b94ae56),
	.w6(32'h39e1e3ea),
	.w7(32'h3b1fa4d0),
	.w8(32'hbad7af5e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b894aef),
	.w1(32'h3ab87ebb),
	.w2(32'h3abf6ad6),
	.w3(32'h3bc859b8),
	.w4(32'h3b9800dc),
	.w5(32'h3b23b552),
	.w6(32'hba152d1c),
	.w7(32'h3ada4efb),
	.w8(32'h3b2fb73f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d0868),
	.w1(32'h3b871c6c),
	.w2(32'h3b309cd9),
	.w3(32'h3b1e922f),
	.w4(32'h3b1c8b64),
	.w5(32'h3b98d889),
	.w6(32'h39bf0843),
	.w7(32'h3b2994a7),
	.w8(32'hbbd7a874),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1e057),
	.w1(32'h3c4c71cf),
	.w2(32'h3c88f08c),
	.w3(32'hbb3a650d),
	.w4(32'h3c02ede8),
	.w5(32'h3c0b6448),
	.w6(32'h3c962908),
	.w7(32'h3c560747),
	.w8(32'h3bdaf6e4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec2f74),
	.w1(32'hbb288652),
	.w2(32'h3b304db6),
	.w3(32'hba694d19),
	.w4(32'hbb5b3e1c),
	.w5(32'h3a627f2c),
	.w6(32'hbb2114df),
	.w7(32'h3b6a7d50),
	.w8(32'h39bc5ec0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2470e),
	.w1(32'hbb876c7b),
	.w2(32'hbc8aa5a3),
	.w3(32'hbb05d632),
	.w4(32'h3b244bde),
	.w5(32'hbbe3f5b3),
	.w6(32'hbc3a5c57),
	.w7(32'hbba7d3b3),
	.w8(32'hbbe09c19),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2460ff),
	.w1(32'h3b713c37),
	.w2(32'hbc6eb18e),
	.w3(32'hbc62ac28),
	.w4(32'h3c3be897),
	.w5(32'hbb7c4497),
	.w6(32'h3930d884),
	.w7(32'h3b0e09e3),
	.w8(32'hbc31a7b6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f83bc),
	.w1(32'h3cb8a9e6),
	.w2(32'hbc138634),
	.w3(32'hbc3e7113),
	.w4(32'h3cad8065),
	.w5(32'h3a8dc278),
	.w6(32'h3c3b1aad),
	.w7(32'hbba864ea),
	.w8(32'hbc3abd7c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21e620),
	.w1(32'h3c031d77),
	.w2(32'hbc280c76),
	.w3(32'hbc04ef79),
	.w4(32'h3baa1afb),
	.w5(32'h3b810e25),
	.w6(32'hbb14f0be),
	.w7(32'hbc223a5f),
	.w8(32'hbc320950),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7efb04),
	.w1(32'hbc290f9a),
	.w2(32'h3c551068),
	.w3(32'hbc141d9d),
	.w4(32'hbbc90077),
	.w5(32'hb94ad39f),
	.w6(32'hbb93a94a),
	.w7(32'hbb7f5bd0),
	.w8(32'h3c5dbcea),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7866a1),
	.w1(32'hbc8b1b6f),
	.w2(32'h3c9c99c1),
	.w3(32'h3cafaba9),
	.w4(32'hbc99feb8),
	.w5(32'h3b5a6575),
	.w6(32'hbc8a42d3),
	.w7(32'h3c8368be),
	.w8(32'h3c14772c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01ba3a),
	.w1(32'hbbf3b7ce),
	.w2(32'h3ca76f17),
	.w3(32'hbb5156ad),
	.w4(32'hbc4702b8),
	.w5(32'h3bd96557),
	.w6(32'hbb5d1e5d),
	.w7(32'h3c3b3524),
	.w8(32'h3b33b5b9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c09f7),
	.w1(32'hbc98bf7e),
	.w2(32'hbbc0f01e),
	.w3(32'h3c4ba6aa),
	.w4(32'hbc35e1c5),
	.w5(32'hbbaa7364),
	.w6(32'hbc4a9327),
	.w7(32'h3aa7b471),
	.w8(32'h3c0a376e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde865a),
	.w1(32'hbb776ceb),
	.w2(32'hbcb2c67a),
	.w3(32'h3ab31bb9),
	.w4(32'h3ba623c7),
	.w5(32'hbc7b4e79),
	.w6(32'h3b68ad32),
	.w7(32'hbc0f493b),
	.w8(32'h3c690724),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1833cd),
	.w1(32'hbbb461ea),
	.w2(32'h3ab54315),
	.w3(32'h3c061ec5),
	.w4(32'hbae862b8),
	.w5(32'h3a9e31c5),
	.w6(32'hbb3fc52c),
	.w7(32'h3b80cf23),
	.w8(32'h3a86f70a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac1271),
	.w1(32'hbb43f5bf),
	.w2(32'hba52eeca),
	.w3(32'hbb16da39),
	.w4(32'hbb7f7628),
	.w5(32'hba4ef200),
	.w6(32'hbb26a4e7),
	.w7(32'h3b7a7e49),
	.w8(32'h3ab7a341),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb667d30),
	.w1(32'hbb8a0fbd),
	.w2(32'hbbbc98f3),
	.w3(32'hbc2a3767),
	.w4(32'hbbac1db5),
	.w5(32'hbc5e955c),
	.w6(32'hbb58f1f9),
	.w7(32'hbc35c2ac),
	.w8(32'hbc0968fe),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a2b6e),
	.w1(32'h3c496d6c),
	.w2(32'h3bff4b93),
	.w3(32'hbbc94f11),
	.w4(32'h3bde7e75),
	.w5(32'h3bdef120),
	.w6(32'h3c64e2e0),
	.w7(32'h3b7ea670),
	.w8(32'h3ab254e1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2dc98),
	.w1(32'h3a3bcabb),
	.w2(32'h3b2f3510),
	.w3(32'h3918d2f3),
	.w4(32'hbabec2ed),
	.w5(32'h3b69ff90),
	.w6(32'h38323b4f),
	.w7(32'h3a6214a0),
	.w8(32'hb911fea8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a836745),
	.w1(32'hbbff0ebd),
	.w2(32'h3cb5e418),
	.w3(32'h3ac39395),
	.w4(32'hbc16613f),
	.w5(32'h3c3bc658),
	.w6(32'h3aa74e75),
	.w7(32'h3bbfbd28),
	.w8(32'hbb2f0a6e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc72251),
	.w1(32'h3b1b0264),
	.w2(32'hb87fac50),
	.w3(32'h3ca78987),
	.w4(32'h39c1467b),
	.w5(32'hbb072c10),
	.w6(32'h3a66e82e),
	.w7(32'h3b4cb366),
	.w8(32'h3b8bd9a9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa278c3),
	.w1(32'h3c00e22c),
	.w2(32'h3c99d2c7),
	.w3(32'hba766e59),
	.w4(32'h3b74c791),
	.w5(32'h3c8c2acc),
	.w6(32'h3bb247e1),
	.w7(32'h3c6dcf98),
	.w8(32'h3b03a372),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5922f),
	.w1(32'hbcacee98),
	.w2(32'hbc5932a2),
	.w3(32'hba9a8472),
	.w4(32'hbc4d91c8),
	.w5(32'hbb884f3f),
	.w6(32'hbc8a1e9d),
	.w7(32'hbb3620c6),
	.w8(32'h3b3096e2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa5bb6),
	.w1(32'hbc00754b),
	.w2(32'hbb71c630),
	.w3(32'hbbd7e51b),
	.w4(32'hbb0eb8a5),
	.w5(32'hbb522818),
	.w6(32'hbb9609d4),
	.w7(32'hbb638a97),
	.w8(32'h3aac3f29),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f8146),
	.w1(32'h3b629c07),
	.w2(32'h3bae03b6),
	.w3(32'h3bc9dc6d),
	.w4(32'h3b2ddda6),
	.w5(32'h3bd06f94),
	.w6(32'h3a83a668),
	.w7(32'h3b07de89),
	.w8(32'h3a63ae0d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad68b),
	.w1(32'h3b1d2756),
	.w2(32'hbbb3e50c),
	.w3(32'h3b227a25),
	.w4(32'h3bd2c6c9),
	.w5(32'hba70ca1b),
	.w6(32'hbb0e3083),
	.w7(32'hbc1148b7),
	.w8(32'h3b73f487),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8db64),
	.w1(32'h3ba31836),
	.w2(32'h3c52281c),
	.w3(32'h3c09533e),
	.w4(32'h3b0c454a),
	.w5(32'h3c3d0a8c),
	.w6(32'h3bfcad37),
	.w7(32'h3bd4245f),
	.w8(32'hbb11ea06),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45d6b1),
	.w1(32'h3b1eade6),
	.w2(32'h3c542055),
	.w3(32'hbba8da64),
	.w4(32'hbc0d2038),
	.w5(32'h3c05bdec),
	.w6(32'hbab05637),
	.w7(32'h3b58cf84),
	.w8(32'hbba5e1f8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab2c87),
	.w1(32'h39ef8324),
	.w2(32'h39dbc04d),
	.w3(32'h3baf6a33),
	.w4(32'hbb248609),
	.w5(32'hbb3713c5),
	.w6(32'h3abe9b45),
	.w7(32'hb8b50e0a),
	.w8(32'h3b2a89b5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb4ffa),
	.w1(32'h3c89c216),
	.w2(32'h3c7d90e2),
	.w3(32'h3b41866b),
	.w4(32'h3b9f22fc),
	.w5(32'h3bc760d5),
	.w6(32'h3ba69a94),
	.w7(32'h3c0946d4),
	.w8(32'hbbb5bb59),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf11f73),
	.w1(32'h3af90b6d),
	.w2(32'hba9d8abc),
	.w3(32'hbb64ce61),
	.w4(32'h3ba467be),
	.w5(32'h3a8cdce8),
	.w6(32'h3a08309f),
	.w7(32'hba379f20),
	.w8(32'hbbd565fd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84d656),
	.w1(32'h3b16185f),
	.w2(32'h3bb394cb),
	.w3(32'hba9e8b49),
	.w4(32'h3ace8bba),
	.w5(32'h3b928692),
	.w6(32'h39908a3d),
	.w7(32'h3b44012e),
	.w8(32'hb9acf2f0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02ab91),
	.w1(32'h3ab02946),
	.w2(32'h3c1750fe),
	.w3(32'h3b4c1f46),
	.w4(32'hbaf2268d),
	.w5(32'h3ba0f14b),
	.w6(32'hbba036df),
	.w7(32'h3bbc3004),
	.w8(32'h3b7cef2b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76699c),
	.w1(32'hbc747717),
	.w2(32'h3c95b727),
	.w3(32'hbb340486),
	.w4(32'hbc2ae4db),
	.w5(32'h3b0e49d9),
	.w6(32'hbc6aa731),
	.w7(32'h3c554c6d),
	.w8(32'h3be15f40),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cce93),
	.w1(32'hbc0905c2),
	.w2(32'hbcd0c4e8),
	.w3(32'h3c1d4eeb),
	.w4(32'hbc0953d0),
	.w5(32'hbc025e5d),
	.w6(32'hbbb64497),
	.w7(32'hbbb48d0a),
	.w8(32'h3c4d1a62),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2eab3),
	.w1(32'hbb0f4357),
	.w2(32'hbbad652f),
	.w3(32'h3a954fea),
	.w4(32'hba2f272b),
	.w5(32'hba5a558c),
	.w6(32'hbb08c78a),
	.w7(32'hbb658526),
	.w8(32'hbaed2c3b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad030d),
	.w1(32'hbbb59f36),
	.w2(32'hbc736c5b),
	.w3(32'h39753ef4),
	.w4(32'h3c1622ff),
	.w5(32'h39cccda6),
	.w6(32'h3a3c768a),
	.w7(32'h3b8dc7ff),
	.w8(32'h3c8c0e75),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule