module layer_8_featuremap_141(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c255ff2),
	.w1(32'h3bd9e329),
	.w2(32'hbb35797a),
	.w3(32'h3c4c92ab),
	.w4(32'h3be630c6),
	.w5(32'h3b6fe252),
	.w6(32'h3c070f05),
	.w7(32'h3be3e57c),
	.w8(32'hbadf3268),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fe381),
	.w1(32'h38ebe264),
	.w2(32'hba699972),
	.w3(32'hbbe5a2ea),
	.w4(32'h3ac9975a),
	.w5(32'h3a08f3f1),
	.w6(32'hbb8998ac),
	.w7(32'h3b798ece),
	.w8(32'h3b6caeec),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb5162),
	.w1(32'h3b441912),
	.w2(32'h3b66fc51),
	.w3(32'hbbaa2113),
	.w4(32'h3b852d12),
	.w5(32'h3b5d5949),
	.w6(32'hbbc48566),
	.w7(32'h3b8bd29f),
	.w8(32'h3ba0368b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb438397),
	.w1(32'h38e30d9b),
	.w2(32'hbc87f676),
	.w3(32'hbb808572),
	.w4(32'h3ae2efab),
	.w5(32'hbbc7511e),
	.w6(32'hbc2b4307),
	.w7(32'hbb39f442),
	.w8(32'hbc730d2f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc906555),
	.w1(32'hbc131606),
	.w2(32'hbbaeacde),
	.w3(32'hbc119193),
	.w4(32'h3ac5e5f1),
	.w5(32'h3b4589c5),
	.w6(32'hbbb7880e),
	.w7(32'h3bf2da48),
	.w8(32'h3bf2e46e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd393ab2),
	.w1(32'hbbf61bea),
	.w2(32'hbba42f3b),
	.w3(32'hbd0215df),
	.w4(32'h3bc40531),
	.w5(32'h3b4e508e),
	.w6(32'hbcf7e7b7),
	.w7(32'h3b9503f0),
	.w8(32'h3a8bdcc8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3bc00),
	.w1(32'h3915f64c),
	.w2(32'h39307811),
	.w3(32'h39cac9ce),
	.w4(32'h37937877),
	.w5(32'h38017578),
	.w6(32'h39be71e6),
	.w7(32'h38037df5),
	.w8(32'h3833e096),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81ba68),
	.w1(32'hbb8d2b90),
	.w2(32'hbc45a6c0),
	.w3(32'hbc205fd4),
	.w4(32'hbb0adca4),
	.w5(32'h380fe6fa),
	.w6(32'hbaa2f0d7),
	.w7(32'h38ea280c),
	.w8(32'hb980fb0d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe64e44),
	.w1(32'hba2bf270),
	.w2(32'h3ad8cc76),
	.w3(32'hbaa63b04),
	.w4(32'h3bb1617a),
	.w5(32'h3bffebbd),
	.w6(32'h3ba69d64),
	.w7(32'h3c5bfa60),
	.w8(32'h3c5427b9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1fda3),
	.w1(32'h3a9bf270),
	.w2(32'hbb9d643a),
	.w3(32'h3ae85788),
	.w4(32'h3b85f4a7),
	.w5(32'h3b05ff10),
	.w6(32'h3bb5da11),
	.w7(32'h3bbbf35a),
	.w8(32'h3b58755d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94df7fe),
	.w1(32'hbb7d3f64),
	.w2(32'hbc54a297),
	.w3(32'h3bcf38e6),
	.w4(32'hbab9ca5c),
	.w5(32'hbb9d1c1e),
	.w6(32'hba4b3d5e),
	.w7(32'h3b03cbc3),
	.w8(32'hbbd737e3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86c5bb),
	.w1(32'hbbbb4ba6),
	.w2(32'hbc83e8ba),
	.w3(32'hbb397c8d),
	.w4(32'h3bd4d1fc),
	.w5(32'hba7a3359),
	.w6(32'hbc00e2c3),
	.w7(32'h3bbd6bf9),
	.w8(32'hbb41513e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94a370),
	.w1(32'hbb39d8a4),
	.w2(32'hbad07eda),
	.w3(32'hbc2d1238),
	.w4(32'h3c1b263f),
	.w5(32'h3a1663ea),
	.w6(32'hbc16e927),
	.w7(32'h3c56c6d2),
	.w8(32'h3c273ebe),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4540dc),
	.w1(32'h3addfaa0),
	.w2(32'hbb50df49),
	.w3(32'hb9d7d3e4),
	.w4(32'hbba3782c),
	.w5(32'hba5425c4),
	.w6(32'h3bcafca1),
	.w7(32'hbbc22f9a),
	.w8(32'h3a961f8b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ad950),
	.w1(32'hbc0c7dda),
	.w2(32'hbbf1a8ff),
	.w3(32'hbbaa6606),
	.w4(32'hbbeaa756),
	.w5(32'hbb29a19c),
	.w6(32'hbc1b04f9),
	.w7(32'hbc0efe9d),
	.w8(32'hb945b5ab),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9183d6b),
	.w1(32'hbb89372e),
	.w2(32'h3c4084a8),
	.w3(32'hbb601f2c),
	.w4(32'h3bcfc56c),
	.w5(32'h3b8fa169),
	.w6(32'hbb7c6bfd),
	.w7(32'h3c881f34),
	.w8(32'hbb8188bd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb821631),
	.w1(32'hbbb10b1c),
	.w2(32'h3c16c7a7),
	.w3(32'hbbd76add),
	.w4(32'h3bf2f5e0),
	.w5(32'hba64b5a8),
	.w6(32'hbc5376a0),
	.w7(32'hbc1831fc),
	.w8(32'hbc5db35f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d0996),
	.w1(32'hbd1c24db),
	.w2(32'hbb4556f8),
	.w3(32'hbcfe1870),
	.w4(32'h3c3067dd),
	.w5(32'h3b236358),
	.w6(32'hbd03f9e8),
	.w7(32'h3c6cca7d),
	.w8(32'h3b855097),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc578c20),
	.w1(32'hbc9c2216),
	.w2(32'hbd1b89f1),
	.w3(32'hbc9aeb6b),
	.w4(32'hbc9dde58),
	.w5(32'hbd0e6f33),
	.w6(32'hbc4b82e3),
	.w7(32'hbca9cef1),
	.w8(32'hbd49723e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9ecd1),
	.w1(32'hbcd50369),
	.w2(32'hbc67c31c),
	.w3(32'hbceb3980),
	.w4(32'h3c94f42c),
	.w5(32'h3b247489),
	.w6(32'hbd2b6bf3),
	.w7(32'h3c0d9ec6),
	.w8(32'h3b9a2eae),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94e0e1),
	.w1(32'hbaaa4062),
	.w2(32'hb9e559c2),
	.w3(32'hbc372945),
	.w4(32'hbc3261d7),
	.w5(32'h3b5248ef),
	.w6(32'hbc695e6a),
	.w7(32'hbd483207),
	.w8(32'h3b748dcf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88b320),
	.w1(32'h3c8eb32e),
	.w2(32'h3cf941ea),
	.w3(32'hbbb53b10),
	.w4(32'hbbd3e371),
	.w5(32'hbb919c5c),
	.w6(32'hbb8e68ab),
	.w7(32'h3c45cc1e),
	.w8(32'hbb83ad4f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d330da8),
	.w1(32'h3acaa945),
	.w2(32'h3bf711a2),
	.w3(32'h3d79af3e),
	.w4(32'h3d20574b),
	.w5(32'h3cb9d2d1),
	.w6(32'h3d38e27f),
	.w7(32'h3d36adbe),
	.w8(32'h3d5c885b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc990976),
	.w1(32'hbbdd2e4a),
	.w2(32'h3c341543),
	.w3(32'hbcbc6220),
	.w4(32'h3c25e105),
	.w5(32'h3c5d8b24),
	.w6(32'hbc03e1b4),
	.w7(32'h3d025238),
	.w8(32'h3c87aa39),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dc672),
	.w1(32'hbbcfd95c),
	.w2(32'hbcbdfe34),
	.w3(32'hbbe888ce),
	.w4(32'hbc229bce),
	.w5(32'hbca5ff43),
	.w6(32'hbbe578db),
	.w7(32'hbcc5fc2b),
	.w8(32'hbca65dd9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6156a),
	.w1(32'hbbb1526b),
	.w2(32'h3beac7f0),
	.w3(32'h3bab4421),
	.w4(32'hba8a35b9),
	.w5(32'h3bb692b4),
	.w6(32'hbbd19aaf),
	.w7(32'hbc08ef2f),
	.w8(32'h3c9081d9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b865b08),
	.w1(32'h3c03e3d9),
	.w2(32'hbbc3c24d),
	.w3(32'h3ad0873c),
	.w4(32'h3c235c2c),
	.w5(32'hbc99de16),
	.w6(32'h3c39cc82),
	.w7(32'h3c01f545),
	.w8(32'hbb8630f0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdcf0ef2),
	.w1(32'h3bc224b6),
	.w2(32'hbd83460c),
	.w3(32'hbc9aed53),
	.w4(32'h3d8515f0),
	.w5(32'h3c12702b),
	.w6(32'hbddb2601),
	.w7(32'hbd20b917),
	.w8(32'hbd85222a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9eb91),
	.w1(32'h3c20bd38),
	.w2(32'hbbf6b440),
	.w3(32'h3c198377),
	.w4(32'hbb1dd0d4),
	.w5(32'h3b4be450),
	.w6(32'h3c11e699),
	.w7(32'hb9ae2b60),
	.w8(32'h3c5c2890),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc582b07),
	.w1(32'hbbade4c6),
	.w2(32'hb9fa49eb),
	.w3(32'hbc27bfc1),
	.w4(32'h3b9bf121),
	.w5(32'hb9d059f3),
	.w6(32'h3c35b136),
	.w7(32'h3c3f41ca),
	.w8(32'hbc945f44),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc25d94),
	.w1(32'hbc656812),
	.w2(32'hbbd6333a),
	.w3(32'hba63fb6c),
	.w4(32'hbb860eb5),
	.w5(32'hbb69c2d2),
	.w6(32'hbc5e5fd8),
	.w7(32'hbc02eab0),
	.w8(32'hbb9416b8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85f8a6),
	.w1(32'hbbb22d53),
	.w2(32'h3ccc771f),
	.w3(32'hbc596d6d),
	.w4(32'h3b21287a),
	.w5(32'hbba9b05d),
	.w6(32'hbc2df4a8),
	.w7(32'h3cfe7f94),
	.w8(32'hbb70504a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23b134),
	.w1(32'hbcf335b3),
	.w2(32'h3bd49d0c),
	.w3(32'hbc5f4e80),
	.w4(32'h3b241d58),
	.w5(32'hbcb9804a),
	.w6(32'hbc962452),
	.w7(32'h3b61fdae),
	.w8(32'h3cb900d1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a7730),
	.w1(32'h3a51926b),
	.w2(32'h3c402814),
	.w3(32'hbbde6966),
	.w4(32'h3c04215a),
	.w5(32'hb9d02822),
	.w6(32'h3c12203d),
	.w7(32'h3c274b57),
	.w8(32'hbcbdd85a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4196ed),
	.w1(32'hbbd6a66b),
	.w2(32'hbbd80935),
	.w3(32'hbcd57e47),
	.w4(32'hbc10e33b),
	.w5(32'h3a82f808),
	.w6(32'hbd2b1fbc),
	.w7(32'hbce821d2),
	.w8(32'hbb26797b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73e16b),
	.w1(32'hbaca5adb),
	.w2(32'hbc1c79d2),
	.w3(32'hbb2bd035),
	.w4(32'hba0cf1db),
	.w5(32'hbbdf57af),
	.w6(32'h3a96432d),
	.w7(32'h3d390736),
	.w8(32'h3d4b9efa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bd457),
	.w1(32'hbc5b65b4),
	.w2(32'h3a466a9f),
	.w3(32'hbb3d1a29),
	.w4(32'h3aa8e7f7),
	.w5(32'hbb1ab479),
	.w6(32'h3b48d7ac),
	.w7(32'hbc5c4758),
	.w8(32'h3bf1be2f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc155345),
	.w1(32'hbc06ac83),
	.w2(32'h3c7e9c43),
	.w3(32'hbbef8a02),
	.w4(32'hbb993fdf),
	.w5(32'hbcec9ddf),
	.w6(32'h3b650441),
	.w7(32'h3d0b9426),
	.w8(32'hbd1f5776),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d5d95),
	.w1(32'hbc7fe825),
	.w2(32'h3cc2337f),
	.w3(32'hbc346958),
	.w4(32'hbad08727),
	.w5(32'hbc827ea2),
	.w6(32'hbc4481a1),
	.w7(32'h3c0cfd8c),
	.w8(32'hbcc1abfb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43b4d3),
	.w1(32'hbca23855),
	.w2(32'h3ac4112d),
	.w3(32'hbc20c5d5),
	.w4(32'h3b9f3f37),
	.w5(32'hbbacab5d),
	.w6(32'hbc902073),
	.w7(32'h3b92aa0d),
	.w8(32'hb9f4276e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8455bb),
	.w1(32'h3c4c757f),
	.w2(32'hbce8fc99),
	.w3(32'hbd3c09ed),
	.w4(32'h3d30ad21),
	.w5(32'h3b9421e8),
	.w6(32'hbd68a6ca),
	.w7(32'h3d00dd59),
	.w8(32'hbc2a6bb7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c8127),
	.w1(32'hbbb3dcc2),
	.w2(32'hbcbd5aff),
	.w3(32'hbc979122),
	.w4(32'hbc0dfdd3),
	.w5(32'h3c0f5cfd),
	.w6(32'hbc74afce),
	.w7(32'hbc93fa87),
	.w8(32'h3c28a7a3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab3628),
	.w1(32'h3c48b14f),
	.w2(32'hbb937a55),
	.w3(32'h3be2a69e),
	.w4(32'hbc552055),
	.w5(32'hbca262a9),
	.w6(32'h3c9aeccf),
	.w7(32'h3c41f951),
	.w8(32'hbb864281),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc736468),
	.w1(32'hbbb7c1c1),
	.w2(32'hbba67176),
	.w3(32'hbc52316d),
	.w4(32'h3bdde4bc),
	.w5(32'hbbca92fd),
	.w6(32'hbbf4f7ef),
	.w7(32'h3bc106ec),
	.w8(32'h3b950885),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b770f89),
	.w1(32'h3a9a9235),
	.w2(32'hbd004b6d),
	.w3(32'h3c01edd6),
	.w4(32'hbbbc1845),
	.w5(32'hbc221d72),
	.w6(32'h3c02bf0e),
	.w7(32'hba056d21),
	.w8(32'hbc3a743e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6a570),
	.w1(32'hbbf434be),
	.w2(32'hbc32804d),
	.w3(32'hbc7d824a),
	.w4(32'h3c092e26),
	.w5(32'hbc3e19ad),
	.w6(32'hbbd890a3),
	.w7(32'h3c297984),
	.w8(32'hbca59855),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5af294),
	.w1(32'hbbf5bcde),
	.w2(32'h3bc83d75),
	.w3(32'hbc508d6c),
	.w4(32'hbba34808),
	.w5(32'h3b74a470),
	.w6(32'hbc37304b),
	.w7(32'hbbfcc2c5),
	.w8(32'hbac933a4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c328d78),
	.w1(32'hb9202309),
	.w2(32'hbc62d659),
	.w3(32'h3c8777ed),
	.w4(32'h3b5484a4),
	.w5(32'hbc6eede2),
	.w6(32'h3c878ce0),
	.w7(32'h3c509e49),
	.w8(32'hbb960108),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a9684),
	.w1(32'hbccb40e8),
	.w2(32'hbaa9ec47),
	.w3(32'hbc35c2da),
	.w4(32'h3cf94f74),
	.w5(32'hbbc8aaee),
	.w6(32'hbc315ec1),
	.w7(32'h3c6f2bcf),
	.w8(32'hbbb861ed),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e5fbc),
	.w1(32'hbc8b6bd7),
	.w2(32'h3cdf5887),
	.w3(32'hbc6c80f6),
	.w4(32'h3d13aaaf),
	.w5(32'hbcbe2033),
	.w6(32'hbcad2892),
	.w7(32'h3d96b699),
	.w8(32'hbcee3b1a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0cfea0),
	.w1(32'hbd22f2d0),
	.w2(32'h3ac5b592),
	.w3(32'hbd71a316),
	.w4(32'h3c005dd2),
	.w5(32'h3d0e84d6),
	.w6(32'hbd8539ec),
	.w7(32'h3cd1a1ec),
	.w8(32'h3cfe6b19),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd92e906),
	.w1(32'hbd14673b),
	.w2(32'hbd7291c8),
	.w3(32'hbd10e389),
	.w4(32'hbd17653f),
	.w5(32'hbbc693ec),
	.w6(32'hbcccb364),
	.w7(32'hbdc86d7e),
	.w8(32'hbd00b14b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc060754),
	.w1(32'h3d2a00c6),
	.w2(32'hba050141),
	.w3(32'h3ce9a17d),
	.w4(32'h394e3b91),
	.w5(32'h3c5a524e),
	.w6(32'h3cee828c),
	.w7(32'h3cc93b36),
	.w8(32'hbc4a7ae8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc241c84),
	.w1(32'hbc4854b0),
	.w2(32'hbbf896ae),
	.w3(32'hbc0c54a4),
	.w4(32'h3b84c474),
	.w5(32'hbb98ff8b),
	.w6(32'hbc5b1803),
	.w7(32'hba38caae),
	.w8(32'hbbc434a8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab93e7c),
	.w1(32'hbb1428b6),
	.w2(32'hbb5c23cc),
	.w3(32'hbba6407b),
	.w4(32'h3c27552c),
	.w5(32'h3a939aca),
	.w6(32'hb960c306),
	.w7(32'h3b847af2),
	.w8(32'h3b0dc2f6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb485e3),
	.w1(32'hbc2415f7),
	.w2(32'hbc0c1b81),
	.w3(32'hbbd8aa85),
	.w4(32'h3d118cc3),
	.w5(32'hbc7c3912),
	.w6(32'hbd06aef7),
	.w7(32'h3d07e872),
	.w8(32'hbcaa0c10),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64f02f),
	.w1(32'hbc894088),
	.w2(32'hbc296ab9),
	.w3(32'hbcce2ec6),
	.w4(32'hbb50a743),
	.w5(32'hb9c69185),
	.w6(32'hbcb7f26d),
	.w7(32'hbb087799),
	.w8(32'hb953e66c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce14512),
	.w1(32'hbc42d25b),
	.w2(32'hbccfd85e),
	.w3(32'hbcff0da6),
	.w4(32'h3b56578c),
	.w5(32'h3cac1d46),
	.w6(32'hbc467bcd),
	.w7(32'hbc3c556d),
	.w8(32'h3bd4a4f6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45c6ac),
	.w1(32'hbb0fa861),
	.w2(32'h3ba503a0),
	.w3(32'h3be852da),
	.w4(32'h3ba9b1cc),
	.w5(32'hbbf93ff1),
	.w6(32'h3c01d4fd),
	.w7(32'h3bfaeb13),
	.w8(32'h3b8c464e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc629444),
	.w1(32'hbb3b8a00),
	.w2(32'hbb2bb742),
	.w3(32'hbc5ade10),
	.w4(32'hb9dd59ba),
	.w5(32'hbc2eca4d),
	.w6(32'hbc186bed),
	.w7(32'hbc79f1d4),
	.w8(32'h3c768fd6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee864b),
	.w1(32'h3c802b0f),
	.w2(32'h3c069fe9),
	.w3(32'hbc446b56),
	.w4(32'hbbf3565e),
	.w5(32'hbc872465),
	.w6(32'h3b385691),
	.w7(32'h3cbd5f2b),
	.w8(32'hbc4ed0d6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc703cdf),
	.w1(32'h3afbb7cf),
	.w2(32'h3b7c0c8f),
	.w3(32'hbca51a2b),
	.w4(32'h3bf24fbd),
	.w5(32'h3c3e4c2d),
	.w6(32'hbc738c25),
	.w7(32'h3bb64609),
	.w8(32'h3b9b972a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd269358),
	.w1(32'hbb643ac1),
	.w2(32'hbbc78d9f),
	.w3(32'hbc8a8f7e),
	.w4(32'h3cfa1af8),
	.w5(32'hbb33606e),
	.w6(32'hbc33c060),
	.w7(32'h3d4d543f),
	.w8(32'hbb799033),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47538b),
	.w1(32'hbb94341c),
	.w2(32'hbb31c514),
	.w3(32'h39cd62b9),
	.w4(32'hbb6e4c61),
	.w5(32'hbc1b52e0),
	.w6(32'hbc0a44d6),
	.w7(32'hbab9ee90),
	.w8(32'hbc6a1bcc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5b0d8),
	.w1(32'hbb45013e),
	.w2(32'h3b844a20),
	.w3(32'h3b7beb5c),
	.w4(32'h39b44cf7),
	.w5(32'h3c27ba85),
	.w6(32'h3b542ec1),
	.w7(32'hbc1cf295),
	.w8(32'h3bba3ea0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7d671),
	.w1(32'h3c21e284),
	.w2(32'hbc2ab030),
	.w3(32'h3ba1c6f6),
	.w4(32'hbc967e64),
	.w5(32'hbc5ec3b3),
	.w6(32'h3b4c1671),
	.w7(32'hbc2bf74b),
	.w8(32'hbc415167),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd47ef2),
	.w1(32'hbb495331),
	.w2(32'h3b5440a6),
	.w3(32'hbc938609),
	.w4(32'h3c896822),
	.w5(32'h3bd9d425),
	.w6(32'hbc73cd2f),
	.w7(32'h3d149964),
	.w8(32'hbb6ca41b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13d834),
	.w1(32'hbb4cad0e),
	.w2(32'h3b01d456),
	.w3(32'hbbb9c594),
	.w4(32'h392f6b8d),
	.w5(32'hb9c3c559),
	.w6(32'hbcbbf309),
	.w7(32'hbca97c0d),
	.w8(32'hbcaa090b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f0e2c),
	.w1(32'h3bfabc85),
	.w2(32'hbbdf0b8d),
	.w3(32'h3a3f7440),
	.w4(32'hbc620047),
	.w5(32'hbc555236),
	.w6(32'hbb343e56),
	.w7(32'hbbed8b79),
	.w8(32'hbc3c7b30),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e0e68),
	.w1(32'hbcbebc18),
	.w2(32'hbc81bcb8),
	.w3(32'h3a9e2000),
	.w4(32'h3ca5bd58),
	.w5(32'h3b3cb595),
	.w6(32'hbd03fc95),
	.w7(32'h3b54eaf0),
	.w8(32'hbc26ec3f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad45ec),
	.w1(32'hbb999059),
	.w2(32'hbc93740a),
	.w3(32'hbc5d5a2e),
	.w4(32'hbbb70dab),
	.w5(32'hbc3ffd7a),
	.w6(32'h3b2694a9),
	.w7(32'hbb1c9f71),
	.w8(32'h3c5226d3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53a756),
	.w1(32'hba40b208),
	.w2(32'hbb911086),
	.w3(32'hbc449f7e),
	.w4(32'h3c6aa66a),
	.w5(32'hbc45224f),
	.w6(32'hbbda424e),
	.w7(32'h3b3741b8),
	.w8(32'hbca37bb7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1d91),
	.w1(32'hbbb9f2fa),
	.w2(32'h3c5bdf09),
	.w3(32'h3c0dfca1),
	.w4(32'h3b444728),
	.w5(32'h3c96eb6f),
	.w6(32'hbaef6d70),
	.w7(32'hbc832945),
	.w8(32'hbc491c0b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd022e2),
	.w1(32'hbcaa1789),
	.w2(32'hbd1cc559),
	.w3(32'h3c1b1174),
	.w4(32'h3ca5c617),
	.w5(32'h3c1231f6),
	.w6(32'hbc08c12d),
	.w7(32'h3b8fd17b),
	.w8(32'h3c9c5642),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc773ed7),
	.w1(32'h3c2ec4dd),
	.w2(32'h3b9ff9da),
	.w3(32'h3c47eba3),
	.w4(32'h3ca827ee),
	.w5(32'hbc9b029d),
	.w6(32'h3c89b97e),
	.w7(32'h3d4acfdc),
	.w8(32'hbc337fa9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc656e0c),
	.w1(32'hbcb5467f),
	.w2(32'hbc5db49f),
	.w3(32'hbcb26f2b),
	.w4(32'h3bb16648),
	.w5(32'hbbf9f294),
	.w6(32'hbcb99a25),
	.w7(32'hbc8bdc5a),
	.w8(32'hbbdc031c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba898df8),
	.w1(32'hb98652a1),
	.w2(32'hbb6c752e),
	.w3(32'hba9e8683),
	.w4(32'hbb116bbd),
	.w5(32'hbaf34c04),
	.w6(32'h3bacf25b),
	.w7(32'hbb13047e),
	.w8(32'h3b516f83),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c06c6),
	.w1(32'h3c13ff0c),
	.w2(32'hbc2648ca),
	.w3(32'hbb842ffb),
	.w4(32'h3bf0df15),
	.w5(32'hb9cefad6),
	.w6(32'hbb928292),
	.w7(32'h3bb41865),
	.w8(32'hba560268),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b83fc),
	.w1(32'hbb4ffb48),
	.w2(32'hbc0199ea),
	.w3(32'hbc038bc3),
	.w4(32'hba826999),
	.w5(32'hbb371e80),
	.w6(32'hbb5132ea),
	.w7(32'hbbe3eb29),
	.w8(32'hbc37b01c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fac8ad),
	.w1(32'h3ac977aa),
	.w2(32'h399d3351),
	.w3(32'hb9bbb92d),
	.w4(32'hbb869500),
	.w5(32'hbb2ca7dc),
	.w6(32'h3a062ff2),
	.w7(32'hbab5eb14),
	.w8(32'hbad0fe19),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb155dfb),
	.w1(32'hbab94ad0),
	.w2(32'hbbdfb7db),
	.w3(32'hbb0099b6),
	.w4(32'hbbf8ac5e),
	.w5(32'hbbad06af),
	.w6(32'hbacd47b9),
	.w7(32'hbc45ad40),
	.w8(32'hbc5e8db8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1794b4),
	.w1(32'hbcb2b133),
	.w2(32'hbc868fb7),
	.w3(32'hbc315e7b),
	.w4(32'hbb0608d0),
	.w5(32'hbb55868b),
	.w6(32'hbca1d1b9),
	.w7(32'hbbb255a8),
	.w8(32'hbb85f88a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce188c3),
	.w1(32'hba71b106),
	.w2(32'hbc09ceab),
	.w3(32'hbc53d9b6),
	.w4(32'h3bb26bf7),
	.w5(32'hbb1c3ad6),
	.w6(32'hbcb00912),
	.w7(32'h3a97b722),
	.w8(32'hbbd23a9b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9a7ddd),
	.w1(32'hbb9ff8b4),
	.w2(32'hba3f0775),
	.w3(32'hbd56a4b9),
	.w4(32'h3ce4b8eb),
	.w5(32'h3c151b91),
	.w6(32'hbd991e5d),
	.w7(32'h3bd3c045),
	.w8(32'h3b622f89),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd64fa),
	.w1(32'h3b37d009),
	.w2(32'hbcb01ec4),
	.w3(32'hbc173ad1),
	.w4(32'h3cf24ce7),
	.w5(32'h3c5f0a4a),
	.w6(32'hbcaa7f80),
	.w7(32'h3c8de24b),
	.w8(32'h3aa04861),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fdb75),
	.w1(32'hbb92cc08),
	.w2(32'hbc942066),
	.w3(32'h3c8a2e16),
	.w4(32'h3c15e46c),
	.w5(32'h3bfbaf0e),
	.w6(32'h3c151360),
	.w7(32'h3b4ff790),
	.w8(32'hbb81a40b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c336a),
	.w1(32'h3ae5dc45),
	.w2(32'h3b0b92a8),
	.w3(32'h3c2bcbfe),
	.w4(32'h3bf7742c),
	.w5(32'h3b0bd8da),
	.w6(32'h3c3df1d6),
	.w7(32'h3c1ab9d1),
	.w8(32'h3b8dc288),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a7968),
	.w1(32'h3bffb688),
	.w2(32'hbb99e2d3),
	.w3(32'h3bc02920),
	.w4(32'hbb314e86),
	.w5(32'h3b17808e),
	.w6(32'h3c1c41e4),
	.w7(32'hbb4c2921),
	.w8(32'hb9a97641),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d69a9a),
	.w1(32'h3a5fe326),
	.w2(32'hbb86fddc),
	.w3(32'hb936df38),
	.w4(32'hbc209ba6),
	.w5(32'hbc608659),
	.w6(32'hb9c916f6),
	.w7(32'hbc39897b),
	.w8(32'hbc97a558),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3a09c),
	.w1(32'hbbc8feb9),
	.w2(32'h3c98b1ef),
	.w3(32'h3aa819c1),
	.w4(32'hbb2a9131),
	.w5(32'hbbb09580),
	.w6(32'hbb77b643),
	.w7(32'h3c2ff7f2),
	.w8(32'h38a18fa1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87c71d),
	.w1(32'h3b8a5e31),
	.w2(32'h3a54df26),
	.w3(32'h3b389ba4),
	.w4(32'hbabe38fb),
	.w5(32'hbb6c81d7),
	.w6(32'h3b05152f),
	.w7(32'h3bb9f6d1),
	.w8(32'hbb4d6000),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06a2be),
	.w1(32'h3b642745),
	.w2(32'h3c1ef058),
	.w3(32'h3af8b2d9),
	.w4(32'hba98a006),
	.w5(32'hbbbba29a),
	.w6(32'hbb9c25c1),
	.w7(32'h3abcebf1),
	.w8(32'hbc1d656e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd072b4b),
	.w1(32'hbc636271),
	.w2(32'hbac86358),
	.w3(32'hbca2447a),
	.w4(32'hbb90757d),
	.w5(32'hbc0c17a1),
	.w6(32'hbce1b403),
	.w7(32'h3af840db),
	.w8(32'h3b61311d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b437b),
	.w1(32'h3b56e873),
	.w2(32'hbc24faab),
	.w3(32'hbba863c5),
	.w4(32'hbaa3c06f),
	.w5(32'h3ae5078c),
	.w6(32'hba8e1fd8),
	.w7(32'h3b064a7d),
	.w8(32'h3adf9c00),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc304b53),
	.w1(32'hbb94267c),
	.w2(32'hbb0f7a06),
	.w3(32'h39aeb5be),
	.w4(32'h3b4cde0e),
	.w5(32'h3b368911),
	.w6(32'hbb0348e5),
	.w7(32'h3b1d6df3),
	.w8(32'h3b2f90d8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57f680),
	.w1(32'hba8b99e0),
	.w2(32'hbc044e89),
	.w3(32'hbb49eb8f),
	.w4(32'h3b0964f7),
	.w5(32'h3b1fb249),
	.w6(32'hbb6a2651),
	.w7(32'hbbed4eac),
	.w8(32'hbb85691c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd39491),
	.w1(32'hbbedec87),
	.w2(32'hbc623535),
	.w3(32'hb977dd82),
	.w4(32'h3ce14fc2),
	.w5(32'h3cf2c491),
	.w6(32'hbb86ef01),
	.w7(32'h3c3ca508),
	.w8(32'h3cd0958b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67729a),
	.w1(32'h3ce569d9),
	.w2(32'hbc492678),
	.w3(32'h3c090393),
	.w4(32'hbbf51ab5),
	.w5(32'hba6f1bb0),
	.w6(32'h3cc76d56),
	.w7(32'hbbd029cc),
	.w8(32'hbc29cf14),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2291ad),
	.w1(32'hbc7b324d),
	.w2(32'h38909ee0),
	.w3(32'h3a9a29e0),
	.w4(32'hbb6cb8b2),
	.w5(32'hbb91f6c8),
	.w6(32'hbc5a66e3),
	.w7(32'hbb80fa60),
	.w8(32'hba9ee498),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eac30),
	.w1(32'h3b8e3aad),
	.w2(32'h3b7b3c54),
	.w3(32'hbac68eae),
	.w4(32'h3c498d79),
	.w5(32'h3b211b7f),
	.w6(32'h3b5c3a76),
	.w7(32'h3cc470f0),
	.w8(32'h3d0562cd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca50acc),
	.w1(32'h3d29eea4),
	.w2(32'h3b298467),
	.w3(32'h3c040cdf),
	.w4(32'h3b977750),
	.w5(32'h3ba54174),
	.w6(32'h3d344b5b),
	.w7(32'hbb93ec62),
	.w8(32'h3b002bcd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c032850),
	.w1(32'h3c185fe0),
	.w2(32'h3b222438),
	.w3(32'h3c322d75),
	.w4(32'h3a7cbfdd),
	.w5(32'hbabbcefe),
	.w6(32'h3c0a589e),
	.w7(32'h3bea2796),
	.w8(32'h3b14d44f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83c984),
	.w1(32'hbac70f9d),
	.w2(32'h3ba72747),
	.w3(32'h3b590b8d),
	.w4(32'h3a4984de),
	.w5(32'hbb518f4a),
	.w6(32'h3b23960e),
	.w7(32'h3b6a2cb6),
	.w8(32'hbb8c272e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1e2db),
	.w1(32'hbc09c428),
	.w2(32'hbb1765c8),
	.w3(32'hbca68c79),
	.w4(32'h3b80b248),
	.w5(32'h3b7c2977),
	.w6(32'hbcb0375d),
	.w7(32'hb9b553de),
	.w8(32'h3acd1a64),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d0e4a),
	.w1(32'h3b4dbedd),
	.w2(32'hbb7afaa1),
	.w3(32'hbbbf20c0),
	.w4(32'hb9a83557),
	.w5(32'hbabd123d),
	.w6(32'hbc0813c6),
	.w7(32'hbb0d68b7),
	.w8(32'hbc0cda41),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96a6f7),
	.w1(32'hbb121f06),
	.w2(32'hbb726ac1),
	.w3(32'h3c05a4bd),
	.w4(32'h3c86c74a),
	.w5(32'h3ba4bc98),
	.w6(32'hbbaadfd8),
	.w7(32'h3b859a2f),
	.w8(32'hbc66bdc4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb36b7f),
	.w1(32'hbb209c22),
	.w2(32'hbc8c0620),
	.w3(32'h3c1eb81b),
	.w4(32'hbc4252bf),
	.w5(32'hbc037c1b),
	.w6(32'hba4e07ff),
	.w7(32'hbb311fd8),
	.w8(32'hbab77f4f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce25c4),
	.w1(32'h3a9d3422),
	.w2(32'hbbddeb35),
	.w3(32'hbc90e407),
	.w4(32'h3bb79160),
	.w5(32'h3ab63e86),
	.w6(32'h3a53c9be),
	.w7(32'h3b91cd5a),
	.w8(32'h3b9953f0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81f95e),
	.w1(32'h3c385230),
	.w2(32'hbb9220ba),
	.w3(32'hbb14b9c3),
	.w4(32'h3a8cb0a6),
	.w5(32'hbb5b02ab),
	.w6(32'h3c0ed92c),
	.w7(32'hba10eebe),
	.w8(32'hbc040b41),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3da642),
	.w1(32'hbc1a93df),
	.w2(32'hbc0ef43a),
	.w3(32'h3c0577c3),
	.w4(32'hbb4ae4c4),
	.w5(32'hbbd65ac0),
	.w6(32'h3c0a378e),
	.w7(32'h3c03426e),
	.w8(32'h3bb2dbc6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd49f930),
	.w1(32'hbc06cb05),
	.w2(32'hbb14f1db),
	.w3(32'hbd031a5b),
	.w4(32'h3bf2d80e),
	.w5(32'h3bfddd8b),
	.w6(32'hbceeddbf),
	.w7(32'h3bb2f272),
	.w8(32'h3c3b3dcd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb333e4),
	.w1(32'h3b19e4c4),
	.w2(32'hbc0186a9),
	.w3(32'hbcb676c2),
	.w4(32'hbb59c31b),
	.w5(32'hbb8d49c5),
	.w6(32'hbca01fae),
	.w7(32'h3bd747bd),
	.w8(32'h3b8709e8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2b3c0),
	.w1(32'h3c9beec0),
	.w2(32'hbc3584f9),
	.w3(32'h3bc08729),
	.w4(32'h3b2d5854),
	.w5(32'hbbc80daa),
	.w6(32'h3c749466),
	.w7(32'hbc24dc81),
	.w8(32'hbcbe54af),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc213c83),
	.w1(32'hbc178d46),
	.w2(32'hbb7909d8),
	.w3(32'hbbca0a0d),
	.w4(32'hbc255a2b),
	.w5(32'hbbb0bf42),
	.w6(32'hbc1ab392),
	.w7(32'hbc3fa084),
	.w8(32'hbc68da6a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b5f3),
	.w1(32'hbbe6fe6f),
	.w2(32'h39df8793),
	.w3(32'h3b1db686),
	.w4(32'h3ac9f59d),
	.w5(32'hba4e121a),
	.w6(32'hbc22e6ad),
	.w7(32'h3baec524),
	.w8(32'h3bd8631a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a2410),
	.w1(32'h3b5043d9),
	.w2(32'hbc406c47),
	.w3(32'h3bccbdef),
	.w4(32'hbc6b69f5),
	.w5(32'hbc77c16f),
	.w6(32'h3c4bce91),
	.w7(32'hbc8b8bb8),
	.w8(32'hbce3975a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd32f088),
	.w1(32'hbd14bf9f),
	.w2(32'hbbdeda39),
	.w3(32'hbcedd869),
	.w4(32'h3b75a742),
	.w5(32'hba969b88),
	.w6(32'hbd35e43b),
	.w7(32'hbb06834f),
	.w8(32'h3a722b8e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f9f0f),
	.w1(32'h3b3a8f5e),
	.w2(32'hbc3cd229),
	.w3(32'hbbb125f7),
	.w4(32'h3b016bfd),
	.w5(32'hbb6782b5),
	.w6(32'hbc666b0a),
	.w7(32'hba877f91),
	.w8(32'hbb2f0508),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30353c),
	.w1(32'h3bb12880),
	.w2(32'h3ba46401),
	.w3(32'hb757a528),
	.w4(32'h3aaf7c38),
	.w5(32'hbaf567fb),
	.w6(32'h3bd5991b),
	.w7(32'h3b97ffd2),
	.w8(32'hbb12ccc6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec9228),
	.w1(32'h3acacfa9),
	.w2(32'hbb2877ef),
	.w3(32'h39d3b0e8),
	.w4(32'hb9449e31),
	.w5(32'h3b070394),
	.w6(32'hbb61040d),
	.w7(32'h3ae7a59e),
	.w8(32'h3ab03d12),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8edad5),
	.w1(32'hbbb8ddb4),
	.w2(32'hbc311925),
	.w3(32'h3bccfcae),
	.w4(32'h3c2ed068),
	.w5(32'h3b98e2be),
	.w6(32'h3b8a43b4),
	.w7(32'h3b02ceb7),
	.w8(32'hb924a0af),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf24ba),
	.w1(32'hbc014543),
	.w2(32'h3c0f031b),
	.w3(32'h3b6ec86a),
	.w4(32'hbc78c177),
	.w5(32'hbc4f66c0),
	.w6(32'hbbd08812),
	.w7(32'hbade8b3d),
	.w8(32'hbb8ec3ae),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaefd7d),
	.w1(32'hbb213894),
	.w2(32'hbbd8c0cf),
	.w3(32'hbb9284cb),
	.w4(32'hbbd36fe2),
	.w5(32'hbbb48d01),
	.w6(32'h3bae3036),
	.w7(32'hbbfa800d),
	.w8(32'hbb027003),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144f2a),
	.w1(32'h3c13d9da),
	.w2(32'hbacc296a),
	.w3(32'h3acef842),
	.w4(32'h3bd21038),
	.w5(32'h3b0e67bf),
	.w6(32'h3c176680),
	.w7(32'h3b784c39),
	.w8(32'h3a4dafc3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bf59d),
	.w1(32'hbb432995),
	.w2(32'hbc3f480a),
	.w3(32'h3ade6367),
	.w4(32'hbb545c30),
	.w5(32'hbadde299),
	.w6(32'h3a717ba9),
	.w7(32'h3b7b2e74),
	.w8(32'h3b2a7314),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70f132),
	.w1(32'h3c029496),
	.w2(32'h385ce3cc),
	.w3(32'hbbaf569a),
	.w4(32'h3b1144b7),
	.w5(32'hbb58b52d),
	.w6(32'h3b987be6),
	.w7(32'hba2f4607),
	.w8(32'hbc0abbad),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17f275),
	.w1(32'hbb689467),
	.w2(32'hbc329615),
	.w3(32'h3b942480),
	.w4(32'hbaf88181),
	.w5(32'hba79c075),
	.w6(32'hbb8c1202),
	.w7(32'hbb428bab),
	.w8(32'h3ae088ee),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac31e1c),
	.w1(32'hb92a7210),
	.w2(32'hbb50ed1d),
	.w3(32'hbb9c6af2),
	.w4(32'hba45f900),
	.w5(32'h3b1e256f),
	.w6(32'hbbde1b5b),
	.w7(32'hbba1edb8),
	.w8(32'hba0f0351),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule