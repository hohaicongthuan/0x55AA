module layer_6_featuremap_61(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3a0205),
	.w1(32'h3b5557dd),
	.w2(32'h3c456be7),
	.w3(32'hbbd6cfaa),
	.w4(32'hbb2efe46),
	.w5(32'hbb8e28ec),
	.w6(32'hbaf3d8d4),
	.w7(32'h3bedbed1),
	.w8(32'h3b6924c5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed41d7),
	.w1(32'hba6bba41),
	.w2(32'hb821a79a),
	.w3(32'h3ab741bd),
	.w4(32'h3b930d66),
	.w5(32'h3b694469),
	.w6(32'h3c374303),
	.w7(32'h3c348699),
	.w8(32'h3c445ecb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17338f),
	.w1(32'hbc219ce5),
	.w2(32'hbc28f0da),
	.w3(32'hbc7c8b65),
	.w4(32'hbc5984d4),
	.w5(32'hbbe65899),
	.w6(32'hbc3edf10),
	.w7(32'hbae18012),
	.w8(32'h3ab95287),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2304bb),
	.w1(32'hbafbe8a1),
	.w2(32'hbc1fbed6),
	.w3(32'h3bad3f19),
	.w4(32'h3ba795be),
	.w5(32'h3b22db73),
	.w6(32'h3b1040d7),
	.w7(32'hbb580341),
	.w8(32'hbbab3f5f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b6874),
	.w1(32'hbbd0ccdc),
	.w2(32'h3bbc6f45),
	.w3(32'hbb48645b),
	.w4(32'h39bba466),
	.w5(32'h3acc8c26),
	.w6(32'hbb4e83e3),
	.w7(32'hbaa0a06b),
	.w8(32'hbc1b0311),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7edb56),
	.w1(32'h3c93d81c),
	.w2(32'h3ce21a80),
	.w3(32'hbbf2f56b),
	.w4(32'hbb7282d4),
	.w5(32'h39c8aaf4),
	.w6(32'h3c072385),
	.w7(32'h3c8f1163),
	.w8(32'h3c99c35a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce7cb54),
	.w1(32'hbce41fe1),
	.w2(32'hbd31210d),
	.w3(32'h3c16c073),
	.w4(32'h3b32b558),
	.w5(32'h3a89c9ee),
	.w6(32'hbc554ffc),
	.w7(32'hbcdf6cb3),
	.w8(32'hbcb6623a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd12e1f9),
	.w1(32'h3bfbb3fb),
	.w2(32'h3bc872cb),
	.w3(32'hbb86ab7e),
	.w4(32'hbc7c710c),
	.w5(32'hbc53862a),
	.w6(32'h3bc07a58),
	.w7(32'h3b529974),
	.w8(32'hbb003d9e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b265307),
	.w1(32'h3c66fc17),
	.w2(32'h3a68cf9d),
	.w3(32'hb9c53c12),
	.w4(32'hbae84bff),
	.w5(32'h3a357742),
	.w6(32'h3c23e22c),
	.w7(32'h3ca762d0),
	.w8(32'h3b615221),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f48d9),
	.w1(32'h3cc12fcf),
	.w2(32'h3cfc102f),
	.w3(32'hb9fa00c3),
	.w4(32'h3b98beed),
	.w5(32'h3b3cd565),
	.w6(32'h3c8726d1),
	.w7(32'h3cc95c15),
	.w8(32'h3c9cba93),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc29383),
	.w1(32'hbbb335ac),
	.w2(32'hbacf9ffa),
	.w3(32'h3b73f8b9),
	.w4(32'h3b64a98a),
	.w5(32'h3be8980d),
	.w6(32'hbbe34217),
	.w7(32'h3b94bfee),
	.w8(32'h3c2b9090),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa9078),
	.w1(32'h3a09ed35),
	.w2(32'h3c0e4026),
	.w3(32'hbbc25ad5),
	.w4(32'hbbba1992),
	.w5(32'hbbf93896),
	.w6(32'hbb5532ce),
	.w7(32'h3a74f979),
	.w8(32'h3b79f739),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33d673),
	.w1(32'hbba4f7b8),
	.w2(32'hbbd6081b),
	.w3(32'h3bec7441),
	.w4(32'h3c0555eb),
	.w5(32'h3b55c803),
	.w6(32'h3b8f0d64),
	.w7(32'h3b81f5e3),
	.w8(32'hb979081e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc179b48),
	.w1(32'h3b38e2b4),
	.w2(32'h3c2c4430),
	.w3(32'h3c617999),
	.w4(32'h3c287352),
	.w5(32'h3be778ea),
	.w6(32'h3c57e82a),
	.w7(32'h3c4bdd2f),
	.w8(32'h3c0ef682),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b7d1b),
	.w1(32'hbbb9e939),
	.w2(32'hbba166f6),
	.w3(32'h393facea),
	.w4(32'h3b9efa63),
	.w5(32'h3babbe0e),
	.w6(32'hbb3df562),
	.w7(32'hbab036f4),
	.w8(32'hbbee382d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfff44d),
	.w1(32'h3b8d9848),
	.w2(32'h3be3f27b),
	.w3(32'hbb1c6097),
	.w4(32'hbb434520),
	.w5(32'hbb35aefa),
	.w6(32'hba2b8623),
	.w7(32'h3a911888),
	.w8(32'h3b02e1ca),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f6095),
	.w1(32'h3bacf1a4),
	.w2(32'hba86731a),
	.w3(32'h3b28e2b9),
	.w4(32'h3b196d74),
	.w5(32'hbb92f251),
	.w6(32'h399df4e0),
	.w7(32'hbb927ff3),
	.w8(32'hbc808ecd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c46c3),
	.w1(32'h3ba5a22d),
	.w2(32'h3c36e9e7),
	.w3(32'hba6a6263),
	.w4(32'h3b96332f),
	.w5(32'h3ac85b77),
	.w6(32'h3ac93661),
	.w7(32'h3c099055),
	.w8(32'h3b9ce5d2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c237152),
	.w1(32'h3b057f3c),
	.w2(32'hbaf4bb52),
	.w3(32'hbb59d545),
	.w4(32'hbbd0aef8),
	.w5(32'hbbbcadc0),
	.w6(32'hb9d02bcc),
	.w7(32'hbba29138),
	.w8(32'hbba8aa32),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49f72b),
	.w1(32'hbb2a2e0f),
	.w2(32'hbbb2a0c8),
	.w3(32'h3b643db4),
	.w4(32'hbbad24d3),
	.w5(32'hbbbe8ee6),
	.w6(32'hba720ad5),
	.w7(32'hbb009651),
	.w8(32'hbb71f04d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e0540),
	.w1(32'hbb6c4305),
	.w2(32'hbbd25c16),
	.w3(32'h3a4e65a7),
	.w4(32'h3b195e45),
	.w5(32'h3b3f3dda),
	.w6(32'hbb3cf131),
	.w7(32'hbb7e57aa),
	.w8(32'hbb365b37),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d4ed),
	.w1(32'h3a4e287e),
	.w2(32'h3a8f86f1),
	.w3(32'h39418e9c),
	.w4(32'h3bcb9e66),
	.w5(32'h3c1283aa),
	.w6(32'h3b1fcb32),
	.w7(32'h3bbb51e3),
	.w8(32'h3b8609a1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a19ac),
	.w1(32'h3b59e745),
	.w2(32'h3bd1f0f1),
	.w3(32'hbc140452),
	.w4(32'h3b1f7220),
	.w5(32'h3b7ef568),
	.w6(32'h3c09f5dc),
	.w7(32'h3c189e07),
	.w8(32'h3b8986d5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb486321),
	.w1(32'h3b8aa89b),
	.w2(32'h3ba457b6),
	.w3(32'hbaba4a33),
	.w4(32'h3b6b263e),
	.w5(32'h3c355b2e),
	.w6(32'h3cb60831),
	.w7(32'h3c9cff4b),
	.w8(32'h3c6289ff),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b078eb1),
	.w1(32'hbbef43ba),
	.w2(32'hbb74691b),
	.w3(32'hbb94c5ab),
	.w4(32'hbb771ae3),
	.w5(32'h3a1cc77f),
	.w6(32'hbc0211e7),
	.w7(32'hbb3aca06),
	.w8(32'hb9e5b463),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba118bbc),
	.w1(32'hbbafe6f8),
	.w2(32'hbab29046),
	.w3(32'h3ab91ec6),
	.w4(32'hbb4be300),
	.w5(32'h3a83278a),
	.w6(32'hbb83be43),
	.w7(32'hba2da240),
	.w8(32'hbb8d3a29),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7146cb),
	.w1(32'hbae6a274),
	.w2(32'h39806815),
	.w3(32'hba0276f3),
	.w4(32'hba9c102d),
	.w5(32'hbb155250),
	.w6(32'hbb597bd3),
	.w7(32'h3961af2b),
	.w8(32'h3b46a15f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37ab90),
	.w1(32'hbc8c42d9),
	.w2(32'hbce813ff),
	.w3(32'h3b63629e),
	.w4(32'hbb3d9205),
	.w5(32'hbafb7e72),
	.w6(32'hbc297187),
	.w7(32'hbcadde88),
	.w8(32'hbc82c9b3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6cb76),
	.w1(32'hbaa8868e),
	.w2(32'hbb33664c),
	.w3(32'h389a70b8),
	.w4(32'hba2ef0e6),
	.w5(32'h39ebd44d),
	.w6(32'hbac19a05),
	.w7(32'hbb25fb22),
	.w8(32'hba8c22d9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4e6f4),
	.w1(32'h3b0874e3),
	.w2(32'h39fef572),
	.w3(32'h3bea7ae8),
	.w4(32'h3c5fe8e8),
	.w5(32'h3b349cf2),
	.w6(32'h3c067a50),
	.w7(32'h3c0b4c68),
	.w8(32'h3c1b10f2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8b66f),
	.w1(32'hbc838593),
	.w2(32'hbcb9a932),
	.w3(32'hbab71ce6),
	.w4(32'hbc8313e9),
	.w5(32'hbc8fc6f5),
	.w6(32'hbc9f2d4a),
	.w7(32'hbd2e75b8),
	.w8(32'hbcf96a10),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3ab3c),
	.w1(32'h3b8adcf0),
	.w2(32'h3c1b913c),
	.w3(32'hbc4d70fb),
	.w4(32'hbc3f74ad),
	.w5(32'hbc29deab),
	.w6(32'hbb16de4f),
	.w7(32'h3b476d47),
	.w8(32'h3b72e88d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c890a),
	.w1(32'hbb814073),
	.w2(32'hbc8b2c60),
	.w3(32'hbb547db2),
	.w4(32'hba6aae07),
	.w5(32'hbbaf04d0),
	.w6(32'hbba58892),
	.w7(32'hbbf589a9),
	.w8(32'hbb8cb430),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44a242),
	.w1(32'h3c243e9f),
	.w2(32'h3bfbae09),
	.w3(32'h3a811728),
	.w4(32'hbb2ef17e),
	.w5(32'h3b370bea),
	.w6(32'h3c11953c),
	.w7(32'h3bee7998),
	.w8(32'hbb8a545e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b47f),
	.w1(32'h3c10ea7d),
	.w2(32'h3c3db6cf),
	.w3(32'hbc0b797f),
	.w4(32'hbbd0c6f2),
	.w5(32'hbbb1bfa4),
	.w6(32'h3b7d6421),
	.w7(32'h3be2aa70),
	.w8(32'h3bc6821d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18fe4a),
	.w1(32'hbc10fb09),
	.w2(32'hbbbe3186),
	.w3(32'hbc0162de),
	.w4(32'hbbbd3204),
	.w5(32'hbb0e3287),
	.w6(32'hbb6ba456),
	.w7(32'hbbda6572),
	.w8(32'hbbc9e89b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb71d61),
	.w1(32'h3b220a43),
	.w2(32'h3c33a5de),
	.w3(32'hbb6879ad),
	.w4(32'hbb5e3ede),
	.w5(32'hbaf91722),
	.w6(32'hb9a6b855),
	.w7(32'h3b94cec3),
	.w8(32'h3b24cbf6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f4ae),
	.w1(32'hbabbd311),
	.w2(32'hbb782b2f),
	.w3(32'h3bab2fd7),
	.w4(32'h3b7f1ee3),
	.w5(32'h3ba2ef4c),
	.w6(32'h3aa20b19),
	.w7(32'hba0d3f04),
	.w8(32'h3aa379fb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1df511),
	.w1(32'h3c0f913e),
	.w2(32'h3b974ca8),
	.w3(32'h3c0860bd),
	.w4(32'h3c71b622),
	.w5(32'h3c737369),
	.w6(32'h3c0ed9d1),
	.w7(32'h3bbc0be6),
	.w8(32'h3c1af0a3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6682),
	.w1(32'h3a457b7f),
	.w2(32'h3bc999b2),
	.w3(32'hbc246098),
	.w4(32'h3bae2810),
	.w5(32'h3c8c34ab),
	.w6(32'hbbc22f69),
	.w7(32'hba8f4683),
	.w8(32'h3bf4b13e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ba253),
	.w1(32'hbb12a36a),
	.w2(32'hbc203a78),
	.w3(32'hbc1cd4cd),
	.w4(32'h36f8eb7a),
	.w5(32'h3a5b3db3),
	.w6(32'hbbd1ad37),
	.w7(32'hbaa57035),
	.w8(32'h3c0c4f29),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3104f),
	.w1(32'hbb3a138a),
	.w2(32'hbc170ea7),
	.w3(32'h3ba36e21),
	.w4(32'h3b81b5c3),
	.w5(32'h3b3ccece),
	.w6(32'h3a503e86),
	.w7(32'hbb81fb8a),
	.w8(32'hbb58235f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be3fd),
	.w1(32'h3bd7767a),
	.w2(32'h3c60690a),
	.w3(32'hbb1cfb9e),
	.w4(32'h3abc2e64),
	.w5(32'h3ab75aee),
	.w6(32'h3b16747f),
	.w7(32'h3c3fdad9),
	.w8(32'h3c0fb042),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ff202),
	.w1(32'hbbc4e562),
	.w2(32'hbbcb481b),
	.w3(32'h3b4895ac),
	.w4(32'hbb9c5804),
	.w5(32'h3a51c934),
	.w6(32'hba224a29),
	.w7(32'hbb8cc5b7),
	.w8(32'h3bd7ef48),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b329d9),
	.w1(32'hbaa95f3b),
	.w2(32'hbad4fb14),
	.w3(32'hbaf2a6be),
	.w4(32'h3aeec90d),
	.w5(32'h3b73c8dd),
	.w6(32'hbab1439e),
	.w7(32'h3ad0fb67),
	.w8(32'h3b39abc0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb5fa6),
	.w1(32'hbbe4ef2c),
	.w2(32'h3b24de14),
	.w3(32'hbc4c33f9),
	.w4(32'h3b7399ac),
	.w5(32'h3c00de2a),
	.w6(32'hbbea2c55),
	.w7(32'h3bb8cf36),
	.w8(32'h3c5540c0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83c957),
	.w1(32'h3bf1603a),
	.w2(32'hbb1d632f),
	.w3(32'h3bc4568e),
	.w4(32'h3c246398),
	.w5(32'h3cb9d971),
	.w6(32'h3c6d65f4),
	.w7(32'h3c2d10fa),
	.w8(32'h3beff063),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc025bcf),
	.w1(32'h3aee0c03),
	.w2(32'hbb924bc2),
	.w3(32'h3ba17f19),
	.w4(32'h3bd222a0),
	.w5(32'h3c04388c),
	.w6(32'h3ba4eed7),
	.w7(32'hba82c511),
	.w8(32'hbb38c323),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda08ef),
	.w1(32'h3ae5d665),
	.w2(32'h3b16adfd),
	.w3(32'h3b270308),
	.w4(32'h3b9b3ac3),
	.w5(32'h3bdd8e3a),
	.w6(32'h3a6db3be),
	.w7(32'h3ada9df5),
	.w8(32'h3b845dc2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ad026),
	.w1(32'hbba82121),
	.w2(32'hbc3f104e),
	.w3(32'hbb540c19),
	.w4(32'hbbdf8887),
	.w5(32'hba748d82),
	.w6(32'hbc2607ab),
	.w7(32'hbc99dd43),
	.w8(32'hbc060976),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58fa95),
	.w1(32'hbb2e9606),
	.w2(32'hbc5b3113),
	.w3(32'h3c163d7f),
	.w4(32'h3c29b291),
	.w5(32'h3bff94ca),
	.w6(32'h3bcacb1c),
	.w7(32'h3a45df53),
	.w8(32'h394ff2f1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20e6a3),
	.w1(32'hbbeacb03),
	.w2(32'hbc6148a5),
	.w3(32'h3aeb72f4),
	.w4(32'hbafd1c20),
	.w5(32'h3ab048b5),
	.w6(32'hbb152d76),
	.w7(32'hbc0960e1),
	.w8(32'hbb95e8a3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36d123),
	.w1(32'hbb9964ca),
	.w2(32'hbc990d5d),
	.w3(32'h3c3dd56c),
	.w4(32'h3c35744a),
	.w5(32'h3c668352),
	.w6(32'hb7c4679c),
	.w7(32'hbc0e2b62),
	.w8(32'hbbb1d165),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f1aaa),
	.w1(32'hbcf0bc5c),
	.w2(32'hbd2a1544),
	.w3(32'h3b976aca),
	.w4(32'h3b8de214),
	.w5(32'h3c1e1954),
	.w6(32'hbc9dbb5d),
	.w7(32'hbcd2b4ab),
	.w8(32'hbc9d199f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07e4e0),
	.w1(32'hbba243f9),
	.w2(32'hbc4de95e),
	.w3(32'h3be28010),
	.w4(32'h3c261281),
	.w5(32'h3be66ff5),
	.w6(32'h3c124151),
	.w7(32'h3bde9176),
	.w8(32'h3ba9c648),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3600fc),
	.w1(32'h3b989d06),
	.w2(32'hbbdac74a),
	.w3(32'hbc5b5758),
	.w4(32'hbbcd695e),
	.w5(32'hbaf3f533),
	.w6(32'hbbbc335e),
	.w7(32'hbc458272),
	.w8(32'hbc69f21b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc052407),
	.w1(32'h3c251afb),
	.w2(32'h3cc45b88),
	.w3(32'h3855e411),
	.w4(32'h3c2a7749),
	.w5(32'hbb6e2d09),
	.w6(32'h3c7211fd),
	.w7(32'h3cffdf79),
	.w8(32'h3c51d498),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12bd69),
	.w1(32'h3ca39ba1),
	.w2(32'h3c1826d6),
	.w3(32'h3b82e915),
	.w4(32'hba4d1de6),
	.w5(32'hbbbf5cdf),
	.w6(32'h3c84d2b1),
	.w7(32'h3c24f490),
	.w8(32'h3bea5bed),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5133e),
	.w1(32'hbaf902c0),
	.w2(32'hbc238a80),
	.w3(32'h3b6e4a13),
	.w4(32'hbaed387b),
	.w5(32'h39c17f86),
	.w6(32'hbb674e61),
	.w7(32'hbc37d98d),
	.w8(32'hbbf7cc91),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99338d),
	.w1(32'hbc84d980),
	.w2(32'hbc214195),
	.w3(32'h3b554482),
	.w4(32'hbbf6ec05),
	.w5(32'hb953e202),
	.w6(32'hbbe8fdd2),
	.w7(32'hbc07b945),
	.w8(32'hbbbba284),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0386bf),
	.w1(32'h3bce8bd0),
	.w2(32'hbb3af1ea),
	.w3(32'h3c1cbb2c),
	.w4(32'h3b72562b),
	.w5(32'h3bc38729),
	.w6(32'h3b8b09f0),
	.w7(32'hbbb10f08),
	.w8(32'hbb0197c1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab881e),
	.w1(32'h3b318f92),
	.w2(32'h3c8483e6),
	.w3(32'h3b016241),
	.w4(32'h3b576c63),
	.w5(32'hbcab18cc),
	.w6(32'h3c491ad5),
	.w7(32'h3bc5f091),
	.w8(32'hbc856152),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb297d5e),
	.w1(32'hbc77d2de),
	.w2(32'hbcaa4856),
	.w3(32'h3a4dae97),
	.w4(32'h3a73c5e5),
	.w5(32'h3c1c5eb1),
	.w6(32'hbcc2d95a),
	.w7(32'hbd12f034),
	.w8(32'hbbb9a9c9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fc5d6),
	.w1(32'hbae15844),
	.w2(32'hbcf3833b),
	.w3(32'hbbc3468b),
	.w4(32'hbcccfb4b),
	.w5(32'hbc8a44b9),
	.w6(32'hbca7c78d),
	.w7(32'hbd61baf0),
	.w8(32'hbd36a583),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule