module layer_8_featuremap_196(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea5c14),
	.w1(32'h3a8d7d97),
	.w2(32'hbbb8225e),
	.w3(32'hbbee5ce7),
	.w4(32'h3bbc2b05),
	.w5(32'h3c3ab506),
	.w6(32'hbad5180c),
	.w7(32'h3bb231e6),
	.w8(32'hbc016c51),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e705d),
	.w1(32'h3ab529a5),
	.w2(32'h3b45d4a9),
	.w3(32'h3b6d6ed7),
	.w4(32'h3ac5ffb6),
	.w5(32'h3a26853a),
	.w6(32'hba9a3a46),
	.w7(32'h397e4401),
	.w8(32'hbb666798),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35a0f3),
	.w1(32'h3a55064f),
	.w2(32'hba31b85b),
	.w3(32'hb984df4f),
	.w4(32'h3a279120),
	.w5(32'h3b96292e),
	.w6(32'hbbf2da3e),
	.w7(32'hbb8b9c0f),
	.w8(32'hbb9b9d42),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9430b),
	.w1(32'hba63c884),
	.w2(32'h3c2d3499),
	.w3(32'h37328e30),
	.w4(32'hbb3d2e39),
	.w5(32'h3c1c3b8c),
	.w6(32'hbb815277),
	.w7(32'hbbd0578d),
	.w8(32'h3a55d132),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3706ad),
	.w1(32'h396411f6),
	.w2(32'hbb37cc07),
	.w3(32'h3c8a996d),
	.w4(32'h3b8db34c),
	.w5(32'h3b0ca285),
	.w6(32'hbb2e1d7a),
	.w7(32'hbb61b255),
	.w8(32'hbb65b608),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7131),
	.w1(32'hbb9f810c),
	.w2(32'hbb4e1974),
	.w3(32'h3b574763),
	.w4(32'h3b240929),
	.w5(32'h3b0a4b03),
	.w6(32'h3ac86e58),
	.w7(32'hbb9916ce),
	.w8(32'hbb0e5d3b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f53f),
	.w1(32'hbbee2bef),
	.w2(32'hbb4f1ea8),
	.w3(32'h3c336112),
	.w4(32'hbb875579),
	.w5(32'h3a0044bc),
	.w6(32'hbc222717),
	.w7(32'hbbe582c2),
	.w8(32'hbbe625d1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee33c),
	.w1(32'hba7803db),
	.w2(32'h39dee793),
	.w3(32'h3b587c49),
	.w4(32'hbc64ac3d),
	.w5(32'hbb54a6d9),
	.w6(32'hbb3dbcdb),
	.w7(32'hbb186fb0),
	.w8(32'h3a7b7be9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd52b39),
	.w1(32'hbb7747f5),
	.w2(32'hba34c06d),
	.w3(32'hbae10d2b),
	.w4(32'h39cf5afa),
	.w5(32'h3ba2173d),
	.w6(32'hbc6981a0),
	.w7(32'hbc54fd44),
	.w8(32'hbc0636da),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86d89),
	.w1(32'h3b00347b),
	.w2(32'h3bdc3455),
	.w3(32'h3c1d1a3d),
	.w4(32'h3baa7707),
	.w5(32'hba3d00c4),
	.w6(32'h3996b153),
	.w7(32'hba4360ae),
	.w8(32'hbbb4ea7a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9aa2a),
	.w1(32'hbb9e7527),
	.w2(32'h3b9035a9),
	.w3(32'hbb13ef54),
	.w4(32'hbb94940f),
	.w5(32'h3c27a055),
	.w6(32'hbc850f45),
	.w7(32'hbc2afec2),
	.w8(32'h3aa03873),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c350265),
	.w1(32'hbc3a6fb8),
	.w2(32'hbbfe8574),
	.w3(32'h3c5f99cb),
	.w4(32'hbc2b0384),
	.w5(32'hbaaa9b14),
	.w6(32'hbafe95cf),
	.w7(32'hbc1b5d92),
	.w8(32'hbc83aac3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90fe1e),
	.w1(32'h3a9a79da),
	.w2(32'hba9069d1),
	.w3(32'h3aaadaec),
	.w4(32'hb9d52861),
	.w5(32'h390d73e1),
	.w6(32'h38466b4e),
	.w7(32'h3b0754a4),
	.w8(32'h3b82ce06),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa77229),
	.w1(32'hba5d731a),
	.w2(32'h3b3f9e15),
	.w3(32'hbb713716),
	.w4(32'hbb2fcb5a),
	.w5(32'h3bd1a3fe),
	.w6(32'h3ab437da),
	.w7(32'hbb0b230a),
	.w8(32'hbba2d1b6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a7374),
	.w1(32'hbc0863ba),
	.w2(32'hbc0cff4f),
	.w3(32'h3c1629d2),
	.w4(32'hbc1788ef),
	.w5(32'hbc254c6f),
	.w6(32'hbbfaea36),
	.w7(32'hbc1cb1c0),
	.w8(32'hbc0a91cd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7e382),
	.w1(32'h3b696ab4),
	.w2(32'h3a94f0b4),
	.w3(32'hbbf7b22c),
	.w4(32'hba84ca96),
	.w5(32'h398ec983),
	.w6(32'hbbdfbbb5),
	.w7(32'hba0aa68b),
	.w8(32'h3a5d7bed),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeaedd),
	.w1(32'hb991b1d4),
	.w2(32'h3a89e9a6),
	.w3(32'h3a3221f4),
	.w4(32'hbb8cde65),
	.w5(32'h3bb41173),
	.w6(32'hb9d5516d),
	.w7(32'hbb9bd63d),
	.w8(32'hb9c382d6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab08ed8),
	.w1(32'h3ba5e031),
	.w2(32'h3aa82d1a),
	.w3(32'hba628dfd),
	.w4(32'hbaab3b9d),
	.w5(32'h3970c244),
	.w6(32'hbc1ad3b7),
	.w7(32'hbbad75bd),
	.w8(32'hbb9e9bd3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c305e34),
	.w1(32'h3bfcc2ef),
	.w2(32'h39fdac6a),
	.w3(32'h3c214d79),
	.w4(32'h3a59c0d5),
	.w5(32'h3a6f3e3c),
	.w6(32'hbba393ef),
	.w7(32'hbb7c82b1),
	.w8(32'hbb948c53),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ffc08),
	.w1(32'hba6bce54),
	.w2(32'hbb7f3b69),
	.w3(32'h3bebcf86),
	.w4(32'h3aa13684),
	.w5(32'h3af5493f),
	.w6(32'hbbabeb1a),
	.w7(32'hbbd57ffa),
	.w8(32'hbb40e596),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e806d),
	.w1(32'hbbc5fba1),
	.w2(32'h3aa0861f),
	.w3(32'h3bdcbbd9),
	.w4(32'h3aa2ea9b),
	.w5(32'h3ab76654),
	.w6(32'hbaecb433),
	.w7(32'hbb30a14a),
	.w8(32'h39912fe4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84aca8),
	.w1(32'h3a1eaa6e),
	.w2(32'h3b9f5b89),
	.w3(32'hb9a6d12f),
	.w4(32'hbaf4ca93),
	.w5(32'h3bd25445),
	.w6(32'h3890e9fd),
	.w7(32'hbb07e70e),
	.w8(32'h3ba96c20),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb47e4a),
	.w1(32'h3b062fbc),
	.w2(32'hbb1c6386),
	.w3(32'h3b65e462),
	.w4(32'h3aaa99a7),
	.w5(32'h3a490833),
	.w6(32'hbc2c3d87),
	.w7(32'hbbb1ecdf),
	.w8(32'hbb9a3162),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c462f1e),
	.w1(32'hba227f04),
	.w2(32'h3bde2581),
	.w3(32'h3c3925ab),
	.w4(32'h3c32d29f),
	.w5(32'h3c09381e),
	.w6(32'hbad0fabe),
	.w7(32'hbbe8a440),
	.w8(32'h3bcf75a0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c250a),
	.w1(32'hba90fbe9),
	.w2(32'h3b1eac9e),
	.w3(32'h3b4f01a7),
	.w4(32'h3c2c96d4),
	.w5(32'h3c5fe9b5),
	.w6(32'h3b8f2d49),
	.w7(32'h3ba44cb2),
	.w8(32'hbae91305),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9330b1),
	.w1(32'h3b4f9b44),
	.w2(32'h3bad6764),
	.w3(32'h3c3377c1),
	.w4(32'h3bfc49cc),
	.w5(32'h3b4b3aa9),
	.w6(32'hba315c6c),
	.w7(32'hbb226833),
	.w8(32'h3b684f6e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cd276),
	.w1(32'h3b804295),
	.w2(32'h3be90219),
	.w3(32'h3b6885fe),
	.w4(32'h3b1fc61a),
	.w5(32'h3bf90f4f),
	.w6(32'h3b47f061),
	.w7(32'hb97cccf6),
	.w8(32'h3b10f8c5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c348037),
	.w1(32'h3b1397b3),
	.w2(32'h3c2ee4f0),
	.w3(32'h3ca5d6d7),
	.w4(32'hbaa6087c),
	.w5(32'h3c11bf9c),
	.w6(32'hbc228150),
	.w7(32'hbbcede9d),
	.w8(32'hbc14b02c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02cdfa),
	.w1(32'h3bb6f13d),
	.w2(32'h3bad2851),
	.w3(32'hba66477f),
	.w4(32'hba139ae9),
	.w5(32'hbaaf402c),
	.w6(32'hbc194f0c),
	.w7(32'hbaf4510f),
	.w8(32'hbbda0b0d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a412c4e),
	.w1(32'hbc78d6ed),
	.w2(32'hbcbf0b62),
	.w3(32'h3a7c60be),
	.w4(32'h3d5ba3ca),
	.w5(32'h3daa97ac),
	.w6(32'hbbb5bba0),
	.w7(32'hbc8371b5),
	.w8(32'h3d6ab725),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db668a9),
	.w1(32'h3bbbe212),
	.w2(32'h3b63523c),
	.w3(32'h3e49263a),
	.w4(32'hbb88c655),
	.w5(32'h3b11cd77),
	.w6(32'hbad4af95),
	.w7(32'h3b45e433),
	.w8(32'h3b68c336),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac86d42),
	.w1(32'h3a956258),
	.w2(32'h3b95a92e),
	.w3(32'h3bb1ed80),
	.w4(32'h3ab32aab),
	.w5(32'h3b805f63),
	.w6(32'hbbd718d7),
	.w7(32'hbb945f6c),
	.w8(32'hbbe76aff),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb17cdf),
	.w1(32'h3b9da7e6),
	.w2(32'h3b3e6a94),
	.w3(32'hba9ce0e0),
	.w4(32'h3b1b2b34),
	.w5(32'h3a2e4aef),
	.w6(32'hba45115a),
	.w7(32'h3b2aa871),
	.w8(32'hbbeb3a79),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad42a6d),
	.w1(32'h3b5ae015),
	.w2(32'h3ba34c0b),
	.w3(32'hb96d73b1),
	.w4(32'hba847380),
	.w5(32'h3a5b6e64),
	.w6(32'hbb7bff05),
	.w7(32'h3b509705),
	.w8(32'h3bb1fc90),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb210),
	.w1(32'hbba337f9),
	.w2(32'hbba590fe),
	.w3(32'h3bbc0763),
	.w4(32'hba932c9a),
	.w5(32'h3b078df6),
	.w6(32'h36eea1b8),
	.w7(32'h39c23404),
	.w8(32'hbb149ea9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a54f1),
	.w1(32'hbbd4ca70),
	.w2(32'hba45598b),
	.w3(32'hbba28193),
	.w4(32'hbb1086ca),
	.w5(32'hbb2c49e2),
	.w6(32'hbbb6ea8d),
	.w7(32'hbc1ec77b),
	.w8(32'hbb6b2ba6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc309e6),
	.w1(32'hbb9f877b),
	.w2(32'hbb14a966),
	.w3(32'hba921328),
	.w4(32'h3a98b88b),
	.w5(32'h3bc3f67d),
	.w6(32'hbb58d009),
	.w7(32'h3b2435d5),
	.w8(32'h3bbc5e72),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8103df),
	.w1(32'hbb4690cf),
	.w2(32'hbbfda792),
	.w3(32'h3a2e023f),
	.w4(32'hbbfe119f),
	.w5(32'hbc6b066c),
	.w6(32'hbb11e76a),
	.w7(32'hbc0121b6),
	.w8(32'hbbd9a068),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1b3f7),
	.w1(32'hbb502a3e),
	.w2(32'h3a1dbac2),
	.w3(32'hbc0df7da),
	.w4(32'h3b8be1c1),
	.w5(32'h3b03c27b),
	.w6(32'hbb325d1e),
	.w7(32'hbbfc8603),
	.w8(32'h3b6a4114),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a491076),
	.w1(32'hba30fc65),
	.w2(32'h3b63e8a6),
	.w3(32'h3be97d84),
	.w4(32'h3afcf08f),
	.w5(32'h3b397d7a),
	.w6(32'hbb19aa10),
	.w7(32'h3a0e35f6),
	.w8(32'h386291dd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caa719),
	.w1(32'hbb710e67),
	.w2(32'h3c06f971),
	.w3(32'h3b53739e),
	.w4(32'hbb8b8682),
	.w5(32'h3c6b4aec),
	.w6(32'h3b28f556),
	.w7(32'h3bd58069),
	.w8(32'hbb1a790e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963322a),
	.w1(32'h3c27986e),
	.w2(32'h3c889035),
	.w3(32'hbaecea3f),
	.w4(32'h3b8322a5),
	.w5(32'h3c7848f2),
	.w6(32'hba71547d),
	.w7(32'h3ab97103),
	.w8(32'hbc24fc0c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76ecb7),
	.w1(32'h3aa45879),
	.w2(32'h3abc0568),
	.w3(32'hbacc94e4),
	.w4(32'h3bb5eaad),
	.w5(32'h3b5dba22),
	.w6(32'hb854f58c),
	.w7(32'h3b9cc679),
	.w8(32'hbb39efd5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda4982),
	.w1(32'hbabb3300),
	.w2(32'h39a553e3),
	.w3(32'h3c08bbc7),
	.w4(32'h3a62d0da),
	.w5(32'hbb1ca5dc),
	.w6(32'hbc208351),
	.w7(32'hbc2fb09e),
	.w8(32'hbc0be058),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc66613),
	.w1(32'h3be4f3f6),
	.w2(32'h3c06d0d0),
	.w3(32'h3bf288f7),
	.w4(32'h3c06bb0a),
	.w5(32'h3c4121d5),
	.w6(32'hbb9e9d0e),
	.w7(32'hbb2bd4d5),
	.w8(32'h3bff25a9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb2c91),
	.w1(32'h3b2957a2),
	.w2(32'h3c828797),
	.w3(32'h3c15d688),
	.w4(32'h3bead80f),
	.w5(32'h3ca93c04),
	.w6(32'hbb35bc6e),
	.w7(32'h3baa30f5),
	.w8(32'h3bb9e057),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c862e6d),
	.w1(32'hbb630daa),
	.w2(32'h3ac3bdb8),
	.w3(32'h3ca1714c),
	.w4(32'hbba559ce),
	.w5(32'hb9ce2218),
	.w6(32'hbc028e64),
	.w7(32'hbba1e2e8),
	.w8(32'hbbd9c706),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb905c96),
	.w1(32'hbbc779af),
	.w2(32'hbb9a837c),
	.w3(32'hbc50b626),
	.w4(32'h3bd00a8a),
	.w5(32'h3be3dc28),
	.w6(32'hba96b583),
	.w7(32'h3b26dc99),
	.w8(32'h3a8f8e17),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12fdc4),
	.w1(32'hbbb841df),
	.w2(32'hbb123ffc),
	.w3(32'h3be37f53),
	.w4(32'h3b85ba14),
	.w5(32'hbadb87c0),
	.w6(32'hbc179684),
	.w7(32'hbbbee7c6),
	.w8(32'h3bad48ea),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd99e2b),
	.w1(32'hbad89fd4),
	.w2(32'h3b993ee0),
	.w3(32'h3bd8bb59),
	.w4(32'h3b18f589),
	.w5(32'h3a46e857),
	.w6(32'hbb107b9d),
	.w7(32'hbb8635a9),
	.w8(32'hbb6351b0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaad99),
	.w1(32'hbbca792f),
	.w2(32'h3c3d797b),
	.w3(32'h3c2b1e83),
	.w4(32'h3a43dac7),
	.w5(32'h3c5be110),
	.w6(32'h3bcd96a8),
	.w7(32'h3c2cefbb),
	.w8(32'h3b569660),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45ae31),
	.w1(32'h3a4d46d9),
	.w2(32'h3b08838f),
	.w3(32'h3b305ca3),
	.w4(32'h3c476c16),
	.w5(32'h3c27cfa4),
	.w6(32'h3b8a95ba),
	.w7(32'h3bba5401),
	.w8(32'h3bc8b51e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7762c2),
	.w1(32'h3b9d166b),
	.w2(32'h3c369799),
	.w3(32'h3ca5e146),
	.w4(32'hbbcaaa30),
	.w5(32'hbaaad7ca),
	.w6(32'hba7f890a),
	.w7(32'h3b0bade9),
	.w8(32'hbbdf6708),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51c6a4),
	.w1(32'h3b1cacb2),
	.w2(32'h3b24d57f),
	.w3(32'hbc281bfc),
	.w4(32'h3abf3801),
	.w5(32'h3c06e522),
	.w6(32'h3c116d29),
	.w7(32'h3b61b8bb),
	.w8(32'h3c11f11c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3946a9),
	.w1(32'h39b638f3),
	.w2(32'h3be8b5be),
	.w3(32'h3c9a63b6),
	.w4(32'h3b762713),
	.w5(32'h3b7f0f72),
	.w6(32'hbadda928),
	.w7(32'h3ac0ba21),
	.w8(32'hbb09579a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94a0f7),
	.w1(32'h3b5f87c2),
	.w2(32'h3c39873a),
	.w3(32'hb9f94ce1),
	.w4(32'h39ae491a),
	.w5(32'h3bf0a341),
	.w6(32'hbc2da749),
	.w7(32'hbba867ed),
	.w8(32'hbbc673aa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab738f7),
	.w1(32'h3c107bf9),
	.w2(32'h3c1a5ad8),
	.w3(32'h3a6d3b6e),
	.w4(32'h3c1f9e62),
	.w5(32'h3b2cfba6),
	.w6(32'hbbc0fc04),
	.w7(32'hba1d1076),
	.w8(32'h39c48530),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09edf8),
	.w1(32'hb9aae51f),
	.w2(32'hbb78e6ad),
	.w3(32'h3a1ac019),
	.w4(32'h3bae70dd),
	.w5(32'hba62af38),
	.w6(32'hbbd9e226),
	.w7(32'hbc2a19cc),
	.w8(32'hbaef5862),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36eb20),
	.w1(32'hba23e2f7),
	.w2(32'hbb03e5c2),
	.w3(32'h3c215429),
	.w4(32'h38d08b68),
	.w5(32'hbb40a001),
	.w6(32'h3a9ff88a),
	.w7(32'hbabd0a19),
	.w8(32'hbbb5702b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cff86),
	.w1(32'hba95bf7e),
	.w2(32'hbaab9fec),
	.w3(32'hbb863af0),
	.w4(32'h3a9d8a7e),
	.w5(32'h3bb5cd73),
	.w6(32'hbac0dfbf),
	.w7(32'hbb87924d),
	.w8(32'h380a8b05),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9d49c),
	.w1(32'hbbc2dc64),
	.w2(32'hbbfe6ba3),
	.w3(32'h3bd1b112),
	.w4(32'hbc1fe8ca),
	.w5(32'hbbe46b61),
	.w6(32'hbb777ffe),
	.w7(32'hbc048230),
	.w8(32'hbbdd35dc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24cf00),
	.w1(32'hbb9a67ba),
	.w2(32'hbbae5ac7),
	.w3(32'hbc07ae61),
	.w4(32'hbc232a44),
	.w5(32'h3a7db7f7),
	.w6(32'hbc15561b),
	.w7(32'hbafebcae),
	.w8(32'hba4ee6ae),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a29b),
	.w1(32'h3a7053c8),
	.w2(32'h3b818cf5),
	.w3(32'h3b35c865),
	.w4(32'h3b823786),
	.w5(32'h3c85ce66),
	.w6(32'hbc1216ad),
	.w7(32'hbbf6dd40),
	.w8(32'h3b104242),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6edfa),
	.w1(32'hbbb8bbb2),
	.w2(32'hbbb8621a),
	.w3(32'h3d048e4d),
	.w4(32'hbbacc310),
	.w5(32'hbbd22ab7),
	.w6(32'h3aa6e529),
	.w7(32'hba3c3827),
	.w8(32'hbc830675),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e77a6),
	.w1(32'h3b00e931),
	.w2(32'h3aec649f),
	.w3(32'hbc720237),
	.w4(32'hba81488d),
	.w5(32'hba88e1a1),
	.w6(32'h3b074fc7),
	.w7(32'h3abbdaf6),
	.w8(32'hbac4f3ee),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b151412),
	.w1(32'hb9a3e56e),
	.w2(32'h3a356cb6),
	.w3(32'hba4b7285),
	.w4(32'h3af00b6a),
	.w5(32'h3b8d7886),
	.w6(32'hbaa52ca9),
	.w7(32'hbb841c4b),
	.w8(32'h3a28f4f0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86f28),
	.w1(32'h3ba4e916),
	.w2(32'h3ac577cd),
	.w3(32'h3bd043af),
	.w4(32'h3b3e11b0),
	.w5(32'h3b9573a4),
	.w6(32'h3b164f3b),
	.w7(32'h3b721402),
	.w8(32'hb7a1976b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39dc77),
	.w1(32'hbc32dacd),
	.w2(32'hbc516006),
	.w3(32'hbbf45ba5),
	.w4(32'h3ac9d6d3),
	.w5(32'h3a63583b),
	.w6(32'hbc31f400),
	.w7(32'hbc51bd8d),
	.w8(32'h39a734cd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcdc2d),
	.w1(32'h3b77de7f),
	.w2(32'h3add8fb3),
	.w3(32'h3bb19ec6),
	.w4(32'hbbcfa41b),
	.w5(32'h3bccdd70),
	.w6(32'hbbd9059f),
	.w7(32'hba92ee9a),
	.w8(32'hb9cf515f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdada66),
	.w1(32'hbb8e2578),
	.w2(32'hbb152943),
	.w3(32'h3bbbd92f),
	.w4(32'h3b408f1b),
	.w5(32'hbb1c8835),
	.w6(32'h3af9da3f),
	.w7(32'hbb94c8bd),
	.w8(32'hbb987270),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ac751),
	.w1(32'hbb3f546b),
	.w2(32'hbb9953f7),
	.w3(32'hba80474b),
	.w4(32'h3b8fccaf),
	.w5(32'hbb3c543f),
	.w6(32'hbbd7397b),
	.w7(32'hbc048781),
	.w8(32'hbc14e556),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6286a),
	.w1(32'hbb926632),
	.w2(32'hbbaa1180),
	.w3(32'h3afba919),
	.w4(32'hbade6582),
	.w5(32'hbaad9e3f),
	.w6(32'hbc074317),
	.w7(32'h392e84f1),
	.w8(32'hbbe42666),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3dbaa),
	.w1(32'hbc2b6dec),
	.w2(32'h3b45c385),
	.w3(32'h3b0040f9),
	.w4(32'hbbda48fb),
	.w5(32'h3b343ded),
	.w6(32'hbc082e73),
	.w7(32'hba8c401d),
	.w8(32'hbb792cf3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b072496),
	.w1(32'h3b0af163),
	.w2(32'h3ae9012f),
	.w3(32'h391f2954),
	.w4(32'hbb19a89c),
	.w5(32'hbba395e8),
	.w6(32'hbb5eb145),
	.w7(32'hbb096c9a),
	.w8(32'h3b144c47),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bd37b),
	.w1(32'h3971ca2c),
	.w2(32'hb9e4f355),
	.w3(32'h3b5dac23),
	.w4(32'hbb864946),
	.w5(32'hbbb996b8),
	.w6(32'h3afd3349),
	.w7(32'hbb31d544),
	.w8(32'hbbd67ef5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc5be1),
	.w1(32'h3b10fd26),
	.w2(32'h3b8a87f7),
	.w3(32'h3bc4338c),
	.w4(32'h3b8999a2),
	.w5(32'h3ad9f112),
	.w6(32'hb9f817a8),
	.w7(32'hbba906b0),
	.w8(32'hbc1df3b9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd269e),
	.w1(32'h3bacc887),
	.w2(32'h3b8b0d86),
	.w3(32'h3a84cbf8),
	.w4(32'h3c0637e7),
	.w5(32'h3b7b4e7c),
	.w6(32'h3a9d76dc),
	.w7(32'h3adc484f),
	.w8(32'h3b24dd83),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2229c),
	.w1(32'h3badb6d5),
	.w2(32'hb9481663),
	.w3(32'h3c152c12),
	.w4(32'h3b8b188e),
	.w5(32'hb9f76e93),
	.w6(32'hba8edcc7),
	.w7(32'hbb56b82e),
	.w8(32'h3c376664),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78977a),
	.w1(32'hbab920e0),
	.w2(32'hbbbc4a7b),
	.w3(32'h3c5c8565),
	.w4(32'h3b97baeb),
	.w5(32'hbae83a5c),
	.w6(32'hbb19ba0c),
	.w7(32'hbb1e51c9),
	.w8(32'hbc0b8ab0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd424e),
	.w1(32'h3b900edc),
	.w2(32'h3c01fea3),
	.w3(32'h3a819ff9),
	.w4(32'h3c11d463),
	.w5(32'h3c386b5b),
	.w6(32'hbc09102f),
	.w7(32'h3b818175),
	.w8(32'hbacfc8e9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42c398),
	.w1(32'hba8719fc),
	.w2(32'hbac2b0d4),
	.w3(32'h3c0c4833),
	.w4(32'hb95dc3cb),
	.w5(32'hbb730302),
	.w6(32'hba9250c7),
	.w7(32'hbb59ed8d),
	.w8(32'hbb8e3889),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9ad8d),
	.w1(32'hba37acf1),
	.w2(32'hba8b2f9b),
	.w3(32'h3a862d93),
	.w4(32'h3a41c955),
	.w5(32'hba23dc2f),
	.w6(32'hbac61984),
	.w7(32'hb9f8d37b),
	.w8(32'hbb37877c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f0634),
	.w1(32'hbbccb5b8),
	.w2(32'hbb6eaa69),
	.w3(32'h3bb1b82b),
	.w4(32'hbb98ba42),
	.w5(32'hbbb195bc),
	.w6(32'hbbce74fe),
	.w7(32'hbc2936a4),
	.w8(32'h3b04759a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed1d29),
	.w1(32'hbc0dc421),
	.w2(32'hbaa74b45),
	.w3(32'h3a918d87),
	.w4(32'hbbadc261),
	.w5(32'hbaaed4b5),
	.w6(32'h3b52abe3),
	.w7(32'hbaa2e111),
	.w8(32'hbb4a0303),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc78ff),
	.w1(32'h3b898a12),
	.w2(32'h3a5e937f),
	.w3(32'h3c0db9f9),
	.w4(32'hbc183690),
	.w5(32'hbb99610d),
	.w6(32'hbbc8bf8c),
	.w7(32'hbbd2786f),
	.w8(32'hbb767075),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9d10c),
	.w1(32'hbb9331a4),
	.w2(32'hbc6e9b8f),
	.w3(32'h3b7c1c36),
	.w4(32'h3b8b1bed),
	.w5(32'h3c132d89),
	.w6(32'hbb11822c),
	.w7(32'hbb518e9a),
	.w8(32'hbc0643be),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0e45e),
	.w1(32'h3b6dd766),
	.w2(32'h3b8a6dad),
	.w3(32'h3c6d512d),
	.w4(32'h3c2736a2),
	.w5(32'h3bc2b22b),
	.w6(32'h3acd41ae),
	.w7(32'h3a023d41),
	.w8(32'h3bb792e8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c610cf3),
	.w1(32'hbb42caaf),
	.w2(32'h3c0b8b49),
	.w3(32'h3bca6598),
	.w4(32'hbbdb8b22),
	.w5(32'hbb0019e6),
	.w6(32'hbbd449a9),
	.w7(32'h3a85cb18),
	.w8(32'hbb19e231),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30720b),
	.w1(32'hbc0d1a59),
	.w2(32'hba835e97),
	.w3(32'h3a840181),
	.w4(32'h3b4edea5),
	.w5(32'h3c9f9559),
	.w6(32'hbbafb188),
	.w7(32'hbb994d71),
	.w8(32'hbb7bcb3b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163d85),
	.w1(32'h3abeade9),
	.w2(32'hb8b13102),
	.w3(32'h3c7140ab),
	.w4(32'hbba7be82),
	.w5(32'h3b264930),
	.w6(32'hbbd1b221),
	.w7(32'hbb40bde3),
	.w8(32'h3afe8afa),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed637),
	.w1(32'hbc37a8f0),
	.w2(32'hbc077804),
	.w3(32'h3b095b86),
	.w4(32'h3ab3bdd2),
	.w5(32'h3c08c94d),
	.w6(32'hbb0120bd),
	.w7(32'hba25b7ff),
	.w8(32'hb9c41420),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42da1f),
	.w1(32'h3abeb6d0),
	.w2(32'h3adee33e),
	.w3(32'h3b3101aa),
	.w4(32'h3b1a7200),
	.w5(32'h3c142a58),
	.w6(32'hbbc6e88d),
	.w7(32'hbb1d10a9),
	.w8(32'h3a3ea6e0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d8964),
	.w1(32'h39f41c49),
	.w2(32'hbaf52891),
	.w3(32'hbad625e5),
	.w4(32'h3b5146a4),
	.w5(32'h3a6879d2),
	.w6(32'h3b2038a1),
	.w7(32'h3a1dd337),
	.w8(32'h3b78c9e2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fd4c0),
	.w1(32'h3b222b6c),
	.w2(32'h3b48d765),
	.w3(32'h3c3230be),
	.w4(32'h3b02ed27),
	.w5(32'h3a0b3050),
	.w6(32'hba1ac658),
	.w7(32'h3a22fb4a),
	.w8(32'hb9224ea2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab81714),
	.w1(32'hbb804729),
	.w2(32'h3a214271),
	.w3(32'hbad089f6),
	.w4(32'hbb03b72a),
	.w5(32'hbb1828a4),
	.w6(32'hbacb08a6),
	.w7(32'hbb185bfc),
	.w8(32'hbc04cc23),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b628617),
	.w1(32'h3a38479d),
	.w2(32'h3c08f795),
	.w3(32'h3bb3d715),
	.w4(32'hba7e0ca4),
	.w5(32'h3b340990),
	.w6(32'hbb7291ca),
	.w7(32'hbab11f37),
	.w8(32'hbb323ff6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e924c),
	.w1(32'h3aab3298),
	.w2(32'hbc092f66),
	.w3(32'hb9882601),
	.w4(32'hbac68b87),
	.w5(32'hbb1e2ede),
	.w6(32'hbba18546),
	.w7(32'hbbf2978c),
	.w8(32'hbb497382),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf4bce),
	.w1(32'hbbe46ee9),
	.w2(32'hbbc3ce1e),
	.w3(32'h39d8f269),
	.w4(32'hbb9e5f41),
	.w5(32'hbb0b9cf5),
	.w6(32'hbb73897b),
	.w7(32'hbb718cfb),
	.w8(32'hbbb0f187),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f6f90),
	.w1(32'hbadd1b09),
	.w2(32'h3c186e75),
	.w3(32'h3b7808f3),
	.w4(32'hbb0d229f),
	.w5(32'h3bbc9a54),
	.w6(32'hbc16e5da),
	.w7(32'hbc21af49),
	.w8(32'h3aecf46b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f22f),
	.w1(32'hbba15048),
	.w2(32'hbb079db9),
	.w3(32'h3c2a5017),
	.w4(32'hbba35500),
	.w5(32'h3aaaa3be),
	.w6(32'hbbc948ef),
	.w7(32'hbb8a6aee),
	.w8(32'hba337ac1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59779b),
	.w1(32'hbba83b91),
	.w2(32'hbba86ca7),
	.w3(32'hbb91a5b4),
	.w4(32'h3b42507a),
	.w5(32'h3696ec36),
	.w6(32'hbc20aba4),
	.w7(32'hbbd0bd91),
	.w8(32'hbbd889aa),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a705eeb),
	.w1(32'hbb789197),
	.w2(32'hbc12a40d),
	.w3(32'h3b075e95),
	.w4(32'hba3d3610),
	.w5(32'hbc79330d),
	.w6(32'h3b5d4445),
	.w7(32'hbb377639),
	.w8(32'hb9ee985f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba84bc5),
	.w1(32'h3ba40c6b),
	.w2(32'h3c29b064),
	.w3(32'h3bfddc67),
	.w4(32'hb98bff4c),
	.w5(32'h3b8bd9cb),
	.w6(32'hbb840b04),
	.w7(32'h3a675343),
	.w8(32'hbb2009ff),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ce550),
	.w1(32'hbc2bc4b7),
	.w2(32'h3a6e0c38),
	.w3(32'h3ae963ea),
	.w4(32'h3b27a430),
	.w5(32'hb70d68cb),
	.w6(32'hbc42aca7),
	.w7(32'hbb1aa4de),
	.w8(32'hb98b2dac),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395bcd87),
	.w1(32'hbbf586ff),
	.w2(32'h3c06f064),
	.w3(32'hbb8c3807),
	.w4(32'hba53debb),
	.w5(32'h3c4afe47),
	.w6(32'hbc0640ae),
	.w7(32'hbb77c6a6),
	.w8(32'hbb45ef72),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46c0c0),
	.w1(32'hb9f0e0ca),
	.w2(32'h3bf6e312),
	.w3(32'h3bfa0f90),
	.w4(32'hbaec0fcd),
	.w5(32'h3bdadf7a),
	.w6(32'hbb795232),
	.w7(32'h3a4290fb),
	.w8(32'h3a13737c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873b4e),
	.w1(32'hbbbd8791),
	.w2(32'h3b50dbed),
	.w3(32'h3b6b09d2),
	.w4(32'hbb90aded),
	.w5(32'hba2e99e3),
	.w6(32'hbbfcf388),
	.w7(32'hb9bfcc31),
	.w8(32'hbb907ced),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6636b5),
	.w1(32'hbb94e41b),
	.w2(32'hbbdbc4a2),
	.w3(32'h3b443347),
	.w4(32'h384862fe),
	.w5(32'h3c52ac4a),
	.w6(32'hbb1195ba),
	.w7(32'hbb1a88f3),
	.w8(32'hbb6584eb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ccb0b),
	.w1(32'hbc9b630f),
	.w2(32'hbca37774),
	.w3(32'hbb8a6a1a),
	.w4(32'hbca45698),
	.w5(32'hbc832b2e),
	.w6(32'hbc933991),
	.w7(32'hbc97dab4),
	.w8(32'hbc98201b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99de6e),
	.w1(32'h3b2d2f95),
	.w2(32'h390dbc58),
	.w3(32'hbc5236d6),
	.w4(32'h3a0d116f),
	.w5(32'hba7a84f0),
	.w6(32'hb93a4830),
	.w7(32'hba318285),
	.w8(32'hbb0aff7d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec373c),
	.w1(32'hbb13386a),
	.w2(32'h3b834c8b),
	.w3(32'hba882d15),
	.w4(32'hb9b284da),
	.w5(32'h3be7cb83),
	.w6(32'hba8a9626),
	.w7(32'h3a399814),
	.w8(32'hbbbef363),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76ecaa),
	.w1(32'hbaddeb06),
	.w2(32'h3babdba9),
	.w3(32'h3c129e64),
	.w4(32'h3b08b8b8),
	.w5(32'h3c1d21c8),
	.w6(32'hbbb2f47f),
	.w7(32'hba2a01cc),
	.w8(32'hbb05c2c3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb09dad),
	.w1(32'hbc5ffbad),
	.w2(32'hbb7bec5b),
	.w3(32'h3c2729f7),
	.w4(32'hbc85a131),
	.w5(32'hbbd81c04),
	.w6(32'hbbf40622),
	.w7(32'hbc233a06),
	.w8(32'hbbe94d41),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c8ff8),
	.w1(32'hbc337558),
	.w2(32'hba61e46f),
	.w3(32'hbbcf5ee7),
	.w4(32'hbb61ebf2),
	.w5(32'hb9dde06a),
	.w6(32'hbc159156),
	.w7(32'hbb085e41),
	.w8(32'hbaf48f96),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39254288),
	.w1(32'h3a8b0db6),
	.w2(32'hb9b94a1f),
	.w3(32'hbb7c509b),
	.w4(32'hbb47de84),
	.w5(32'h3c438fec),
	.w6(32'h3b40c840),
	.w7(32'h3b43c66e),
	.w8(32'h3ba94bb2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcf061),
	.w1(32'h3ba39efc),
	.w2(32'h3b878ee1),
	.w3(32'h3c83f876),
	.w4(32'h3b20a171),
	.w5(32'h3ab4596b),
	.w6(32'h3b8136a2),
	.w7(32'h3b86340f),
	.w8(32'h3a9a6ad2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b84e7),
	.w1(32'hba354a2d),
	.w2(32'h3a8ad6ec),
	.w3(32'h3a864459),
	.w4(32'h3b75e6ff),
	.w5(32'h3c9b6ee6),
	.w6(32'h3b27d8b6),
	.w7(32'hbaa18e13),
	.w8(32'h399ced2a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ee1ad),
	.w1(32'hbb21100a),
	.w2(32'hbbac3499),
	.w3(32'h3d01a349),
	.w4(32'hbc05647d),
	.w5(32'hbae9901f),
	.w6(32'hbb9e3333),
	.w7(32'hbbf951ca),
	.w8(32'hbc0df245),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5410f),
	.w1(32'h3b6b6f32),
	.w2(32'h3bf74b32),
	.w3(32'hbb87134c),
	.w4(32'hbb06dbb0),
	.w5(32'h3ab18aee),
	.w6(32'hbbe58d1f),
	.w7(32'h3a35dcc2),
	.w8(32'h3b8d7be1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13b05d),
	.w1(32'h3a5f6724),
	.w2(32'h3b0e14d9),
	.w3(32'h3ba340e2),
	.w4(32'h3bf5d49d),
	.w5(32'h3be7d8cd),
	.w6(32'h3a4ec3a4),
	.w7(32'h3a7a66aa),
	.w8(32'h3bb2f6d7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1eb6d5),
	.w1(32'h3b8e0b98),
	.w2(32'h3baebdd0),
	.w3(32'h3c961467),
	.w4(32'h3b65a710),
	.w5(32'h3c01e31e),
	.w6(32'hbc03729b),
	.w7(32'hbb2beb62),
	.w8(32'hbba055b6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad222b7),
	.w1(32'h3b8874a9),
	.w2(32'h3bbd7a2c),
	.w3(32'h3b2d2b09),
	.w4(32'hbb0175c5),
	.w5(32'hbadf1c6e),
	.w6(32'hb9b27966),
	.w7(32'h3c06b5a7),
	.w8(32'hb9bbb044),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5b32),
	.w1(32'h38f295bc),
	.w2(32'h3b9cdbe9),
	.w3(32'hbc3b30bc),
	.w4(32'hb9ab9edf),
	.w5(32'h3ba1fc46),
	.w6(32'hbacb2b8b),
	.w7(32'h3b629b2c),
	.w8(32'hb9b4a253),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5453e),
	.w1(32'hbb41f2da),
	.w2(32'hbb901b19),
	.w3(32'h3b008ecc),
	.w4(32'hbbe314e0),
	.w5(32'hbbce94d8),
	.w6(32'hbc00aebf),
	.w7(32'hbbe8223e),
	.w8(32'hbc4c9dcd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1cf11),
	.w1(32'hbaaa919c),
	.w2(32'h3b85e832),
	.w3(32'hbbc55be6),
	.w4(32'hba83b772),
	.w5(32'h3ba4806f),
	.w6(32'hba71c673),
	.w7(32'hbb455480),
	.w8(32'h3bd917d4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05355e),
	.w1(32'h3a719f5a),
	.w2(32'h3bb8c135),
	.w3(32'h3c763553),
	.w4(32'h3b925b59),
	.w5(32'h3b1b03c8),
	.w6(32'hbb9dcdc8),
	.w7(32'hbb0e27d8),
	.w8(32'h39494a0d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c429),
	.w1(32'hba167b34),
	.w2(32'hbaa8714a),
	.w3(32'h3a6ebd6a),
	.w4(32'hba2c44b9),
	.w5(32'hba926d0a),
	.w6(32'hb927db14),
	.w7(32'hb986a6e0),
	.w8(32'h39d59229),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399979b1),
	.w1(32'h3b4df115),
	.w2(32'h3c6e2b81),
	.w3(32'hb95013bf),
	.w4(32'hbb95d501),
	.w5(32'h3a86249c),
	.w6(32'h3ac86ff9),
	.w7(32'hbaefeaf8),
	.w8(32'h3bbeb523),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule