module layer_8_featuremap_140(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01e430),
	.w1(32'hb9f3abfe),
	.w2(32'h3aa057bd),
	.w3(32'hba9a035a),
	.w4(32'hb8ed6d94),
	.w5(32'hb9170550),
	.w6(32'hbadf1e8b),
	.w7(32'hb9995225),
	.w8(32'hba659f36),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88b0ea),
	.w1(32'hb9c0064a),
	.w2(32'hb9c9dab8),
	.w3(32'hba394098),
	.w4(32'hb91136cc),
	.w5(32'hba5e5e09),
	.w6(32'hbab31899),
	.w7(32'hbaa6662b),
	.w8(32'hbb316d7e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac08c21),
	.w1(32'hb9dd1f04),
	.w2(32'hb9a38202),
	.w3(32'hba8f6547),
	.w4(32'hba81553e),
	.w5(32'h3a65953a),
	.w6(32'hbb2eb0f7),
	.w7(32'hbb29b2e2),
	.w8(32'h3a735c93),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce9542),
	.w1(32'h3a9d8b55),
	.w2(32'hbabd2402),
	.w3(32'h3b011ab7),
	.w4(32'h392e8a42),
	.w5(32'hba1d3401),
	.w6(32'h3b061fcf),
	.w7(32'hbad5534a),
	.w8(32'hbb1cdddd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dfaec),
	.w1(32'hbb1cd41a),
	.w2(32'h39242329),
	.w3(32'hbb0f7626),
	.w4(32'hb9931284),
	.w5(32'hba44aeac),
	.w6(32'hbb2fe92b),
	.w7(32'h38e6bf81),
	.w8(32'hba954ecc),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5f9e0),
	.w1(32'h39f8b76c),
	.w2(32'hb8566b7a),
	.w3(32'hba89aa39),
	.w4(32'h3a313a90),
	.w5(32'h39f6ce14),
	.w6(32'hba34804e),
	.w7(32'h37bcdeda),
	.w8(32'hb9d0ccc0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9905896),
	.w1(32'hb8455eb2),
	.w2(32'h39007aac),
	.w3(32'h38148fd1),
	.w4(32'h3ab6034b),
	.w5(32'hba4edc0d),
	.w6(32'hb9f91532),
	.w7(32'hb84b2e90),
	.w8(32'hbb222d73),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcfecd),
	.w1(32'hb923ab08),
	.w2(32'h3a540790),
	.w3(32'hba96e097),
	.w4(32'hb9ab998d),
	.w5(32'h39b2cf0f),
	.w6(32'hbb0c0d21),
	.w7(32'hb990cabd),
	.w8(32'hb9e2188e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac13100),
	.w1(32'hbb1fcfa9),
	.w2(32'hba79db88),
	.w3(32'hbb6c36e4),
	.w4(32'hbb7f3989),
	.w5(32'hbb11d1e8),
	.w6(32'hbb6716ba),
	.w7(32'hbb80bd9e),
	.w8(32'hbb309a0e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb868abe9),
	.w1(32'hb98c0a63),
	.w2(32'hbaaf8499),
	.w3(32'hbaa15486),
	.w4(32'h3a905738),
	.w5(32'h39de2128),
	.w6(32'hba9005b2),
	.w7(32'h396c9d4c),
	.w8(32'hbafab51a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae751c1),
	.w1(32'hba537a3c),
	.w2(32'hbb3d7e1f),
	.w3(32'hb9b96ec8),
	.w4(32'hbb8953b5),
	.w5(32'hbb43015a),
	.w6(32'hba445235),
	.w7(32'hbb773c86),
	.w8(32'hba5b2af2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b3ca9),
	.w1(32'hbaca5a9b),
	.w2(32'h38acb13c),
	.w3(32'hbaac624a),
	.w4(32'hb6d61f1a),
	.w5(32'h39470754),
	.w6(32'hbaa32cc4),
	.w7(32'hb9aac3f5),
	.w8(32'hba14db96),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a803378),
	.w1(32'h3a28df0f),
	.w2(32'h3a3e3400),
	.w3(32'hb82c793e),
	.w4(32'hba79408c),
	.w5(32'hb946141e),
	.w6(32'h388dc2a5),
	.w7(32'hb9afad62),
	.w8(32'hb94291a6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880f7fd),
	.w1(32'h39588e08),
	.w2(32'h39c7856f),
	.w3(32'hb8635ee3),
	.w4(32'h39b784ed),
	.w5(32'h39f6f91f),
	.w6(32'h3971b945),
	.w7(32'h39e597a7),
	.w8(32'h3a06af5a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944167a),
	.w1(32'h379c2f6c),
	.w2(32'h390fc0e2),
	.w3(32'hb82a287b),
	.w4(32'h3964c0fe),
	.w5(32'h39a941a5),
	.w6(32'h3944538f),
	.w7(32'h392e4ba0),
	.w8(32'h39c30c6d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952d765),
	.w1(32'hb96f5790),
	.w2(32'hbac40584),
	.w3(32'hb9aeedc1),
	.w4(32'hbadead0d),
	.w5(32'hbac34de9),
	.w6(32'hb95e455e),
	.w7(32'hbacdcff6),
	.w8(32'hbaa1e530),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66428d),
	.w1(32'hba39b725),
	.w2(32'hb9abc3bc),
	.w3(32'hbadfd9b7),
	.w4(32'hb9e4c396),
	.w5(32'hba977c32),
	.w6(32'hbaa5e0f4),
	.w7(32'hba1b3991),
	.w8(32'hbab31f08),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f568cc),
	.w1(32'h39ef790e),
	.w2(32'h3a6c8911),
	.w3(32'hbaaaa11f),
	.w4(32'hbaa3224c),
	.w5(32'hba490567),
	.w6(32'hba8aca2a),
	.w7(32'hba8d5a20),
	.w8(32'hb98afcdf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50e9b0),
	.w1(32'hbb3f3075),
	.w2(32'hbb3fa1d0),
	.w3(32'hbb2f15f3),
	.w4(32'hbb225840),
	.w5(32'hbb32991d),
	.w6(32'hbb20873b),
	.w7(32'hbb28ed33),
	.w8(32'hbb1e2d13),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e29e3c),
	.w1(32'hb8caa6dc),
	.w2(32'hbab7d3c0),
	.w3(32'hbae7670b),
	.w4(32'hba9781d1),
	.w5(32'hbb7a6f85),
	.w6(32'hba11cddc),
	.w7(32'hba2fda03),
	.w8(32'hbae2bafa),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908b51f),
	.w1(32'hba678db7),
	.w2(32'hbb0102ea),
	.w3(32'hbadeaf01),
	.w4(32'hbab60482),
	.w5(32'hba315184),
	.w6(32'hb8d8a998),
	.w7(32'hba8cf362),
	.w8(32'hb9b9b08c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8b65f),
	.w1(32'h3b4aaba3),
	.w2(32'h3a13aed3),
	.w3(32'h3aabf037),
	.w4(32'h3b0cc2c1),
	.w5(32'h3b0e373f),
	.w6(32'h3ad7e423),
	.w7(32'h3a1690cb),
	.w8(32'h3a094d5a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba946ec7),
	.w1(32'hbb35839c),
	.w2(32'hbb5a3782),
	.w3(32'hbab89dd8),
	.w4(32'hbb8b5632),
	.w5(32'hbb51db2f),
	.w6(32'hba256783),
	.w7(32'hbb88143b),
	.w8(32'hbb2454d6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b069de3),
	.w1(32'h3ad2d745),
	.w2(32'hba5d191a),
	.w3(32'h39d9805b),
	.w4(32'hbad249ca),
	.w5(32'hba8cbad0),
	.w6(32'h3a29c7d4),
	.w7(32'hbb102119),
	.w8(32'hbac82ddc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06c5cd),
	.w1(32'hbaea2c63),
	.w2(32'hbab64d8a),
	.w3(32'hbaff5c66),
	.w4(32'hbaadffa8),
	.w5(32'hbb09949b),
	.w6(32'hbb0f7052),
	.w7(32'hbaf5cfb4),
	.w8(32'hbb094363),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f100ca),
	.w1(32'hb90dae3b),
	.w2(32'h3acbd7a4),
	.w3(32'hb9f10159),
	.w4(32'h3a1de21a),
	.w5(32'hba7b82f4),
	.w6(32'hba1ffdb3),
	.w7(32'hba84b814),
	.w8(32'hbb21e1e3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80b147),
	.w1(32'hba984406),
	.w2(32'hba10f0db),
	.w3(32'hb8c96893),
	.w4(32'h39e38571),
	.w5(32'h397b1a53),
	.w6(32'hba122933),
	.w7(32'hb932364c),
	.w8(32'hb9651743),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fd0dd),
	.w1(32'hbc1ce854),
	.w2(32'hbc66bd22),
	.w3(32'hbc40090d),
	.w4(32'hbbe7c622),
	.w5(32'hbc412a8b),
	.w6(32'hbbc55286),
	.w7(32'hbbc5f415),
	.w8(32'hbbf2b92d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf14b9),
	.w1(32'hbaf7d35d),
	.w2(32'hbabbce52),
	.w3(32'hba105093),
	.w4(32'hba839543),
	.w5(32'hba3589f4),
	.w6(32'hba9cc607),
	.w7(32'hba8290fe),
	.w8(32'hbaa4f3eb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819048),
	.w1(32'hb97616bc),
	.w2(32'h3aa85eb2),
	.w3(32'h37d9d9fa),
	.w4(32'h395e171f),
	.w5(32'h39cec1e7),
	.w6(32'hba04147f),
	.w7(32'h3a7fe307),
	.w8(32'h39ec5827),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a4ec7),
	.w1(32'h3b334d1b),
	.w2(32'h3ac2d33d),
	.w3(32'h3b74bda5),
	.w4(32'h3af221c5),
	.w5(32'h3ae047ff),
	.w6(32'h3b6208e9),
	.w7(32'h3b27db44),
	.w8(32'h3b042289),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee8e4d),
	.w1(32'h392da642),
	.w2(32'hbabe278a),
	.w3(32'h3964b218),
	.w4(32'hbab00f87),
	.w5(32'hbaa9db21),
	.w6(32'h3a3b27d9),
	.w7(32'hba3a288a),
	.w8(32'hb9e06aa6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac64107),
	.w1(32'hbaa4eff6),
	.w2(32'h3aa674c4),
	.w3(32'hbaada294),
	.w4(32'hb95f8a1e),
	.w5(32'hb8e0ab1d),
	.w6(32'hba634161),
	.w7(32'h39ebe480),
	.w8(32'h3a97d4e0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eaeef),
	.w1(32'h3b1d17fa),
	.w2(32'h39bfea1b),
	.w3(32'hb8234a44),
	.w4(32'h395d7d5c),
	.w5(32'hb9f227e2),
	.w6(32'h3aba40b5),
	.w7(32'h398b8db1),
	.w8(32'hb9f29a3c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831df9b),
	.w1(32'h3a7a4e25),
	.w2(32'hb7c55c90),
	.w3(32'h3ab53e83),
	.w4(32'h3aa54f7a),
	.w5(32'hb97c29b7),
	.w6(32'h3aabe622),
	.w7(32'h3a884e73),
	.w8(32'hba263f89),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b534b),
	.w1(32'hbaadac09),
	.w2(32'hba37d7e2),
	.w3(32'hb8b6ef4f),
	.w4(32'hbad60362),
	.w5(32'hba951615),
	.w6(32'hb9538987),
	.w7(32'hba098035),
	.w8(32'h3924f7fc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984b5e4),
	.w1(32'h3a498c46),
	.w2(32'hba3ce04b),
	.w3(32'h3a658a86),
	.w4(32'hba34d518),
	.w5(32'hba0c4987),
	.w6(32'h3aa31e8b),
	.w7(32'hba9ac923),
	.w8(32'hba8d0069),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39579847),
	.w1(32'h3a2605fc),
	.w2(32'hba8e59a9),
	.w3(32'h39ae3b74),
	.w4(32'hba2b1eb8),
	.w5(32'hb9f89916),
	.w6(32'h3a665add),
	.w7(32'hba0657e5),
	.w8(32'hba91d7e9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b82ef),
	.w1(32'hba21669e),
	.w2(32'hba2b5f1a),
	.w3(32'hba47af37),
	.w4(32'hba8cd726),
	.w5(32'hbae75804),
	.w6(32'hba635a09),
	.w7(32'hba718d06),
	.w8(32'hbad3d66e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba781d52),
	.w1(32'hba60c0e6),
	.w2(32'h3a193060),
	.w3(32'hbab82d81),
	.w4(32'hba0b7285),
	.w5(32'hba3f4d13),
	.w6(32'hbaaf74d1),
	.w7(32'hb936ec27),
	.w8(32'hb96a0f1b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fea4c),
	.w1(32'hbaae85cd),
	.w2(32'hbb02e6d2),
	.w3(32'hbb0018c1),
	.w4(32'hba997f4f),
	.w5(32'hbae75a63),
	.w6(32'hba4abb45),
	.w7(32'hba6b4ee8),
	.w8(32'hbabf1e8b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47b972),
	.w1(32'hba231586),
	.w2(32'hb8396f5e),
	.w3(32'hbacac303),
	.w4(32'hb9028b3b),
	.w5(32'h39b0e0d4),
	.w6(32'hba20b675),
	.w7(32'hb9e4e61f),
	.w8(32'hb91a0fab),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba521e01),
	.w1(32'hba16d6b1),
	.w2(32'h399af900),
	.w3(32'h3a173a8f),
	.w4(32'h37e3ea27),
	.w5(32'hb7b5aa59),
	.w6(32'hb9c43fa8),
	.w7(32'h3903dfd0),
	.w8(32'h394088db),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a72e5),
	.w1(32'h389b6a21),
	.w2(32'hba2f8f56),
	.w3(32'hba224a4f),
	.w4(32'hba437902),
	.w5(32'hba6f14a8),
	.w6(32'h394465e1),
	.w7(32'hba1aaf4b),
	.w8(32'hba46fc94),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d342f),
	.w1(32'h3a74ae4b),
	.w2(32'h3aa0d9f7),
	.w3(32'hb6c273b5),
	.w4(32'hb82c077e),
	.w5(32'h39e627dd),
	.w6(32'h39b9ceeb),
	.w7(32'hba02fb2f),
	.w8(32'hb9b26a07),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba196895),
	.w1(32'hb96d81a9),
	.w2(32'h390378d9),
	.w3(32'hb83dc512),
	.w4(32'hb937e6a6),
	.w5(32'hba4ee433),
	.w6(32'hb904ba66),
	.w7(32'hb966b1f5),
	.w8(32'hba5e537f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820c97),
	.w1(32'hbb005c54),
	.w2(32'hb6e5fcc9),
	.w3(32'hba4ab065),
	.w4(32'h39a65650),
	.w5(32'h398c5633),
	.w6(32'hba8e1383),
	.w7(32'h38ebff1d),
	.w8(32'h39e27769),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992e655),
	.w1(32'hbabc763c),
	.w2(32'hbb1f7149),
	.w3(32'hbaa44aa9),
	.w4(32'hbaf48bde),
	.w5(32'hbafe4c9a),
	.w6(32'hba1833e4),
	.w7(32'hbb0a70a7),
	.w8(32'hbae89480),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba666301),
	.w1(32'hba98b53f),
	.w2(32'hbb00ce43),
	.w3(32'hba358d39),
	.w4(32'hbad7ca09),
	.w5(32'hbaec2ba0),
	.w6(32'hb9610697),
	.w7(32'hbadbc01e),
	.w8(32'hbaec46e6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03223b),
	.w1(32'hbab64cc4),
	.w2(32'hba6f2f44),
	.w3(32'hbab2a5f2),
	.w4(32'hbb15b4d3),
	.w5(32'hba88182c),
	.w6(32'hba7f1cd1),
	.w7(32'hbb26eeba),
	.w8(32'hbb07224b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb8f8b),
	.w1(32'hb87727fd),
	.w2(32'hba86b0b4),
	.w3(32'hba188f21),
	.w4(32'h3a5a4fb8),
	.w5(32'h3a16247c),
	.w6(32'h382a1ebe),
	.w7(32'h3ad357df),
	.w8(32'h39d1f02d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba980da1),
	.w1(32'h390df143),
	.w2(32'hbb384c2e),
	.w3(32'hbb198440),
	.w4(32'hbaa936c4),
	.w5(32'hbb888aa1),
	.w6(32'hbafae211),
	.w7(32'hbadfbc52),
	.w8(32'hbb016e51),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399670d9),
	.w1(32'h3943d2fd),
	.w2(32'h3a2c3723),
	.w3(32'hbb181024),
	.w4(32'hbb3fee20),
	.w5(32'hbb11b549),
	.w6(32'hbab30dc4),
	.w7(32'hbb425981),
	.w8(32'hbace4369),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a93fc6),
	.w1(32'hba7e295b),
	.w2(32'hb8c12e2c),
	.w3(32'hba84405b),
	.w4(32'hba40ef1f),
	.w5(32'hb9d47cd0),
	.w6(32'hba9098d6),
	.w7(32'hb9f7a1a2),
	.w8(32'hb98ed720),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3833f61b),
	.w1(32'h38aef1d8),
	.w2(32'hba1bca87),
	.w3(32'h38480c48),
	.w4(32'h39099f28),
	.w5(32'hb93d076b),
	.w6(32'h396f0124),
	.w7(32'hb9973be6),
	.w8(32'hb9c94ac2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fd1b7),
	.w1(32'hba1329e6),
	.w2(32'hba8ff1a3),
	.w3(32'hb887d187),
	.w4(32'hba38b9fa),
	.w5(32'hb9bc00dd),
	.w6(32'h395c642d),
	.w7(32'hba3dcf47),
	.w8(32'hba5dd22b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9a7ca),
	.w1(32'hb9de24d0),
	.w2(32'h39bec7d1),
	.w3(32'hba9fe781),
	.w4(32'h39aa527f),
	.w5(32'h39996144),
	.w6(32'hba5327ce),
	.w7(32'h39aaed61),
	.w8(32'h399a4d83),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9e638),
	.w1(32'h399b3bdd),
	.w2(32'hba428853),
	.w3(32'hb9950cde),
	.w4(32'h3a325237),
	.w5(32'h3a8e2108),
	.w6(32'hba471cb8),
	.w7(32'hb9b8b054),
	.w8(32'h3832b245),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0699c5),
	.w1(32'hb8f54095),
	.w2(32'hb7e9876f),
	.w3(32'h3a4d500a),
	.w4(32'hb91485c3),
	.w5(32'hb9a7986e),
	.w6(32'hb5b6553d),
	.w7(32'h38f0be16),
	.w8(32'hb8a950bd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c83517),
	.w1(32'hb92b02eb),
	.w2(32'hb7ac75c1),
	.w3(32'hb95f6d3a),
	.w4(32'hb986aa43),
	.w5(32'hba3a3c3e),
	.w6(32'hb953973c),
	.w7(32'hba6507c9),
	.w8(32'hbb12db27),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf80238),
	.w1(32'hbb3f9a92),
	.w2(32'hb7a20a07),
	.w3(32'hbb23e56a),
	.w4(32'hba54fc26),
	.w5(32'hba66b952),
	.w6(32'hbb64758a),
	.w7(32'hba1964c0),
	.w8(32'hba52a25a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a669fe6),
	.w1(32'h3a268848),
	.w2(32'hba2e83f5),
	.w3(32'h3a0860f1),
	.w4(32'h3953158f),
	.w5(32'h39fefb35),
	.w6(32'hb8e0b950),
	.w7(32'hba0e4169),
	.w8(32'hb8670686),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eac863),
	.w1(32'hb912250e),
	.w2(32'hba60e11d),
	.w3(32'h3905947f),
	.w4(32'hbab190aa),
	.w5(32'hbae3f12d),
	.w6(32'h38081387),
	.w7(32'hba81e3b7),
	.w8(32'hbaabd5aa),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f40b72),
	.w1(32'hbaac265b),
	.w2(32'h38ffed71),
	.w3(32'hbaf5d346),
	.w4(32'hba9f4c86),
	.w5(32'hbadb9fd7),
	.w6(32'hbb16ce6b),
	.w7(32'hbabdc173),
	.w8(32'hbab40bd0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c2cf43),
	.w1(32'h395b9b21),
	.w2(32'hb73a3d05),
	.w3(32'hb9ca8561),
	.w4(32'hb9a88472),
	.w5(32'hba0e54a2),
	.w6(32'hb9259f10),
	.w7(32'hb9b3c2a4),
	.w8(32'hb95e5ab3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ae118),
	.w1(32'hba30eb75),
	.w2(32'hbafedfa2),
	.w3(32'hba80c7e6),
	.w4(32'hbb1e5299),
	.w5(32'hba876b40),
	.w6(32'hba9dbdce),
	.w7(32'hbb274a30),
	.w8(32'hba87c9b5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba378e4e),
	.w1(32'hba8777d4),
	.w2(32'hbae11081),
	.w3(32'hbab20c37),
	.w4(32'hbb11fa4a),
	.w5(32'hbb1d878c),
	.w6(32'hbabbdf6d),
	.w7(32'hbb198103),
	.w8(32'hbb418f35),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb5ffd),
	.w1(32'hbacb5ce1),
	.w2(32'h3ab73494),
	.w3(32'hba9e74ca),
	.w4(32'h39052698),
	.w5(32'hb7ceaa94),
	.w6(32'hbafe2a8b),
	.w7(32'h3a756f37),
	.w8(32'h3a2d3652),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99810a),
	.w1(32'h3a27ba87),
	.w2(32'hba582858),
	.w3(32'hb9d6538d),
	.w4(32'hba894296),
	.w5(32'hba1f86d4),
	.w6(32'h38e631ca),
	.w7(32'hba8884d9),
	.w8(32'hba817679),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfdbac),
	.w1(32'hbb5c4b68),
	.w2(32'hbb324de2),
	.w3(32'hbaee1f98),
	.w4(32'hbb019097),
	.w5(32'hbb508e68),
	.w6(32'hbb3f26a5),
	.w7(32'hbb420814),
	.w8(32'hbb79663b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9735847),
	.w1(32'h39deb082),
	.w2(32'hba638487),
	.w3(32'h38d58bd4),
	.w4(32'hba99822c),
	.w5(32'hba62bea3),
	.w6(32'hb8618536),
	.w7(32'hba686f64),
	.w8(32'hba010687),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadcccd),
	.w1(32'hba52c7ff),
	.w2(32'hbac5b223),
	.w3(32'hbad30a23),
	.w4(32'hba9c894e),
	.w5(32'hbaff40c7),
	.w6(32'hbac7e6e9),
	.w7(32'hbb0a92b2),
	.w8(32'hbb0b104d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad05a25),
	.w1(32'hba763323),
	.w2(32'hb98b3180),
	.w3(32'hba559656),
	.w4(32'hb981cb6c),
	.w5(32'hb95705c2),
	.w6(32'hbaa8d60c),
	.w7(32'hb9c4ed1b),
	.w8(32'hb7f3cb2b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba167264),
	.w1(32'hba406525),
	.w2(32'hba8bab8e),
	.w3(32'hbaa60e51),
	.w4(32'h39b8648d),
	.w5(32'h39f01711),
	.w6(32'hba038fb5),
	.w7(32'hb87f7516),
	.w8(32'hb6d1d93b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9288996),
	.w1(32'h390c77cd),
	.w2(32'hba9651ef),
	.w3(32'hbaa61c45),
	.w4(32'hba9ce8ae),
	.w5(32'hba8c6b26),
	.w6(32'h390b9140),
	.w7(32'hba8c24dd),
	.w8(32'hbac9d92a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb428d1e),
	.w1(32'hbb3b529c),
	.w2(32'hbaccf84a),
	.w3(32'hbad18879),
	.w4(32'hbaaf4f57),
	.w5(32'hbac2422b),
	.w6(32'hbaa975c5),
	.w7(32'hba210fcf),
	.w8(32'hba68f2e1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef85d6),
	.w1(32'hba0a4382),
	.w2(32'hb84aca83),
	.w3(32'hba4b25ab),
	.w4(32'hb87a1b0b),
	.w5(32'hb79ee854),
	.w6(32'hba1b6378),
	.w7(32'hb7990886),
	.w8(32'hb5f155d3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66e756),
	.w1(32'hba8727eb),
	.w2(32'hba785c2a),
	.w3(32'hba671cfc),
	.w4(32'hbad209d4),
	.w5(32'hbacc6722),
	.w6(32'hba4f6ce2),
	.w7(32'hbac1e348),
	.w8(32'hbab04ca8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba759ecc),
	.w1(32'hba73c54f),
	.w2(32'hba3ad4df),
	.w3(32'hba881ffb),
	.w4(32'hb9c9e9eb),
	.w5(32'hba278439),
	.w6(32'hba643c4d),
	.w7(32'hba52453c),
	.w8(32'hb9a3833d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971a9f4),
	.w1(32'hb980180f),
	.w2(32'hb90821ce),
	.w3(32'hb9e57ea9),
	.w4(32'hba0fef1a),
	.w5(32'hb9b41583),
	.w6(32'hb9edc549),
	.w7(32'hb8f4e5eb),
	.w8(32'hb9d46e1d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eeb7ad),
	.w1(32'h37e33b39),
	.w2(32'h388c0e3b),
	.w3(32'h37ae76c6),
	.w4(32'h37d8e13c),
	.w5(32'h38944fde),
	.w6(32'h376f70f8),
	.w7(32'h380be676),
	.w8(32'h389e82a5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c0bd84),
	.w1(32'h3a10f23a),
	.w2(32'h3a43d278),
	.w3(32'hb9309ea1),
	.w4(32'h39e4b385),
	.w5(32'h3a3f2528),
	.w6(32'hb8893e26),
	.w7(32'h39c907c8),
	.w8(32'h3a1f34cf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a326956),
	.w1(32'h3aa4ef32),
	.w2(32'h3a64d628),
	.w3(32'hb9f366c2),
	.w4(32'hb9279eb0),
	.w5(32'h376f4fc0),
	.w6(32'hb981d2e1),
	.w7(32'hba2051f5),
	.w8(32'hba14f401),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3db7e0),
	.w1(32'hb6cc6f4d),
	.w2(32'hb9247c37),
	.w3(32'hba694df5),
	.w4(32'h39dc1b02),
	.w5(32'h394a977e),
	.w6(32'hba2f0a79),
	.w7(32'h3a069df2),
	.w8(32'h392a00d4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6de4c),
	.w1(32'hbaa1768e),
	.w2(32'hba7b9127),
	.w3(32'hbb414c7f),
	.w4(32'hbb3ce369),
	.w5(32'hbb3a0c18),
	.w6(32'hbaf206bc),
	.w7(32'hbb68b14b),
	.w8(32'hbb1cf460),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2003f0),
	.w1(32'hba0d3044),
	.w2(32'hb9ec98ad),
	.w3(32'hbadd3d2c),
	.w4(32'hbb07ed1b),
	.w5(32'hbb02a730),
	.w6(32'hba5d06d0),
	.w7(32'hba9959ec),
	.w8(32'hbab8a6b1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a7ade4),
	.w1(32'h389bf010),
	.w2(32'h38c9ba14),
	.w3(32'h38e38b22),
	.w4(32'h3898f038),
	.w5(32'h38d7e253),
	.w6(32'h391373c1),
	.w7(32'h38d8d3a9),
	.w8(32'h38fa3fb9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5cd9953),
	.w1(32'hb70fbecc),
	.w2(32'h34943141),
	.w3(32'h36c4dae9),
	.w4(32'hb68279cc),
	.w5(32'h35c4b709),
	.w6(32'h36e358af),
	.w7(32'hb65456c9),
	.w8(32'h35909f82),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6232c11),
	.w1(32'h38b5c9c0),
	.w2(32'h3899b0fe),
	.w3(32'h36ee90df),
	.w4(32'h389619ec),
	.w5(32'h38a64aba),
	.w6(32'h38a50756),
	.w7(32'h380d09da),
	.w8(32'h385abf28),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7057c8),
	.w1(32'hb7c2e422),
	.w2(32'hb9d1109e),
	.w3(32'hb8866da2),
	.w4(32'hbaa196c6),
	.w5(32'hbab2139a),
	.w6(32'h3948e109),
	.w7(32'hba538b55),
	.w8(32'hba6851ea),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904b70c),
	.w1(32'hb8255823),
	.w2(32'h38ffe117),
	.w3(32'hba13e343),
	.w4(32'hba202cf0),
	.w5(32'hb99f0883),
	.w6(32'hba097eca),
	.w7(32'hba21be20),
	.w8(32'hb9ba2738),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2826b),
	.w1(32'hb96a6702),
	.w2(32'hb9ee27e7),
	.w3(32'h396ad53e),
	.w4(32'hb8ba9cc0),
	.w5(32'hb9b87904),
	.w6(32'h39a32fed),
	.w7(32'h3806847b),
	.w8(32'hb9b0b315),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fbd068),
	.w1(32'h38d8b02d),
	.w2(32'h39e16304),
	.w3(32'hba0b8c7a),
	.w4(32'hba29170f),
	.w5(32'hb912c8f0),
	.w6(32'hb96c9bed),
	.w7(32'hb9575c42),
	.w8(32'h39fdb752),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09ad19),
	.w1(32'h39d2eb49),
	.w2(32'h3888f392),
	.w3(32'hb949128f),
	.w4(32'hb9cc68d1),
	.w5(32'hba3947e4),
	.w6(32'hb8e96851),
	.w7(32'hba2276ed),
	.w8(32'hba6d3f91),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4abef3),
	.w1(32'h3a952c24),
	.w2(32'h3a5e0eaa),
	.w3(32'h3a2aa73c),
	.w4(32'h3a029750),
	.w5(32'h3a7151b6),
	.w6(32'h3a6bf31f),
	.w7(32'h3984541a),
	.w8(32'h3a05ceb0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9514df),
	.w1(32'h3a009685),
	.w2(32'h3a50d3c3),
	.w3(32'h3a0da077),
	.w4(32'hb9d9111c),
	.w5(32'hb84535cc),
	.w6(32'h3a9b4a2f),
	.w7(32'h39845eed),
	.w8(32'h3a05533d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d243d5),
	.w1(32'hb73fd103),
	.w2(32'hba8d8b3a),
	.w3(32'hbb1390f2),
	.w4(32'hbb2a5fe6),
	.w5(32'hbb1e3c14),
	.w6(32'hb9ba74a7),
	.w7(32'hbae79a83),
	.w8(32'hbac58dde),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3671a528),
	.w1(32'hb6ef22e5),
	.w2(32'h369d3579),
	.w3(32'hb7479712),
	.w4(32'hb789fd41),
	.w5(32'hb5ae7dde),
	.w6(32'h365ef7de),
	.w7(32'hb74d0fba),
	.w8(32'hb5ecc84e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3769e4e9),
	.w1(32'hb7a9bd89),
	.w2(32'h378ee9e0),
	.w3(32'h372aa494),
	.w4(32'hb7f4c650),
	.w5(32'h37585f22),
	.w6(32'h35e9282f),
	.w7(32'hb7e50057),
	.w8(32'h37820835),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379c5e07),
	.w1(32'hb6d2f146),
	.w2(32'h3719480e),
	.w3(32'h378c9784),
	.w4(32'hb676680d),
	.w5(32'h372215e4),
	.w6(32'h378d9f77),
	.w7(32'hb4b11637),
	.w8(32'h378168e9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e70196),
	.w1(32'h368a34ea),
	.w2(32'hb8830c15),
	.w3(32'h38ea7506),
	.w4(32'h3780ec14),
	.w5(32'hb899011e),
	.w6(32'h38c0cd2f),
	.w7(32'hb553cba4),
	.w8(32'hb87514d4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2182b8),
	.w1(32'h39f15279),
	.w2(32'hb8b8f301),
	.w3(32'h38efec96),
	.w4(32'hb92543b4),
	.w5(32'hb9602d42),
	.w6(32'h3a911a62),
	.w7(32'h3a0f0060),
	.w8(32'hb942e74a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4d3b0),
	.w1(32'hba888dfe),
	.w2(32'hba833f2a),
	.w3(32'hbaab0f35),
	.w4(32'hba991f6e),
	.w5(32'hba9da3f6),
	.w6(32'hba55754c),
	.w7(32'hba36157b),
	.w8(32'hb99fd523),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2bccc),
	.w1(32'h398b9717),
	.w2(32'hb990f83c),
	.w3(32'hb816a408),
	.w4(32'h3a396cb6),
	.w5(32'h398794e8),
	.w6(32'hba135d3d),
	.w7(32'hb6342758),
	.w8(32'h389288c8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dc0408),
	.w1(32'h37b0846c),
	.w2(32'hb903761c),
	.w3(32'h38906c47),
	.w4(32'h387bcc35),
	.w5(32'hb87562c8),
	.w6(32'hb8e72aef),
	.w7(32'hb7529070),
	.w8(32'h37ac8773),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8f861),
	.w1(32'hba6b7cb5),
	.w2(32'hba838507),
	.w3(32'hbb632964),
	.w4(32'hbb19bad7),
	.w5(32'hbb03e162),
	.w6(32'hbb4d98fd),
	.w7(32'hbb397684),
	.w8(32'hbaef777d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a2a74),
	.w1(32'h3a0bd100),
	.w2(32'h38cc85f5),
	.w3(32'h399814ff),
	.w4(32'hb9d7e1a3),
	.w5(32'hb963641c),
	.w6(32'h3a23e5de),
	.w7(32'hba41291c),
	.w8(32'hba0d9d17),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cc2ac),
	.w1(32'h39991e54),
	.w2(32'hb90dafe7),
	.w3(32'hb8c586eb),
	.w4(32'hb94226c4),
	.w5(32'hb950c401),
	.w6(32'h3917aab7),
	.w7(32'hb8b74058),
	.w8(32'hb9c3612f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6abc84),
	.w1(32'h3a7df396),
	.w2(32'h3a008c2e),
	.w3(32'h3a9174ab),
	.w4(32'h3ab60ea2),
	.w5(32'h3a874484),
	.w6(32'h3a8c5684),
	.w7(32'h3abe30c2),
	.w8(32'h3a9f2d82),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d68518),
	.w1(32'hba8654f0),
	.w2(32'hba4a9878),
	.w3(32'hbac86187),
	.w4(32'hbb0fbe4a),
	.w5(32'hba90654f),
	.w6(32'hba165730),
	.w7(32'hba904fd7),
	.w8(32'hba66f95d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993269f),
	.w1(32'h39ceb521),
	.w2(32'h3976330f),
	.w3(32'hb897c9da),
	.w4(32'h39f65de9),
	.w5(32'h39f330a7),
	.w6(32'h3a49aa9a),
	.w7(32'h3aa7f6df),
	.w8(32'h3a133a8d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ec972),
	.w1(32'hb9183a84),
	.w2(32'hba16371c),
	.w3(32'hba34166b),
	.w4(32'h374a3d6b),
	.w5(32'hba36acf6),
	.w6(32'hb96e9461),
	.w7(32'h39c9349e),
	.w8(32'hb909b829),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0d247),
	.w1(32'h3956835f),
	.w2(32'hb98c10f6),
	.w3(32'h3a008cd2),
	.w4(32'h3a471650),
	.w5(32'h3815e8f5),
	.w6(32'h38a76bb5),
	.w7(32'h39af34ff),
	.w8(32'h389e509a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb792b59e),
	.w1(32'hb9103d57),
	.w2(32'hb88882f8),
	.w3(32'hb8664ac4),
	.w4(32'hb9690001),
	.w5(32'hb8a1463a),
	.w6(32'hb80c4d4f),
	.w7(32'hb91e5279),
	.w8(32'hb860fd1a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e292c),
	.w1(32'hb86e7eea),
	.w2(32'h388d0475),
	.w3(32'hb89ea041),
	.w4(32'hb9536a2b),
	.w5(32'hb8b1959a),
	.w6(32'h37eccb78),
	.w7(32'hb90827fe),
	.w8(32'hb6042012),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a780d),
	.w1(32'hba31d2f0),
	.w2(32'hba6b1b35),
	.w3(32'hba3c42a8),
	.w4(32'hba7e55d0),
	.w5(32'hba86db4c),
	.w6(32'hb9661692),
	.w7(32'hba0e5ad0),
	.w8(32'hba0d2db4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9905fa1),
	.w1(32'hb8ed4c45),
	.w2(32'hb93fff41),
	.w3(32'hb967501f),
	.w4(32'h39de2d74),
	.w5(32'h37fbaa8c),
	.w6(32'h392fb42c),
	.w7(32'h3a3e99ef),
	.w8(32'h3948a5ff),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2de0f1),
	.w1(32'hb9a37cdb),
	.w2(32'hba08c187),
	.w3(32'hb9918cb6),
	.w4(32'h38bac4c0),
	.w5(32'hb889f92c),
	.w6(32'hb9239955),
	.w7(32'h3985380f),
	.w8(32'hb8ab4ad3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35aae324),
	.w1(32'hb6c328d2),
	.w2(32'h3638c3f6),
	.w3(32'h36cabf3a),
	.w4(32'hb5fba171),
	.w5(32'h3719c995),
	.w6(32'h36da8873),
	.w7(32'h36121a3d),
	.w8(32'h3779b475),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85f9e82),
	.w1(32'hb8285e0b),
	.w2(32'hb82cb771),
	.w3(32'hb5caa902),
	.w4(32'hb7b52131),
	.w5(32'hb7160f3c),
	.w6(32'h3711db3a),
	.w7(32'hb6c7813c),
	.w8(32'hb6e83f9e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ecc8b),
	.w1(32'h39013336),
	.w2(32'h3963e8d4),
	.w3(32'hb9f3aa45),
	.w4(32'hba26ed50),
	.w5(32'hba194637),
	.w6(32'h38ec49bc),
	.w7(32'hb9607564),
	.w8(32'hba275d38),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ac3be),
	.w1(32'hbad65abb),
	.w2(32'hbb0f404d),
	.w3(32'hba8d3f4a),
	.w4(32'hbaebdee8),
	.w5(32'hbadffaf3),
	.w6(32'hb944d3c0),
	.w7(32'hba3516c7),
	.w8(32'hbab03c14),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b45d1),
	.w1(32'hb8cbedc4),
	.w2(32'hb9870ee9),
	.w3(32'hb9062994),
	.w4(32'hb7c19c53),
	.w5(32'hb808c0c9),
	.w6(32'hb88e2db5),
	.w7(32'h38d39b4c),
	.w8(32'h399013cb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b31b73),
	.w1(32'h3995d24b),
	.w2(32'hb9d8f7d1),
	.w3(32'h3a18da0b),
	.w4(32'h3a5278db),
	.w5(32'h396f552b),
	.w6(32'h3a3b83b0),
	.w7(32'h3aaa78d6),
	.w8(32'h3a124c15),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998bff6),
	.w1(32'h39dcdccf),
	.w2(32'hb877f162),
	.w3(32'h39949ad0),
	.w4(32'h39f63b5a),
	.w5(32'h39ef9807),
	.w6(32'h3a928767),
	.w7(32'h3a5ff559),
	.w8(32'h39677dba),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9265f),
	.w1(32'hb9ffdd5e),
	.w2(32'hb8ceecf4),
	.w3(32'hba0c0ef1),
	.w4(32'hb9f1fc79),
	.w5(32'hb88e730d),
	.w6(32'hb9a0dab6),
	.w7(32'hb99ce99d),
	.w8(32'hb9482236),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933b300),
	.w1(32'hb9c1f536),
	.w2(32'hba552808),
	.w3(32'hb9c77fc3),
	.w4(32'h3821faa0),
	.w5(32'h38036d55),
	.w6(32'h3a2c5c0e),
	.w7(32'h38a1ca4d),
	.w8(32'h3967b2c6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9179e),
	.w1(32'hb9c472c1),
	.w2(32'hb9e2f659),
	.w3(32'hb8a9b07d),
	.w4(32'h361648e2),
	.w5(32'hb933fb8c),
	.w6(32'h39199e85),
	.w7(32'hb846a07d),
	.w8(32'h38581222),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule