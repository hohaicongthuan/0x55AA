module layer_8_featuremap_247(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80e6d8),
	.w1(32'hba03abce),
	.w2(32'h3ac8ac22),
	.w3(32'hbb34d6e4),
	.w4(32'hbbe12554),
	.w5(32'hb9c22019),
	.w6(32'hbab016cf),
	.w7(32'h3a404a96),
	.w8(32'h3b2b1104),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb222a1),
	.w1(32'hbad82e5a),
	.w2(32'hbb915458),
	.w3(32'hbbd24ea9),
	.w4(32'hbac6cf89),
	.w5(32'hbba6513b),
	.w6(32'hba6504f6),
	.w7(32'hba8c7d7b),
	.w8(32'h3b710819),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ae2a95),
	.w1(32'h3c363dae),
	.w2(32'h3c2d8d51),
	.w3(32'hbb2629eb),
	.w4(32'h3c5352af),
	.w5(32'h3c4f4cff),
	.w6(32'h3a04efd1),
	.w7(32'hbafa2098),
	.w8(32'h39b8d770),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ece06),
	.w1(32'h3b960e1c),
	.w2(32'h3c77e614),
	.w3(32'h3c19080e),
	.w4(32'h3bca7aae),
	.w5(32'h3c2d9cbc),
	.w6(32'h3b19db23),
	.w7(32'h3bf64511),
	.w8(32'h3b95e0c3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b0a70),
	.w1(32'h3a323901),
	.w2(32'h39870d24),
	.w3(32'h3c6993d7),
	.w4(32'hbb482134),
	.w5(32'h3abd10be),
	.w6(32'hba3321fd),
	.w7(32'hbb0d6d71),
	.w8(32'hbb93836a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b3f83),
	.w1(32'hbc630b63),
	.w2(32'hbcf0686d),
	.w3(32'h3aa5f733),
	.w4(32'hbc57e6e6),
	.w5(32'hbcd946b3),
	.w6(32'hbb9a9fa0),
	.w7(32'hbc38b793),
	.w8(32'hbbe39b04),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5a6ec),
	.w1(32'h3b9b6884),
	.w2(32'h3bd5c30a),
	.w3(32'hbce348c1),
	.w4(32'h3b4fd266),
	.w5(32'h3c09525e),
	.w6(32'h3a9154cc),
	.w7(32'h3b842ec1),
	.w8(32'h39e3a4fd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa2277),
	.w1(32'h3a96cce4),
	.w2(32'hbb6ad832),
	.w3(32'h3c1482dd),
	.w4(32'hbbafadc3),
	.w5(32'hbc1d0563),
	.w6(32'hbbf2c426),
	.w7(32'h3a083214),
	.w8(32'hbb111373),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ab87f),
	.w1(32'h3ab451a3),
	.w2(32'h3bb87566),
	.w3(32'h3b74cd7b),
	.w4(32'hba7ae327),
	.w5(32'h3ac5197b),
	.w6(32'hbb118f8d),
	.w7(32'h398dc860),
	.w8(32'hb96f97aa),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56a27f),
	.w1(32'h3b7c827e),
	.w2(32'h3c14d06b),
	.w3(32'hb98db954),
	.w4(32'h3bdd42f8),
	.w5(32'h3b39f2a4),
	.w6(32'h3b2b1bd6),
	.w7(32'h3be1efa1),
	.w8(32'h3a7aee68),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b6867f),
	.w1(32'hbc1303ab),
	.w2(32'hbaccc556),
	.w3(32'h3ac72f54),
	.w4(32'h3b905c87),
	.w5(32'hb9c2c622),
	.w6(32'hbc00197f),
	.w7(32'h3b548c71),
	.w8(32'h3c61769b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aa261),
	.w1(32'h3c0c8ee5),
	.w2(32'h3becff00),
	.w3(32'h3baa138b),
	.w4(32'h3b360182),
	.w5(32'h3bec0bf7),
	.w6(32'h3c25150b),
	.w7(32'h3b4bae3c),
	.w8(32'h3c02e940),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c132b6d),
	.w1(32'h3beeb980),
	.w2(32'h3be97b01),
	.w3(32'h3c0fd299),
	.w4(32'h3c014b93),
	.w5(32'h3bd78bb8),
	.w6(32'h3c440850),
	.w7(32'h3c122c28),
	.w8(32'h3c13ed43),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18e5cd),
	.w1(32'h3b2cbea9),
	.w2(32'h3b9ac3bf),
	.w3(32'h3c1fb802),
	.w4(32'h39891139),
	.w5(32'h3c0fc00c),
	.w6(32'hbb53d648),
	.w7(32'hbbfef595),
	.w8(32'hbb9fef7f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb50f90),
	.w1(32'hbb5f0c42),
	.w2(32'h3add3272),
	.w3(32'h3a74d16b),
	.w4(32'hbb6dba94),
	.w5(32'h391fb746),
	.w6(32'hbb10358d),
	.w7(32'h3ab01fa3),
	.w8(32'hbb31fc7d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbdefd),
	.w1(32'hbb97d08d),
	.w2(32'hbc2bc201),
	.w3(32'h3adeee38),
	.w4(32'h3bdc6fa2),
	.w5(32'h3b84afce),
	.w6(32'hb8b987e1),
	.w7(32'hbb9ec821),
	.w8(32'h3c26fe03),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8987cf),
	.w1(32'hbc113865),
	.w2(32'hbcab1a7a),
	.w3(32'h3c0d70bb),
	.w4(32'hbc8b7bfb),
	.w5(32'hbc7a3722),
	.w6(32'hbbacd212),
	.w7(32'hbc3b1a28),
	.w8(32'hbcb52efb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca42a1a),
	.w1(32'h3c29c032),
	.w2(32'h3bf952c9),
	.w3(32'hbb3d5e9b),
	.w4(32'h3c2093d3),
	.w5(32'h3c3580dc),
	.w6(32'h3c837945),
	.w7(32'h3c2ad912),
	.w8(32'h3bedc0f7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf69a12),
	.w1(32'h3c21cb6d),
	.w2(32'h3b675f3a),
	.w3(32'h3a07c9b6),
	.w4(32'h3bb17efc),
	.w5(32'h3b9a4a9f),
	.w6(32'h3b86695e),
	.w7(32'hbbd3b54a),
	.w8(32'h3bf6327d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bfd9d),
	.w1(32'h3a9245d2),
	.w2(32'h3b88adfd),
	.w3(32'hbba0bee5),
	.w4(32'h3abcf65a),
	.w5(32'h3aaa1dfa),
	.w6(32'hbaed7db2),
	.w7(32'h3aa2cc59),
	.w8(32'h3a899d6f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d8f75),
	.w1(32'h3b9a512f),
	.w2(32'hbb19f1ca),
	.w3(32'h3b8b8f8c),
	.w4(32'h3ad8250f),
	.w5(32'h3b1b72c4),
	.w6(32'h3b85deb1),
	.w7(32'h3bda9680),
	.w8(32'h3be620ad),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63be50),
	.w1(32'hbcb4f194),
	.w2(32'hbd27d7cb),
	.w3(32'hba70ea64),
	.w4(32'hbc789e97),
	.w5(32'hbc9f5356),
	.w6(32'hbc01912b),
	.w7(32'hbcd21dd6),
	.w8(32'hbc71b3ad),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce531a4),
	.w1(32'hbc3e1803),
	.w2(32'hbccad614),
	.w3(32'hbcde4f9a),
	.w4(32'hbb90146b),
	.w5(32'hbcd9cc37),
	.w6(32'hbc2c9dcb),
	.w7(32'hbc7684c1),
	.w8(32'hba1017e4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80a295),
	.w1(32'hbc46892c),
	.w2(32'hbcd982ae),
	.w3(32'hbc3567c8),
	.w4(32'hbb394678),
	.w5(32'hbc29d181),
	.w6(32'hbbd634e5),
	.w7(32'hbc4ccc7d),
	.w8(32'hba769ece),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb043e7),
	.w1(32'hba6a0de7),
	.w2(32'h398b2ce8),
	.w3(32'hbc088aa8),
	.w4(32'h3bc43246),
	.w5(32'h3c0be881),
	.w6(32'h3a7e7aa7),
	.w7(32'h3b65429b),
	.w8(32'h3aeb79ab),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b244229),
	.w1(32'hbacb46bf),
	.w2(32'hbb966ef6),
	.w3(32'h3a86f219),
	.w4(32'hbb8a3974),
	.w5(32'hb9ee3642),
	.w6(32'hbc0b6f74),
	.w7(32'hba88981f),
	.w8(32'h3b629b52),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c378d),
	.w1(32'hb9531821),
	.w2(32'h3b9362c9),
	.w3(32'hbc03d50f),
	.w4(32'h3bbeaa99),
	.w5(32'h3b82dcf8),
	.w6(32'h3be4959f),
	.w7(32'h3bec0b85),
	.w8(32'h3b1c8768),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9f94),
	.w1(32'h3b9d7f23),
	.w2(32'h3bbd3a87),
	.w3(32'h3a810df2),
	.w4(32'h3c03db48),
	.w5(32'hbab6d76b),
	.w6(32'h3ba0bfd7),
	.w7(32'h3ba02a4d),
	.w8(32'h3c4bab51),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beee69c),
	.w1(32'hbb440c4f),
	.w2(32'hbb1e36f6),
	.w3(32'h3a0c46a3),
	.w4(32'h3abcc8c7),
	.w5(32'h39d66eb0),
	.w6(32'hbbb6dea9),
	.w7(32'hba124690),
	.w8(32'hba8f84a8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43f413),
	.w1(32'h3ac9951b),
	.w2(32'h3b065d2a),
	.w3(32'hbaa42e67),
	.w4(32'hbb5163ce),
	.w5(32'h3ab76f0b),
	.w6(32'h39a9b679),
	.w7(32'h3aba014d),
	.w8(32'h3c76ea2b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccb1941),
	.w1(32'h3b486940),
	.w2(32'h3afc5bf7),
	.w3(32'h3cd39fbd),
	.w4(32'h3b498d03),
	.w5(32'h3b9f9cf2),
	.w6(32'hb7145809),
	.w7(32'h3abd47d3),
	.w8(32'h3a8bc6b1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75e660),
	.w1(32'h39bca44d),
	.w2(32'h39ced886),
	.w3(32'h3bbe71de),
	.w4(32'hba0f7d4c),
	.w5(32'h3b9936f5),
	.w6(32'h3aa189d3),
	.w7(32'h3b906602),
	.w8(32'h3c0fe3c2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be445f9),
	.w1(32'hbc06cd78),
	.w2(32'hbc0d5a26),
	.w3(32'h3b72ad2d),
	.w4(32'h3b766b50),
	.w5(32'hbc1ca247),
	.w6(32'hbb9059c4),
	.w7(32'h3a20bbd0),
	.w8(32'h3c0c0ed3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0da739),
	.w1(32'hbb16a630),
	.w2(32'hbc17c5ac),
	.w3(32'hbc218cf0),
	.w4(32'h3bdca274),
	.w5(32'hbb1ec1c8),
	.w6(32'hbbfd9645),
	.w7(32'hbbbf458e),
	.w8(32'h3c597422),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc7f24),
	.w1(32'h3bfcc5d0),
	.w2(32'h3c1b9ec6),
	.w3(32'hbbb6a553),
	.w4(32'h3c4c8a71),
	.w5(32'h3c691562),
	.w6(32'h3c640dd9),
	.w7(32'h3c80b5c0),
	.w8(32'h3c54f208),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ecadd),
	.w1(32'h3c0a9a54),
	.w2(32'hb91087aa),
	.w3(32'h3c707e64),
	.w4(32'h3b26fbcf),
	.w5(32'hbb1d686f),
	.w6(32'h3c000f98),
	.w7(32'h3c11ad63),
	.w8(32'hbae595f5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea1759),
	.w1(32'hbab60c9c),
	.w2(32'h393e3c1f),
	.w3(32'h3b274ede),
	.w4(32'hbb1dbc3c),
	.w5(32'hba0ba5bd),
	.w6(32'h3b42d783),
	.w7(32'h3ae8624a),
	.w8(32'hbbcb02f5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba638c29),
	.w1(32'hba873b18),
	.w2(32'h3930a76d),
	.w3(32'h3a3bb301),
	.w4(32'hba15c79b),
	.w5(32'h3a9a4f95),
	.w6(32'h3a7e6530),
	.w7(32'hb8e4c4f6),
	.w8(32'hb9f6b363),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0859),
	.w1(32'hbcb3b23b),
	.w2(32'hbd361be0),
	.w3(32'h3b009752),
	.w4(32'hbc1c94c6),
	.w5(32'hbd04d8cb),
	.w6(32'hbc8af57d),
	.w7(32'hbcf28021),
	.w8(32'hbcb59beb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0fe5ef),
	.w1(32'hbb84113c),
	.w2(32'hbc839721),
	.w3(32'hbcef620c),
	.w4(32'hbb0c8d87),
	.w5(32'hbbe3b873),
	.w6(32'h393be11c),
	.w7(32'hbb8201a9),
	.w8(32'h3b705175),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba173db),
	.w1(32'h39c73398),
	.w2(32'h3bec01ba),
	.w3(32'h3b8ba2c4),
	.w4(32'h3b1a5eb5),
	.w5(32'h3c14af5e),
	.w6(32'h3b94e94e),
	.w7(32'h3c09b2bc),
	.w8(32'h3b0ad4d2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab590fe),
	.w1(32'h3c162be1),
	.w2(32'h3a55fb53),
	.w3(32'h3bd0721f),
	.w4(32'h3b7bc6ce),
	.w5(32'h3bed1556),
	.w6(32'h3b26f63e),
	.w7(32'hbbf4bab2),
	.w8(32'hbc13bde9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dda8c),
	.w1(32'h3b952a0a),
	.w2(32'hb9e1f26b),
	.w3(32'hbbb85d98),
	.w4(32'hbb674eac),
	.w5(32'hbb027720),
	.w6(32'h3c120c30),
	.w7(32'h3c0628b9),
	.w8(32'h3b81c21a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70f178),
	.w1(32'h3c5e3816),
	.w2(32'h3cca7312),
	.w3(32'hbaba8c4b),
	.w4(32'h3b82c364),
	.w5(32'h3c6916a2),
	.w6(32'h3c82bfce),
	.w7(32'h3c70e27b),
	.w8(32'h3c11b2be),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e2faf),
	.w1(32'hbbe960c9),
	.w2(32'hbc7b059b),
	.w3(32'h3c4b01a7),
	.w4(32'hbbe80f10),
	.w5(32'hbc9b5344),
	.w6(32'hbc136be6),
	.w7(32'hbc5239cd),
	.w8(32'hbbe123f8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ec7ef),
	.w1(32'h3ab540d3),
	.w2(32'hbab2b315),
	.w3(32'hbc987ad0),
	.w4(32'h3b00eca5),
	.w5(32'hba9d37fd),
	.w6(32'hbb95e55a),
	.w7(32'hbb7a009f),
	.w8(32'h3b0f35ba),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf0d22),
	.w1(32'h3a2e320a),
	.w2(32'h3bb25709),
	.w3(32'h3bcc59be),
	.w4(32'hbacf16e6),
	.w5(32'h3bf8075e),
	.w6(32'h3b41465e),
	.w7(32'h3c1d5ab2),
	.w8(32'h3b8a262b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd45a21),
	.w1(32'hbcf05c02),
	.w2(32'hbd57fccd),
	.w3(32'h3c151fde),
	.w4(32'hbca07a98),
	.w5(32'hbd241337),
	.w6(32'hbc3c4212),
	.w7(32'hbc8f170f),
	.w8(32'hbc856218),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd38b235),
	.w1(32'hbce03e9d),
	.w2(32'hbd5db68b),
	.w3(32'hbce86f18),
	.w4(32'hbcc426c3),
	.w5(32'hbd387f47),
	.w6(32'hbc25907a),
	.w7(32'hbca0e19e),
	.w8(32'hbc34c90b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06b478),
	.w1(32'h3aeaa13e),
	.w2(32'h3aa3df5c),
	.w3(32'hbcfa4a2c),
	.w4(32'h3ad5d355),
	.w5(32'h3a47772d),
	.w6(32'hbb9d23aa),
	.w7(32'hbb681d61),
	.w8(32'h3ab6effa),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917cc7),
	.w1(32'hbaa0ebc9),
	.w2(32'h3ade5886),
	.w3(32'hbb5e68d2),
	.w4(32'h3abdab43),
	.w5(32'h3bfab0ab),
	.w6(32'h3b3c9af2),
	.w7(32'h3bb683a1),
	.w8(32'h399e5cb1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9862f2),
	.w1(32'h3b99808d),
	.w2(32'h3af16869),
	.w3(32'h3af23f13),
	.w4(32'h3aec24e9),
	.w5(32'h3b6892f7),
	.w6(32'h3bcb999a),
	.w7(32'hb9cf57cd),
	.w8(32'h3a6740bd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36004e),
	.w1(32'hbaa2847f),
	.w2(32'hba4f7cc8),
	.w3(32'h3b62a862),
	.w4(32'hba7b5ccd),
	.w5(32'h39768189),
	.w6(32'h3b366814),
	.w7(32'h3b5bb24b),
	.w8(32'h3b929fd7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b927cc7),
	.w1(32'hbb5c0992),
	.w2(32'h3ad2db58),
	.w3(32'h3bc0b614),
	.w4(32'h3aac4659),
	.w5(32'h39ee9401),
	.w6(32'hbb89a609),
	.w7(32'hbc120261),
	.w8(32'hb95c257e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdc365),
	.w1(32'h3b93d0f3),
	.w2(32'h3b69d672),
	.w3(32'hbbef0225),
	.w4(32'hba72082e),
	.w5(32'hbb9549df),
	.w6(32'h3b81fca6),
	.w7(32'h3947d68b),
	.w8(32'hbad1921b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee16eb),
	.w1(32'h3cad93e0),
	.w2(32'h3d0c0d9a),
	.w3(32'h3a139c83),
	.w4(32'h3cb67968),
	.w5(32'h3cf46c60),
	.w6(32'h3c90fb44),
	.w7(32'h3cbd0999),
	.w8(32'h3cccd56c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce6cd44),
	.w1(32'hbbd0a02e),
	.w2(32'hbcd5e99f),
	.w3(32'h3c9f884a),
	.w4(32'hbb8fd70d),
	.w5(32'hbce4c5ac),
	.w6(32'hbbdea2a0),
	.w7(32'hbc3e2051),
	.w8(32'hb9b27df2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6637c1),
	.w1(32'h3b770703),
	.w2(32'hbadc60e1),
	.w3(32'hbc88c345),
	.w4(32'h3b308ded),
	.w5(32'hbb99defa),
	.w6(32'h3b91952b),
	.w7(32'h3b254d0c),
	.w8(32'h3b016d57),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affed1f),
	.w1(32'h3a2b2054),
	.w2(32'h38bdc579),
	.w3(32'hbb3455ca),
	.w4(32'hbab55d90),
	.w5(32'h3b16f8e3),
	.w6(32'h3ba15562),
	.w7(32'h3b8a4486),
	.w8(32'h3a4752e0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b5598),
	.w1(32'hbca840d2),
	.w2(32'hbd3a608d),
	.w3(32'h3b37d765),
	.w4(32'hbc58d981),
	.w5(32'hbcd54ca4),
	.w6(32'hbc2d40e7),
	.w7(32'hbcaa7311),
	.w8(32'h3a456842),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd11617),
	.w1(32'h3b3eea6c),
	.w2(32'h3bcce9d1),
	.w3(32'hbcacfb9e),
	.w4(32'hb9a02979),
	.w5(32'h3b848a6f),
	.w6(32'h3c05c172),
	.w7(32'h3b786259),
	.w8(32'h3b4840fe),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c171973),
	.w1(32'hbbf118a8),
	.w2(32'hbb311b69),
	.w3(32'hba1c0155),
	.w4(32'h3a647281),
	.w5(32'h3be1eff3),
	.w6(32'hbb7eab47),
	.w7(32'h3b170911),
	.w8(32'hbadb388d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b980b20),
	.w1(32'hbb4e241e),
	.w2(32'h3bcd81ea),
	.w3(32'h3bd63ce8),
	.w4(32'hba1a6c5e),
	.w5(32'h39361254),
	.w6(32'hbbde8997),
	.w7(32'hb93c3053),
	.w8(32'h3bc797a2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54e935),
	.w1(32'hbab85a9b),
	.w2(32'h3b10d73e),
	.w3(32'h3b81ad49),
	.w4(32'hbba2f33e),
	.w5(32'hb99759f9),
	.w6(32'h3ae9b335),
	.w7(32'h3ba30c48),
	.w8(32'h3aef815c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39578ba4),
	.w1(32'hbb0dce02),
	.w2(32'hb9aa6828),
	.w3(32'h3b22e81c),
	.w4(32'hbb30d42b),
	.w5(32'hbabbb2d5),
	.w6(32'hbad60bd7),
	.w7(32'h3b523588),
	.w8(32'h3bb354cf),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f311e),
	.w1(32'hbb2d095f),
	.w2(32'hbc266cb1),
	.w3(32'h3a04def0),
	.w4(32'h3bee8d22),
	.w5(32'h3b36019b),
	.w6(32'hba8ca649),
	.w7(32'hbb898e1b),
	.w8(32'hbbb032ae),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2e0c3),
	.w1(32'h3a658791),
	.w2(32'h3b399933),
	.w3(32'hbbc11d6e),
	.w4(32'h3a72a8c3),
	.w5(32'hba8a074d),
	.w6(32'h3b9520f1),
	.w7(32'h3bde3ed8),
	.w8(32'h3c22de49),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fbed2),
	.w1(32'h3bbcd17a),
	.w2(32'h3c18038e),
	.w3(32'hbbe2f6b1),
	.w4(32'h3bad6f5c),
	.w5(32'h3b9e7e6a),
	.w6(32'h3be703ed),
	.w7(32'h3c00b01b),
	.w8(32'h3beef74d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48136f),
	.w1(32'hbc0f908f),
	.w2(32'hbc945e50),
	.w3(32'h3aa313b4),
	.w4(32'h3bd08436),
	.w5(32'hbbf6fc21),
	.w6(32'hbcc9f84d),
	.w7(32'hbba16cdd),
	.w8(32'h3c67286c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4297f5),
	.w1(32'hbc5e2556),
	.w2(32'hbcbcc063),
	.w3(32'hbc99e2ab),
	.w4(32'hbb2a7185),
	.w5(32'hbcb6c4b7),
	.w6(32'hbbee892c),
	.w7(32'hbc2ee463),
	.w8(32'hbb9d02ec),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d8ed0),
	.w1(32'hbb3c0b4d),
	.w2(32'hba8476ff),
	.w3(32'hbccafbc0),
	.w4(32'hbbbe65ff),
	.w5(32'h3acfcda0),
	.w6(32'hba03004a),
	.w7(32'hba28d5bc),
	.w8(32'h3be8981b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c016369),
	.w1(32'h3ce7619d),
	.w2(32'h3d226293),
	.w3(32'h3c0e6217),
	.w4(32'h3c139236),
	.w5(32'h3cdf79b6),
	.w6(32'h3ca8db02),
	.w7(32'h3cbda26d),
	.w8(32'h3ca822d6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc56b07),
	.w1(32'h3cbaf6c8),
	.w2(32'h3c9f5cc1),
	.w3(32'h3ce07187),
	.w4(32'h3be30531),
	.w5(32'h3bfb6257),
	.w6(32'h3ca22f51),
	.w7(32'h3c4f6de7),
	.w8(32'h3b9c5921),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d068f),
	.w1(32'h3b567653),
	.w2(32'h3bfaf6f9),
	.w3(32'h3c8dd388),
	.w4(32'h3b992336),
	.w5(32'h39a5d6dd),
	.w6(32'h3b6813ce),
	.w7(32'h3b38fca0),
	.w8(32'h3b2255f7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18067b),
	.w1(32'hbb8e6fa1),
	.w2(32'hbbd6a33a),
	.w3(32'h3abe7d43),
	.w4(32'h3ba49e3e),
	.w5(32'h3aee5894),
	.w6(32'h3b837345),
	.w7(32'h39a16d7a),
	.w8(32'h3b91f39b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ff21),
	.w1(32'hbbafc5d2),
	.w2(32'hbccc5c02),
	.w3(32'hbb3d9a81),
	.w4(32'hbb0ec79a),
	.w5(32'hbc9c7db3),
	.w6(32'hbb1901b4),
	.w7(32'hbb8e7c85),
	.w8(32'hb94da1bc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83f680),
	.w1(32'hbaa7a7fb),
	.w2(32'hbbe7e124),
	.w3(32'hbc8ec054),
	.w4(32'h3b379f1c),
	.w5(32'hbb3f6cc1),
	.w6(32'hba2b45d9),
	.w7(32'hbb47e000),
	.w8(32'hba5a80dd),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31fa2f),
	.w1(32'h3ad275a9),
	.w2(32'h3a24f90a),
	.w3(32'hbab00916),
	.w4(32'h36a517d6),
	.w5(32'hbb2c2e58),
	.w6(32'h3bb8e7bf),
	.w7(32'h3b8851e0),
	.w8(32'h3b866c29),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a7e7f),
	.w1(32'h3bbd6b6c),
	.w2(32'h3b49bd97),
	.w3(32'hba0586aa),
	.w4(32'h3b192d3a),
	.w5(32'h3b7db3bb),
	.w6(32'h3be528b0),
	.w7(32'h3b27fbd7),
	.w8(32'hbbd1b78c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76cb66),
	.w1(32'h3cbb8988),
	.w2(32'h3cfd1f3d),
	.w3(32'h3b94667b),
	.w4(32'h3c8b1096),
	.w5(32'h3ca2a48d),
	.w6(32'h3cb78c15),
	.w7(32'h3c585d0b),
	.w8(32'h3c8a6b19),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdfb822),
	.w1(32'h3bcd02a7),
	.w2(32'h3c57453b),
	.w3(32'h3c4af562),
	.w4(32'h3a6e3f49),
	.w5(32'h3c1dcf47),
	.w6(32'hbb82e7e4),
	.w7(32'hb91284dc),
	.w8(32'h3bf4e423),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b5d82),
	.w1(32'hbcbc93b6),
	.w2(32'hbce2096e),
	.w3(32'h3c063c2c),
	.w4(32'hbaa88d86),
	.w5(32'hbc8d37f0),
	.w6(32'hbcd2cce2),
	.w7(32'hbcc4305b),
	.w8(32'h39c508fd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6112f4),
	.w1(32'hbc085fc3),
	.w2(32'hbc56e931),
	.w3(32'hbcdb5909),
	.w4(32'hbb89fe0a),
	.w5(32'hbc40fff5),
	.w6(32'hb9477837),
	.w7(32'hbbaae7c3),
	.w8(32'h3b116894),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52f2c9),
	.w1(32'hbaafc782),
	.w2(32'hbaaf50da),
	.w3(32'hbc9544bf),
	.w4(32'hbba0fad6),
	.w5(32'hbbe4cbf3),
	.w6(32'h3bd6d667),
	.w7(32'hbbe31bf7),
	.w8(32'hbb2fe341),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc217ec),
	.w1(32'h3c03411f),
	.w2(32'h3bb7d11b),
	.w3(32'hbbadd02e),
	.w4(32'h3be7e81e),
	.w5(32'h3c32a210),
	.w6(32'hbbffa900),
	.w7(32'hba0669c0),
	.w8(32'h39d9911c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46959a),
	.w1(32'h3ac8803f),
	.w2(32'hb8cf6b3a),
	.w3(32'h3c2b057b),
	.w4(32'h3b285365),
	.w5(32'hbbd0abc8),
	.w6(32'h3b9eb823),
	.w7(32'h3ac23b82),
	.w8(32'hba307a2c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb2993),
	.w1(32'h392d2228),
	.w2(32'h3b3ac36d),
	.w3(32'hbb93d41e),
	.w4(32'hbb631deb),
	.w5(32'hbb37d139),
	.w6(32'h3ab69ca9),
	.w7(32'h3b4c7679),
	.w8(32'h3b9cefab),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12293f),
	.w1(32'hbbdec1bc),
	.w2(32'h39564a27),
	.w3(32'hbb13cabb),
	.w4(32'hbb2af6cf),
	.w5(32'hbae73680),
	.w6(32'h3b1ca131),
	.w7(32'h3b8c6a6c),
	.w8(32'h3b2b32c9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc66fd4),
	.w1(32'hbb9fa0de),
	.w2(32'hb9a92657),
	.w3(32'h3968e7b6),
	.w4(32'h3b0d62b7),
	.w5(32'h3b3474bf),
	.w6(32'hb998da57),
	.w7(32'hb9fae1dd),
	.w8(32'h3ae1cac9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4e616),
	.w1(32'h3a58dd49),
	.w2(32'hbc286551),
	.w3(32'h3b41fe9e),
	.w4(32'h3babefe2),
	.w5(32'hbb9e42a8),
	.w6(32'hbb9c26f8),
	.w7(32'hbc497ab8),
	.w8(32'hbb3bf87d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6f67e),
	.w1(32'h3cede1b7),
	.w2(32'h3d0644b9),
	.w3(32'hbb0011c4),
	.w4(32'h3c686f05),
	.w5(32'h3ca89b1d),
	.w6(32'h3cd80882),
	.w7(32'h3cb39e89),
	.w8(32'h3bde6ddf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0251dd),
	.w1(32'hbc085655),
	.w2(32'hbc7e05ad),
	.w3(32'h3c9150e8),
	.w4(32'hbb6e49b2),
	.w5(32'hbba91cda),
	.w6(32'hbbc99166),
	.w7(32'hbb79c65e),
	.w8(32'h3b3ac3f0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2be0b2),
	.w1(32'hba836946),
	.w2(32'hb94702bf),
	.w3(32'hbc2823a9),
	.w4(32'h3ae15749),
	.w5(32'h38259e87),
	.w6(32'hbb32af66),
	.w7(32'hba7fafcd),
	.w8(32'h3abb504f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff4e94),
	.w1(32'hba8ec766),
	.w2(32'hbb12a50a),
	.w3(32'hba2234bf),
	.w4(32'hba7e4139),
	.w5(32'hba182570),
	.w6(32'hba57e18a),
	.w7(32'hbacb7ed3),
	.w8(32'h3af93c7b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98c1ee),
	.w1(32'h3b2f81c7),
	.w2(32'hba51f0e1),
	.w3(32'h3b2259a1),
	.w4(32'hbb3ee751),
	.w5(32'h3b651465),
	.w6(32'h3bc637eb),
	.w7(32'h3b231dae),
	.w8(32'hbb08acd4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912f29),
	.w1(32'h3c0076bb),
	.w2(32'h3c1b7b58),
	.w3(32'hbb9c82c2),
	.w4(32'h3c529d21),
	.w5(32'h3c095fc9),
	.w6(32'h3ac02111),
	.w7(32'h3bd9759c),
	.w8(32'h3c0db2c1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5063e),
	.w1(32'hbce2c7c3),
	.w2(32'hbd57f71f),
	.w3(32'h3b615188),
	.w4(32'hbc797cd8),
	.w5(32'hbd025b8a),
	.w6(32'hbc0ee395),
	.w7(32'hbd02afe7),
	.w8(32'hbc82b2d1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd32f195),
	.w1(32'hbc3cab42),
	.w2(32'hbd102fd5),
	.w3(32'hbcfb6352),
	.w4(32'hbc4aced9),
	.w5(32'hbc8555a5),
	.w6(32'hbc48b9ad),
	.w7(32'hbccc740f),
	.w8(32'hbc6032c9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd169034),
	.w1(32'hbbd7e996),
	.w2(32'hbcd64c3c),
	.w3(32'hbd083085),
	.w4(32'hbbba4eb1),
	.w5(32'hbc4e050d),
	.w6(32'hbb13ec3d),
	.w7(32'hbce25d35),
	.w8(32'hbc98b252),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc935a9),
	.w1(32'hbb4d95de),
	.w2(32'hbaee5de3),
	.w3(32'hbc8acfa6),
	.w4(32'hba3b59a2),
	.w5(32'hbb52bddb),
	.w6(32'h3bad0424),
	.w7(32'h3b7f80d0),
	.w8(32'h3b9aaa1a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3ad87),
	.w1(32'hbab8c741),
	.w2(32'hbc42f581),
	.w3(32'h3baf5724),
	.w4(32'h3c02f893),
	.w5(32'h3b8ec215),
	.w6(32'hbc216079),
	.w7(32'hbbfe6f78),
	.w8(32'h3c02d46b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87039f),
	.w1(32'h3b16a189),
	.w2(32'h3ca5151f),
	.w3(32'hbc6af27f),
	.w4(32'hbb920aee),
	.w5(32'h3b8b6f7f),
	.w6(32'h3b204feb),
	.w7(32'h3c0864df),
	.w8(32'h3bd08e32),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c164667),
	.w1(32'hbc2f44c3),
	.w2(32'hbc63ba63),
	.w3(32'h3c24f7aa),
	.w4(32'hbaa3aa0d),
	.w5(32'hbb663742),
	.w6(32'hbc6d37cf),
	.w7(32'hbc07f9cb),
	.w8(32'hbbe66e49),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fbfbf),
	.w1(32'hbc4743a4),
	.w2(32'hbc70cd6b),
	.w3(32'hbb68bcb3),
	.w4(32'h3bc68eab),
	.w5(32'hbc087801),
	.w6(32'hbc2b8c1c),
	.w7(32'hbbe094e1),
	.w8(32'hbb8aefd2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84ddb5),
	.w1(32'h3c386ecb),
	.w2(32'h3b0d29ba),
	.w3(32'hbbedf93d),
	.w4(32'h3c37f20f),
	.w5(32'hbbab39f6),
	.w6(32'h3ab5b8f0),
	.w7(32'h3bcc208d),
	.w8(32'h3bd1c817),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be24c60),
	.w1(32'hbb82b32b),
	.w2(32'hbb838175),
	.w3(32'h3c2fa2b8),
	.w4(32'hbb315a0e),
	.w5(32'hbbde604f),
	.w6(32'hbbb55643),
	.w7(32'hbb871009),
	.w8(32'h38de8fe3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af68b36),
	.w1(32'hbb187ec7),
	.w2(32'h3a5723bd),
	.w3(32'h3a53ac74),
	.w4(32'h3b8f453d),
	.w5(32'h3b73d53e),
	.w6(32'hbb902f80),
	.w7(32'h39889771),
	.w8(32'h3b4b03e3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd72da),
	.w1(32'hbb26aa7f),
	.w2(32'h3b278eac),
	.w3(32'hba4f6478),
	.w4(32'hbb3b8515),
	.w5(32'h3b99e521),
	.w6(32'h3bce83f8),
	.w7(32'h3c153557),
	.w8(32'hbb195153),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4051d2),
	.w1(32'h3be8f0d5),
	.w2(32'h3c8c166b),
	.w3(32'h395e57d6),
	.w4(32'hbab6105b),
	.w5(32'h3c6d40eb),
	.w6(32'h3be8290a),
	.w7(32'h3c38c0ca),
	.w8(32'h3b670a29),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c752717),
	.w1(32'h3aa63d49),
	.w2(32'h3a902f35),
	.w3(32'h3c91bf17),
	.w4(32'h3ae240b6),
	.w5(32'h3b0e5b92),
	.w6(32'h3aac49f9),
	.w7(32'h3ace19c9),
	.w8(32'h3b8d029c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a7728),
	.w1(32'hba738a63),
	.w2(32'h3aba8eb9),
	.w3(32'h3b03f8aa),
	.w4(32'hba4af346),
	.w5(32'h3b623728),
	.w6(32'hbba20eee),
	.w7(32'hbb401e0f),
	.w8(32'h3bb050c1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c4b26),
	.w1(32'h3b996536),
	.w2(32'h3c05e04c),
	.w3(32'hbb66bc7e),
	.w4(32'h3b1d012d),
	.w5(32'h3b928dfe),
	.w6(32'hba9ca0a3),
	.w7(32'h3b5a10c8),
	.w8(32'h3b8eec73),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd72aa5),
	.w1(32'h3c21c409),
	.w2(32'h3c9e08f2),
	.w3(32'h3bf52ff7),
	.w4(32'h3c308832),
	.w5(32'h3c753d6e),
	.w6(32'h3c1217be),
	.w7(32'h3c7bfc6c),
	.w8(32'h3c11da2f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c404b0e),
	.w1(32'h3c2af026),
	.w2(32'h3c28eb09),
	.w3(32'h3b85c03d),
	.w4(32'h3bc8b729),
	.w5(32'h3b352c36),
	.w6(32'h3c14a3e2),
	.w7(32'h3bb62965),
	.w8(32'h3b5487dd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f18f52),
	.w1(32'h3b25eb7a),
	.w2(32'h3baac5fc),
	.w3(32'hbaf28dc8),
	.w4(32'h3b12eee3),
	.w5(32'h3c156d62),
	.w6(32'hbab1ad79),
	.w7(32'hbb364b21),
	.w8(32'hbb90479b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d302b),
	.w1(32'h3a874e14),
	.w2(32'h3b2f3bcc),
	.w3(32'h3c5a4711),
	.w4(32'h3b14b8cd),
	.w5(32'h3b1e411c),
	.w6(32'h3ae4561f),
	.w7(32'h3b8f0005),
	.w8(32'h3ba8820c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ff9d9),
	.w1(32'h3c17b2e2),
	.w2(32'h3c28580c),
	.w3(32'h3b58b764),
	.w4(32'h3be4ebea),
	.w5(32'h3bb187f0),
	.w6(32'h3b555472),
	.w7(32'h3b90b49e),
	.w8(32'h3c41cf6d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c769c23),
	.w1(32'h3c27eab5),
	.w2(32'h3c812aa4),
	.w3(32'h3c0f56b0),
	.w4(32'h3c0e1aa7),
	.w5(32'h3c43d297),
	.w6(32'h3b65a897),
	.w7(32'h3c68e54a),
	.w8(32'h3c3e4018),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e15f5),
	.w1(32'hbbb2e5a6),
	.w2(32'hbbdd60b8),
	.w3(32'h3c43cb2d),
	.w4(32'hbb4858d9),
	.w5(32'hbbbeed09),
	.w6(32'hbc874b97),
	.w7(32'hbc4a5345),
	.w8(32'hbb4f2e33),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fc46c),
	.w1(32'hbb47663a),
	.w2(32'h3abccece),
	.w3(32'hbbd08f0f),
	.w4(32'h3b9f15aa),
	.w5(32'h3bb6b573),
	.w6(32'h3b73e819),
	.w7(32'h3afb9a22),
	.w8(32'h3bf6cc5c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e7dd5),
	.w1(32'h3bab9823),
	.w2(32'hbb346d58),
	.w3(32'h3bffd0e7),
	.w4(32'h3bf47c5e),
	.w5(32'hb8b9616b),
	.w6(32'hbc09dabe),
	.w7(32'h3aec7cf0),
	.w8(32'h3c552d2a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fda10),
	.w1(32'hbbcf4b6f),
	.w2(32'hbbe89b94),
	.w3(32'hbbde7a6e),
	.w4(32'hbc232df1),
	.w5(32'hbbd6eceb),
	.w6(32'hbb9e6751),
	.w7(32'hbc111ef5),
	.w8(32'hbc3a8e93),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc582c1c),
	.w1(32'h3b94f8d7),
	.w2(32'h3bf9762b),
	.w3(32'hbb43284e),
	.w4(32'h3b6450a6),
	.w5(32'h3b9e4639),
	.w6(32'h3b43a04a),
	.w7(32'h3b80b96c),
	.w8(32'h3b5e559c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbabd54),
	.w1(32'h3b66a5c9),
	.w2(32'h3c0e63b5),
	.w3(32'h3b97d066),
	.w4(32'h3c3eb068),
	.w5(32'h3c60e57a),
	.w6(32'h3ad4daa7),
	.w7(32'h3c07db0f),
	.w8(32'hbb16aec8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1fa24),
	.w1(32'h3bff83c5),
	.w2(32'h3c767ffe),
	.w3(32'h3bb8f870),
	.w4(32'h3b7da052),
	.w5(32'hba0858b4),
	.w6(32'h3a757239),
	.w7(32'h3bce4cb5),
	.w8(32'h3c0917b2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b997736),
	.w1(32'hbcde0d53),
	.w2(32'hbd5edf16),
	.w3(32'h3a531861),
	.w4(32'hbcadffc4),
	.w5(32'hbd0e2d83),
	.w6(32'hbbdd0426),
	.w7(32'hbcb55594),
	.w8(32'hbc640cab),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd08072d),
	.w1(32'h3b7436f7),
	.w2(32'h3ab54b41),
	.w3(32'hbd023e30),
	.w4(32'hb9e60824),
	.w5(32'hbae1811f),
	.w6(32'hb9e8eba2),
	.w7(32'hbadc0009),
	.w8(32'hb89d1fcb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48ad71),
	.w1(32'h3b55c4d8),
	.w2(32'h3c96c0e9),
	.w3(32'hb8283a99),
	.w4(32'h3bd5a624),
	.w5(32'h3c611f21),
	.w6(32'hbb4376aa),
	.w7(32'h3c0a8469),
	.w8(32'h3c172948),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule