module layer_6_featuremap_44(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2bf25),
	.w1(32'h3b9e4225),
	.w2(32'h3b27e2cb),
	.w3(32'h3b9459ea),
	.w4(32'h3bdbc51c),
	.w5(32'h3ac7c043),
	.w6(32'h3b806616),
	.w7(32'h3bd289a0),
	.w8(32'h3b6c3a29),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb63b6d),
	.w1(32'h3b5c10cc),
	.w2(32'hba37d684),
	.w3(32'hbb258c0c),
	.w4(32'hbb4ee58a),
	.w5(32'hbb9ffbe5),
	.w6(32'h3be1d202),
	.w7(32'h3bdd8eaa),
	.w8(32'h3c24ce2b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc499b5d),
	.w1(32'hbcb779b5),
	.w2(32'hbc8c5629),
	.w3(32'hbc1f8b4b),
	.w4(32'hb8bf41c4),
	.w5(32'hbc29b4d5),
	.w6(32'h3a9367e6),
	.w7(32'h3c34eba1),
	.w8(32'h3be3538d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6735d1),
	.w1(32'hbb8065c5),
	.w2(32'hbbd07c20),
	.w3(32'hbb908bf4),
	.w4(32'hbc1009d0),
	.w5(32'hbc454a19),
	.w6(32'hb7c78d4b),
	.w7(32'hbbb991ee),
	.w8(32'hbbaa1f38),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff6149),
	.w1(32'hbd40fe1b),
	.w2(32'hbc9c4db1),
	.w3(32'hbb69f3c4),
	.w4(32'hbc821d23),
	.w5(32'hbc12b886),
	.w6(32'h3d75c60e),
	.w7(32'h3d773c98),
	.w8(32'h3caaae99),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d280dfe),
	.w1(32'hbbaaf12b),
	.w2(32'hbb840fc8),
	.w3(32'hbb89e437),
	.w4(32'hbb6e8461),
	.w5(32'hbb07c1e3),
	.w6(32'hba9a023e),
	.w7(32'hbb712590),
	.w8(32'hbc032969),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad906),
	.w1(32'h3bb496c5),
	.w2(32'h3b895475),
	.w3(32'hbbb54072),
	.w4(32'hba259d99),
	.w5(32'h3b057a84),
	.w6(32'hbc4bfbbf),
	.w7(32'hbbdfc97e),
	.w8(32'h392c2acf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe4e90),
	.w1(32'h3c2d5785),
	.w2(32'h3cfeeaf2),
	.w3(32'hbb08ed22),
	.w4(32'h3b6e617f),
	.w5(32'hbc836f4a),
	.w6(32'h3cf88826),
	.w7(32'h3d1dfe4d),
	.w8(32'h3d0fdd5c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b2a85),
	.w1(32'hbd60c371),
	.w2(32'hbde4d6af),
	.w3(32'h3caeb813),
	.w4(32'h3c5da28c),
	.w5(32'hbc7e6c55),
	.w6(32'hbc359d7d),
	.w7(32'h3d2a2b31),
	.w8(32'h3d2b181b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3d13f4),
	.w1(32'hbb4b598f),
	.w2(32'hbbbc2575),
	.w3(32'h3ba50159),
	.w4(32'h3a946749),
	.w5(32'hbb8e8884),
	.w6(32'h3ace28f3),
	.w7(32'h3b081d87),
	.w8(32'hbb44e09e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1992c8),
	.w1(32'hbb824fd3),
	.w2(32'hbc6c4066),
	.w3(32'hbb115dda),
	.w4(32'h3b242b8d),
	.w5(32'hbc290a4c),
	.w6(32'h3b181f68),
	.w7(32'hbc17061f),
	.w8(32'h3bbc1140),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc110d21),
	.w1(32'hbbf6669c),
	.w2(32'hbc8df5e9),
	.w3(32'hbb1aff5b),
	.w4(32'h3a2fbe07),
	.w5(32'hbba9b74b),
	.w6(32'hbc58f260),
	.w7(32'hbb385724),
	.w8(32'h3badd769),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5d8a0),
	.w1(32'h3a004e41),
	.w2(32'h399e53c1),
	.w3(32'hbb11c386),
	.w4(32'h3b9084a5),
	.w5(32'h3a8151e4),
	.w6(32'hbb13da84),
	.w7(32'h38d59ee3),
	.w8(32'h399858c7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22226d),
	.w1(32'hbd14fd64),
	.w2(32'hbbef4200),
	.w3(32'hbca695fc),
	.w4(32'hbc601201),
	.w5(32'hbb9a9d32),
	.w6(32'hba9aee9e),
	.w7(32'h3c3d1044),
	.w8(32'h3b4549ca),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1420b1),
	.w1(32'hbb1e26d4),
	.w2(32'hbac8037b),
	.w3(32'h3ba2269d),
	.w4(32'hb9b75144),
	.w5(32'hbb3a59fe),
	.w6(32'h3be53099),
	.w7(32'h3bab8154),
	.w8(32'h3ba9838c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd549f4),
	.w1(32'hba5db184),
	.w2(32'h3b28d5e5),
	.w3(32'h3b3854ac),
	.w4(32'h3ba07db4),
	.w5(32'h3ab75188),
	.w6(32'hba4b918c),
	.w7(32'h3b39714e),
	.w8(32'h3b3f46dd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8829d6),
	.w1(32'hbce7a31c),
	.w2(32'hbcac5812),
	.w3(32'hbc083cdd),
	.w4(32'hbc79072d),
	.w5(32'hbbd0546d),
	.w6(32'h3a6aebd6),
	.w7(32'h3c841b69),
	.w8(32'h3c4007cf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba546123),
	.w1(32'h3b97f268),
	.w2(32'h3b1fcc34),
	.w3(32'h3b9fa84a),
	.w4(32'h3ba68573),
	.w5(32'h3a776d83),
	.w6(32'hbbc60648),
	.w7(32'hbb841acd),
	.w8(32'h3a61b829),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bb126),
	.w1(32'h3b1f0d78),
	.w2(32'h3b13bd93),
	.w3(32'h3af244d5),
	.w4(32'h3850037c),
	.w5(32'h3b6c004a),
	.w6(32'hba94ceee),
	.w7(32'hbb8add64),
	.w8(32'hbb133077),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85b252),
	.w1(32'hbb960858),
	.w2(32'hbca68483),
	.w3(32'h3bc65ad0),
	.w4(32'h3baea30c),
	.w5(32'hbaf6e684),
	.w6(32'hbbe0a048),
	.w7(32'h3c696336),
	.w8(32'h3bdfc663),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc982e9c),
	.w1(32'hba9a0a95),
	.w2(32'hb97be7a1),
	.w3(32'hbb0ac09c),
	.w4(32'hbbc52f23),
	.w5(32'hbad3ff6b),
	.w6(32'hba9b2847),
	.w7(32'hbb830253),
	.w8(32'h3a4acc02),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d13b0),
	.w1(32'hbca5ddf4),
	.w2(32'hbc9cac76),
	.w3(32'hbb169988),
	.w4(32'hbb9162b2),
	.w5(32'hbb773e60),
	.w6(32'h3986cc2b),
	.w7(32'hba914111),
	.w8(32'h3c06bbfb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1c08e),
	.w1(32'h3c977bce),
	.w2(32'h3cdadf26),
	.w3(32'hbca20bd9),
	.w4(32'hbc000d42),
	.w5(32'hbc06af2f),
	.w6(32'h3bd7cc07),
	.w7(32'hbbc1827b),
	.w8(32'hbcba3196),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d230bc9),
	.w1(32'h3ca3f8d9),
	.w2(32'hbccb6855),
	.w3(32'hbc945edd),
	.w4(32'h3c89589e),
	.w5(32'h3caaba9c),
	.w6(32'hbd90a931),
	.w7(32'hbd983474),
	.w8(32'hbbd3033f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce371b2),
	.w1(32'hbd3013af),
	.w2(32'hbc4a9361),
	.w3(32'hbc0f7d79),
	.w4(32'hbcc07366),
	.w5(32'hbd19c94f),
	.w6(32'hbc03fa23),
	.w7(32'h3bf23536),
	.w8(32'h3b8e6a9f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbff049),
	.w1(32'hbcef974d),
	.w2(32'hbcfd3161),
	.w3(32'hbc34adc7),
	.w4(32'hbd0bf2d1),
	.w5(32'hbcf37024),
	.w6(32'hbcc229fc),
	.w7(32'hbca9513e),
	.w8(32'hbcb4c2ed),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78bee0),
	.w1(32'h3adbf003),
	.w2(32'hbbd9c6fa),
	.w3(32'h3b110382),
	.w4(32'hb94e4a1d),
	.w5(32'hbad9c96e),
	.w6(32'hbb88214c),
	.w7(32'hbc5a42c9),
	.w8(32'hbbc90d1a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd31af8),
	.w1(32'hbbc8a28a),
	.w2(32'hba997036),
	.w3(32'h3aa42ac7),
	.w4(32'h3bb754f5),
	.w5(32'h3aceddfa),
	.w6(32'hba9eafec),
	.w7(32'h379b1177),
	.w8(32'h3bcb13c0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a6b0d),
	.w1(32'hbb2fb296),
	.w2(32'hbb365b6c),
	.w3(32'hb9beaf23),
	.w4(32'hbb15d214),
	.w5(32'hbb5a3fa4),
	.w6(32'h39e24d71),
	.w7(32'hb9ae6550),
	.w8(32'h3a8fc3a2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfd91e),
	.w1(32'h3cca68cc),
	.w2(32'h3c450a2e),
	.w3(32'hbbbbaddd),
	.w4(32'hbc8a6880),
	.w5(32'hbcc20db1),
	.w6(32'hbc3e7574),
	.w7(32'hbcb34eeb),
	.w8(32'hbc8db588),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb51b33),
	.w1(32'h3b4972e4),
	.w2(32'h3d1c94f6),
	.w3(32'hbcd6b21b),
	.w4(32'hbc6cadae),
	.w5(32'h3c08d353),
	.w6(32'h3c021206),
	.w7(32'hbcb5aa3e),
	.w8(32'hbd053216),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a9d89),
	.w1(32'hbbc57fb8),
	.w2(32'h3c1dc8fa),
	.w3(32'h3c0568d3),
	.w4(32'h3ad01b1c),
	.w5(32'hbb6fa4f7),
	.w6(32'h3b9d622e),
	.w7(32'h3c0b19ed),
	.w8(32'h3b48c0ab),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6a4e1),
	.w1(32'hbbf24a2c),
	.w2(32'hbc393628),
	.w3(32'h3c095224),
	.w4(32'h3bdb214a),
	.w5(32'h3be61b58),
	.w6(32'hbbe5848c),
	.w7(32'hbbc51e6b),
	.w8(32'hbade15d4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce079f3),
	.w1(32'hbcbc21b0),
	.w2(32'hbc89d729),
	.w3(32'hbba620ea),
	.w4(32'hbc83e924),
	.w5(32'hbc1b5ee4),
	.w6(32'hbc88ee8a),
	.w7(32'hba2a3de4),
	.w8(32'hbcae94ca),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb081712),
	.w1(32'hbb355099),
	.w2(32'hbb0598a4),
	.w3(32'hbaab1b96),
	.w4(32'hbb6c5ccc),
	.w5(32'hbb6ccf30),
	.w6(32'h3b94bcc5),
	.w7(32'h3b30e670),
	.w8(32'hb694cefb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0fbed),
	.w1(32'hbbded494),
	.w2(32'hbbc836fb),
	.w3(32'hbc04c789),
	.w4(32'hbcae8c8a),
	.w5(32'hbc7757aa),
	.w6(32'hbc48948e),
	.w7(32'hbcf1668a),
	.w8(32'hbcec53b5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5c273),
	.w1(32'hbb1c18a7),
	.w2(32'h3aab823e),
	.w3(32'h39e70606),
	.w4(32'hb9e96c01),
	.w5(32'h3b2a1175),
	.w6(32'h3b891c8f),
	.w7(32'h3a0fd1cb),
	.w8(32'hbc34cd7d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c69a1),
	.w1(32'hbbd2eeda),
	.w2(32'hbb4212fd),
	.w3(32'hbbfa631f),
	.w4(32'hbc3ef02a),
	.w5(32'hbbc99ca5),
	.w6(32'hbb004e46),
	.w7(32'hbab3e734),
	.w8(32'hba7a5fb8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eba8c),
	.w1(32'hbc97bb0a),
	.w2(32'hbc5e8b67),
	.w3(32'h3c06723b),
	.w4(32'h3c89c97a),
	.w5(32'hbb959617),
	.w6(32'hbbc8b708),
	.w7(32'hbc7b7e19),
	.w8(32'hbc3ed898),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47040f),
	.w1(32'hbdb777de),
	.w2(32'hbdd038a7),
	.w3(32'h3cc3d1db),
	.w4(32'h3c277afc),
	.w5(32'hbb1dfcc7),
	.w6(32'hbc974ec5),
	.w7(32'h3d2d1201),
	.w8(32'h3d22845b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd49480e),
	.w1(32'hbc57114c),
	.w2(32'hbca618c9),
	.w3(32'h3c3090c8),
	.w4(32'hbc383ec7),
	.w5(32'hbcbe088c),
	.w6(32'h3d0d0d8b),
	.w7(32'h3cda684a),
	.w8(32'h3cbcb53f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12327c),
	.w1(32'hbaa2300e),
	.w2(32'h3968a0b0),
	.w3(32'hbb8391ce),
	.w4(32'hbbe4e346),
	.w5(32'hbb737cc9),
	.w6(32'hbb6421f6),
	.w7(32'hbc076e3c),
	.w8(32'hbbb69366),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7b4ca),
	.w1(32'hbbe9331b),
	.w2(32'hbc06620b),
	.w3(32'h3bce5280),
	.w4(32'h3ae6a24a),
	.w5(32'hbbb87cc9),
	.w6(32'hb9ea328c),
	.w7(32'h3ad28ee1),
	.w8(32'hbb5058a7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc204d56),
	.w1(32'hbc3ccf73),
	.w2(32'h3bbd1d0c),
	.w3(32'hbc81c20a),
	.w4(32'hbd518271),
	.w5(32'hbce0cade),
	.w6(32'h3b998cef),
	.w7(32'hbcf5ef32),
	.w8(32'hbd0e9147),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74f58c),
	.w1(32'hbcd864b9),
	.w2(32'hbcd2d29c),
	.w3(32'hbc3f00b2),
	.w4(32'hbbc89cba),
	.w5(32'hbb9e2269),
	.w6(32'hbc52e8b0),
	.w7(32'hbc14d633),
	.w8(32'h3ba14695),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f8d58),
	.w1(32'hbc9067f9),
	.w2(32'hbc434cf6),
	.w3(32'hbc22bf40),
	.w4(32'hbc8ec676),
	.w5(32'hbbc8e4e8),
	.w6(32'hbb473138),
	.w7(32'hbcdf846b),
	.w8(32'hbcb3db20),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc832709),
	.w1(32'h3c4296ad),
	.w2(32'h3c97f661),
	.w3(32'hbbab6552),
	.w4(32'hbb86dd74),
	.w5(32'h3b49fca1),
	.w6(32'hbb9b1aa8),
	.w7(32'hbb837268),
	.w8(32'h3c05e4e6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1371da),
	.w1(32'h3b7ad696),
	.w2(32'h3bb7cf28),
	.w3(32'hbaa8d646),
	.w4(32'h39d09651),
	.w5(32'h3c41220a),
	.w6(32'hbadd3503),
	.w7(32'hbbd2b11d),
	.w8(32'h3b8c0fb7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff7beb),
	.w1(32'h3b5b7634),
	.w2(32'h3ac3e480),
	.w3(32'hbadb9737),
	.w4(32'h3acfe381),
	.w5(32'h3bc03256),
	.w6(32'hbaffba67),
	.w7(32'h37e28749),
	.w8(32'h3b72ecf5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d3431),
	.w1(32'h3c954a08),
	.w2(32'h3d6cbef9),
	.w3(32'hbcc7a6d6),
	.w4(32'hbc4f5a6d),
	.w5(32'hbb4e290b),
	.w6(32'h3c2399f0),
	.w7(32'hbcbb141a),
	.w8(32'hbd4b6ee1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e2922),
	.w1(32'hbb3188f0),
	.w2(32'hbb6e8fa3),
	.w3(32'hbc14c958),
	.w4(32'hbc4d6a39),
	.w5(32'hbc348a0e),
	.w6(32'hbaca5848),
	.w7(32'hbbad7a8c),
	.w8(32'hbb582f09),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad144ed),
	.w1(32'hbb44a16f),
	.w2(32'hbc351fab),
	.w3(32'hbb6d4409),
	.w4(32'hbc4ad287),
	.w5(32'hbc842283),
	.w6(32'hb8a515f4),
	.w7(32'hbb5eec6c),
	.w8(32'hbc1d8ecf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc94dde),
	.w1(32'hbc09d296),
	.w2(32'hba5a0ab8),
	.w3(32'hbbcd7db6),
	.w4(32'h3b822724),
	.w5(32'h3c829a50),
	.w6(32'hbb82dc0f),
	.w7(32'h3be8c579),
	.w8(32'h3d00abd3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25728d),
	.w1(32'h3c8361f6),
	.w2(32'h3c854393),
	.w3(32'h3a15f5dc),
	.w4(32'h3c4a410d),
	.w5(32'h3c0b4e5b),
	.w6(32'h3c371b2e),
	.w7(32'h3cc004b5),
	.w8(32'h3cd7093f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc205e1),
	.w1(32'h3b9f3459),
	.w2(32'h3b256e00),
	.w3(32'hb91bff5c),
	.w4(32'hba340a7f),
	.w5(32'h3a908ab3),
	.w6(32'hbbb7c3d3),
	.w7(32'hbbd31f86),
	.w8(32'h3adcc8ca),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7af196),
	.w1(32'hbc504b7f),
	.w2(32'hbbd0f004),
	.w3(32'hbc126e72),
	.w4(32'hbcb0acd0),
	.w5(32'hbc867664),
	.w6(32'hb9ee445c),
	.w7(32'hbb577b00),
	.w8(32'hbbe7e481),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c313fbd),
	.w1(32'hbd279f4e),
	.w2(32'hbda0505c),
	.w3(32'hbcc49b5f),
	.w4(32'hbd7768e1),
	.w5(32'hbd4376fc),
	.w6(32'hbd6a2e43),
	.w7(32'hbdc7c49d),
	.w8(32'hbda36f45),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd978f52),
	.w1(32'hbbb12105),
	.w2(32'hbb918d62),
	.w3(32'hba4ea46b),
	.w4(32'h3ae85a9d),
	.w5(32'h399125fb),
	.w6(32'hbb13f455),
	.w7(32'hbb5d337b),
	.w8(32'h38cbd63b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd61dc3),
	.w1(32'h3bd7c408),
	.w2(32'h3c34f526),
	.w3(32'h3bed4b86),
	.w4(32'h3c23ad81),
	.w5(32'h3c1f29ac),
	.w6(32'h3c162f38),
	.w7(32'h3c666583),
	.w8(32'h3c6548a3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19d9bf),
	.w1(32'hbd32e21b),
	.w2(32'hbd53bd9b),
	.w3(32'hbba0f300),
	.w4(32'hbc764499),
	.w5(32'hbd015b18),
	.w6(32'hbc643c44),
	.w7(32'hbc200e24),
	.w8(32'hbc888cf9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22bc1b),
	.w1(32'hbbfd62e5),
	.w2(32'hbbaf2212),
	.w3(32'hbb5aa71a),
	.w4(32'hbc181bd3),
	.w5(32'hbbc9e809),
	.w6(32'hbc2d1a13),
	.w7(32'hbc49e111),
	.w8(32'hbc032e25),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad97dc7),
	.w1(32'hbc1957a3),
	.w2(32'hbc8988db),
	.w3(32'hbb06750d),
	.w4(32'hbcacf8f5),
	.w5(32'hbca1b0fb),
	.w6(32'h3b04cb87),
	.w7(32'hbc47cf41),
	.w8(32'hbc621926),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ed803),
	.w1(32'h3d072dbb),
	.w2(32'hbc06ef0e),
	.w3(32'h3c9fc179),
	.w4(32'h3b930294),
	.w5(32'hbb6067fe),
	.w6(32'hba28da04),
	.w7(32'hbd89bd7e),
	.w8(32'hbd36f543),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba18db2),
	.w1(32'hbcfae6bd),
	.w2(32'hbd430d6e),
	.w3(32'hbcb2d34c),
	.w4(32'hbd13d366),
	.w5(32'hbcda9fb2),
	.w6(32'hbd2dc26c),
	.w7(32'hbd84ab88),
	.w8(32'hbd4468c9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule