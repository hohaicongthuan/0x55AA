module layer_10_featuremap_229(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e7c62),
	.w1(32'hbb2f0069),
	.w2(32'hba4545dd),
	.w3(32'h3a3a7bad),
	.w4(32'hbbb5a5f1),
	.w5(32'hbaae6ede),
	.w6(32'hbb5771c6),
	.w7(32'hbb1ff18d),
	.w8(32'hbbac44c9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1359fc),
	.w1(32'hbbddc05e),
	.w2(32'hbb12238d),
	.w3(32'hbc069b3c),
	.w4(32'h3bf5ed9a),
	.w5(32'h3ab30017),
	.w6(32'h3b8a626e),
	.w7(32'hb98add38),
	.w8(32'hbb55973a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4e0e3),
	.w1(32'hbb9eb3cb),
	.w2(32'hbb862bf6),
	.w3(32'h3b5c8192),
	.w4(32'h3c278b0e),
	.w5(32'hbafedbd6),
	.w6(32'hbcc350fb),
	.w7(32'h39abf4c6),
	.w8(32'h38f5aa5f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8256fb),
	.w1(32'hbc77ed23),
	.w2(32'hbb60f6b1),
	.w3(32'hbc1e73df),
	.w4(32'hba819cc1),
	.w5(32'hbb8afbd6),
	.w6(32'hba22fae6),
	.w7(32'h3aea755d),
	.w8(32'h3c575ec7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c216e),
	.w1(32'h3a1acbd2),
	.w2(32'h395f54e8),
	.w3(32'hbb0badfa),
	.w4(32'hbb8ed7f6),
	.w5(32'hba0c48ab),
	.w6(32'hbb5e402b),
	.w7(32'h3c1509d1),
	.w8(32'h3cef8369),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e1377),
	.w1(32'h3a96cca6),
	.w2(32'h3bc5c573),
	.w3(32'hbad318d5),
	.w4(32'h3b02d395),
	.w5(32'hbb911cb2),
	.w6(32'h3b75e011),
	.w7(32'hba8572a2),
	.w8(32'h3bb8880a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bbbeb),
	.w1(32'h38711dce),
	.w2(32'h3b295c57),
	.w3(32'h3b390b8a),
	.w4(32'hbd03551a),
	.w5(32'h3bca0030),
	.w6(32'h3b3fc1bf),
	.w7(32'h3b7bae11),
	.w8(32'hba2bdf4c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb53d59),
	.w1(32'hbc581d63),
	.w2(32'h3c05fb10),
	.w3(32'h3b821014),
	.w4(32'h3b844abb),
	.w5(32'hbbaad3ca),
	.w6(32'hbbabe2ed),
	.w7(32'hbbe602aa),
	.w8(32'h3b1f4ada),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4940c1),
	.w1(32'hbc547cd5),
	.w2(32'h3aeb0b68),
	.w3(32'h3af44051),
	.w4(32'hbb857ba2),
	.w5(32'h3b67e486),
	.w6(32'hbb45983c),
	.w7(32'hbbc39e5a),
	.w8(32'h3a9a8744),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5fc143),
	.w1(32'hba06dc92),
	.w2(32'hbbef6ac7),
	.w3(32'h3c0d8a45),
	.w4(32'h3b60befb),
	.w5(32'h3a34c5f8),
	.w6(32'hbc9b0efc),
	.w7(32'hbc4888d3),
	.w8(32'hbc7e48d7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd5856),
	.w1(32'hbb684c1e),
	.w2(32'h3b693e73),
	.w3(32'hbb473e83),
	.w4(32'hbbfd076b),
	.w5(32'h39709506),
	.w6(32'h3bb82bb0),
	.w7(32'hbb11789b),
	.w8(32'h39b51a4d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967549),
	.w1(32'hbbc93348),
	.w2(32'h3bac1cc4),
	.w3(32'hbadd6ad5),
	.w4(32'hbac8f25d),
	.w5(32'hba2ddf6b),
	.w6(32'hba22d766),
	.w7(32'hb8c9df56),
	.w8(32'hbbc99c3f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16db9e),
	.w1(32'hbbb73a31),
	.w2(32'hba902add),
	.w3(32'hbb513696),
	.w4(32'hbb92298e),
	.w5(32'hbbdf7d3c),
	.w6(32'h3b7e8ef3),
	.w7(32'hbbc3f6f9),
	.w8(32'h3c0cdda1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b7abd),
	.w1(32'hbbc90cb2),
	.w2(32'h3c192a36),
	.w3(32'hbb2aa10c),
	.w4(32'hbc30041c),
	.w5(32'hbba97383),
	.w6(32'hbc4b84c1),
	.w7(32'hbb128103),
	.w8(32'hb990a465),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc23c11),
	.w1(32'h3ba08080),
	.w2(32'h3b69bf5a),
	.w3(32'hbbbf7036),
	.w4(32'hbc2d54e6),
	.w5(32'hbb036a41),
	.w6(32'hbaeee489),
	.w7(32'h3aa6c435),
	.w8(32'h3b775f1a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc093914),
	.w1(32'hbb3bfc8d),
	.w2(32'h3b62cf0f),
	.w3(32'hbbde681f),
	.w4(32'hba4d3380),
	.w5(32'hba4b1007),
	.w6(32'hbbb3f539),
	.w7(32'h3aa92ef0),
	.w8(32'hbcd60e17),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f157),
	.w1(32'hba9e726f),
	.w2(32'hbc0a4178),
	.w3(32'hbb98dba3),
	.w4(32'hb95263a3),
	.w5(32'hbc0520d8),
	.w6(32'hbb15d6eb),
	.w7(32'hbc144f46),
	.w8(32'h3a8d2524),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01a798),
	.w1(32'hbc46f9bb),
	.w2(32'hbb9d5eb5),
	.w3(32'h3912c5a9),
	.w4(32'hbb7fe743),
	.w5(32'hb8abc94b),
	.w6(32'hbbee56ae),
	.w7(32'h3d4b7aa5),
	.w8(32'h3afe562c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d5cd2),
	.w1(32'h3c0acf30),
	.w2(32'hbb29533e),
	.w3(32'hbc04a373),
	.w4(32'h3b24459c),
	.w5(32'hbc12007b),
	.w6(32'hbb66a486),
	.w7(32'hba8e7fe9),
	.w8(32'hbb62bc19),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba983cf),
	.w1(32'h3b580c7e),
	.w2(32'hbc026114),
	.w3(32'h3b653d11),
	.w4(32'hbd4ef6d5),
	.w5(32'h3b1bd2d5),
	.w6(32'h3a9792a3),
	.w7(32'h3ac5c457),
	.w8(32'hbb215028),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92425b),
	.w1(32'hbb68c1ad),
	.w2(32'hbd544748),
	.w3(32'hbb5f9606),
	.w4(32'h3b642f65),
	.w5(32'h3ad193d7),
	.w6(32'h3bef228c),
	.w7(32'hbb68988f),
	.w8(32'hbc25ed87),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b01d6),
	.w1(32'h3aab71e1),
	.w2(32'h3996130b),
	.w3(32'h38e526c5),
	.w4(32'hbb8e42f0),
	.w5(32'hbb81d8da),
	.w6(32'h3ccfb14e),
	.w7(32'hb993a523),
	.w8(32'hbb3caad5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba362a7),
	.w1(32'h38abbf6b),
	.w2(32'h3c63cd31),
	.w3(32'h39b89862),
	.w4(32'h3ad1ea45),
	.w5(32'h3c03b75f),
	.w6(32'h38f0955b),
	.w7(32'hbb93f82e),
	.w8(32'hbc20c9f9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a244d),
	.w1(32'hbc1ecda7),
	.w2(32'h3b968b13),
	.w3(32'h3b2428e7),
	.w4(32'h3aa35458),
	.w5(32'h3a220a46),
	.w6(32'h3b77b05c),
	.w7(32'hbc5e5e1a),
	.w8(32'hbb9dccc6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b7ff5),
	.w1(32'hbb000f3d),
	.w2(32'h3b82b5d8),
	.w3(32'hba967f57),
	.w4(32'h3a1dd69a),
	.w5(32'hbc1a68a3),
	.w6(32'h3bca0000),
	.w7(32'hbbd36914),
	.w8(32'hbcb47b23),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc136285),
	.w1(32'hb78f9a4d),
	.w2(32'h3b282062),
	.w3(32'hbbbe84ca),
	.w4(32'hb8ee782b),
	.w5(32'hbc0a3633),
	.w6(32'hbbcac928),
	.w7(32'hbaebf05c),
	.w8(32'hbaa7aa8e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd0c0),
	.w1(32'hbc300ba7),
	.w2(32'h3abfbcb9),
	.w3(32'hbadcc223),
	.w4(32'hbbd57eb1),
	.w5(32'hbb2a6676),
	.w6(32'hbb4f8926),
	.w7(32'hba82510f),
	.w8(32'h3b134c7a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba87c06),
	.w1(32'h3b3d58b4),
	.w2(32'h3a084450),
	.w3(32'h3aa42adc),
	.w4(32'h3bc342d0),
	.w5(32'hbb046737),
	.w6(32'hbb74c0dd),
	.w7(32'h3c11358c),
	.w8(32'h3bf8b9d9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77c86f),
	.w1(32'h3b5f7abf),
	.w2(32'h3a99b2f9),
	.w3(32'h3c19b9e8),
	.w4(32'hb863d063),
	.w5(32'h3c1d14de),
	.w6(32'hbbfb7945),
	.w7(32'hbb16cf9d),
	.w8(32'h3c399447),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6365b3),
	.w1(32'h3b87fa12),
	.w2(32'hbb9338c8),
	.w3(32'hbbc1256c),
	.w4(32'h3c0ced9c),
	.w5(32'h3bbc2710),
	.w6(32'h3ccd5220),
	.w7(32'hba48ec45),
	.w8(32'h39d6477e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a3ddf),
	.w1(32'hbb416fde),
	.w2(32'h3b7491c5),
	.w3(32'hbbfa0ec6),
	.w4(32'hbaebb869),
	.w5(32'h3b76c6f2),
	.w6(32'h3bb1d5ba),
	.w7(32'h3b91d225),
	.w8(32'hbc496824),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafea3a1),
	.w1(32'h39c6845c),
	.w2(32'hbbf0ed7a),
	.w3(32'hbc2ecbc4),
	.w4(32'hbb835293),
	.w5(32'hbb89c3e9),
	.w6(32'h3c264323),
	.w7(32'h3bd95ec4),
	.w8(32'h3b739988),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83a935),
	.w1(32'h3b613f71),
	.w2(32'h3bb58283),
	.w3(32'h3c0371ad),
	.w4(32'hba8947fb),
	.w5(32'h3bdc73bf),
	.w6(32'hbadd0877),
	.w7(32'h3a4d4966),
	.w8(32'hbbc8311e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912149),
	.w1(32'h3b433d8a),
	.w2(32'hbb6bb87e),
	.w3(32'hba0a364f),
	.w4(32'hbafa73cc),
	.w5(32'hba99c3bf),
	.w6(32'h3b633ce7),
	.w7(32'h3b59461e),
	.w8(32'h3b814463),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52eb15),
	.w1(32'hbb33e422),
	.w2(32'h3b6836f1),
	.w3(32'h3c2ded40),
	.w4(32'hba918866),
	.w5(32'hbb8b2fce),
	.w6(32'h3b71d218),
	.w7(32'h3c6646a6),
	.w8(32'hbc0fa805),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5db37),
	.w1(32'hbafe5147),
	.w2(32'hbba0cec9),
	.w3(32'hbc3ddf3a),
	.w4(32'h3c784d6a),
	.w5(32'h3c878452),
	.w6(32'hba289cfb),
	.w7(32'h3b6a23f2),
	.w8(32'h3b052938),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54e867),
	.w1(32'h3be09dda),
	.w2(32'h3b92ae1c),
	.w3(32'hbc1cce28),
	.w4(32'hbbf08621),
	.w5(32'hbc2b2c23),
	.w6(32'h3b1466d5),
	.w7(32'h3cbafcd2),
	.w8(32'hbb759ff2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b521e6f),
	.w1(32'h3aa29bef),
	.w2(32'h3b0f5486),
	.w3(32'hb9c9d0e9),
	.w4(32'h3be11367),
	.w5(32'hb94b79cc),
	.w6(32'hbbbdccaf),
	.w7(32'h3b99b415),
	.w8(32'hbaf3c308),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17b182),
	.w1(32'h3cf9f20b),
	.w2(32'hb8b8c3d1),
	.w3(32'hbc9bfc8a),
	.w4(32'h3ccb5e6a),
	.w5(32'h3a140f07),
	.w6(32'h3a27e7c3),
	.w7(32'h3cc55ac6),
	.w8(32'hbc04de79),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38baa7ad),
	.w1(32'hbb9258f8),
	.w2(32'h3b8b91a2),
	.w3(32'hbb6c3e04),
	.w4(32'h3bd72b80),
	.w5(32'hbb839ef6),
	.w6(32'h3be063d6),
	.w7(32'h3ca5369a),
	.w8(32'h3b09c51f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902c2f6),
	.w1(32'h3bd48af9),
	.w2(32'h3b451b95),
	.w3(32'h3ae7201d),
	.w4(32'hbb2f4e50),
	.w5(32'hbb299f56),
	.w6(32'h38a680ec),
	.w7(32'h3b46b09f),
	.w8(32'hba7c4ec4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babfad5),
	.w1(32'h3b901b1d),
	.w2(32'h3bf12fce),
	.w3(32'h3b716256),
	.w4(32'hbc8aeb69),
	.w5(32'h3bdc574a),
	.w6(32'h3c0c5688),
	.w7(32'hbb0e48fa),
	.w8(32'h3b741149),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89d07d),
	.w1(32'h3c12751e),
	.w2(32'hbb2c17f7),
	.w3(32'hbbc382c9),
	.w4(32'h3b12eb4e),
	.w5(32'hbbd612d4),
	.w6(32'h3c2b2eaa),
	.w7(32'hbb94d83c),
	.w8(32'h3a8a2178),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf446f),
	.w1(32'h3b006cc0),
	.w2(32'hbb870206),
	.w3(32'h3ba46320),
	.w4(32'h3b6d55a5),
	.w5(32'hbb108d14),
	.w6(32'h3bb2b8bc),
	.w7(32'h3af3c25d),
	.w8(32'h3b0951e7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a09c1),
	.w1(32'hbc3b41d3),
	.w2(32'h3bd9a391),
	.w3(32'hbbe68179),
	.w4(32'h3b6015aa),
	.w5(32'hbbd24005),
	.w6(32'hba788709),
	.w7(32'hbb55549f),
	.w8(32'h397d4378),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82c5a6),
	.w1(32'h3acc3447),
	.w2(32'h3b9f30d7),
	.w3(32'h3c4c40aa),
	.w4(32'hbaaa496d),
	.w5(32'h3b7ce819),
	.w6(32'hbbc4c894),
	.w7(32'h351f3432),
	.w8(32'hbb2b3966),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae89f87),
	.w1(32'h3b3e4f3b),
	.w2(32'h3b06818e),
	.w3(32'h3ad24080),
	.w4(32'h3bb89404),
	.w5(32'h3bf36dd8),
	.w6(32'h39e1d7b5),
	.w7(32'hbaa8827a),
	.w8(32'h3bbf8ea7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27cc4b),
	.w1(32'h3bc61451),
	.w2(32'hbb7b9d88),
	.w3(32'hbb99b673),
	.w4(32'h3b50b235),
	.w5(32'h3bd52d30),
	.w6(32'h3c18af27),
	.w7(32'h3b1f4769),
	.w8(32'h3b088f9e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aade324),
	.w1(32'hb8b5e721),
	.w2(32'hbbdae422),
	.w3(32'h3bcbd094),
	.w4(32'h3c3bc46c),
	.w5(32'hbab936b0),
	.w6(32'h39bc97b1),
	.w7(32'hbbc22991),
	.w8(32'hbb34f334),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eb2e0),
	.w1(32'hbac9ab19),
	.w2(32'hbb4d8954),
	.w3(32'h3b4f1c19),
	.w4(32'hbc1b76c4),
	.w5(32'h3c09563c),
	.w6(32'hbbbf808b),
	.w7(32'hbb051578),
	.w8(32'h3c2366fb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f3d5bd),
	.w1(32'h3ba0c059),
	.w2(32'h3a8da60d),
	.w3(32'hbba33368),
	.w4(32'h3a2957c6),
	.w5(32'hb9dde201),
	.w6(32'h38dd1ae3),
	.w7(32'h39ce092f),
	.w8(32'h3a6a46c8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4aa0f),
	.w1(32'h3bc4d583),
	.w2(32'hbc3fd263),
	.w3(32'h3baeacc0),
	.w4(32'hbb312ff9),
	.w5(32'h3be01fdf),
	.w6(32'hbbf43b58),
	.w7(32'hba47a3f7),
	.w8(32'hbb6de2a3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba853ff9),
	.w1(32'h3b003400),
	.w2(32'hbc266edb),
	.w3(32'hbbdc6d69),
	.w4(32'h3a0f8a0b),
	.w5(32'h3c2cce07),
	.w6(32'hbc128865),
	.w7(32'h3c0204d4),
	.w8(32'hbabf24ad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ff035),
	.w1(32'hbc508966),
	.w2(32'h3b5b493d),
	.w3(32'hb522b48a),
	.w4(32'hbc672097),
	.w5(32'h3c237277),
	.w6(32'h3acc60e8),
	.w7(32'hbb2faa29),
	.w8(32'hbc40c55c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1852a9),
	.w1(32'h3bd5bc48),
	.w2(32'h3c861f7d),
	.w3(32'h3caca961),
	.w4(32'h3badd582),
	.w5(32'hbc46577e),
	.w6(32'h3c86ad4e),
	.w7(32'h3b09367a),
	.w8(32'h3af9a112),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23cfe7),
	.w1(32'hbb6c4161),
	.w2(32'hbbaadd16),
	.w3(32'hbca914e3),
	.w4(32'hbc9f306f),
	.w5(32'hbb5aa671),
	.w6(32'h3a726dcb),
	.w7(32'h388d5d7d),
	.w8(32'h3c0924de),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe23268),
	.w1(32'hb97709e4),
	.w2(32'h3b7c9a32),
	.w3(32'h3c9660af),
	.w4(32'hbc2cecbd),
	.w5(32'hba315d33),
	.w6(32'hbb5f6db7),
	.w7(32'hbb1c686f),
	.w8(32'hbac5aa0d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad693cb),
	.w1(32'hb8ae2c4a),
	.w2(32'hbca439c0),
	.w3(32'h3a24676e),
	.w4(32'h3b80801b),
	.w5(32'hbc47190f),
	.w6(32'hbc789372),
	.w7(32'hbc30e33c),
	.w8(32'hbb916b53),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79a5eb),
	.w1(32'h3d31d350),
	.w2(32'hbbe91321),
	.w3(32'hbbe388ad),
	.w4(32'hbc30d4ed),
	.w5(32'h3bf104b5),
	.w6(32'h396cab0a),
	.w7(32'hba00b498),
	.w8(32'h3a46de36),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12c0cf),
	.w1(32'hba28caa1),
	.w2(32'hbca275d6),
	.w3(32'h3a0a472e),
	.w4(32'hbb15a693),
	.w5(32'h3af87415),
	.w6(32'hbbc40c38),
	.w7(32'hbb1f41b8),
	.w8(32'h3a58bb38),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8425c),
	.w1(32'h3b1b86e6),
	.w2(32'hbc4c212d),
	.w3(32'h3b963e5a),
	.w4(32'hbb31466b),
	.w5(32'hbcbb4fc5),
	.w6(32'h3c8ad4ce),
	.w7(32'hbb1fe257),
	.w8(32'h3b2ca9c4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44bb75),
	.w1(32'hbbaeccec),
	.w2(32'hba564d64),
	.w3(32'h3b7c5d47),
	.w4(32'hbc32d724),
	.w5(32'h39cc6884),
	.w6(32'h3bf2fc86),
	.w7(32'h3a55b245),
	.w8(32'hbc3960a4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08a570),
	.w1(32'h3a130f60),
	.w2(32'hbc7a2b6b),
	.w3(32'hbb7fdf25),
	.w4(32'h3b23c531),
	.w5(32'h3a9283e7),
	.w6(32'hbb06d13b),
	.w7(32'h3bf30947),
	.w8(32'hbb8a8e3b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9f042),
	.w1(32'h3bbc0c84),
	.w2(32'h3c05ea38),
	.w3(32'h3bc22700),
	.w4(32'h3c59b7ee),
	.w5(32'hbbc9fc95),
	.w6(32'h3bf1de1d),
	.w7(32'h3c28b4d8),
	.w8(32'h37fab8f6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5a000),
	.w1(32'hbb967f43),
	.w2(32'hbb4b5813),
	.w3(32'h3c23afcf),
	.w4(32'hbc01f9e8),
	.w5(32'hbbfa33ec),
	.w6(32'hbb8d9a4c),
	.w7(32'h38d4514d),
	.w8(32'h39bf4e73),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca033a4),
	.w1(32'hbbc78e4d),
	.w2(32'h3b485c90),
	.w3(32'hbbf4b66b),
	.w4(32'h3b5bbb90),
	.w5(32'h391500e3),
	.w6(32'hba155a27),
	.w7(32'hbc44a10a),
	.w8(32'h3bd88b96),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04fe86),
	.w1(32'hbbe3a1d8),
	.w2(32'hbc1e399f),
	.w3(32'h3beaef5d),
	.w4(32'h3bdcb575),
	.w5(32'hbc4282a6),
	.w6(32'h3a023829),
	.w7(32'h3a4f0f41),
	.w8(32'h3c571da1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf05c6),
	.w1(32'hbbb5e7c7),
	.w2(32'hbb595864),
	.w3(32'h3bfdcf19),
	.w4(32'h3b782ad8),
	.w5(32'h3c0578f7),
	.w6(32'h3b19fb71),
	.w7(32'hbb04b38f),
	.w8(32'h39c48011),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05f983),
	.w1(32'hbc81ff2f),
	.w2(32'hb9a7737c),
	.w3(32'hbc749f59),
	.w4(32'hb9263b4c),
	.w5(32'hbc6396ee),
	.w6(32'hb92ffc1b),
	.w7(32'h3ab01a11),
	.w8(32'hbb112f23),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15df09),
	.w1(32'h3b391270),
	.w2(32'hbc012713),
	.w3(32'h3acbb9cc),
	.w4(32'hbc8957ea),
	.w5(32'h3aa5c384),
	.w6(32'hbb921e94),
	.w7(32'hbc1dc70d),
	.w8(32'hbc20b3b5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba939e0e),
	.w1(32'hbaca4ffc),
	.w2(32'h3b121ff2),
	.w3(32'h3b1ceb20),
	.w4(32'hbba01e8a),
	.w5(32'hbb9c58f9),
	.w6(32'h39d1e1d7),
	.w7(32'h3aa17228),
	.w8(32'h3c41bd5f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbb4c1),
	.w1(32'h3ba53d30),
	.w2(32'h3c87efa1),
	.w3(32'h3c6d5106),
	.w4(32'h3d516e81),
	.w5(32'hb9141792),
	.w6(32'hbcb59dcf),
	.w7(32'hbb87ee26),
	.w8(32'h3b5127e1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66df51),
	.w1(32'hbb17d59f),
	.w2(32'hbb786297),
	.w3(32'h3ba84561),
	.w4(32'hbb844694),
	.w5(32'hbc34aef8),
	.w6(32'hbaf50f74),
	.w7(32'h3c701942),
	.w8(32'h3c051c38),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a8eba),
	.w1(32'hb8b97959),
	.w2(32'hbb921dae),
	.w3(32'hbbb6d7e8),
	.w4(32'h3b440ff3),
	.w5(32'h3adf99ff),
	.w6(32'h38b98d15),
	.w7(32'hbc455c2c),
	.w8(32'hbc06aac1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3d762),
	.w1(32'h39f31212),
	.w2(32'h39736ffe),
	.w3(32'hbb5866e1),
	.w4(32'hbb35f7dd),
	.w5(32'h3b92db59),
	.w6(32'hbbe61718),
	.w7(32'hbc0fbdbf),
	.w8(32'hbbd15df7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1ff0e),
	.w1(32'h39d15279),
	.w2(32'h3bd63fbf),
	.w3(32'h3c580e9b),
	.w4(32'hbc38a539),
	.w5(32'hbc95c59d),
	.w6(32'hbaa0a49f),
	.w7(32'h3b4633fb),
	.w8(32'h3a92f0e7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3ac3d),
	.w1(32'hbb33fa66),
	.w2(32'h39f5afdb),
	.w3(32'h3c20991c),
	.w4(32'h3cb46561),
	.w5(32'hbaf650be),
	.w6(32'hbc391fc8),
	.w7(32'h3a093ba8),
	.w8(32'hba9c1d27),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073336),
	.w1(32'hbbe08b4c),
	.w2(32'h3beea4b0),
	.w3(32'h3aae3566),
	.w4(32'hbbeda0af),
	.w5(32'hbb7c4f8d),
	.w6(32'hbbd01195),
	.w7(32'h3aec4a13),
	.w8(32'h3ad4d1c1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f3c1c),
	.w1(32'hb60225ec),
	.w2(32'hbac86190),
	.w3(32'h3b0a11f4),
	.w4(32'h38ce09e3),
	.w5(32'hbb8d8f3b),
	.w6(32'h3b8cf65f),
	.w7(32'hbc21de48),
	.w8(32'hba083e57),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b0e6a),
	.w1(32'h3ab1daae),
	.w2(32'hba8d1314),
	.w3(32'hbaf94922),
	.w4(32'h38100d0a),
	.w5(32'hbb96005e),
	.w6(32'h3a2ea216),
	.w7(32'hbc1bb6b1),
	.w8(32'h3a1fdd42),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c503e3f),
	.w1(32'h3bce851e),
	.w2(32'hbc393116),
	.w3(32'h3c324fc8),
	.w4(32'h3babf5dc),
	.w5(32'hbb354de6),
	.w6(32'hbc79cef7),
	.w7(32'h3b1adc27),
	.w8(32'h3c23a459),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbabcc5),
	.w1(32'h3a2563a8),
	.w2(32'h3a247c3a),
	.w3(32'hbbfc62cd),
	.w4(32'hbb640c28),
	.w5(32'h3b7570ac),
	.w6(32'hbb5ea43e),
	.w7(32'hbb0c8ecd),
	.w8(32'hbc8aebc9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc002fca),
	.w1(32'hba1bc920),
	.w2(32'hbc637f57),
	.w3(32'hbae68943),
	.w4(32'hbb380d1b),
	.w5(32'hbc1d9bba),
	.w6(32'h3af78cf9),
	.w7(32'hbbeb96e0),
	.w8(32'h3bac5fd5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a595),
	.w1(32'hbb0fe929),
	.w2(32'hbb519554),
	.w3(32'h3c215544),
	.w4(32'hbb8518c3),
	.w5(32'h3cbad155),
	.w6(32'hbb8708eb),
	.w7(32'h3b97577d),
	.w8(32'h3c20fd27),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3832b1),
	.w1(32'h3bf3f1b1),
	.w2(32'hbbed5bdd),
	.w3(32'h3bfc6c22),
	.w4(32'hbc28a525),
	.w5(32'hba1f48d0),
	.w6(32'h3b9658f7),
	.w7(32'h3b323710),
	.w8(32'h3cccaf31),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad14ceb),
	.w1(32'h3c3bb763),
	.w2(32'hbc564451),
	.w3(32'h3cb25bad),
	.w4(32'h3c2aeef4),
	.w5(32'hbc751470),
	.w6(32'hbc8bc69f),
	.w7(32'h3b244aa2),
	.w8(32'h3bee6273),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42183c),
	.w1(32'h3bacf9ea),
	.w2(32'hbc70753d),
	.w3(32'hbc8bcaa8),
	.w4(32'hbbb9885c),
	.w5(32'h3ccd9eed),
	.w6(32'h3c36226c),
	.w7(32'hbc547476),
	.w8(32'hbc93ff9e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990df4e),
	.w1(32'hbbdcfd10),
	.w2(32'h3ca200c0),
	.w3(32'hbb1df2f8),
	.w4(32'hbb8b0f11),
	.w5(32'h3ba3a118),
	.w6(32'h3ca49e1e),
	.w7(32'h3b4cf8d5),
	.w8(32'h3c199efc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e2b72),
	.w1(32'h3945008f),
	.w2(32'h3be235ab),
	.w3(32'h3b3a2752),
	.w4(32'h3c6e6129),
	.w5(32'h3bc319df),
	.w6(32'h3c4a1689),
	.w7(32'hbbc3b88a),
	.w8(32'hbbd99263),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba96dba),
	.w1(32'hbc827fc9),
	.w2(32'h3befbd12),
	.w3(32'h3c25da02),
	.w4(32'h3b54dea2),
	.w5(32'h3c0056b0),
	.w6(32'h3cf781e0),
	.w7(32'h3b8e134e),
	.w8(32'h3c3aa381),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1110bf),
	.w1(32'h3b7d524e),
	.w2(32'hbc306a70),
	.w3(32'hbacbde34),
	.w4(32'h3c849c98),
	.w5(32'hbb5e683c),
	.w6(32'h3ac05a04),
	.w7(32'hbb8fa082),
	.w8(32'h3c769b68),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77a651),
	.w1(32'h3a2af1e3),
	.w2(32'hbd242b76),
	.w3(32'hbb4deb00),
	.w4(32'hbb7d0b8e),
	.w5(32'h3b6b995a),
	.w6(32'h3c0603f1),
	.w7(32'hbc30536c),
	.w8(32'hbc47f48e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9421be),
	.w1(32'hbbe5c5a5),
	.w2(32'h3b2ae8d2),
	.w3(32'hbbc44099),
	.w4(32'h3c4795df),
	.w5(32'h3acf3b9d),
	.w6(32'h3bc48712),
	.w7(32'h3b87b5ef),
	.w8(32'hbcba9522),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12ea61),
	.w1(32'h3c09107c),
	.w2(32'hbb9b9801),
	.w3(32'hbbac4315),
	.w4(32'h3b0d3856),
	.w5(32'hbc980942),
	.w6(32'hbbec3bfc),
	.w7(32'hbcc48b6d),
	.w8(32'h3cac5f16),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb406ad4),
	.w1(32'hbbeec6a3),
	.w2(32'h39bf8e48),
	.w3(32'h3c83c81e),
	.w4(32'h3b0f90fe),
	.w5(32'h3b298a67),
	.w6(32'hbb52befe),
	.w7(32'h3bd317da),
	.w8(32'h3c83bc86),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb74f72),
	.w1(32'hbca4edfb),
	.w2(32'hbc34741b),
	.w3(32'h3c3c69ab),
	.w4(32'hbab48a39),
	.w5(32'hbb76617c),
	.w6(32'h3c80631c),
	.w7(32'hbb84800c),
	.w8(32'h3c820271),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4727a2),
	.w1(32'hbb23f138),
	.w2(32'h3c5259b9),
	.w3(32'hb986a39a),
	.w4(32'hbab723e0),
	.w5(32'h3bc3ecdb),
	.w6(32'hbbd730ea),
	.w7(32'h3c49e52d),
	.w8(32'hba3139e9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8498ee),
	.w1(32'hbc4e6f97),
	.w2(32'h3c777805),
	.w3(32'h3a57abf3),
	.w4(32'h3c7a3751),
	.w5(32'h3b5b0b8d),
	.w6(32'hbd28aa94),
	.w7(32'hbbe5735d),
	.w8(32'h3bfbed60),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6361bc),
	.w1(32'h3b104f26),
	.w2(32'h3c20bdc5),
	.w3(32'hbc4bd210),
	.w4(32'hbc2c9692),
	.w5(32'h3c0d27bb),
	.w6(32'h3c96d0f0),
	.w7(32'h3a671213),
	.w8(32'h3abeb33d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0d06d),
	.w1(32'hbab9f0a8),
	.w2(32'h3c6a3880),
	.w3(32'h3c7a2593),
	.w4(32'h3bf1e8ce),
	.w5(32'h3cc25212),
	.w6(32'h3c2938ff),
	.w7(32'h3c566b4f),
	.w8(32'h3c68a040),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e1407),
	.w1(32'h3c2785a9),
	.w2(32'h3ce8ede6),
	.w3(32'h3baf890a),
	.w4(32'h3adf52c2),
	.w5(32'h3cb73ec4),
	.w6(32'h3c1ae0bc),
	.w7(32'h3bc7a9de),
	.w8(32'h3c1ffb11),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1982b),
	.w1(32'h3c1b8449),
	.w2(32'h3c8ccf08),
	.w3(32'h3c8ca59e),
	.w4(32'hbb1356eb),
	.w5(32'h395957c6),
	.w6(32'h3b877cd3),
	.w7(32'h3c68dd4b),
	.w8(32'h3c575fde),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e0003),
	.w1(32'h3c00a915),
	.w2(32'h3bba0000),
	.w3(32'hbc65f9fc),
	.w4(32'h3ca7f512),
	.w5(32'h3caf63b6),
	.w6(32'hbc1952b3),
	.w7(32'hba247e91),
	.w8(32'h3c4a2903),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66faad),
	.w1(32'h39edaa35),
	.w2(32'hbc0616eb),
	.w3(32'h3ad17855),
	.w4(32'h3d024594),
	.w5(32'h3c3b4610),
	.w6(32'h3c0ed1f1),
	.w7(32'h3ca1851f),
	.w8(32'hbbb5b426),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e2162),
	.w1(32'h37be7c68),
	.w2(32'h3c468680),
	.w3(32'h3c2ee24f),
	.w4(32'h3c207df7),
	.w5(32'h3bbe9f31),
	.w6(32'h3cad471a),
	.w7(32'h3c56b5e0),
	.w8(32'h3c1aa18d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc653992),
	.w1(32'hbc64aaa2),
	.w2(32'h3c89bb91),
	.w3(32'hbc1872ac),
	.w4(32'hbbc983bc),
	.w5(32'h3c3eb0db),
	.w6(32'h3ab49449),
	.w7(32'hbb45eeb5),
	.w8(32'h3b23aaeb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30b52e),
	.w1(32'h3c0775cb),
	.w2(32'hbc259904),
	.w3(32'hbce6b663),
	.w4(32'h3ae4ee0e),
	.w5(32'h3bebaac3),
	.w6(32'h3b392f5d),
	.w7(32'h3b73958e),
	.w8(32'hb9f6e19f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3df944),
	.w1(32'h3c8e1791),
	.w2(32'hb9048480),
	.w3(32'h3bf91e60),
	.w4(32'h3c8d11f2),
	.w5(32'h3c5ce4fa),
	.w6(32'h3c624abf),
	.w7(32'h3ae733a0),
	.w8(32'h3c82222d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f20f3),
	.w1(32'h3c07ccbd),
	.w2(32'h3cd3bee0),
	.w3(32'h3c810376),
	.w4(32'h3c61ac53),
	.w5(32'h3c091d63),
	.w6(32'h3b26124e),
	.w7(32'h3bdf1797),
	.w8(32'h3a5087f3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba744e1d),
	.w1(32'h3b262005),
	.w2(32'hbb106cbe),
	.w3(32'h3c3985bc),
	.w4(32'h3ca32c1a),
	.w5(32'h3cc8855b),
	.w6(32'h3c5298b1),
	.w7(32'h3b9d4138),
	.w8(32'hbc012912),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6ee00),
	.w1(32'hbaaba1e9),
	.w2(32'h3cc64a9d),
	.w3(32'h3c6c12ba),
	.w4(32'hba7825a0),
	.w5(32'hbc0ab1d9),
	.w6(32'h3a559f0c),
	.w7(32'h3b4bbb5c),
	.w8(32'h3bccc121),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8434f6),
	.w1(32'h3d33cd16),
	.w2(32'h3a8ce0dc),
	.w3(32'hbb07ef22),
	.w4(32'h3c869b16),
	.w5(32'h3bc5c3cb),
	.w6(32'h3c989075),
	.w7(32'h3c88715b),
	.w8(32'hbb4897cf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c474a7f),
	.w1(32'hbcbb02c4),
	.w2(32'hbbaa9e36),
	.w3(32'h3bb63a91),
	.w4(32'h3b08a861),
	.w5(32'h3ab8d627),
	.w6(32'h3be8c474),
	.w7(32'h3cb56370),
	.w8(32'hbc25b21e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec0d2d),
	.w1(32'h3c1fe59b),
	.w2(32'hb905c241),
	.w3(32'h3bb4dcc5),
	.w4(32'h3a76851e),
	.w5(32'hbba5b7e2),
	.w6(32'hbb6a6444),
	.w7(32'h3ba81a53),
	.w8(32'hbba9d6d9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2ad2f),
	.w1(32'hbc4f12e6),
	.w2(32'h3c2d79bd),
	.w3(32'h3b654699),
	.w4(32'hbc1c9bd8),
	.w5(32'h3c107ebb),
	.w6(32'hba1fa9b6),
	.w7(32'h3d1cf643),
	.w8(32'h3d202078),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc7c9),
	.w1(32'hbc167b03),
	.w2(32'hba353e74),
	.w3(32'hbbab9ec6),
	.w4(32'h3addffbe),
	.w5(32'hbb78ef4e),
	.w6(32'hba5f577c),
	.w7(32'hbb5c08f9),
	.w8(32'h3bffc989),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c3b92),
	.w1(32'h3cc8d0fa),
	.w2(32'h3c3d76a6),
	.w3(32'h3c804e3a),
	.w4(32'hbce03917),
	.w5(32'h3cef5107),
	.w6(32'h3bf30176),
	.w7(32'h3bf2a08d),
	.w8(32'h3b907913),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c741deb),
	.w1(32'h3c0af142),
	.w2(32'hbceef335),
	.w3(32'h3b43be3b),
	.w4(32'hbb722288),
	.w5(32'hbbf5c7cf),
	.w6(32'hbc7cdc90),
	.w7(32'h3bb96c6e),
	.w8(32'h395f4fc7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac06c1f),
	.w1(32'h3c205409),
	.w2(32'h3b962c7d),
	.w3(32'h3c545c21),
	.w4(32'h3c05d62b),
	.w5(32'h3888942e),
	.w6(32'h3c8e194e),
	.w7(32'h3b2d12a1),
	.w8(32'h3c04b450),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa70441),
	.w1(32'hbc5306ef),
	.w2(32'hbac328ea),
	.w3(32'h3c261c52),
	.w4(32'hba80643c),
	.w5(32'h3a809cf4),
	.w6(32'hbb19d866),
	.w7(32'hbcf9d179),
	.w8(32'hbc07c842),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0da639),
	.w1(32'h3b8ad59a),
	.w2(32'hbc63e6a2),
	.w3(32'h3d7dd503),
	.w4(32'h3c1e4008),
	.w5(32'hbbe87390),
	.w6(32'h3c0b6f2d),
	.w7(32'hbc8c5d90),
	.w8(32'h3bb9e21e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd066e3e),
	.w1(32'hbc6992b1),
	.w2(32'hbc6e4aa8),
	.w3(32'h3c28450f),
	.w4(32'h3c55d940),
	.w5(32'hbaf3997e),
	.w6(32'hbc07a1cf),
	.w7(32'h3be8f327),
	.w8(32'h3cb97f69),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae788c),
	.w1(32'h39beab74),
	.w2(32'hbaae7743),
	.w3(32'hba8cb461),
	.w4(32'h3c391b1a),
	.w5(32'hba19229b),
	.w6(32'h3c4bf5a3),
	.w7(32'hbbfe47fc),
	.w8(32'h3bd6a516),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21df69),
	.w1(32'h3a3104dc),
	.w2(32'h3ce7bdde),
	.w3(32'hb9ede450),
	.w4(32'h3c9c90bf),
	.w5(32'h3b068079),
	.w6(32'hbbf99ff5),
	.w7(32'hbb6b63c1),
	.w8(32'h3c68629d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad17fcd),
	.w1(32'h3a80d9aa),
	.w2(32'h3c8a1f9c),
	.w3(32'h3be21fb2),
	.w4(32'h3a15deda),
	.w5(32'hbbed71e6),
	.w6(32'hbc25d8a8),
	.w7(32'h3c78aeee),
	.w8(32'h3ca972ee),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afea1c),
	.w1(32'h378617bd),
	.w2(32'hbc945cf5),
	.w3(32'h3ba272e9),
	.w4(32'h3adaeffb),
	.w5(32'hbbb57f9d),
	.w6(32'hbb259ab8),
	.w7(32'h3ace069b),
	.w8(32'h3bfa6edc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd17315),
	.w1(32'hbbee13c5),
	.w2(32'hbbc5a4c9),
	.w3(32'h3adb9f7c),
	.w4(32'hbb79fb1d),
	.w5(32'hbba6db8d),
	.w6(32'h3bf1e243),
	.w7(32'hbc05faac),
	.w8(32'hbac40840),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01b3ea),
	.w1(32'hbce22f02),
	.w2(32'h3a7471ef),
	.w3(32'h3afd5937),
	.w4(32'hbcd47d59),
	.w5(32'h3bc32b54),
	.w6(32'h3b47fe66),
	.w7(32'hbb9be8a7),
	.w8(32'h3a6e8ebf),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0881b1),
	.w1(32'hbc145a8b),
	.w2(32'hbc0d0430),
	.w3(32'h3c6130a2),
	.w4(32'h3c828f2f),
	.w5(32'h3bbfd09b),
	.w6(32'h3b2bde09),
	.w7(32'h3c4fe530),
	.w8(32'hbc60da8b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89f48c),
	.w1(32'hbc5394c8),
	.w2(32'hbb60b0f9),
	.w3(32'h3b3fd742),
	.w4(32'h3b9371e1),
	.w5(32'h3c847920),
	.w6(32'h3b68bc27),
	.w7(32'h3b171039),
	.w8(32'h3ce53f88),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80724e),
	.w1(32'h3c24d6d7),
	.w2(32'h3bc74736),
	.w3(32'hbc4a7123),
	.w4(32'hb9787614),
	.w5(32'hbc38ea90),
	.w6(32'h389a4034),
	.w7(32'hbba440c5),
	.w8(32'h3be51622),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9328e),
	.w1(32'hba675b42),
	.w2(32'h3bb338b6),
	.w3(32'h3bc283d6),
	.w4(32'hbb599f6f),
	.w5(32'h3bc0a9cb),
	.w6(32'h3ac5e87c),
	.w7(32'h3a197ea8),
	.w8(32'h3acf2fe8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c4e15),
	.w1(32'h3acef634),
	.w2(32'h3c8ddbb0),
	.w3(32'hbb4ab120),
	.w4(32'h3c7a5390),
	.w5(32'hbae047ba),
	.w6(32'h3c3efea6),
	.w7(32'h3bc53eda),
	.w8(32'h3bec1dfb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3af693),
	.w1(32'h3b1696a7),
	.w2(32'hbb470a11),
	.w3(32'h3c670e8d),
	.w4(32'h3c198b6b),
	.w5(32'h3bb2127a),
	.w6(32'h3c1b8c0f),
	.w7(32'h3bacd546),
	.w8(32'hbc85a6da),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a20da),
	.w1(32'hbb8bb23e),
	.w2(32'h3b507177),
	.w3(32'h3c3bd23a),
	.w4(32'hbbd24bf4),
	.w5(32'hbb9717b7),
	.w6(32'h3a96a07a),
	.w7(32'hbcc9858a),
	.w8(32'h3bd934c0),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eac26),
	.w1(32'h386ba8bd),
	.w2(32'h3c1964b5),
	.w3(32'h3a862e17),
	.w4(32'hba12f47b),
	.w5(32'h3c0bd9e2),
	.w6(32'h3a7757d0),
	.w7(32'h3a87b8cf),
	.w8(32'hbb99d8ed),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfb3e9),
	.w1(32'hbc49ebd9),
	.w2(32'h3c032cfd),
	.w3(32'hb902277b),
	.w4(32'h3c080b7f),
	.w5(32'h3b47db01),
	.w6(32'h3b8a16d6),
	.w7(32'hbd149d8d),
	.w8(32'hbb993a1f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a578cd6),
	.w1(32'hba837880),
	.w2(32'h3c213526),
	.w3(32'hbbef030b),
	.w4(32'h3a1e855a),
	.w5(32'h3b951690),
	.w6(32'hbbdfeb83),
	.w7(32'hbbd7a4c0),
	.w8(32'hbc2ef17b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cd885),
	.w1(32'hba2041f7),
	.w2(32'hbc646f13),
	.w3(32'hbb6b2881),
	.w4(32'h3c5107d1),
	.w5(32'h3bb9e69a),
	.w6(32'h3c1c35c8),
	.w7(32'h3bf385b9),
	.w8(32'hb9459d6b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ee4be),
	.w1(32'h3b936fee),
	.w2(32'h3b489cd7),
	.w3(32'hbd0e776a),
	.w4(32'h3d7b77a2),
	.w5(32'hbd016f75),
	.w6(32'h3c349607),
	.w7(32'h3bf6282d),
	.w8(32'hbb393345),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85c4fe),
	.w1(32'h3c2d0704),
	.w2(32'h3b3b770b),
	.w3(32'h3ac8478e),
	.w4(32'h3b8ebaeb),
	.w5(32'h3ce1c532),
	.w6(32'hb8d26af3),
	.w7(32'hb85ef450),
	.w8(32'hbb98b6b0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6f732),
	.w1(32'hbc2677ac),
	.w2(32'h3a10af4c),
	.w3(32'hbb8bad66),
	.w4(32'hbafee3ed),
	.w5(32'hbb8e5de0),
	.w6(32'h3c84c7f0),
	.w7(32'h3a962d8f),
	.w8(32'h3c4bc615),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc18b9),
	.w1(32'hbb1afab1),
	.w2(32'h3b351acb),
	.w3(32'hb8ed8dfc),
	.w4(32'hbb6fb9c3),
	.w5(32'h3b8fea05),
	.w6(32'hbade9b06),
	.w7(32'h3c8ed490),
	.w8(32'h3b622dce),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48d186),
	.w1(32'h3bba09a3),
	.w2(32'hbc46f99f),
	.w3(32'hba1673a0),
	.w4(32'hbbeb88d0),
	.w5(32'h3b5b48b8),
	.w6(32'hbb2b3b95),
	.w7(32'h3bd98931),
	.w8(32'h3a3ddefe),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4f035),
	.w1(32'h3c91f2a5),
	.w2(32'hbc5a8a35),
	.w3(32'hbb4ef1e8),
	.w4(32'h3a8f5da2),
	.w5(32'hb8c25f99),
	.w6(32'hbc2a895a),
	.w7(32'hbb249af5),
	.w8(32'h3af7f22c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8afb51),
	.w1(32'hba82ec23),
	.w2(32'hbc9098b9),
	.w3(32'hbab50a27),
	.w4(32'hbad69e4c),
	.w5(32'h3b62d448),
	.w6(32'h38f341d7),
	.w7(32'hbc3afdf2),
	.w8(32'hbc1cf353),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ab0c1),
	.w1(32'hbc72c063),
	.w2(32'h3b3f4008),
	.w3(32'h3d22a862),
	.w4(32'h3c9829a2),
	.w5(32'hbb9fd311),
	.w6(32'hbba8474b),
	.w7(32'hbc875aeb),
	.w8(32'h3b8356ab),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4240b),
	.w1(32'hbbeabef5),
	.w2(32'hbb79df60),
	.w3(32'hbc86c3ba),
	.w4(32'hba641cb1),
	.w5(32'h3b166eaf),
	.w6(32'hbb77ab78),
	.w7(32'h3bd8cb46),
	.w8(32'h3c55b745),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10985e),
	.w1(32'hbb782f39),
	.w2(32'hbbfc13ce),
	.w3(32'h3bd98e89),
	.w4(32'hbbbb8666),
	.w5(32'h3c77b044),
	.w6(32'hbab36f55),
	.w7(32'h396c73cc),
	.w8(32'h3c5186f6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3145),
	.w1(32'hba22f0fd),
	.w2(32'hbb33aabe),
	.w3(32'hbc0ccb9b),
	.w4(32'hbc5a91a2),
	.w5(32'h3bb68834),
	.w6(32'h3d5142a2),
	.w7(32'hbc540f8d),
	.w8(32'hbb1cc891),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af84ad7),
	.w1(32'hbc153ea0),
	.w2(32'hbbefc1b1),
	.w3(32'hbb61aac4),
	.w4(32'h3c0fa86a),
	.w5(32'hbb9dc8ec),
	.w6(32'hbb7ee386),
	.w7(32'h3b1ef1e6),
	.w8(32'h3c00a161),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ca709),
	.w1(32'hbc333492),
	.w2(32'hbbbd257a),
	.w3(32'h3ab684fb),
	.w4(32'hbbe62ab2),
	.w5(32'hbc521784),
	.w6(32'h3b8c002a),
	.w7(32'h3886f8c1),
	.w8(32'hbb395930),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa82949),
	.w1(32'hbca4016f),
	.w2(32'hbc1f80dd),
	.w3(32'h3cdb0b93),
	.w4(32'hbc59efa2),
	.w5(32'h3c403d28),
	.w6(32'hbbb17254),
	.w7(32'hbb288197),
	.w8(32'hbb3a83ee),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa08d14),
	.w1(32'h3b305843),
	.w2(32'hbbaee1f5),
	.w3(32'h3b2dbfe0),
	.w4(32'h3c129d0b),
	.w5(32'h37bdbdb2),
	.w6(32'hbb823c88),
	.w7(32'h3bd22504),
	.w8(32'h3acb6601),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982b2af),
	.w1(32'h3be1a502),
	.w2(32'h3b88f15f),
	.w3(32'hbbc4a4ad),
	.w4(32'h3bb4a65b),
	.w5(32'hbb4f2d9a),
	.w6(32'hbb267321),
	.w7(32'hbb97b22e),
	.w8(32'hbcbed51a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9888f4),
	.w1(32'hbc7a6690),
	.w2(32'h3b958f80),
	.w3(32'h3bea4913),
	.w4(32'h3c449f43),
	.w5(32'hbb37960f),
	.w6(32'hbbb22488),
	.w7(32'hba1896f0),
	.w8(32'h3c1acc1a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b138bf5),
	.w1(32'h3b50a5d9),
	.w2(32'hbbd54fac),
	.w3(32'hbbc74cd7),
	.w4(32'hbbfc6e1f),
	.w5(32'hbd193a62),
	.w6(32'h3b7f82a7),
	.w7(32'h3a01c837),
	.w8(32'h3b751b14),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc668a08),
	.w1(32'hb964ec89),
	.w2(32'h39e51317),
	.w3(32'h3ab387eb),
	.w4(32'h3b8edfc3),
	.w5(32'hbbc61008),
	.w6(32'hbc8081bf),
	.w7(32'h3b4a0228),
	.w8(32'hbb942caa),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff9b62),
	.w1(32'hbae70950),
	.w2(32'hb8475ddc),
	.w3(32'hbbeb9b84),
	.w4(32'hbb85d3a3),
	.w5(32'h3bf6acba),
	.w6(32'h3c28b144),
	.w7(32'hbc0491ea),
	.w8(32'h3cf40df0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefe5ad),
	.w1(32'h3b3dd598),
	.w2(32'hbc21996d),
	.w3(32'h3c79991e),
	.w4(32'h3bcc1525),
	.w5(32'h3a93c117),
	.w6(32'hbc32a34f),
	.w7(32'hbbd85d6b),
	.w8(32'hbbf07552),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba813552),
	.w1(32'hb9ec119d),
	.w2(32'h3c576e24),
	.w3(32'h3aa5c324),
	.w4(32'hbb0ecade),
	.w5(32'hbc80a436),
	.w6(32'h3c12e8af),
	.w7(32'hbbc416af),
	.w8(32'hbbc6d061),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7057f),
	.w1(32'hbc4b156e),
	.w2(32'hbba8ef41),
	.w3(32'hb9cc430f),
	.w4(32'hbbc26897),
	.w5(32'h3c48bd56),
	.w6(32'h38d3f8f9),
	.w7(32'h3bc6c181),
	.w8(32'hb894182e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba698e39),
	.w1(32'h3aaa98f1),
	.w2(32'h3b2691c8),
	.w3(32'hbaee0ae4),
	.w4(32'h3aa1d84a),
	.w5(32'hbb7ac96a),
	.w6(32'h3c071439),
	.w7(32'hbbf78629),
	.w8(32'h3bd809ea),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be794e6),
	.w1(32'h38d26403),
	.w2(32'h38df8849),
	.w3(32'h3b4c927f),
	.w4(32'hbb5450d6),
	.w5(32'h392a94df),
	.w6(32'hbc96b367),
	.w7(32'hb9a015b7),
	.w8(32'hbb6b8b3e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5708a1),
	.w1(32'hba987ea9),
	.w2(32'h3be77767),
	.w3(32'hba91f664),
	.w4(32'hba5310c0),
	.w5(32'h3a8e0c56),
	.w6(32'h3b899d5a),
	.w7(32'h38fcb1c3),
	.w8(32'hbbe07e82),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fade),
	.w1(32'h3a0d8298),
	.w2(32'hbb80e48b),
	.w3(32'hbb9a01f6),
	.w4(32'h3c09053d),
	.w5(32'hbb806d8f),
	.w6(32'hbc6ccd21),
	.w7(32'h3c4b0618),
	.w8(32'h3b995252),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e5324),
	.w1(32'h3ca02d0d),
	.w2(32'hbc51f981),
	.w3(32'hbc2a2f7a),
	.w4(32'h39f2b4cf),
	.w5(32'hbc9d04f3),
	.w6(32'h3c417d5a),
	.w7(32'h3991abc1),
	.w8(32'h3bec4ff4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31da90),
	.w1(32'hbc4c6f19),
	.w2(32'h3ca8964b),
	.w3(32'hba5d243d),
	.w4(32'h3be66415),
	.w5(32'h3caf419b),
	.w6(32'hbc985723),
	.w7(32'hbc27b70d),
	.w8(32'h3c165d58),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00a370),
	.w1(32'hbb6eccba),
	.w2(32'h3bc88a0b),
	.w3(32'hbbadda13),
	.w4(32'hbb787307),
	.w5(32'hbbb47ba4),
	.w6(32'hbbd92591),
	.w7(32'h3bceedb4),
	.w8(32'h3c2018dc),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af83670),
	.w1(32'hbbf480b0),
	.w2(32'hbb5b57a3),
	.w3(32'h3b874b3b),
	.w4(32'h3bedccca),
	.w5(32'h3c51d2ff),
	.w6(32'h3b806a68),
	.w7(32'hbc1138c2),
	.w8(32'hbb50b417),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c59c2),
	.w1(32'hbb9f8bfe),
	.w2(32'hbc2688aa),
	.w3(32'hbc1b6577),
	.w4(32'hba9506ba),
	.w5(32'hbadf4df3),
	.w6(32'h3a0ef2d2),
	.w7(32'h3ad9c2e6),
	.w8(32'hbbd1511f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c578de3),
	.w1(32'hba8dec71),
	.w2(32'h3934b730),
	.w3(32'hbc029d7a),
	.w4(32'h3c1bc0a7),
	.w5(32'h3cb42311),
	.w6(32'hbc000fe0),
	.w7(32'h3ba68148),
	.w8(32'hbc2feea9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8024a8),
	.w1(32'hbb3b860b),
	.w2(32'h3c2fe2c7),
	.w3(32'hbc6624a7),
	.w4(32'hbb21df2f),
	.w5(32'h3b91cd90),
	.w6(32'hb994c97c),
	.w7(32'h3b9ab470),
	.w8(32'h3a5d3d83),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816b02),
	.w1(32'hbc9a756c),
	.w2(32'h3cab7fca),
	.w3(32'h3c6d0067),
	.w4(32'h3c0ec1ab),
	.w5(32'h3c48fc6a),
	.w6(32'h3befba7e),
	.w7(32'hbbcaf9b1),
	.w8(32'h3c4e9f93),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac58579),
	.w1(32'hbb8f4596),
	.w2(32'hbba6c94c),
	.w3(32'hb9c75746),
	.w4(32'hbbaad2be),
	.w5(32'hb9ffd28b),
	.w6(32'h3bdef2d3),
	.w7(32'h3cbb1282),
	.w8(32'h3a9eea0e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25f05d),
	.w1(32'hbb29ef70),
	.w2(32'hbbcc603f),
	.w3(32'hb8e44a26),
	.w4(32'hbaed258b),
	.w5(32'hba512ab5),
	.w6(32'h3b291546),
	.w7(32'h3a8c9946),
	.w8(32'h3b936341),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fe051),
	.w1(32'h3a073496),
	.w2(32'hbbcab613),
	.w3(32'hb9eb4ab8),
	.w4(32'hbc43fc8d),
	.w5(32'h3be658f4),
	.w6(32'hbbe8be3e),
	.w7(32'h3a7632b9),
	.w8(32'h3b819e69),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1d19e),
	.w1(32'hbb5bdc28),
	.w2(32'hb84dd837),
	.w3(32'hbc48a5b7),
	.w4(32'hbc4772f5),
	.w5(32'h3bd82888),
	.w6(32'hbb6d944c),
	.w7(32'h3b28a6d5),
	.w8(32'hbcb9a8c1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63e6ec),
	.w1(32'hbae70b0a),
	.w2(32'hbb92850c),
	.w3(32'hbad349b4),
	.w4(32'h3a995777),
	.w5(32'h3cb05e60),
	.w6(32'hbc3966ce),
	.w7(32'h39486022),
	.w8(32'hbb60e999),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09675a),
	.w1(32'h3b728675),
	.w2(32'hbad9f576),
	.w3(32'h3bf0460b),
	.w4(32'hbbabd242),
	.w5(32'h3baca17d),
	.w6(32'h3c5f410e),
	.w7(32'h3b318711),
	.w8(32'hbb39cd5e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9372316),
	.w1(32'hbbf5e514),
	.w2(32'hbc6bc228),
	.w3(32'hbb9deaa5),
	.w4(32'hbc2b602f),
	.w5(32'h3c02277a),
	.w6(32'hbc340484),
	.w7(32'h3d2a5cb9),
	.w8(32'hbc2c4f3d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4c84b),
	.w1(32'h3bf4bdb5),
	.w2(32'hbac198b2),
	.w3(32'hbadef1e0),
	.w4(32'h3a01415c),
	.w5(32'hbb89874e),
	.w6(32'h3b1816b1),
	.w7(32'h3c056719),
	.w8(32'hbaf3cb73),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeffed),
	.w1(32'hbc063809),
	.w2(32'h3b37736e),
	.w3(32'h3ae20785),
	.w4(32'h39b073bc),
	.w5(32'h3ad60dd0),
	.w6(32'h3768d45a),
	.w7(32'hbd015067),
	.w8(32'h3bbc3295),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d825),
	.w1(32'hbbe20681),
	.w2(32'hbc2c128a),
	.w3(32'hba0df3ae),
	.w4(32'hbaed7193),
	.w5(32'hbc0fce44),
	.w6(32'hbb0a68c7),
	.w7(32'hbb0ec1b4),
	.w8(32'h3be8fbcc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986a9d3),
	.w1(32'hbb84f109),
	.w2(32'hbc1a0f79),
	.w3(32'h3b8ba8d9),
	.w4(32'h3b817b63),
	.w5(32'h3c1dc2e7),
	.w6(32'h38690a08),
	.w7(32'h3a7dfb32),
	.w8(32'hbb379e90),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba419d9),
	.w1(32'h3c11481a),
	.w2(32'hbc10d0e2),
	.w3(32'h3bd766ff),
	.w4(32'h3b5f5cd7),
	.w5(32'hbb0f8a7c),
	.w6(32'hbc00d25c),
	.w7(32'h3a98cbaf),
	.w8(32'h3c2935a3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c388228),
	.w1(32'hba205761),
	.w2(32'h3b93b401),
	.w3(32'h3a582cbf),
	.w4(32'hb9e4b746),
	.w5(32'h3bdc3efc),
	.w6(32'hbbbb5b24),
	.w7(32'hbb5ae733),
	.w8(32'h3bea40b8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc037711),
	.w1(32'h3c9951f0),
	.w2(32'hbc469f00),
	.w3(32'h37fcfdc7),
	.w4(32'h3b639fd5),
	.w5(32'h3c325898),
	.w6(32'h3bc00ce0),
	.w7(32'hbb9bf863),
	.w8(32'hbcdb1abd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af28ff7),
	.w1(32'hb92d69a7),
	.w2(32'h3ba75469),
	.w3(32'hbc2c1a29),
	.w4(32'h39a27f36),
	.w5(32'h3b253ee2),
	.w6(32'h3be9643d),
	.w7(32'hbb7c7079),
	.w8(32'hbb927dab),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec48c4),
	.w1(32'h3ba745c6),
	.w2(32'hbb7f0c06),
	.w3(32'hbacecf42),
	.w4(32'h3c577adb),
	.w5(32'hbaeaea16),
	.w6(32'hbb4303b2),
	.w7(32'h3bb564dc),
	.w8(32'h3c4ab238),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbfb3c),
	.w1(32'hbb98584c),
	.w2(32'hbbceeee9),
	.w3(32'h3b7e347b),
	.w4(32'h3bc8c74d),
	.w5(32'h3ae89b68),
	.w6(32'hba9f422e),
	.w7(32'h3acefaf0),
	.w8(32'hbb477fcf),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08d394),
	.w1(32'h3c9ed0cb),
	.w2(32'hbc21be56),
	.w3(32'hb9d0e615),
	.w4(32'hbc0bea29),
	.w5(32'h3b52ee2b),
	.w6(32'hbb739774),
	.w7(32'hbb862bd5),
	.w8(32'h3afba487),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be050c2),
	.w1(32'h3bb35be7),
	.w2(32'h3bb48c5f),
	.w3(32'h3aa2beb6),
	.w4(32'hbb8a2bf9),
	.w5(32'h3af79517),
	.w6(32'h3815f723),
	.w7(32'h3ba19b4c),
	.w8(32'h3baa0a75),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367ccdff),
	.w1(32'hbb92a767),
	.w2(32'hbaa1d671),
	.w3(32'hbb047344),
	.w4(32'h3bf98dbe),
	.w5(32'hbb802d04),
	.w6(32'hbc394a59),
	.w7(32'hbc2140e9),
	.w8(32'h3b8d84e5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb94ead),
	.w1(32'hbc978975),
	.w2(32'h3af57df3),
	.w3(32'h3b8e4ae9),
	.w4(32'h3b06dd85),
	.w5(32'h3c085c10),
	.w6(32'hbc001c63),
	.w7(32'h3affffba),
	.w8(32'h3a63e990),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb284203),
	.w1(32'h3b9db2fc),
	.w2(32'hbc57e963),
	.w3(32'hbb892760),
	.w4(32'hbbbe4011),
	.w5(32'hbb032563),
	.w6(32'hbc1107cf),
	.w7(32'h39d610cf),
	.w8(32'hb9eda21c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9bd6b),
	.w1(32'h3c5307e0),
	.w2(32'hbcf1d37d),
	.w3(32'hbd090f3b),
	.w4(32'hbb49bcfe),
	.w5(32'h3bd61bb1),
	.w6(32'h3ae81ca3),
	.w7(32'hba952952),
	.w8(32'h3b1840c0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd96f3e),
	.w1(32'hbbd0e766),
	.w2(32'hbc0b8a0d),
	.w3(32'h3b2b2fe6),
	.w4(32'hbb7178d2),
	.w5(32'h3bd1ddff),
	.w6(32'hbac61444),
	.w7(32'hbbda1d64),
	.w8(32'hbc863a80),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2be646),
	.w1(32'hbc6e1273),
	.w2(32'hbc299c5c),
	.w3(32'hb90eb23b),
	.w4(32'hbb5e6807),
	.w5(32'h3b715900),
	.w6(32'hbb41518a),
	.w7(32'h3c0eb3c4),
	.w8(32'hbc478fe8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41723f),
	.w1(32'h3bb5795e),
	.w2(32'h3a59b31f),
	.w3(32'h3a786da6),
	.w4(32'hbc567d90),
	.w5(32'h3af1956d),
	.w6(32'hbbbcf3ea),
	.w7(32'hbc327715),
	.w8(32'h3c80fa68),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabbf2c),
	.w1(32'h3c19eaf3),
	.w2(32'hbb77afac),
	.w3(32'h386e982f),
	.w4(32'hbab9e883),
	.w5(32'h39d240b8),
	.w6(32'hbc3bf31c),
	.w7(32'hbc5fe5cc),
	.w8(32'hbb07c76d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e50a4),
	.w1(32'hbc050ba8),
	.w2(32'hbb9b322d),
	.w3(32'h3c095c78),
	.w4(32'hbc6ee983),
	.w5(32'hbbe63ea1),
	.w6(32'hbafa1f65),
	.w7(32'h3cd34c6a),
	.w8(32'hbc4e1726),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8237f1),
	.w1(32'hbcde586e),
	.w2(32'hbc85ce25),
	.w3(32'hbcce43b6),
	.w4(32'hbc3e2ea8),
	.w5(32'hb96b2dc2),
	.w6(32'hbbffbf04),
	.w7(32'h3bdb8cf9),
	.w8(32'hbc025120),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12afd6),
	.w1(32'hbc1a8578),
	.w2(32'h3b5fd3b7),
	.w3(32'h3c331656),
	.w4(32'hbc1d51fe),
	.w5(32'hbbcc5172),
	.w6(32'hbbad9a1d),
	.w7(32'hbc3a96c4),
	.w8(32'h3b662b61),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38abffcc),
	.w1(32'h3c24cec2),
	.w2(32'h3bd18020),
	.w3(32'h3a4f60f4),
	.w4(32'hba04942b),
	.w5(32'hbbbfc69b),
	.w6(32'hbc0daa5f),
	.w7(32'h3a8cbf49),
	.w8(32'h3d68eb9f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b6962),
	.w1(32'h3c9553f4),
	.w2(32'hbc4124e3),
	.w3(32'hb9d28cd5),
	.w4(32'hbd66f690),
	.w5(32'h3aad9c0e),
	.w6(32'h3b97417f),
	.w7(32'h3b673c04),
	.w8(32'h3b94e496),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10d1e7),
	.w1(32'h3be60d08),
	.w2(32'hbb30f634),
	.w3(32'hba89a1d4),
	.w4(32'hbc0ca7fd),
	.w5(32'hba66528b),
	.w6(32'hbc18f999),
	.w7(32'h3c48741f),
	.w8(32'hbb81a432),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88c57b),
	.w1(32'h3b327118),
	.w2(32'hbb603ae4),
	.w3(32'h3b0c2f6c),
	.w4(32'hba7fe528),
	.w5(32'h3b69f4da),
	.w6(32'hbcaab496),
	.w7(32'hbd39bc3f),
	.w8(32'h3b077e35),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4255fa),
	.w1(32'hba9f8157),
	.w2(32'h3a12928a),
	.w3(32'hbba22f15),
	.w4(32'hb926cc28),
	.w5(32'hbd0d608c),
	.w6(32'hbbd00be7),
	.w7(32'h3bb8d2e4),
	.w8(32'hbb8344c7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabade3),
	.w1(32'h3c4a6baa),
	.w2(32'hbbe2d9da),
	.w3(32'hbb72e258),
	.w4(32'hbb6f1c40),
	.w5(32'hbc2469a1),
	.w6(32'hbc67fb9c),
	.w7(32'hba9b0d07),
	.w8(32'hbbbe4550),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3700b),
	.w1(32'h3a72f7d8),
	.w2(32'hb6865d21),
	.w3(32'h3b06152f),
	.w4(32'hba16bf36),
	.w5(32'hbb53ae64),
	.w6(32'h3a1f02a2),
	.w7(32'hba3dfec9),
	.w8(32'hbb48edf0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca34535),
	.w1(32'h3beef990),
	.w2(32'h3a8a3d0e),
	.w3(32'hbc7e8650),
	.w4(32'hbc12f944),
	.w5(32'h3cabe2f9),
	.w6(32'hbb898f35),
	.w7(32'hbc0d71d0),
	.w8(32'h3c881c85),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b76c8),
	.w1(32'hbbe85ecc),
	.w2(32'h3bbf6bbf),
	.w3(32'hbb332e9e),
	.w4(32'hbc16c83e),
	.w5(32'h3b585ecd),
	.w6(32'h3ac273a7),
	.w7(32'h3bcef200),
	.w8(32'hbb830bed),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28cf4f),
	.w1(32'h3c5e43c1),
	.w2(32'hbc17c5d3),
	.w3(32'hbb1f5876),
	.w4(32'hbbb93fb4),
	.w5(32'hbc70cc8d),
	.w6(32'hbb9b7b7e),
	.w7(32'hbc884a73),
	.w8(32'h3af5e0e7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac4c76),
	.w1(32'hbbf57db9),
	.w2(32'hbb6e4405),
	.w3(32'hbc865619),
	.w4(32'hbc221bff),
	.w5(32'h3c145c16),
	.w6(32'h3c0ce236),
	.w7(32'hbb87e76d),
	.w8(32'hb9c1c96f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedd78e),
	.w1(32'hbba806bc),
	.w2(32'hbbf13bf8),
	.w3(32'hbbf347f3),
	.w4(32'h3c3846c0),
	.w5(32'hbc683ee1),
	.w6(32'h3b93fb9b),
	.w7(32'hb6b44ef7),
	.w8(32'hbb911edf),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef8630),
	.w1(32'h3c4db82a),
	.w2(32'h3b969404),
	.w3(32'h3c47954d),
	.w4(32'h3b15314c),
	.w5(32'h3b197176),
	.w6(32'hbc6fcb53),
	.w7(32'h3b039576),
	.w8(32'h390b6418),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba45f2),
	.w1(32'hbc0d299e),
	.w2(32'h3caefbd9),
	.w3(32'hba836d51),
	.w4(32'h3b081f2a),
	.w5(32'hbb84b931),
	.w6(32'hbc1a6502),
	.w7(32'hbb17adf8),
	.w8(32'hbc189b45),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc598bb1),
	.w1(32'hbb9b316b),
	.w2(32'hbb2bcb7e),
	.w3(32'hba79dd78),
	.w4(32'hbc4142b0),
	.w5(32'hbadc47d9),
	.w6(32'hbbf41ec6),
	.w7(32'hbc2e7ab5),
	.w8(32'hbaead912),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb568da6),
	.w1(32'hbb8dca7d),
	.w2(32'h3ae71a1f),
	.w3(32'h3b3d6070),
	.w4(32'hbc87775d),
	.w5(32'h3c17e4c3),
	.w6(32'hbbea6fac),
	.w7(32'h3bdba153),
	.w8(32'hbc08be97),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42819a),
	.w1(32'hba00926e),
	.w2(32'hb8915520),
	.w3(32'h39b557fa),
	.w4(32'h3c225511),
	.w5(32'hba6331cb),
	.w6(32'hbb4e7a63),
	.w7(32'hbb9a98ae),
	.w8(32'h38ab19d5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ca9dc),
	.w1(32'hba796e31),
	.w2(32'h3a494742),
	.w3(32'hbc0b2eb2),
	.w4(32'h39a5b5bf),
	.w5(32'hbbac1d68),
	.w6(32'hbc2e7170),
	.w7(32'hbbc76566),
	.w8(32'h3c1f1265),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b08ce),
	.w1(32'hbb82c7ad),
	.w2(32'hbb415b1d),
	.w3(32'hbb1ba366),
	.w4(32'h3a4e6bd2),
	.w5(32'h3c505d6a),
	.w6(32'h3bd61ea6),
	.w7(32'h3b3accc3),
	.w8(32'h3b949c51),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ca2dc),
	.w1(32'hbc72c73a),
	.w2(32'h3b12b2de),
	.w3(32'hba5d71ea),
	.w4(32'h3b6b7ffe),
	.w5(32'hbbb7532c),
	.w6(32'hb89547a3),
	.w7(32'h3bef6015),
	.w8(32'h3a8d26d3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9454f),
	.w1(32'h3b50cbb7),
	.w2(32'hbb192323),
	.w3(32'hbb95a35a),
	.w4(32'h3bfd2a20),
	.w5(32'hbcb61013),
	.w6(32'hb9c54a00),
	.w7(32'hbd0de2ce),
	.w8(32'hbbbc7e94),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc374f59),
	.w1(32'h3ae8ca20),
	.w2(32'hbb8e0b7c),
	.w3(32'h3c1f91fc),
	.w4(32'hbbdfce2c),
	.w5(32'h3bc610bf),
	.w6(32'hbb3bdd04),
	.w7(32'hba15311b),
	.w8(32'hbb8b1b3e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc313bd9),
	.w1(32'hbc7d36a7),
	.w2(32'hbb995a51),
	.w3(32'h3c3352f3),
	.w4(32'h3ad96899),
	.w5(32'h3c4fcb15),
	.w6(32'h3b1e3ffd),
	.w7(32'hbc1c7b63),
	.w8(32'hbb3f1304),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d11632),
	.w1(32'h3b9e5206),
	.w2(32'hba3bb560),
	.w3(32'h3be30484),
	.w4(32'h3c51a18c),
	.w5(32'hbb2511d8),
	.w6(32'hba46fdc1),
	.w7(32'h399bb72f),
	.w8(32'hbb96de80),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c599b80),
	.w1(32'hbd31a1b5),
	.w2(32'h3c4b1809),
	.w3(32'h3a68f364),
	.w4(32'h3aa250a7),
	.w5(32'hbad738fc),
	.w6(32'h3ba92577),
	.w7(32'h3b26bcd7),
	.w8(32'hbb5d3bb6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d2545),
	.w1(32'h3c269c21),
	.w2(32'hbb8f9807),
	.w3(32'h3b21bbb6),
	.w4(32'hbb7e7c2b),
	.w5(32'hbc507ca2),
	.w6(32'h3b5b6536),
	.w7(32'h3bc6aa51),
	.w8(32'hbba020be),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc262d84),
	.w1(32'hbbef19e2),
	.w2(32'hbb4aa8b7),
	.w3(32'hbb0059bb),
	.w4(32'h3bee377e),
	.w5(32'hbc869dfa),
	.w6(32'h3cdd4e1b),
	.w7(32'hbc892b7b),
	.w8(32'h3be66659),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca51251),
	.w1(32'h3c47bb3e),
	.w2(32'h3c796d32),
	.w3(32'hba2e2e84),
	.w4(32'hbb7501d2),
	.w5(32'hb9ed0fbf),
	.w6(32'h3b3b9657),
	.w7(32'hbbbb1b38),
	.w8(32'h3b9f33f4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4f6a1),
	.w1(32'hba3ac85e),
	.w2(32'hbb66462b),
	.w3(32'h3bbadf01),
	.w4(32'hbbd14e63),
	.w5(32'hbb48fb5f),
	.w6(32'h3c1b14b7),
	.w7(32'h3c9a61a4),
	.w8(32'h3ac24aba),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81446a),
	.w1(32'h3cba637f),
	.w2(32'hbc09e059),
	.w3(32'hb8a75342),
	.w4(32'hbb8cec18),
	.w5(32'hbc13232b),
	.w6(32'h3b947a77),
	.w7(32'h3923b69a),
	.w8(32'hbcb0fcea),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe5997),
	.w1(32'hbb0d3d67),
	.w2(32'h3b27eb8c),
	.w3(32'h3b30f16e),
	.w4(32'hbb8e5194),
	.w5(32'h3cc15d11),
	.w6(32'h3aca9a6c),
	.w7(32'h3be153e5),
	.w8(32'hbbc988a0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8439),
	.w1(32'hba7e6b2f),
	.w2(32'hbc2dccc3),
	.w3(32'h3be171ce),
	.w4(32'h3be8a6f4),
	.w5(32'h3bc48dff),
	.w6(32'hbb52f1d7),
	.w7(32'h3b5f98e9),
	.w8(32'h3b165058),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd098502),
	.w1(32'h3c1ce1b0),
	.w2(32'h3a840855),
	.w3(32'hbbd7184b),
	.w4(32'hba03bdaa),
	.w5(32'h3ba51ef9),
	.w6(32'hbc3589ea),
	.w7(32'hbb94d5f0),
	.w8(32'h39c7c45a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06ef26),
	.w1(32'h398507b6),
	.w2(32'h3b80b424),
	.w3(32'h3bd69193),
	.w4(32'hbbd8979f),
	.w5(32'h3c4864a7),
	.w6(32'hbb65507a),
	.w7(32'hbb0c08b3),
	.w8(32'hb8a12924),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c973d1c),
	.w1(32'hbab2baa1),
	.w2(32'h3c31de1d),
	.w3(32'h3be078f6),
	.w4(32'h3be9de65),
	.w5(32'hba43abb5),
	.w6(32'hbbb1bfb7),
	.w7(32'hbaccabb2),
	.w8(32'hbc32c19f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39677877),
	.w1(32'hbb034f25),
	.w2(32'h3bac6ca5),
	.w3(32'h38fffe9b),
	.w4(32'h3d02ef0c),
	.w5(32'hbc3e6a30),
	.w6(32'hbc21ccc0),
	.w7(32'h3c2bba24),
	.w8(32'h3bf573cc),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb570c7e),
	.w1(32'h3baaeb85),
	.w2(32'h3c40a8b1),
	.w3(32'h3bd003b0),
	.w4(32'h3c2928bc),
	.w5(32'hbb9ea66f),
	.w6(32'h3c50a209),
	.w7(32'h3b28dd92),
	.w8(32'h3c93b530),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0715d2),
	.w1(32'h3b279ff5),
	.w2(32'h3bb4c2f7),
	.w3(32'h3bee6790),
	.w4(32'hbb409f76),
	.w5(32'h3d07672a),
	.w6(32'hb9444da0),
	.w7(32'h3bccc82d),
	.w8(32'h3c06d8c6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e3b1),
	.w1(32'h3c2b9a10),
	.w2(32'hbb8237ae),
	.w3(32'hbb52f70c),
	.w4(32'h3b04a150),
	.w5(32'hbbe4d0c2),
	.w6(32'hbbe62573),
	.w7(32'hb9a886ab),
	.w8(32'hbc0e1ecc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb519baf),
	.w1(32'hbc0c95de),
	.w2(32'h3b514254),
	.w3(32'hba89c764),
	.w4(32'hbb1dee6b),
	.w5(32'hbbff9984),
	.w6(32'hbae22b77),
	.w7(32'hbc0d4f35),
	.w8(32'hbbf0c52f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376884b8),
	.w1(32'h3c1dda7f),
	.w2(32'h3aaec17c),
	.w3(32'hbb4e1bde),
	.w4(32'hbaf3ae24),
	.w5(32'h3cc11704),
	.w6(32'h3a766196),
	.w7(32'h3cd321dd),
	.w8(32'hbbd1ba55),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8322d3),
	.w1(32'hb822e156),
	.w2(32'hbab3037b),
	.w3(32'hba03ecd1),
	.w4(32'h3bca6de4),
	.w5(32'h3afe228b),
	.w6(32'hbb0499ab),
	.w7(32'hba3672ef),
	.w8(32'hbc0bf9b7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc4d1b),
	.w1(32'h3aebc51f),
	.w2(32'h3c0430fe),
	.w3(32'h3b8d4438),
	.w4(32'hbc88df33),
	.w5(32'hba058a98),
	.w6(32'hbb9dc98c),
	.w7(32'hbc03625e),
	.w8(32'hbae163db),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31f731),
	.w1(32'hbc03bac8),
	.w2(32'hbc4cb8e8),
	.w3(32'h3a7b21b2),
	.w4(32'h3b58971e),
	.w5(32'h39a5210e),
	.w6(32'hbbbee713),
	.w7(32'h3ba1267e),
	.w8(32'hbbe27d90),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745eb0),
	.w1(32'h3cef5797),
	.w2(32'hba5b4714),
	.w3(32'h3c600994),
	.w4(32'h3b79dba4),
	.w5(32'hbb9fcf15),
	.w6(32'h3c551895),
	.w7(32'hbc0650e5),
	.w8(32'hbc1dfe01),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1620ba),
	.w1(32'h3b9370f8),
	.w2(32'hbbe11031),
	.w3(32'hb9de36a1),
	.w4(32'hbc262791),
	.w5(32'hbb7355d5),
	.w6(32'hb7dd8fe8),
	.w7(32'hbc2ed1f6),
	.w8(32'h3a786377),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d2cd7),
	.w1(32'h3ce814df),
	.w2(32'h3b8e2569),
	.w3(32'h3c933fbf),
	.w4(32'h3c157544),
	.w5(32'hbbbe5fbb),
	.w6(32'h3bf12913),
	.w7(32'h3b10cd52),
	.w8(32'h3cd44c5d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c322bca),
	.w1(32'h3bf4210c),
	.w2(32'hbc02ae72),
	.w3(32'h3bb576ac),
	.w4(32'hbba698f4),
	.w5(32'h3beab267),
	.w6(32'h3ba27ed7),
	.w7(32'hbb838dbf),
	.w8(32'hbb9089c6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9410c),
	.w1(32'hbac55f1a),
	.w2(32'h3c3efce7),
	.w3(32'h3b4ff8c7),
	.w4(32'h3a88088b),
	.w5(32'hbb0a4766),
	.w6(32'hbc097953),
	.w7(32'hbc376984),
	.w8(32'h3cd1d8ee),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91cf3d),
	.w1(32'hb9faddac),
	.w2(32'h3b9f6abe),
	.w3(32'hbb1343fa),
	.w4(32'h3aad9c7b),
	.w5(32'hbc1a5100),
	.w6(32'hbb8bb845),
	.w7(32'h3cf7c40b),
	.w8(32'h3b128924),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37697731),
	.w1(32'hbbad5ce8),
	.w2(32'hbb2fa6e4),
	.w3(32'h3b4368cc),
	.w4(32'hbbfa461a),
	.w5(32'hbb758e1f),
	.w6(32'hbb14ea50),
	.w7(32'hba21895f),
	.w8(32'hbb964402),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe0de7),
	.w1(32'hba9362c3),
	.w2(32'h3bbf0a0f),
	.w3(32'hbb873c74),
	.w4(32'h3bafd206),
	.w5(32'hbc2cc53c),
	.w6(32'hbc4343b6),
	.w7(32'h3ba43fb3),
	.w8(32'h3bd9f0d4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule