module layer_8_featuremap_107(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beda812),
	.w1(32'h3b8ab751),
	.w2(32'hbb697108),
	.w3(32'h3b6bbe04),
	.w4(32'h3cb00f63),
	.w5(32'h3c3d3b43),
	.w6(32'hbb08f796),
	.w7(32'h3c6d93a1),
	.w8(32'h3c8f320b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf5bd77),
	.w1(32'hbc9d7049),
	.w2(32'h3bec6f86),
	.w3(32'h39e584c7),
	.w4(32'h3c642ec7),
	.w5(32'h3c604ed9),
	.w6(32'h3c5eca21),
	.w7(32'h3c8e49d4),
	.w8(32'hbc36afbc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2e162),
	.w1(32'h3c963727),
	.w2(32'h3ba512bb),
	.w3(32'h3bd30331),
	.w4(32'h3ba66253),
	.w5(32'hbbb60642),
	.w6(32'h3aeca79d),
	.w7(32'h3c27d26d),
	.w8(32'hbca50e63),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a19df),
	.w1(32'h3d0032dc),
	.w2(32'h3a6eae41),
	.w3(32'hbc49c595),
	.w4(32'hbb04150f),
	.w5(32'h3b5d37ca),
	.w6(32'hbc7c143e),
	.w7(32'h3c1cbf0e),
	.w8(32'h3c829ee5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07b1b3),
	.w1(32'hbb838dbe),
	.w2(32'hbbf3d2dc),
	.w3(32'h3c097513),
	.w4(32'hbab508ec),
	.w5(32'hbc1adcc5),
	.w6(32'h3bbd2a4d),
	.w7(32'hbc265910),
	.w8(32'hbc947f41),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75d0e4),
	.w1(32'hbb2beac5),
	.w2(32'h3bd1ce2e),
	.w3(32'hbc6dff01),
	.w4(32'h3bb7c47d),
	.w5(32'h3bedc575),
	.w6(32'hbc71b867),
	.w7(32'h3bc7d67a),
	.w8(32'hbc21c0b4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a01cb),
	.w1(32'hbb55daf5),
	.w2(32'h3cb027d3),
	.w3(32'h3bf5d228),
	.w4(32'h3c2a5892),
	.w5(32'h3ce01d52),
	.w6(32'hbc38d134),
	.w7(32'h3c76625a),
	.w8(32'hbb2ce1ae),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd46e16),
	.w1(32'hbc554739),
	.w2(32'h3cc2b7b7),
	.w3(32'h3c704a88),
	.w4(32'hbc3b4bf4),
	.w5(32'hbcda0721),
	.w6(32'hbc68921b),
	.w7(32'hbc43e2c7),
	.w8(32'hbc672bbe),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d86f4a3),
	.w1(32'hbc46f020),
	.w2(32'h3c7a4a5d),
	.w3(32'hbb53ad02),
	.w4(32'hbc05adc2),
	.w5(32'hbbcba0e5),
	.w6(32'h3a9583f0),
	.w7(32'h3cccb40a),
	.w8(32'h3cb5c607),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50ef19),
	.w1(32'hbc6b5801),
	.w2(32'hbbd0eb26),
	.w3(32'hba4374ce),
	.w4(32'h3a5f2d73),
	.w5(32'h3ca8587d),
	.w6(32'h3c02218e),
	.w7(32'h3b92b33d),
	.w8(32'h3ca88496),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd29e9fe),
	.w1(32'hba33cb99),
	.w2(32'h3bca1a24),
	.w3(32'h3ba9b2da),
	.w4(32'hbbf0594a),
	.w5(32'hbcd0d51f),
	.w6(32'h3ba65f24),
	.w7(32'hbcbf6bbe),
	.w8(32'hbcf7347d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d730b38),
	.w1(32'h3c3bbe9d),
	.w2(32'h3c7da75b),
	.w3(32'hbcbe7986),
	.w4(32'hb97bf435),
	.w5(32'hbc70618e),
	.w6(32'hbc90edf7),
	.w7(32'hb9905fc4),
	.w8(32'hbcbe57fa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becf08e),
	.w1(32'hbbf91d95),
	.w2(32'h3ad218b9),
	.w3(32'h3a3b648a),
	.w4(32'hba29f2c4),
	.w5(32'h3c020ebb),
	.w6(32'h3b906d66),
	.w7(32'hbb88ca07),
	.w8(32'hbc226b49),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2cc72),
	.w1(32'h3b5b0ced),
	.w2(32'h3ab227ce),
	.w3(32'h3ba3f283),
	.w4(32'hbbf94dcd),
	.w5(32'h3af2c9cd),
	.w6(32'hbbb7543b),
	.w7(32'hbb7e4c28),
	.w8(32'hb994eb10),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b212d),
	.w1(32'h38f210d3),
	.w2(32'h3ae602c4),
	.w3(32'h399bd759),
	.w4(32'hbbbfb9c3),
	.w5(32'hbb3e3b4d),
	.w6(32'hbaa205d1),
	.w7(32'hbae98b7a),
	.w8(32'hbb197dc8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6c800),
	.w1(32'hbb4ad9d5),
	.w2(32'hbc80deca),
	.w3(32'hba9c1fcb),
	.w4(32'hbc03f67f),
	.w5(32'hbc21c499),
	.w6(32'hbb4b034e),
	.w7(32'h3c35e52a),
	.w8(32'h3c5b4a4c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51d8a2),
	.w1(32'hbb9ae574),
	.w2(32'h3c3dc8cd),
	.w3(32'hbab0ac16),
	.w4(32'hbc9d4c6c),
	.w5(32'hbc93e329),
	.w6(32'hbbaba488),
	.w7(32'hbabcae93),
	.w8(32'h3c466715),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde61d0),
	.w1(32'hbbd920ce),
	.w2(32'hbb9b6025),
	.w3(32'h3b3544c3),
	.w4(32'hbbfc0260),
	.w5(32'h3beec9c8),
	.w6(32'h3ac0ad06),
	.w7(32'h3c3b10b3),
	.w8(32'h3adc93b3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaeabf),
	.w1(32'hbc3f2d72),
	.w2(32'hbc4ffaa8),
	.w3(32'h3c91f3f5),
	.w4(32'h3b8f00b1),
	.w5(32'hbc3dca31),
	.w6(32'hbc988921),
	.w7(32'h3a83db03),
	.w8(32'h3981cfbf),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e72a),
	.w1(32'hbb3a1bb8),
	.w2(32'hba21b3ce),
	.w3(32'hbb7081e3),
	.w4(32'h3c9963cc),
	.w5(32'h3d4d0cea),
	.w6(32'hbc41ff4f),
	.w7(32'hbcc0a0c3),
	.w8(32'hbcd439c2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c05cd),
	.w1(32'hbb86f9fc),
	.w2(32'hbb900b03),
	.w3(32'h3bbb3338),
	.w4(32'h3ba00144),
	.w5(32'h3c36e3cc),
	.w6(32'hbcb2ead0),
	.w7(32'hbbb1e03e),
	.w8(32'h3c042e5f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbe21c),
	.w1(32'h3b883fa7),
	.w2(32'hbbf9d4db),
	.w3(32'hbc095e22),
	.w4(32'hbaac1d44),
	.w5(32'hbca11f23),
	.w6(32'h3b494864),
	.w7(32'hbb54f23a),
	.w8(32'h3ba5cea7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60dc8a),
	.w1(32'hbbc7988f),
	.w2(32'hbac4dd17),
	.w3(32'hbb338845),
	.w4(32'h3bb0983e),
	.w5(32'hbc190a8a),
	.w6(32'h3c9bc83a),
	.w7(32'h3b9a73fb),
	.w8(32'h3c2a9523),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7a964),
	.w1(32'hbb74c8b4),
	.w2(32'h3c83632b),
	.w3(32'hbc9cb508),
	.w4(32'h3b9985e5),
	.w5(32'hbbdd4703),
	.w6(32'hbb4028b4),
	.w7(32'h3c936ec3),
	.w8(32'h3bd88625),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b833df7),
	.w1(32'hbba61ea6),
	.w2(32'h3b5af458),
	.w3(32'hbb96a18d),
	.w4(32'h3a8813aa),
	.w5(32'hbb7f8821),
	.w6(32'hba9c5dad),
	.w7(32'h3aa65736),
	.w8(32'h3c3005bf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2cc90),
	.w1(32'hbb9d0a74),
	.w2(32'h3bc2e494),
	.w3(32'hbb2f8d5a),
	.w4(32'hbc4714b1),
	.w5(32'hbccf67fb),
	.w6(32'h3bd9ead0),
	.w7(32'hba3b6a34),
	.w8(32'h3cee3ca5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba677eec),
	.w1(32'h3b63f6e6),
	.w2(32'hbad1083b),
	.w3(32'hbc59b223),
	.w4(32'hb9a4c221),
	.w5(32'h3cd70778),
	.w6(32'h3cabd818),
	.w7(32'hbbde89c2),
	.w8(32'hbc74bbdd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d203733),
	.w1(32'h3cd2360c),
	.w2(32'hbd276936),
	.w3(32'h3c05d293),
	.w4(32'h3d014fdb),
	.w5(32'h3d5c5492),
	.w6(32'hbd29a7e7),
	.w7(32'hbc87b54a),
	.w8(32'hbc85de85),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a26c5),
	.w1(32'hbc99da7c),
	.w2(32'h3c85e139),
	.w3(32'h3bfd77b5),
	.w4(32'h3cf0858c),
	.w5(32'h3cad4d36),
	.w6(32'hbcd5ba8b),
	.w7(32'hbbd6b135),
	.w8(32'hbc062fe0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc80f0f),
	.w1(32'h3c0c8966),
	.w2(32'h3b3eb79c),
	.w3(32'hbbc25594),
	.w4(32'hbba401b2),
	.w5(32'hbca3d4d9),
	.w6(32'h3c4cd42d),
	.w7(32'h3c02b10e),
	.w8(32'h3ce7e7a2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed7116),
	.w1(32'hbbd8ffbc),
	.w2(32'h3c3b2f09),
	.w3(32'hbc0b44a2),
	.w4(32'h3a8b0135),
	.w5(32'h3bb6c0fc),
	.w6(32'h3c4771f0),
	.w7(32'h3bdce7ed),
	.w8(32'h3c34b0e6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66a3e3),
	.w1(32'h3c8a1b15),
	.w2(32'hbcd103b1),
	.w3(32'h3bc09259),
	.w4(32'h3d00ad69),
	.w5(32'h3d3d117d),
	.w6(32'h3c5f6ab6),
	.w7(32'hbc38b74a),
	.w8(32'hbccbd169),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcef9931),
	.w1(32'hbcf847ca),
	.w2(32'h3cf3f51b),
	.w3(32'h3cb9a3f3),
	.w4(32'hbcb59f3c),
	.w5(32'hbd3eac4b),
	.w6(32'hbd13c28c),
	.w7(32'hbc7c1597),
	.w8(32'hbc355758),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd75e52),
	.w1(32'h3c9b1b32),
	.w2(32'h3aff158b),
	.w3(32'hbbaa1d29),
	.w4(32'hbc21893b),
	.w5(32'hbcc5ab80),
	.w6(32'h3cd7ea92),
	.w7(32'h3b994418),
	.w8(32'h3b7f5974),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a4698),
	.w1(32'h3b942acb),
	.w2(32'h3bea851b),
	.w3(32'hbc87bd45),
	.w4(32'hbb92dcf4),
	.w5(32'h3a1a9525),
	.w6(32'h3c8214e1),
	.w7(32'h3bc4aadf),
	.w8(32'h3c40c7a6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5597d7),
	.w1(32'h3c110f4f),
	.w2(32'hbafa53e1),
	.w3(32'hb9ab1e29),
	.w4(32'hbc2d6649),
	.w5(32'h3accdd57),
	.w6(32'h3b69a429),
	.w7(32'hbba73ee2),
	.w8(32'hbc291dcf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc625b),
	.w1(32'hbc0edf1e),
	.w2(32'hbbe88af4),
	.w3(32'h3c02456c),
	.w4(32'h3c4a64a2),
	.w5(32'h3cab4a0f),
	.w6(32'hbb270e1b),
	.w7(32'hbc88c5d1),
	.w8(32'hbcf1e7de),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b241f),
	.w1(32'hbd042720),
	.w2(32'h3a61fa5c),
	.w3(32'h3b567de1),
	.w4(32'hbc5551f1),
	.w5(32'hbcf92a47),
	.w6(32'hbcdb4497),
	.w7(32'hbb6fe564),
	.w8(32'h3c07e134),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e2c3c),
	.w1(32'h3c25735e),
	.w2(32'hbc096db0),
	.w3(32'hbc16beed),
	.w4(32'h3c880640),
	.w5(32'h3d02a601),
	.w6(32'h3c249ce0),
	.w7(32'hbb4851fb),
	.w8(32'hbc751eba),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52c21f),
	.w1(32'hbc910ed8),
	.w2(32'hbb290d02),
	.w3(32'h3c61f5a6),
	.w4(32'hbc1763b7),
	.w5(32'hbc0d2e8d),
	.w6(32'hbc5077e5),
	.w7(32'h3b4e5f16),
	.w8(32'hbb125dd8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe41b6),
	.w1(32'hbbbae5ab),
	.w2(32'hbba17a76),
	.w3(32'hbbd68ebb),
	.w4(32'h3c99176d),
	.w5(32'h3c319ea8),
	.w6(32'hbadc162f),
	.w7(32'hb9b34a46),
	.w8(32'hbba0ab52),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c690ed5),
	.w1(32'h3bbd3375),
	.w2(32'hbc2486bf),
	.w3(32'hbbd40871),
	.w4(32'hbbcd714e),
	.w5(32'h3caa442a),
	.w6(32'hbc82577f),
	.w7(32'h3bf59a8b),
	.w8(32'hbaca0060),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48c8c5),
	.w1(32'h39c613bc),
	.w2(32'h38177250),
	.w3(32'hba539850),
	.w4(32'hbce23762),
	.w5(32'hbd3f7efe),
	.w6(32'hbd017fff),
	.w7(32'h3c9e29cb),
	.w8(32'h3d605dba),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a2128),
	.w1(32'h3bf4dea4),
	.w2(32'h3b569d4b),
	.w3(32'hbc319b2e),
	.w4(32'h3aa95111),
	.w5(32'h3c0f8900),
	.w6(32'h3d2210b8),
	.w7(32'hbb830f84),
	.w8(32'hbc193706),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8af73e),
	.w1(32'h3bf16e75),
	.w2(32'hbc26e492),
	.w3(32'h3bd6b1b2),
	.w4(32'h3c60423b),
	.w5(32'h3bf4b352),
	.w6(32'hbc0a5dc9),
	.w7(32'h3c5906e0),
	.w8(32'h3c19f734),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69265b),
	.w1(32'hbbbceaf3),
	.w2(32'hbb884da2),
	.w3(32'h3c3ac3b4),
	.w4(32'hbbe250f2),
	.w5(32'h3b80dadc),
	.w6(32'h3a580051),
	.w7(32'hbbc2ef99),
	.w8(32'hbb446d66),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70105f),
	.w1(32'h3b9542f9),
	.w2(32'h3b06daa3),
	.w3(32'h3b44bb0c),
	.w4(32'h3cc2f766),
	.w5(32'h3c0bfb73),
	.w6(32'hbb928a0e),
	.w7(32'hbc8a8c6b),
	.w8(32'hbc20a389),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ed90d),
	.w1(32'hbc2be649),
	.w2(32'hbc837100),
	.w3(32'hbbc270a0),
	.w4(32'hbbb51638),
	.w5(32'hbd07d8b2),
	.w6(32'h3b986021),
	.w7(32'hbc3ce455),
	.w8(32'h3cb70a67),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d6dce),
	.w1(32'h3bc0790e),
	.w2(32'hbd0322a8),
	.w3(32'hbc18903e),
	.w4(32'h3ca24c46),
	.w5(32'h3d03d046),
	.w6(32'h3d0ea743),
	.w7(32'h3c66e25b),
	.w8(32'hbc269993),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd16fdcb),
	.w1(32'hbca995a3),
	.w2(32'hbd0f1502),
	.w3(32'h3ccc1b4e),
	.w4(32'h3d0a0224),
	.w5(32'h3ceb2767),
	.w6(32'hbcffd3ce),
	.w7(32'hbbd12f52),
	.w8(32'hbca62416),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd28441a),
	.w1(32'hbd53dbca),
	.w2(32'hba745b7c),
	.w3(32'hbbe55a53),
	.w4(32'hbc85ce94),
	.w5(32'hbd0d0979),
	.w6(32'hbd1c928e),
	.w7(32'h3cb3635e),
	.w8(32'h3d2b4a78),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d332),
	.w1(32'hbbd002fa),
	.w2(32'hbcdf3505),
	.w3(32'hbbeefe9f),
	.w4(32'h3c3fc6b4),
	.w5(32'h3b2e1df5),
	.w6(32'h3cf87a7a),
	.w7(32'hbccd00fd),
	.w8(32'h3b85b46e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fe51b),
	.w1(32'hbb8c4366),
	.w2(32'hbb896752),
	.w3(32'h3c88278c),
	.w4(32'h3c47bf6c),
	.w5(32'h3bdcee3c),
	.w6(32'h3c8014f1),
	.w7(32'h3c275b64),
	.w8(32'hbb031164),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4670d),
	.w1(32'h3bfbb26c),
	.w2(32'h3ab18f24),
	.w3(32'h3c83bab7),
	.w4(32'hba0836cc),
	.w5(32'h3be6d858),
	.w6(32'h3bc3885a),
	.w7(32'hbb203794),
	.w8(32'hbbd2b26e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb805cb40),
	.w1(32'h3a97c697),
	.w2(32'hbb1fcff1),
	.w3(32'h3ad678ae),
	.w4(32'h3c1d6987),
	.w5(32'h3c9541d3),
	.w6(32'hbba1484a),
	.w7(32'hbc3e8c8c),
	.w8(32'hbc1c81a0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bb5e4),
	.w1(32'hbc22155b),
	.w2(32'hbc634ecf),
	.w3(32'hb95cd458),
	.w4(32'h3c3d1466),
	.w5(32'h3b837415),
	.w6(32'hbc27cc8c),
	.w7(32'hbaa902db),
	.w8(32'hbc3b01a1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a5892),
	.w1(32'hbc647f77),
	.w2(32'hb7fc8e05),
	.w3(32'h3b3fcfee),
	.w4(32'hbc36a1b7),
	.w5(32'hbbe18480),
	.w6(32'hbae28960),
	.w7(32'hbaca1df0),
	.w8(32'h3b78fcc3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9201e),
	.w1(32'h3b35122b),
	.w2(32'h3b3fe012),
	.w3(32'hbbfb4b26),
	.w4(32'hbc1ad0a3),
	.w5(32'hbcbb930f),
	.w6(32'h3a89686c),
	.w7(32'h3c7fb05e),
	.w8(32'h3d4d6f0e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9288ea),
	.w1(32'h3c0b23c2),
	.w2(32'h3b7cbe67),
	.w3(32'hbc87ead3),
	.w4(32'h3a3e244d),
	.w5(32'h3c007675),
	.w6(32'h3cc74a51),
	.w7(32'hbbb2c6c4),
	.w8(32'hbc18c942),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81c384),
	.w1(32'h3b84b5a7),
	.w2(32'hbbafe57c),
	.w3(32'h3b772fcc),
	.w4(32'h3bf920fa),
	.w5(32'h3c813225),
	.w6(32'hbbb2ee45),
	.w7(32'h3b33e73a),
	.w8(32'hbc92cb6a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37c220),
	.w1(32'hba690cd2),
	.w2(32'h3c2de674),
	.w3(32'h39c3c641),
	.w4(32'hbab895b0),
	.w5(32'h3c9c4e33),
	.w6(32'hbc3d4fc9),
	.w7(32'h3c630bb7),
	.w8(32'h3bd57ad7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcedce),
	.w1(32'hbbb15dfb),
	.w2(32'h3c173d0f),
	.w3(32'hbc14ec29),
	.w4(32'h3b575242),
	.w5(32'h3bd2ae13),
	.w6(32'hbc99fdaf),
	.w7(32'h3c4a3e5c),
	.w8(32'h3c11e29c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be68be7),
	.w1(32'h3aac8404),
	.w2(32'hbca07b4c),
	.w3(32'h3ba6b1f1),
	.w4(32'h3c7860cc),
	.w5(32'hbc45a95f),
	.w6(32'h3bef0082),
	.w7(32'h39f9ac53),
	.w8(32'h3bb0f479),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe528ff),
	.w1(32'hbc3f4fc3),
	.w2(32'h3c53657a),
	.w3(32'hbb9bcc29),
	.w4(32'h3cb7f281),
	.w5(32'h3c9f69f3),
	.w6(32'hb987998a),
	.w7(32'hbbcd8922),
	.w8(32'hbc9ab3cb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e5054),
	.w1(32'h3c47d42c),
	.w2(32'hba7a134c),
	.w3(32'h3b81f001),
	.w4(32'h3b397e29),
	.w5(32'hbaa165fe),
	.w6(32'hbb035762),
	.w7(32'hbb1041b6),
	.w8(32'hbb4dd6e7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beff1a4),
	.w1(32'h391932e8),
	.w2(32'h3c9fcc69),
	.w3(32'hbcf2f3fd),
	.w4(32'hbcf797f6),
	.w5(32'hbd40c421),
	.w6(32'hbc551714),
	.w7(32'h3c1f8757),
	.w8(32'h3cf0713e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e9586),
	.w1(32'h3b0170ca),
	.w2(32'h3c2e7231),
	.w3(32'hbca3c6ab),
	.w4(32'hbc22ca7f),
	.w5(32'hbbaa6fbc),
	.w6(32'h3ca78910),
	.w7(32'h3c30deb8),
	.w8(32'h3af9bb36),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14106b),
	.w1(32'h3abee62b),
	.w2(32'hbb919f92),
	.w3(32'h3bd1067e),
	.w4(32'hbc193d57),
	.w5(32'h3c91baf3),
	.w6(32'h39168a8c),
	.w7(32'hbbdb8aa3),
	.w8(32'hbcc811e3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc418881),
	.w1(32'h3c16f613),
	.w2(32'hbb7b3cbf),
	.w3(32'h3c7de283),
	.w4(32'h3ce58832),
	.w5(32'h3d2291cf),
	.w6(32'hbc9a1ca9),
	.w7(32'hbbf4d9b9),
	.w8(32'hbc6b4bb6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c297fa9),
	.w1(32'h3bf87858),
	.w2(32'h3c4798b8),
	.w3(32'h3c94553e),
	.w4(32'hbbbca5c2),
	.w5(32'hbc902931),
	.w6(32'hbcbed28b),
	.w7(32'h3c5c1974),
	.w8(32'h3a7af19a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60289a),
	.w1(32'h3c09362a),
	.w2(32'hbb94351b),
	.w3(32'hbc8b9c32),
	.w4(32'hbceeba3d),
	.w5(32'hbc07ebe5),
	.w6(32'h3c855437),
	.w7(32'hbb3447d2),
	.w8(32'h3c4f6d29),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66f003),
	.w1(32'h3c68de2c),
	.w2(32'hbb9e1e58),
	.w3(32'hbb6ec92d),
	.w4(32'h3bd450a5),
	.w5(32'h3b32afa4),
	.w6(32'hbb921e1d),
	.w7(32'h3b564664),
	.w8(32'hbb704f12),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4be4f9),
	.w1(32'h3c715874),
	.w2(32'hbab1df96),
	.w3(32'hbba97826),
	.w4(32'hbb17e35a),
	.w5(32'h3c4652e8),
	.w6(32'hba2ef696),
	.w7(32'hbc12a039),
	.w8(32'hbc6a8572),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb022e09),
	.w1(32'hbc41f083),
	.w2(32'hbbca94d0),
	.w3(32'h3adac2d5),
	.w4(32'hbc2e2fba),
	.w5(32'h3a229371),
	.w6(32'hbc50c4ef),
	.w7(32'h3bf4606c),
	.w8(32'h3c28aa9a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30094e),
	.w1(32'hbb84da87),
	.w2(32'hbc03fb99),
	.w3(32'h3bb06291),
	.w4(32'h3b99f2c5),
	.w5(32'hbaf0f04d),
	.w6(32'h39ff5401),
	.w7(32'hbc0ede34),
	.w8(32'hbbad2518),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbcfbe),
	.w1(32'hbccd871b),
	.w2(32'hbb13d858),
	.w3(32'h3bd996cd),
	.w4(32'hbb2af046),
	.w5(32'h3c2b6760),
	.w6(32'hbc4aed37),
	.w7(32'h3c34521f),
	.w8(32'hba6b8f69),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ee84e),
	.w1(32'hbc007dac),
	.w2(32'h3aaa5484),
	.w3(32'h3b48814d),
	.w4(32'h3b94db15),
	.w5(32'h3abd4cff),
	.w6(32'h3b09fc7b),
	.w7(32'h3ac41cf2),
	.w8(32'hbb1e4aca),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a234e),
	.w1(32'h3bd0be17),
	.w2(32'hbb39b6bb),
	.w3(32'h3c469af6),
	.w4(32'h3b5fd040),
	.w5(32'h3bd6ddcd),
	.w6(32'hb8e609ef),
	.w7(32'h39e59162),
	.w8(32'hbb4988fd),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3703e2),
	.w1(32'h3be0d64d),
	.w2(32'hbbd59d0a),
	.w3(32'h3c09bb8f),
	.w4(32'hbb7aa4e1),
	.w5(32'hbba64504),
	.w6(32'h3c274023),
	.w7(32'hbb4fcb45),
	.w8(32'hbbf43665),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9fa37),
	.w1(32'hbae545eb),
	.w2(32'hbade4af8),
	.w3(32'hbbaf2e28),
	.w4(32'hbc0f21d6),
	.w5(32'hbb1ae4d8),
	.w6(32'hbbe3f04f),
	.w7(32'hba5732e2),
	.w8(32'h3b2c1d53),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2cb67),
	.w1(32'h3b7ba61b),
	.w2(32'hbb8408e4),
	.w3(32'h3c509449),
	.w4(32'hbcb59503),
	.w5(32'hba47edf1),
	.w6(32'hbaf44dbd),
	.w7(32'hbae45c77),
	.w8(32'h3c638ef2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f5ded),
	.w1(32'h3cd431a7),
	.w2(32'hbb661bdb),
	.w3(32'h3b40f832),
	.w4(32'h3b20d34a),
	.w5(32'hbc07a304),
	.w6(32'h3c37a98c),
	.w7(32'hbb09dfac),
	.w8(32'hbc35371d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc230094),
	.w1(32'hbc60a14e),
	.w2(32'hbad4df4f),
	.w3(32'h3aaa2344),
	.w4(32'h3baeb19a),
	.w5(32'hba7721f1),
	.w6(32'hbc90a306),
	.w7(32'h3c653f07),
	.w8(32'h3aef5890),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387084fc),
	.w1(32'hbcac4620),
	.w2(32'h3c02c466),
	.w3(32'h3c80bc65),
	.w4(32'hba83f682),
	.w5(32'hbbb7d8a2),
	.w6(32'h3cc4f776),
	.w7(32'h3cd75aea),
	.w8(32'h3b345b6b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc18690),
	.w1(32'hbc1dc229),
	.w2(32'hbcba9161),
	.w3(32'h3b4655d0),
	.w4(32'h3c80e729),
	.w5(32'h3bfb5176),
	.w6(32'hbcc0504c),
	.w7(32'h3be8d297),
	.w8(32'h3d5d3b68),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4bd3a),
	.w1(32'h3bcdc0c1),
	.w2(32'hbbcf3140),
	.w3(32'hbcb39b49),
	.w4(32'h397ac5dd),
	.w5(32'h3c52f2b7),
	.w6(32'hbb57d6b3),
	.w7(32'hbc7e806f),
	.w8(32'hb97e6918),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc473a7),
	.w1(32'h3d1b78c3),
	.w2(32'hbc35147c),
	.w3(32'hbcb48b22),
	.w4(32'hba8fb3fd),
	.w5(32'hbc8381c1),
	.w6(32'h3c84cbe7),
	.w7(32'h3c075e36),
	.w8(32'h3c3d9f2d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a4b19),
	.w1(32'h3b1b855e),
	.w2(32'hbbd8dc95),
	.w3(32'h3b813274),
	.w4(32'hbb89c505),
	.w5(32'hbbfbbd5a),
	.w6(32'hbc8d84f8),
	.w7(32'hbbbde1cf),
	.w8(32'hbbf903e3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7ebd8),
	.w1(32'hba359947),
	.w2(32'h3bf9f797),
	.w3(32'hbaae8a13),
	.w4(32'h3ad4a3e6),
	.w5(32'hbbc74c96),
	.w6(32'hbae5638f),
	.w7(32'h3c137c4b),
	.w8(32'h3b0dfd5e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94c922),
	.w1(32'hb9443cff),
	.w2(32'hbc4c87e6),
	.w3(32'hbbe89828),
	.w4(32'hbc82f01b),
	.w5(32'hbbef5ad9),
	.w6(32'h39b50227),
	.w7(32'h3b7a6b81),
	.w8(32'hbbe980a2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c7904),
	.w1(32'h3b874847),
	.w2(32'h3bd77fbc),
	.w3(32'h3c82e41d),
	.w4(32'hbaa2a62f),
	.w5(32'h3bc8800e),
	.w6(32'h3c806692),
	.w7(32'hba65ff2e),
	.w8(32'hbb763585),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1de960),
	.w1(32'hbb7e3481),
	.w2(32'hbb9c0661),
	.w3(32'h3c9d6eef),
	.w4(32'h3bbb6ddc),
	.w5(32'h3c8106fe),
	.w6(32'h3c104e59),
	.w7(32'hbc386f3d),
	.w8(32'hbba4adae),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdfdf87),
	.w1(32'h3cbd6cb3),
	.w2(32'hbb2d279f),
	.w3(32'h3ae2db32),
	.w4(32'hbba4dcbf),
	.w5(32'h3b8505cb),
	.w6(32'h3ce7ce58),
	.w7(32'hbc3949ee),
	.w8(32'hbce3ad2d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19acb0),
	.w1(32'hbd133f3a),
	.w2(32'hbc8b9cd0),
	.w3(32'h3c33c86b),
	.w4(32'hba87f7ed),
	.w5(32'hbb58b0d1),
	.w6(32'h3b85cd08),
	.w7(32'hba9ae299),
	.w8(32'h3a70df84),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7981c8),
	.w1(32'h3be212cc),
	.w2(32'h3a8e2e0c),
	.w3(32'h3c5263ff),
	.w4(32'h3941eba2),
	.w5(32'hb65cd436),
	.w6(32'h3c3ee0cb),
	.w7(32'hb92bcf25),
	.w8(32'hbb456078),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00b286),
	.w1(32'h3b3c4f90),
	.w2(32'hbc9773ec),
	.w3(32'hba4359bc),
	.w4(32'hbb87c90d),
	.w5(32'h3c368a0d),
	.w6(32'hbabf70cc),
	.w7(32'hbcbbd26c),
	.w8(32'h3be782c1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4011a6),
	.w1(32'h3c87130e),
	.w2(32'h3b982e17),
	.w3(32'h3c1098b0),
	.w4(32'hbb62351b),
	.w5(32'h3c6365e2),
	.w6(32'h3c8e36b6),
	.w7(32'h3bc89125),
	.w8(32'h3c9a6507),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d131b58),
	.w1(32'hbc46461d),
	.w2(32'hbbdb4755),
	.w3(32'hbc035920),
	.w4(32'h3b32001c),
	.w5(32'hbc9a4722),
	.w6(32'hbd06bee2),
	.w7(32'h3b6d9c5f),
	.w8(32'hbc2402df),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cb541),
	.w1(32'h3c34d26f),
	.w2(32'h3b61bf52),
	.w3(32'hbb8d7d4b),
	.w4(32'h3c20d833),
	.w5(32'h3ad7505f),
	.w6(32'h3c746f22),
	.w7(32'h3bc9fac1),
	.w8(32'h3c279e10),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bc228),
	.w1(32'h3af8e154),
	.w2(32'hbbd57c55),
	.w3(32'hbbc7a2a4),
	.w4(32'hbc2e868e),
	.w5(32'h3bedb511),
	.w6(32'hbc4bc30f),
	.w7(32'hbca11379),
	.w8(32'hbbaa0d6e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc996f27),
	.w1(32'hbbe2dd50),
	.w2(32'hbc4d2bee),
	.w3(32'h3cb95106),
	.w4(32'h3bf46475),
	.w5(32'h3c6aacc8),
	.w6(32'hba8ddf37),
	.w7(32'hbc03662f),
	.w8(32'h3c0b5dac),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6926cc),
	.w1(32'hbbd51c2f),
	.w2(32'h3a2782ca),
	.w3(32'h3c7385c6),
	.w4(32'hbbe8de28),
	.w5(32'hbc29f116),
	.w6(32'h397809b3),
	.w7(32'hbb1ff3f0),
	.w8(32'hbb13e25b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b861e01),
	.w1(32'h3bda1ce4),
	.w2(32'hbc662247),
	.w3(32'hb942320c),
	.w4(32'hbc052741),
	.w5(32'h3b32b53d),
	.w6(32'h3ce0acbe),
	.w7(32'hbbdab2f1),
	.w8(32'hbc1c9b79),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc529424),
	.w1(32'hbca1106b),
	.w2(32'h3b74b71e),
	.w3(32'h3c37fa6f),
	.w4(32'hbb87767b),
	.w5(32'hbc2b5be7),
	.w6(32'h3bac3158),
	.w7(32'h3b7deafa),
	.w8(32'hb9e41ad4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93bc6ed),
	.w1(32'hbba99fa4),
	.w2(32'hbc1e5997),
	.w3(32'hbc29a005),
	.w4(32'hbc31895d),
	.w5(32'hbbefd826),
	.w6(32'hba641c0f),
	.w7(32'hbc48064b),
	.w8(32'hbc8ef1d8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b384fac),
	.w1(32'h3b644e65),
	.w2(32'h39516b92),
	.w3(32'h3c804738),
	.w4(32'h3c297545),
	.w5(32'h3b40e952),
	.w6(32'hbc053fb8),
	.w7(32'h3bcf4ecf),
	.w8(32'hbaeb59ad),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46d005),
	.w1(32'hbc10fb3b),
	.w2(32'h3b5f6b7e),
	.w3(32'hbb91bb97),
	.w4(32'hbc069deb),
	.w5(32'h3c031a04),
	.w6(32'hbc660df4),
	.w7(32'hbc4c2dbb),
	.w8(32'h3c12e106),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdb0c2),
	.w1(32'hbabf94f7),
	.w2(32'h3b58295b),
	.w3(32'hbb551c20),
	.w4(32'h3b0926ab),
	.w5(32'h384062fa),
	.w6(32'hbbffbe1b),
	.w7(32'hba353699),
	.w8(32'hbc2a77ed),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f4b69),
	.w1(32'hbb2ac049),
	.w2(32'hbb4d6873),
	.w3(32'h3c6c5b0d),
	.w4(32'hbc77252f),
	.w5(32'h3ce378df),
	.w6(32'hba57f18f),
	.w7(32'hbc3573c3),
	.w8(32'h3acc1416),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3c41c),
	.w1(32'h3bdce7a5),
	.w2(32'h3b341c6e),
	.w3(32'h3bff56df),
	.w4(32'h3bb8f59d),
	.w5(32'hbc3cef03),
	.w6(32'h3cb12588),
	.w7(32'h3b10a2ec),
	.w8(32'hbbe0b460),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1242c),
	.w1(32'hbc746e5d),
	.w2(32'hbaa24963),
	.w3(32'h3bdaebd4),
	.w4(32'hbc24c1d5),
	.w5(32'h3b63882c),
	.w6(32'hbca2cf93),
	.w7(32'hbbf25cf2),
	.w8(32'hbc88ed53),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cc1c9),
	.w1(32'hbcbe623c),
	.w2(32'hba25b056),
	.w3(32'h3b2d03db),
	.w4(32'hbbcee412),
	.w5(32'h3cb820a6),
	.w6(32'h3c793134),
	.w7(32'h3b5407cb),
	.w8(32'h3b7bee04),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdc0761),
	.w1(32'hbb84f56c),
	.w2(32'hbc925be6),
	.w3(32'hbc0136e1),
	.w4(32'hbc2d2894),
	.w5(32'h3c08ccbd),
	.w6(32'h3ad3595f),
	.w7(32'hbc5b37f7),
	.w8(32'hbba56118),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac1ecc),
	.w1(32'hbc2453c6),
	.w2(32'hbd1f0a23),
	.w3(32'h3a879288),
	.w4(32'hbd1deb51),
	.w5(32'hba8ec63d),
	.w6(32'hbb130e18),
	.w7(32'hbd23650c),
	.w8(32'hbca3501d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a7900),
	.w1(32'hbbdb73ff),
	.w2(32'h3c1d77a9),
	.w3(32'h3cca2767),
	.w4(32'hbb1b1eed),
	.w5(32'hbcbf1620),
	.w6(32'h3d2cd519),
	.w7(32'hbb3d7770),
	.w8(32'hba6506eb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadb57c),
	.w1(32'hbbd490c7),
	.w2(32'h3bc6002e),
	.w3(32'h3cc47456),
	.w4(32'h3c425ecd),
	.w5(32'hbc6026fc),
	.w6(32'hbcec7829),
	.w7(32'h3d107d5c),
	.w8(32'h3d14c650),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf0c26d),
	.w1(32'h3b8ad583),
	.w2(32'h3cb94e31),
	.w3(32'hbd5a5dfd),
	.w4(32'hbaf746a3),
	.w5(32'hbb32fc3d),
	.w6(32'hbd37dc2b),
	.w7(32'h3a89fb0b),
	.w8(32'h3a8f2946),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0e20e),
	.w1(32'h39f9dcf3),
	.w2(32'hbb2f1f4f),
	.w3(32'h3c1c2432),
	.w4(32'h3bb2e619),
	.w5(32'h3bb6062b),
	.w6(32'h3c6f0f42),
	.w7(32'h39929389),
	.w8(32'hbb3dca46),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9456a98),
	.w1(32'h3b9f1861),
	.w2(32'hbc13b990),
	.w3(32'h3c5ded00),
	.w4(32'hbbfc807b),
	.w5(32'h3a90769d),
	.w6(32'h3c33606d),
	.w7(32'h3b495876),
	.w8(32'h3ba4ff1d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1bb39),
	.w1(32'hbc27d9ba),
	.w2(32'hbab782af),
	.w3(32'h3b92a953),
	.w4(32'hbc059fcb),
	.w5(32'hb8b409cf),
	.w6(32'h3bd042f2),
	.w7(32'hbb32635e),
	.w8(32'hbc8187ec),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc836c5e),
	.w1(32'hba8e1cd0),
	.w2(32'h3b445959),
	.w3(32'h3d0f0632),
	.w4(32'hbac6ebe5),
	.w5(32'h3b0bb72e),
	.w6(32'h3cf358e8),
	.w7(32'hb9a9fe3c),
	.w8(32'h3b699640),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1eb99d),
	.w1(32'hbb92505a),
	.w2(32'hbc13f9b9),
	.w3(32'hbc150242),
	.w4(32'hbb4b916e),
	.w5(32'hbc5bec65),
	.w6(32'hbbb527d2),
	.w7(32'hbb4e9d89),
	.w8(32'h3b160356),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc464b41),
	.w1(32'hbb2a777d),
	.w2(32'h39c61ace),
	.w3(32'h3c7c2e96),
	.w4(32'h3a974789),
	.w5(32'h3ad981d5),
	.w6(32'hbc5eece3),
	.w7(32'hbab701ce),
	.w8(32'hbc0be07e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad1458),
	.w1(32'h3a2d6eb4),
	.w2(32'hbb55aa2c),
	.w3(32'h3c724555),
	.w4(32'h3c22994b),
	.w5(32'h3afde22c),
	.w6(32'h3bb091af),
	.w7(32'hb9615ea6),
	.w8(32'h3c596c52),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a9498),
	.w1(32'hb9a9a3ca),
	.w2(32'hbc3cf6d7),
	.w3(32'h3bff0305),
	.w4(32'hbbd42013),
	.w5(32'h3cad23e0),
	.w6(32'hbb470e71),
	.w7(32'hbcf3de94),
	.w8(32'hbc390a95),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf96bf5),
	.w1(32'h3c211ce4),
	.w2(32'hbc4239d0),
	.w3(32'h3d0a3b43),
	.w4(32'hbc2bb17f),
	.w5(32'h3b406474),
	.w6(32'h3c5e9a31),
	.w7(32'hbc7babf7),
	.w8(32'hbc116168),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c3a68),
	.w1(32'hbc22bec5),
	.w2(32'h3b5df092),
	.w3(32'h39642ed0),
	.w4(32'hbbfe8ac6),
	.w5(32'h3ca25ca6),
	.w6(32'h3b413541),
	.w7(32'h3b296e7a),
	.w8(32'hbcc05439),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7e27e),
	.w1(32'h3c60e2fa),
	.w2(32'hbbc0935d),
	.w3(32'hbb953810),
	.w4(32'h3c0cab89),
	.w5(32'hbb078447),
	.w6(32'h3d1667fe),
	.w7(32'hb857cb58),
	.w8(32'hbb33b166),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule