module layer_10_featuremap_241(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e1fa4),
	.w1(32'hbb93787c),
	.w2(32'hbbaa852b),
	.w3(32'hbba94697),
	.w4(32'hbbaeb17c),
	.w5(32'h3bacc9f0),
	.w6(32'hbbc50366),
	.w7(32'hbbf0956e),
	.w8(32'h397b679a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2c219),
	.w1(32'h3aa48791),
	.w2(32'h3a3f984c),
	.w3(32'h3a3c3f92),
	.w4(32'h3b7c2e67),
	.w5(32'hbbaf3e8e),
	.w6(32'hbb4291b0),
	.w7(32'h3b27f379),
	.w8(32'hbb8b7ab5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8720e1),
	.w1(32'hbbffca70),
	.w2(32'h3b8a61bf),
	.w3(32'hb7c44aa2),
	.w4(32'h3bffce82),
	.w5(32'hbb8be795),
	.w6(32'hbba3acc7),
	.w7(32'h3b8e9581),
	.w8(32'hbb97c10e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aa0ef),
	.w1(32'hbb123008),
	.w2(32'h3b0c1f6a),
	.w3(32'h3a529f1f),
	.w4(32'h3b00008a),
	.w5(32'hbba9a217),
	.w6(32'hba087f0b),
	.w7(32'hb936e563),
	.w8(32'hbb955c1d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3af35d),
	.w1(32'h3c744d36),
	.w2(32'hbc0b51be),
	.w3(32'h3c503421),
	.w4(32'hbc72a4fb),
	.w5(32'hbb6cc356),
	.w6(32'h3cc5f96e),
	.w7(32'hbc31e0f0),
	.w8(32'hbb0c1d3f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bede2),
	.w1(32'h3acfe7c5),
	.w2(32'h3b632264),
	.w3(32'h3af41d35),
	.w4(32'h3b9d3555),
	.w5(32'hba912c0f),
	.w6(32'h3b55df18),
	.w7(32'h3ba2b4d2),
	.w8(32'hb9e4c521),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852ae4),
	.w1(32'hbab34939),
	.w2(32'hbaa51cc5),
	.w3(32'h3abe7334),
	.w4(32'h3b164a9b),
	.w5(32'hbb40d6cc),
	.w6(32'h3a24d450),
	.w7(32'h396548d2),
	.w8(32'hba4766a8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7f6bb),
	.w1(32'h3b2c0074),
	.w2(32'hbb12ed87),
	.w3(32'hbb558421),
	.w4(32'hbb8de501),
	.w5(32'hb9c8b0f8),
	.w6(32'h3b0ba2fc),
	.w7(32'hbb73c51a),
	.w8(32'hb99e8977),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad26469),
	.w1(32'h39e351f1),
	.w2(32'hba6c574e),
	.w3(32'h3a76fdcd),
	.w4(32'h3a0d80be),
	.w5(32'hbb434a42),
	.w6(32'h3ae7d2e2),
	.w7(32'h391cd0df),
	.w8(32'hb94d92b8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba552a21),
	.w1(32'h3af649dc),
	.w2(32'h3b57d6fa),
	.w3(32'h3a373409),
	.w4(32'h3b27ff86),
	.w5(32'hbb543ffb),
	.w6(32'h3b57ff84),
	.w7(32'h3b61ad7b),
	.w8(32'h39c86847),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cf81f),
	.w1(32'hbabcf875),
	.w2(32'h3b611caf),
	.w3(32'h3ba0687e),
	.w4(32'h3b5e14be),
	.w5(32'hb7d9ac3a),
	.w6(32'h3ba7da67),
	.w7(32'h3b1df6cc),
	.w8(32'hba7b698a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd651c5),
	.w1(32'hba0e1879),
	.w2(32'hbba8b31e),
	.w3(32'hbb837c70),
	.w4(32'hbbd63a29),
	.w5(32'h3a8190a4),
	.w6(32'hbbf34e3a),
	.w7(32'hbbdad4ac),
	.w8(32'hb8ba7e5d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9792c9),
	.w1(32'h3c01db47),
	.w2(32'hbb09be87),
	.w3(32'h3c1e5767),
	.w4(32'hbbab6f91),
	.w5(32'h3acc7fb6),
	.w6(32'h3b68ff9d),
	.w7(32'h3866c297),
	.w8(32'hbc1dd9d1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a702ebc),
	.w1(32'hbd0161fc),
	.w2(32'hbaba8de0),
	.w3(32'hbd0f7fd0),
	.w4(32'hbbb1827b),
	.w5(32'hbb1fd7b1),
	.w6(32'hbce70a67),
	.w7(32'hbc3ce101),
	.w8(32'hbb08625c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7a2ee),
	.w1(32'h3b219147),
	.w2(32'h3b3f0993),
	.w3(32'hbb033deb),
	.w4(32'h3b5a90b1),
	.w5(32'hbbef40a4),
	.w6(32'hbb082668),
	.w7(32'h3add8903),
	.w8(32'hbc1b77bc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156aad),
	.w1(32'hbb99ecc0),
	.w2(32'hb9639b97),
	.w3(32'hbb3af25c),
	.w4(32'hbab52c8f),
	.w5(32'hbb31341d),
	.w6(32'hbb1346d7),
	.w7(32'hbadecf45),
	.w8(32'hbbe73ca7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27caa8),
	.w1(32'h3ab59de4),
	.w2(32'h3a0277d6),
	.w3(32'hbb5a5c86),
	.w4(32'h3a8b1aa3),
	.w5(32'hba68d924),
	.w6(32'hbbc4d077),
	.w7(32'hb99d5aec),
	.w8(32'h3914adc9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a1c35),
	.w1(32'h3ade518d),
	.w2(32'h3a3f30df),
	.w3(32'hbb03a9ba),
	.w4(32'hbbd77c1b),
	.w5(32'h3a0f7c97),
	.w6(32'hbac7b44f),
	.w7(32'hba76cca7),
	.w8(32'hbaede68f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5389df),
	.w1(32'hbb85e1e9),
	.w2(32'hba0b20f5),
	.w3(32'h3a7471c0),
	.w4(32'hbac4ed17),
	.w5(32'hbbdb285b),
	.w6(32'hbb008230),
	.w7(32'h3a473e78),
	.w8(32'hbc02ae88),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5de224),
	.w1(32'hbacf5ed2),
	.w2(32'h398a1591),
	.w3(32'hbb2fe450),
	.w4(32'hbc9abac5),
	.w5(32'hbbaee7ae),
	.w6(32'h3c6c205e),
	.w7(32'hbbaa2086),
	.w8(32'hbbef2c28),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec413b),
	.w1(32'hbb0118a3),
	.w2(32'h3b0ac63c),
	.w3(32'h3ac024c5),
	.w4(32'h3bc33374),
	.w5(32'hb8c79677),
	.w6(32'hba867d68),
	.w7(32'h3c023f14),
	.w8(32'h3a7853c4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc0120),
	.w1(32'hba1fdfde),
	.w2(32'hb9359333),
	.w3(32'hbab9b33c),
	.w4(32'h3af2c215),
	.w5(32'hbc63a5b2),
	.w6(32'hbae85a28),
	.w7(32'hbb0f4205),
	.w8(32'hbc41b241),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b0557),
	.w1(32'hbc1ea929),
	.w2(32'h3c83af06),
	.w3(32'hbc0a62e1),
	.w4(32'h3cd257c6),
	.w5(32'hbb640826),
	.w6(32'hbc9401b5),
	.w7(32'h3c7dcaff),
	.w8(32'h3b3f7594),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba36841),
	.w1(32'hbb48448a),
	.w2(32'hbbb31c93),
	.w3(32'h3bb6b1b2),
	.w4(32'hbba283a0),
	.w5(32'hbb8ee729),
	.w6(32'h3b561d00),
	.w7(32'hbbb3d552),
	.w8(32'hbb45a0a6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43b141),
	.w1(32'hbc279c0a),
	.w2(32'hbc43971a),
	.w3(32'hbc128d7c),
	.w4(32'hbbb90843),
	.w5(32'hbabb48af),
	.w6(32'hbc1b22aa),
	.w7(32'hbc38550d),
	.w8(32'hbb60ed2a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82e75ea),
	.w1(32'h3b3e10a9),
	.w2(32'h3a84c24e),
	.w3(32'h3a5deb66),
	.w4(32'hbacbed2d),
	.w5(32'hbabcf50f),
	.w6(32'hbb421ae0),
	.w7(32'h3b334ea2),
	.w8(32'hbb62e32b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb166483),
	.w1(32'h3b460fe0),
	.w2(32'hba388103),
	.w3(32'h39b0a5e9),
	.w4(32'hba750153),
	.w5(32'hbb19c8b4),
	.w6(32'h3a967b35),
	.w7(32'hba939f6f),
	.w8(32'hbb8a9cc8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4c738),
	.w1(32'hbab9d29f),
	.w2(32'hbb5062b7),
	.w3(32'hbb7f242e),
	.w4(32'hba51cc43),
	.w5(32'hbb90d996),
	.w6(32'hbb4e9cbb),
	.w7(32'hbb46248d),
	.w8(32'hbc2bc6d3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6eaf47),
	.w1(32'hbc8667c7),
	.w2(32'hbc3f0671),
	.w3(32'hbca506f0),
	.w4(32'hbc64bedb),
	.w5(32'h3a2536fd),
	.w6(32'hbc515c34),
	.w7(32'hbcc62ae9),
	.w8(32'h3b927c55),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea233a),
	.w1(32'h3a89e359),
	.w2(32'h3bd3a033),
	.w3(32'h3bdf79ca),
	.w4(32'h3bb2cbad),
	.w5(32'h3ba8da24),
	.w6(32'h3bc2d1d8),
	.w7(32'h3be20a55),
	.w8(32'h3ad3bfea),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc933b),
	.w1(32'hbb2f89df),
	.w2(32'hbb55db51),
	.w3(32'h3a252544),
	.w4(32'hbba03208),
	.w5(32'hbaa8ce4f),
	.w6(32'h3a2137da),
	.w7(32'hbbf3f0e1),
	.w8(32'h3c1e1135),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96467b),
	.w1(32'h3be4a5a5),
	.w2(32'h3b313c22),
	.w3(32'hbb9eadde),
	.w4(32'hbb6ca75c),
	.w5(32'h3bf452f1),
	.w6(32'hbb331b4b),
	.w7(32'hbb1798dc),
	.w8(32'h3a2786a9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3b14e),
	.w1(32'h3add98ae),
	.w2(32'hba6642d3),
	.w3(32'hb8830fb8),
	.w4(32'h3b5db7b8),
	.w5(32'h3a9ccd29),
	.w6(32'h3a8b988c),
	.w7(32'h3b8f4bf4),
	.w8(32'hba1a7c38),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f15a3),
	.w1(32'hb9b1eeaf),
	.w2(32'hbb924501),
	.w3(32'hbbd74527),
	.w4(32'hbc22d993),
	.w5(32'hbbc51509),
	.w6(32'hbbbf761b),
	.w7(32'hbbf89a49),
	.w8(32'h3a911e64),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4509d9),
	.w1(32'h3b02cddf),
	.w2(32'h3b728ce4),
	.w3(32'h3c1e048d),
	.w4(32'h3cc7ce60),
	.w5(32'hbaff2c78),
	.w6(32'h3b5d978d),
	.w7(32'h3cd0d945),
	.w8(32'h3babffe8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad89a7e),
	.w1(32'hbb88b2e4),
	.w2(32'hbb64846e),
	.w3(32'hbace105c),
	.w4(32'h3b0d2c21),
	.w5(32'hbb211158),
	.w6(32'hbb3cd6b3),
	.w7(32'h3b870d44),
	.w8(32'hbb839f99),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6e45c),
	.w1(32'h3b6192d5),
	.w2(32'hbbce0e78),
	.w3(32'h3b97948d),
	.w4(32'h3c2e5904),
	.w5(32'h3a61fbcc),
	.w6(32'h3983cd92),
	.w7(32'h3bd6d61a),
	.w8(32'hbada4967),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10e9a9),
	.w1(32'hbb5b0869),
	.w2(32'hbaf0de5d),
	.w3(32'h3ac36a51),
	.w4(32'hbbbb821b),
	.w5(32'hba53f6d1),
	.w6(32'h3a18d491),
	.w7(32'hbae6606c),
	.w8(32'hbb92f292),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48ca6c),
	.w1(32'hbae12774),
	.w2(32'hbc02d841),
	.w3(32'hbad2a713),
	.w4(32'hbc1f6625),
	.w5(32'hbbdc9d4f),
	.w6(32'hbb97a158),
	.w7(32'hbc03addd),
	.w8(32'hbc00b440),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec929d),
	.w1(32'hbb6701fa),
	.w2(32'hbb99fb7c),
	.w3(32'hbb421c1b),
	.w4(32'h3bbbce8d),
	.w5(32'hbb133eec),
	.w6(32'hbbd8574c),
	.w7(32'hbbe18c0d),
	.w8(32'hbb28bf31),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ef8e4),
	.w1(32'hba1f84fd),
	.w2(32'hbc113bff),
	.w3(32'hbbf812de),
	.w4(32'hbc4a0b87),
	.w5(32'hbb2e5ba8),
	.w6(32'h3ae8138d),
	.w7(32'hbc3c3e89),
	.w8(32'hbba28c83),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b0643),
	.w1(32'hb9b147f6),
	.w2(32'hbaba2582),
	.w3(32'hb9d6faad),
	.w4(32'hbbc59bfc),
	.w5(32'h3ac107a5),
	.w6(32'hbb3f1a6c),
	.w7(32'hba8a9765),
	.w8(32'h3b0e8e0d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad125de),
	.w1(32'hbaeee2b2),
	.w2(32'hba2e49b1),
	.w3(32'hb837a04c),
	.w4(32'hbbf7d1d7),
	.w5(32'hbb52ff90),
	.w6(32'h3a9d6740),
	.w7(32'hba8a138e),
	.w8(32'hbb6907a1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71972a),
	.w1(32'h3b226872),
	.w2(32'h3af2de4d),
	.w3(32'hbb20ee59),
	.w4(32'hba5c26f2),
	.w5(32'hbb119fa2),
	.w6(32'hbb12fa5b),
	.w7(32'hbab59e37),
	.w8(32'hbba51184),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e0ed5),
	.w1(32'hbab44715),
	.w2(32'h3ac1389d),
	.w3(32'hbb13556e),
	.w4(32'h3ae545d1),
	.w5(32'h3b74b177),
	.w6(32'hbb8f682c),
	.w7(32'h3b89c38e),
	.w8(32'h3b8418c8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4efb2),
	.w1(32'hb9a27881),
	.w2(32'h3aec87d7),
	.w3(32'h39ba96af),
	.w4(32'hbb1cbb0a),
	.w5(32'h3b2d9c26),
	.w6(32'hba6aa89f),
	.w7(32'hbb45cc29),
	.w8(32'h3a917e28),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47ea13),
	.w1(32'h3bf935ae),
	.w2(32'h3ae5b925),
	.w3(32'h3ba3e1e2),
	.w4(32'hbacda167),
	.w5(32'h39dfd745),
	.w6(32'h3b62badb),
	.w7(32'hb9931ff3),
	.w8(32'h3a656cd4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1dbb6),
	.w1(32'h3b576483),
	.w2(32'hbb900393),
	.w3(32'h3adbd325),
	.w4(32'hbb02eac6),
	.w5(32'h39d49910),
	.w6(32'h3935fbf8),
	.w7(32'hbba81ef1),
	.w8(32'hbb0e97ef),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb7d9),
	.w1(32'hbb4a9bc1),
	.w2(32'hb9fe9bd1),
	.w3(32'hbb46a4c9),
	.w4(32'hbb911015),
	.w5(32'hba04b654),
	.w6(32'hbbb3d774),
	.w7(32'h3b2a0ad3),
	.w8(32'hbb351d5a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba639f55),
	.w1(32'h3b8f15a3),
	.w2(32'hbb7cdfd1),
	.w3(32'h3ad74dd7),
	.w4(32'hbb003a24),
	.w5(32'hba81d3f7),
	.w6(32'h3acca4a8),
	.w7(32'hbbdc0419),
	.w8(32'hbc840729),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc1fcd),
	.w1(32'h3bf39387),
	.w2(32'h3b7128ee),
	.w3(32'h3c09c3bb),
	.w4(32'h3b4ad89d),
	.w5(32'hbb0f2756),
	.w6(32'h3b8f2e37),
	.w7(32'h3bafdfa2),
	.w8(32'h3b266d31),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec1ad5),
	.w1(32'h3b35f4d6),
	.w2(32'h3a1f727c),
	.w3(32'h3ab214b5),
	.w4(32'hba0e3e40),
	.w5(32'h3aebefad),
	.w6(32'h3a11c8d6),
	.w7(32'h3aab614a),
	.w8(32'hbad47a72),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47ded7),
	.w1(32'hbc8d33d1),
	.w2(32'hbb9ebd41),
	.w3(32'hbca7c734),
	.w4(32'hbc8de162),
	.w5(32'hbb2b2a7b),
	.w6(32'hbc986e88),
	.w7(32'hbc7a029d),
	.w8(32'h3a496973),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95cae8),
	.w1(32'h3b26d7b4),
	.w2(32'h3bacf596),
	.w3(32'hbb86d686),
	.w4(32'h3c090fdb),
	.w5(32'hbb824691),
	.w6(32'hba2ef8fe),
	.w7(32'h3b8570fd),
	.w8(32'h3c00f348),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e0ea1),
	.w1(32'h3c83299e),
	.w2(32'h3c33bfac),
	.w3(32'h3babfb30),
	.w4(32'hbb8abb7b),
	.w5(32'hbc025000),
	.w6(32'h3c8e2fc0),
	.w7(32'h3c6f575b),
	.w8(32'hbb1520a2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9643d),
	.w1(32'h3c11cca5),
	.w2(32'h3b508368),
	.w3(32'hbb415e21),
	.w4(32'hbc4de858),
	.w5(32'hbb7cd72a),
	.w6(32'h3c8a2dc7),
	.w7(32'h3ae11359),
	.w8(32'hba17a14d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983f3ed),
	.w1(32'h3a4fdbb7),
	.w2(32'hbc34b2f2),
	.w3(32'hbbc953ae),
	.w4(32'hbc4afde4),
	.w5(32'hbb82d492),
	.w6(32'h3a82f315),
	.w7(32'hbc66eb8f),
	.w8(32'hbb157d8c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c3c0),
	.w1(32'hbb75834e),
	.w2(32'h3b2d5a2b),
	.w3(32'hbb81efa0),
	.w4(32'h3bcfd5c1),
	.w5(32'hba4cfeb6),
	.w6(32'h3b84f8f7),
	.w7(32'h3bd2e873),
	.w8(32'hbb563a52),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba812ec6),
	.w1(32'h3b066a16),
	.w2(32'hbb928e93),
	.w3(32'h39dff8de),
	.w4(32'hbb97ca9a),
	.w5(32'hb8cb0505),
	.w6(32'h38738769),
	.w7(32'hbc024c5c),
	.w8(32'hbbb1aed1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49788d),
	.w1(32'hbbe97654),
	.w2(32'h38f03382),
	.w3(32'hbb2e1732),
	.w4(32'hbc1e7db5),
	.w5(32'hb951a6c8),
	.w6(32'hbb8177e3),
	.w7(32'h3b3c72cd),
	.w8(32'hba5ad723),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f82f2),
	.w1(32'h3a075c87),
	.w2(32'hbb32e225),
	.w3(32'hba4d647d),
	.w4(32'hbb883e96),
	.w5(32'hbaf5ccc5),
	.w6(32'hba6bb65f),
	.w7(32'hbb415c49),
	.w8(32'hbbd517c7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba29a0a),
	.w1(32'hbb39d444),
	.w2(32'hbb9a16ae),
	.w3(32'h3ac54f55),
	.w4(32'hbb052207),
	.w5(32'hbbed75d9),
	.w6(32'hbb7da54b),
	.w7(32'hbaf4b389),
	.w8(32'hbb61f97f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc004d4b),
	.w1(32'h3bd529b3),
	.w2(32'h3c0c91c0),
	.w3(32'h3c60a31c),
	.w4(32'h3cafc292),
	.w5(32'hbc2527dc),
	.w6(32'h3bba07ea),
	.w7(32'h3cda0ad6),
	.w8(32'hbc0f2cec),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25a495),
	.w1(32'h3bbe63af),
	.w2(32'hbb23c102),
	.w3(32'h3ba96cd5),
	.w4(32'h3a287dd1),
	.w5(32'h3bfa2546),
	.w6(32'h3bd239a5),
	.w7(32'h3b865cf6),
	.w8(32'h3cd54a1a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9675c8),
	.w1(32'h3cec4340),
	.w2(32'h3c5fcaf2),
	.w3(32'h3ce33f68),
	.w4(32'h3cfc692e),
	.w5(32'hbbb024cd),
	.w6(32'h3ca28cb0),
	.w7(32'h3d11ea62),
	.w8(32'h3ba9b547),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb65dc8),
	.w1(32'h3bcb162d),
	.w2(32'h3c305bfd),
	.w3(32'hbbf7a0cc),
	.w4(32'hbc4977eb),
	.w5(32'hbb9d0ce3),
	.w6(32'hb98010fc),
	.w7(32'h3c026f21),
	.w8(32'hbbc80da0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cd708),
	.w1(32'hba670c8b),
	.w2(32'hba85a012),
	.w3(32'hba5b8ed9),
	.w4(32'h3b2df0d5),
	.w5(32'hb8e659e7),
	.w6(32'hba912662),
	.w7(32'hbb0c6b0b),
	.w8(32'hbaa0f32d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba705cf6),
	.w1(32'hba9ed3df),
	.w2(32'h3b816848),
	.w3(32'hbb302337),
	.w4(32'h3bb40044),
	.w5(32'h3ba8e388),
	.w6(32'hbada138a),
	.w7(32'h3b41fad1),
	.w8(32'h3cbfc0b1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c859ffa),
	.w1(32'h3c978d38),
	.w2(32'hbc4e50e8),
	.w3(32'h3c4f4764),
	.w4(32'h3ab15362),
	.w5(32'h3b9a4d79),
	.w6(32'h3c86404c),
	.w7(32'hbba13cf9),
	.w8(32'h3a6e73e3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68aca4),
	.w1(32'h3b62c79c),
	.w2(32'hbb0b07c7),
	.w3(32'hbb3093f6),
	.w4(32'hbba07a3b),
	.w5(32'hba0d3ce3),
	.w6(32'hbbe2ca6b),
	.w7(32'hbba84ad2),
	.w8(32'hbb3835e6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bf0dc),
	.w1(32'hbadd4b7a),
	.w2(32'hbb2a4788),
	.w3(32'hbb44af62),
	.w4(32'h393f527d),
	.w5(32'h3ad709b3),
	.w6(32'hbb8608ae),
	.w7(32'hbb136322),
	.w8(32'hba8bc9d2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb584a7f),
	.w1(32'hba5f0c24),
	.w2(32'h38e52284),
	.w3(32'hb98d4f0d),
	.w4(32'hba8c468e),
	.w5(32'h3b047d02),
	.w6(32'hbb3ea16a),
	.w7(32'hbb2b30c7),
	.w8(32'h3a9d046b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb893c98),
	.w1(32'hbb1325e8),
	.w2(32'hbb820b2b),
	.w3(32'hbb085294),
	.w4(32'hbba40c9e),
	.w5(32'hbadbf317),
	.w6(32'hbb229c7a),
	.w7(32'hbba8b737),
	.w8(32'hbb90bbee),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb462e08),
	.w1(32'h3acb2185),
	.w2(32'h3b481e73),
	.w3(32'h3bc47b7d),
	.w4(32'h3bc6e73a),
	.w5(32'hbb667e65),
	.w6(32'h39d96383),
	.w7(32'h3c2c3c18),
	.w8(32'hbb9642e0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacbfdb),
	.w1(32'hbbd29b4c),
	.w2(32'h38199dd5),
	.w3(32'hbb4b2ea1),
	.w4(32'h3a54d540),
	.w5(32'hba0f4942),
	.w6(32'hbb873fc2),
	.w7(32'hbb3ce018),
	.w8(32'hb988d75f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fa275),
	.w1(32'hb91a55fe),
	.w2(32'h3a902eda),
	.w3(32'h3871ae2d),
	.w4(32'hbc0629af),
	.w5(32'hbc35ca83),
	.w6(32'h3b084950),
	.w7(32'hbb164dc8),
	.w8(32'hbc0fa312),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0121f5),
	.w1(32'hbbc10666),
	.w2(32'hbc2221c6),
	.w3(32'hbb9cc34e),
	.w4(32'hbc22b422),
	.w5(32'h3b84979d),
	.w6(32'hbbb2b675),
	.w7(32'hbc5f5647),
	.w8(32'h3b3ba507),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f6158),
	.w1(32'h3b23eedb),
	.w2(32'hbaac0ab5),
	.w3(32'hba5c8196),
	.w4(32'hbb99c1e3),
	.w5(32'hba86387c),
	.w6(32'h3b336d7c),
	.w7(32'hbc0e7b02),
	.w8(32'h3b1a9d95),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be317c1),
	.w1(32'hbb3ac7c2),
	.w2(32'h3a4de312),
	.w3(32'hbb801c04),
	.w4(32'hbb1046f4),
	.w5(32'hbb818f07),
	.w6(32'hbb85f0d9),
	.w7(32'hbb63d8dd),
	.w8(32'hbbcae972),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdba7e2),
	.w1(32'hba9db85e),
	.w2(32'hb9f87084),
	.w3(32'hbac26120),
	.w4(32'h3b8c2705),
	.w5(32'hbb54536b),
	.w6(32'hbb42d459),
	.w7(32'hba795f80),
	.w8(32'hba957803),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15f2cd),
	.w1(32'hbb6489ef),
	.w2(32'hbab00b25),
	.w3(32'hba63c4aa),
	.w4(32'h3a9b1732),
	.w5(32'h3a5d725f),
	.w6(32'h3aa5a94d),
	.w7(32'hba24fe98),
	.w8(32'hbaee66bb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfa472),
	.w1(32'hbaa8f3f3),
	.w2(32'hbb3f0720),
	.w3(32'hb985dac4),
	.w4(32'hbc2241b8),
	.w5(32'h3c9e3772),
	.w6(32'hb933da91),
	.w7(32'hbba3a271),
	.w8(32'h3cf9afff),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a32cf),
	.w1(32'h3b9e7f39),
	.w2(32'h3c035868),
	.w3(32'h3cbc3156),
	.w4(32'h3d0473a2),
	.w5(32'h3b912d72),
	.w6(32'h3c95166a),
	.w7(32'h3c5e3bfb),
	.w8(32'h3a96d642),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac41f63),
	.w1(32'h3b3911a5),
	.w2(32'h3bbd49c0),
	.w3(32'h3ad975c8),
	.w4(32'h3bac7b90),
	.w5(32'h3c281cd2),
	.w6(32'hbaf9ac2c),
	.w7(32'h3b4e275f),
	.w8(32'h3c25c453),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62ffe1),
	.w1(32'hbb04eea5),
	.w2(32'h3c9b3a80),
	.w3(32'h3b6b663e),
	.w4(32'h3d05e834),
	.w5(32'hbb68a199),
	.w6(32'hbb10cee5),
	.w7(32'h3c56afb6),
	.w8(32'hb8a164cd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef8bcb),
	.w1(32'hbb938f2c),
	.w2(32'hbb865095),
	.w3(32'hbbbf540d),
	.w4(32'hbc169e5a),
	.w5(32'h3b046e95),
	.w6(32'hbae3fb3e),
	.w7(32'hbbe4e49e),
	.w8(32'hba40cc9f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b522c24),
	.w1(32'hba0f57d2),
	.w2(32'hbb7a8f52),
	.w3(32'h3b3eafc4),
	.w4(32'hbb6b5eb0),
	.w5(32'hbc2268c9),
	.w6(32'h3b1a3b71),
	.w7(32'hbba27945),
	.w8(32'hbc84b42b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc390a7),
	.w1(32'hbbbc576a),
	.w2(32'h3b7df3f8),
	.w3(32'hbc3cef8e),
	.w4(32'hbca16b9c),
	.w5(32'hbb2846d7),
	.w6(32'hbb627586),
	.w7(32'hbc203e07),
	.w8(32'hbacf4736),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e5f78),
	.w1(32'hba98f0f1),
	.w2(32'hb8b25f04),
	.w3(32'hba66040a),
	.w4(32'h3b3a10b9),
	.w5(32'h3a03eafd),
	.w6(32'hbaeb575f),
	.w7(32'hb9db67c3),
	.w8(32'h3b7cee41),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74b5c6),
	.w1(32'h3b9898f9),
	.w2(32'h3b477b6b),
	.w3(32'hbb1dff37),
	.w4(32'hbc1cecb0),
	.w5(32'h3b1ec9c5),
	.w6(32'h3b73d1ae),
	.w7(32'hbbcdee1f),
	.w8(32'h3b3ed00f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4c9da),
	.w1(32'hbba2f944),
	.w2(32'hba8ed334),
	.w3(32'hbac7a192),
	.w4(32'hbaad4bac),
	.w5(32'hbb46b6e2),
	.w6(32'hbb928d27),
	.w7(32'hbbbc63db),
	.w8(32'h3a550c3c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17e69d),
	.w1(32'h3bc4d6d1),
	.w2(32'h3b313f4d),
	.w3(32'h39d297f1),
	.w4(32'hbc0a2c0f),
	.w5(32'hbb9fa761),
	.w6(32'h3c5af7d0),
	.w7(32'h3a751bad),
	.w8(32'hbc4bcc7b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9671e2),
	.w1(32'h3704fc3c),
	.w2(32'hbbf4a482),
	.w3(32'h39cad559),
	.w4(32'hbbf7f44c),
	.w5(32'hbb2520dc),
	.w6(32'hb9a34684),
	.w7(32'hbc48f87a),
	.w8(32'hbb968773),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74cfc7),
	.w1(32'h3a47b7c4),
	.w2(32'h3c0c92d8),
	.w3(32'h3aba7900),
	.w4(32'h3c608d7a),
	.w5(32'h39a7b246),
	.w6(32'hba33f69e),
	.w7(32'h3c29e240),
	.w8(32'hba2c57f5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56930c),
	.w1(32'h3ab1e8e6),
	.w2(32'hbb033ec1),
	.w3(32'h3aec0bdb),
	.w4(32'hbbb7a09f),
	.w5(32'h3b898de7),
	.w6(32'h3b09ed63),
	.w7(32'hbb18d43f),
	.w8(32'hba8d1312),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b896b1),
	.w1(32'hbbc6ae45),
	.w2(32'hbb82b333),
	.w3(32'hba405602),
	.w4(32'hbbd742ab),
	.w5(32'hb8a644c2),
	.w6(32'hbb978401),
	.w7(32'hbc04c551),
	.w8(32'hb724821f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a878ab5),
	.w1(32'h3b11540d),
	.w2(32'hbb27840a),
	.w3(32'h3b3007ef),
	.w4(32'h3a7f6c8f),
	.w5(32'h3ae53128),
	.w6(32'h3b0fd4a0),
	.w7(32'hbb9f8563),
	.w8(32'hba1724d5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d5a0d),
	.w1(32'h3b369447),
	.w2(32'hbbf8555d),
	.w3(32'hbbb2e1f8),
	.w4(32'hbc3bc4d9),
	.w5(32'h3a8f29b0),
	.w6(32'h3ab27b67),
	.w7(32'hbc517cc1),
	.w8(32'h381f9d30),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a517d59),
	.w1(32'h3b281bba),
	.w2(32'h3b17205e),
	.w3(32'h3abfeea7),
	.w4(32'h3af6ff61),
	.w5(32'hba7c0cb0),
	.w6(32'h3b806b3a),
	.w7(32'h3a94a609),
	.w8(32'hbb2dd2a8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81a001),
	.w1(32'hba0f2bd9),
	.w2(32'hbb0824f5),
	.w3(32'h3a2fe5d0),
	.w4(32'h393828e3),
	.w5(32'hbabff389),
	.w6(32'h3c13cc9b),
	.w7(32'hbaa41fad),
	.w8(32'hb9b71588),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5de2d),
	.w1(32'h3bb4ef20),
	.w2(32'h3b294b69),
	.w3(32'h3a7fa5e9),
	.w4(32'hbb049167),
	.w5(32'hb9a72bf8),
	.w6(32'h39a4f7f5),
	.w7(32'hba3a072e),
	.w8(32'hbb8bd21c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a385c28),
	.w1(32'hbaaae315),
	.w2(32'h3a346c66),
	.w3(32'h3942fc80),
	.w4(32'h3b02d055),
	.w5(32'h3af3cb59),
	.w6(32'hbb36c40b),
	.w7(32'hbb03ff29),
	.w8(32'h3ac4267d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aa022),
	.w1(32'hba104191),
	.w2(32'h3b0be273),
	.w3(32'h3903f170),
	.w4(32'h3b02f4c8),
	.w5(32'hbad7c3e8),
	.w6(32'hba821a07),
	.w7(32'h3b178f66),
	.w8(32'h3b1add5f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dfdb1),
	.w1(32'h3a92c412),
	.w2(32'hba1ac7ca),
	.w3(32'hba829301),
	.w4(32'hba6ab3a0),
	.w5(32'hbb823716),
	.w6(32'h3c3ef6be),
	.w7(32'h3bcc2c6d),
	.w8(32'hbb253528),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21d231),
	.w1(32'h3b093014),
	.w2(32'h3aae1c86),
	.w3(32'hbb02e8c4),
	.w4(32'hbb1403ef),
	.w5(32'hbadc1e4a),
	.w6(32'hbbbadeed),
	.w7(32'hbbc42739),
	.w8(32'hbb415f63),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03d377),
	.w1(32'hb9117b6f),
	.w2(32'hba4a6fdf),
	.w3(32'hbab630f7),
	.w4(32'hbb3d5f06),
	.w5(32'h3bb5be6f),
	.w6(32'h3a26ad38),
	.w7(32'hbadfb6a7),
	.w8(32'hb9eaf534),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd841d),
	.w1(32'h3c08257e),
	.w2(32'h3b2e2a83),
	.w3(32'h3a1e6e3e),
	.w4(32'h3b8783ab),
	.w5(32'h39ebb5bc),
	.w6(32'h3b17939a),
	.w7(32'h3ba8e62a),
	.w8(32'h3a6e9f94),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62c25fd),
	.w1(32'h3a1195d3),
	.w2(32'h3ac80fa0),
	.w3(32'hb995d637),
	.w4(32'h3a947edd),
	.w5(32'h3b1a2f19),
	.w6(32'hb888f58e),
	.w7(32'h3a866963),
	.w8(32'h3b07da17),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b106293),
	.w1(32'h3b87545e),
	.w2(32'h3b867903),
	.w3(32'h3b86106f),
	.w4(32'h3b9e279d),
	.w5(32'hba8c8057),
	.w6(32'h3bc7ea13),
	.w7(32'h3b8950a4),
	.w8(32'hbaf46c01),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985c0ef),
	.w1(32'h3a66457b),
	.w2(32'h3a550d77),
	.w3(32'hb9a37e0b),
	.w4(32'hba4914b0),
	.w5(32'h3b6795ed),
	.w6(32'hba726160),
	.w7(32'hb97834df),
	.w8(32'hba364806),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3c5e3),
	.w1(32'h3b3783d1),
	.w2(32'hba3a0824),
	.w3(32'h3afcdb25),
	.w4(32'h3a6bec0c),
	.w5(32'h3aa9c182),
	.w6(32'hba8361fa),
	.w7(32'hbb27733e),
	.w8(32'h3a1bc007),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960c5ba),
	.w1(32'hb9f8ba4f),
	.w2(32'hb8c92540),
	.w3(32'h372bd391),
	.w4(32'h3b02b90b),
	.w5(32'h37f025a7),
	.w6(32'hba8b86eb),
	.w7(32'h3b0f0301),
	.w8(32'hbb2ec96a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bb8389),
	.w1(32'h3a0ef426),
	.w2(32'hb96bc39d),
	.w3(32'hba1f616b),
	.w4(32'hb9999905),
	.w5(32'hbade5885),
	.w6(32'hbb1997f9),
	.w7(32'hbb158a02),
	.w8(32'h378dec91),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee3f9d),
	.w1(32'h3aa40b7c),
	.w2(32'h3aeed540),
	.w3(32'hbad9bad8),
	.w4(32'hb9026983),
	.w5(32'hb8ebffe7),
	.w6(32'h3978baa9),
	.w7(32'hb8e79e38),
	.w8(32'hba37ae10),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7c89e),
	.w1(32'h3ba4ade9),
	.w2(32'h3b4774c6),
	.w3(32'h3921c9e2),
	.w4(32'h3af711b7),
	.w5(32'h3b19ab2f),
	.w6(32'h3b3b45aa),
	.w7(32'hbb5a4848),
	.w8(32'hb9a109c5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a637096),
	.w1(32'hbb1ff13a),
	.w2(32'hbafc9748),
	.w3(32'hb9623e52),
	.w4(32'h3abc5349),
	.w5(32'hba73241f),
	.w6(32'hba72a205),
	.w7(32'h3a77cfc2),
	.w8(32'h396c34fd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f1883e),
	.w1(32'hbaa4021c),
	.w2(32'hb83c25d4),
	.w3(32'hbaba1f2a),
	.w4(32'hb934bca7),
	.w5(32'hb9b25b72),
	.w6(32'hba8d03cb),
	.w7(32'h39c2d646),
	.w8(32'h3b5bf62f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a653364),
	.w1(32'h398c64ce),
	.w2(32'h3b210c2c),
	.w3(32'h3acb46f5),
	.w4(32'hbb07736d),
	.w5(32'hba3bd3dd),
	.w6(32'h3c004546),
	.w7(32'h3aa9592c),
	.w8(32'hbb74df5e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c9f0e),
	.w1(32'hba12f83c),
	.w2(32'h39f8945c),
	.w3(32'h3adfe31b),
	.w4(32'h3a1ac0ee),
	.w5(32'h3ae07884),
	.w6(32'h3998880e),
	.w7(32'h3a1b89b4),
	.w8(32'h3ad076cf),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d42eb),
	.w1(32'h3b00982c),
	.w2(32'h3a6eac77),
	.w3(32'h3b4e98de),
	.w4(32'h3b830992),
	.w5(32'h3a530775),
	.w6(32'h3b76ec14),
	.w7(32'h3b065036),
	.w8(32'h3b02e281),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7fc04),
	.w1(32'h3a8afac7),
	.w2(32'h3abb657f),
	.w3(32'h39a67f81),
	.w4(32'h3ae26354),
	.w5(32'h3993015b),
	.w6(32'h39de199a),
	.w7(32'h3b170f4e),
	.w8(32'h3a91a86f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f70b9),
	.w1(32'h3a10a4d7),
	.w2(32'h3a697a3f),
	.w3(32'h3a4f6b6a),
	.w4(32'h3a8eb19c),
	.w5(32'h3ba7f3d6),
	.w6(32'hba8ac7b6),
	.w7(32'hba4ea342),
	.w8(32'h3a8970cc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6befea),
	.w1(32'h3b3ae85d),
	.w2(32'h3b180b98),
	.w3(32'h3b87a000),
	.w4(32'h3b4b54a3),
	.w5(32'h3aa0fac6),
	.w6(32'h3b4ef93d),
	.w7(32'h3a28c091),
	.w8(32'h3aa6eac4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d574e),
	.w1(32'hb752b6e1),
	.w2(32'hb93f7d23),
	.w3(32'h399a342d),
	.w4(32'hb9590319),
	.w5(32'h3b1f9af2),
	.w6(32'h3a086489),
	.w7(32'hb90a4761),
	.w8(32'h3b36aa93),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadafb2c),
	.w1(32'hba7a1b36),
	.w2(32'hb9ded936),
	.w3(32'h3b213815),
	.w4(32'h3aa11c38),
	.w5(32'hb9f37589),
	.w6(32'h3b33dc98),
	.w7(32'h3b15cde2),
	.w8(32'hb9b3676e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23b95f),
	.w1(32'hba75901d),
	.w2(32'h3a41441a),
	.w3(32'hbafe143e),
	.w4(32'hbb37c9eb),
	.w5(32'hb9f50aec),
	.w6(32'hba690867),
	.w7(32'hb9a403b9),
	.w8(32'hb981a2a2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e836d),
	.w1(32'h3a059822),
	.w2(32'h3a99de01),
	.w3(32'hba29e1bb),
	.w4(32'h39793707),
	.w5(32'hbad1fd0f),
	.w6(32'h3a84bb3e),
	.w7(32'h3a9587ad),
	.w8(32'h3b34561a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b808569),
	.w1(32'h3ba660b5),
	.w2(32'h3b89df50),
	.w3(32'h3a57606d),
	.w4(32'h3a5e3ccf),
	.w5(32'hbb063748),
	.w6(32'hb9ad742e),
	.w7(32'hb96c8b14),
	.w8(32'hbb5b68cd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0096de),
	.w1(32'hbad70702),
	.w2(32'h3a2613a1),
	.w3(32'hbaf45679),
	.w4(32'hba1c4f58),
	.w5(32'h39de814e),
	.w6(32'hbb69c28f),
	.w7(32'h392402f0),
	.w8(32'hb9392614),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e411d),
	.w1(32'h3a515e57),
	.w2(32'h3abdcc5f),
	.w3(32'hb93dea80),
	.w4(32'h391bb1b2),
	.w5(32'h3b3ea8f5),
	.w6(32'hba939505),
	.w7(32'hba0bb5b8),
	.w8(32'hba43b056),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912352e),
	.w1(32'hbaf1576d),
	.w2(32'hbb022ccc),
	.w3(32'h3b2771fa),
	.w4(32'h3abfba63),
	.w5(32'h3a44dbd3),
	.w6(32'hbb79e1dc),
	.w7(32'hbb5f842e),
	.w8(32'hb893baad),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9443a84),
	.w1(32'h39b1c7e7),
	.w2(32'hb893040e),
	.w3(32'h39382b56),
	.w4(32'hb9947600),
	.w5(32'h3be26397),
	.w6(32'h3a2d039c),
	.w7(32'hba0b42a6),
	.w8(32'h3b23066c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9855f1),
	.w1(32'h3b7072e5),
	.w2(32'h3be2a100),
	.w3(32'h3b76d2ed),
	.w4(32'h3bcba934),
	.w5(32'hba4bb79c),
	.w6(32'h3ab44986),
	.w7(32'h3b18480b),
	.w8(32'hbb0155c7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec7d0d),
	.w1(32'hb87d1ae3),
	.w2(32'h3a1a6281),
	.w3(32'hba32e4b6),
	.w4(32'hb987cf5b),
	.w5(32'hb9f0044a),
	.w6(32'hba148d62),
	.w7(32'hb96feef0),
	.w8(32'hb8ca42a4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a579d56),
	.w1(32'h39d2bcb9),
	.w2(32'h3aa8ec7a),
	.w3(32'hb9d870e8),
	.w4(32'h3a5cd8de),
	.w5(32'hba90d5a8),
	.w6(32'hb887c3ad),
	.w7(32'h39a5a36a),
	.w8(32'hbb06bb3d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1eada),
	.w1(32'h3a6629f5),
	.w2(32'h3a21d806),
	.w3(32'hba48c095),
	.w4(32'h3aa0df47),
	.w5(32'hbabfa0d8),
	.w6(32'h39ea4414),
	.w7(32'h3a1ed308),
	.w8(32'hbb226e9c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0b92b),
	.w1(32'hb7c80153),
	.w2(32'h397615fb),
	.w3(32'hba51a00d),
	.w4(32'hb891eea1),
	.w5(32'h3a4e5184),
	.w6(32'hbb0e3313),
	.w7(32'hba77c7c2),
	.w8(32'hbaab5055),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8e8ed),
	.w1(32'h39e71cb6),
	.w2(32'h3a867e23),
	.w3(32'h39037d22),
	.w4(32'hb910a1d5),
	.w5(32'h3a680df5),
	.w6(32'hb7ab4bb4),
	.w7(32'hb954ce63),
	.w8(32'hb971dd98),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a6d25),
	.w1(32'hb7b9fd8e),
	.w2(32'h39fdab20),
	.w3(32'h3a0b2e72),
	.w4(32'h3a30c125),
	.w5(32'h3a034778),
	.w6(32'h3a86ce14),
	.w7(32'hb8a2cd7b),
	.w8(32'h39a8f714),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b9c94),
	.w1(32'h3bea0615),
	.w2(32'h3b3b06bf),
	.w3(32'h3b03d942),
	.w4(32'h3b444b6e),
	.w5(32'hba091a54),
	.w6(32'h39ef8938),
	.w7(32'h3a5f2c38),
	.w8(32'hba176959),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f294b),
	.w1(32'hbaf32c31),
	.w2(32'hbad6c7f2),
	.w3(32'hbad09abf),
	.w4(32'hb90ae6ca),
	.w5(32'h3b75f9ad),
	.w6(32'h3a9358ec),
	.w7(32'hbaa233c3),
	.w8(32'h3b7b7d66),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7d7c8),
	.w1(32'hba228f21),
	.w2(32'h3a37241c),
	.w3(32'hba82147c),
	.w4(32'h3a57c075),
	.w5(32'h3ad05795),
	.w6(32'hbb44ec5e),
	.w7(32'h39c71284),
	.w8(32'h397e2c87),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39766d47),
	.w1(32'hb902a7cb),
	.w2(32'hb990da23),
	.w3(32'h3ad1fb34),
	.w4(32'h39a323d1),
	.w5(32'h3b1d592b),
	.w6(32'h3934351f),
	.w7(32'hba382080),
	.w8(32'h3adec27c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c993b),
	.w1(32'h3b0b78a2),
	.w2(32'h3b6c7f5d),
	.w3(32'h3a7b21e1),
	.w4(32'hb833ac22),
	.w5(32'hba558840),
	.w6(32'hba25971e),
	.w7(32'hb921d0a9),
	.w8(32'hbaa99f88),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab34de3),
	.w1(32'h3a7c5d92),
	.w2(32'h3ab5c125),
	.w3(32'hba99de11),
	.w4(32'hba47015c),
	.w5(32'h3a29123b),
	.w6(32'hbacbbabe),
	.w7(32'hba4a7fed),
	.w8(32'hb9cf0f81),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383b9746),
	.w1(32'hba24ad9f),
	.w2(32'hba62ddfb),
	.w3(32'hb9507f4f),
	.w4(32'hb99be4f2),
	.w5(32'hbb4e1347),
	.w6(32'h3a72070e),
	.w7(32'hb95abc38),
	.w8(32'hbb3c9b71),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0709a),
	.w1(32'h3986d6e3),
	.w2(32'hbae0e086),
	.w3(32'hba80a367),
	.w4(32'hbb8ae9f7),
	.w5(32'h3a09cd43),
	.w6(32'h3bad8339),
	.w7(32'hba8ca4fe),
	.w8(32'h3a3ed9d8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafe11b),
	.w1(32'h3a1276db),
	.w2(32'h3baca9e1),
	.w3(32'hba18be49),
	.w4(32'hb7ff5411),
	.w5(32'h3a87def9),
	.w6(32'hb7b3f36c),
	.w7(32'h3b066d3b),
	.w8(32'h3a4f36da),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a832e17),
	.w1(32'h3a774c84),
	.w2(32'h3ac5d62a),
	.w3(32'hb403f03c),
	.w4(32'hbabb98cf),
	.w5(32'h3a2895be),
	.w6(32'hba1aac58),
	.w7(32'hba822bc9),
	.w8(32'h3aa2a38c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b0ca3),
	.w1(32'h3a03ab64),
	.w2(32'h3aa3e003),
	.w3(32'h39d0788d),
	.w4(32'h3a915dc3),
	.w5(32'hb9e5b793),
	.w6(32'h3a1ffff2),
	.w7(32'h3ab0d288),
	.w8(32'hba5c0b61),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74d7a7),
	.w1(32'h38706888),
	.w2(32'h3a7a629a),
	.w3(32'hbaf3d622),
	.w4(32'hba3c3e07),
	.w5(32'h3b739c8a),
	.w6(32'hbaff4b43),
	.w7(32'h3a02d1c1),
	.w8(32'h3b108ac7),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b918c89),
	.w1(32'h3abfa8aa),
	.w2(32'h3b3c2729),
	.w3(32'h36fbc796),
	.w4(32'h3889fb98),
	.w5(32'hba19e4e1),
	.w6(32'hba2cafc4),
	.w7(32'hbadca317),
	.w8(32'hb7eb48e2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4597ac),
	.w1(32'hbb5f24e4),
	.w2(32'hbb14245c),
	.w3(32'hbae22353),
	.w4(32'h3a083e98),
	.w5(32'h3a8859ec),
	.w6(32'h399eac2d),
	.w7(32'hba878db1),
	.w8(32'h39c475eb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a20d3f),
	.w1(32'h3b0efcd7),
	.w2(32'h3b1ff4f7),
	.w3(32'h39d96e46),
	.w4(32'hb692f8cd),
	.w5(32'h3a378c53),
	.w6(32'h3921afe9),
	.w7(32'h39d046ca),
	.w8(32'h3af1f5c5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b346edf),
	.w1(32'h3b12d44e),
	.w2(32'h3b5fd872),
	.w3(32'h3a061eb8),
	.w4(32'h3acf7c99),
	.w5(32'hbaa8ec96),
	.w6(32'hbac826c3),
	.w7(32'h390c6855),
	.w8(32'hbb27121f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa40c87),
	.w1(32'hba681655),
	.w2(32'hb9b2b4b2),
	.w3(32'hba96888e),
	.w4(32'hbac13461),
	.w5(32'hba788a42),
	.w6(32'hbb17fbe3),
	.w7(32'hba6c25dc),
	.w8(32'hba12977f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc12a9),
	.w1(32'h398be1ed),
	.w2(32'h3a82b311),
	.w3(32'hbab6297a),
	.w4(32'hbadc823a),
	.w5(32'h3abb1b05),
	.w6(32'hbb09a13d),
	.w7(32'h39cfb1c0),
	.w8(32'h3a96dcc4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceebba),
	.w1(32'h3a5c5bf3),
	.w2(32'h3b274d0b),
	.w3(32'h398df475),
	.w4(32'h3afc18a6),
	.w5(32'hba8073c1),
	.w6(32'hbb01e2aa),
	.w7(32'h39c62342),
	.w8(32'h3b8c94c4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4c0b1),
	.w1(32'hbb2ebf17),
	.w2(32'hba48d126),
	.w3(32'h3b61fd22),
	.w4(32'h3ae74124),
	.w5(32'h3b976604),
	.w6(32'h3c1af619),
	.w7(32'h3b61e30c),
	.w8(32'hba258fa3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c3fba),
	.w1(32'h3bd709ed),
	.w2(32'h3b72f381),
	.w3(32'h3b735805),
	.w4(32'h3b7becc2),
	.w5(32'hbb994e09),
	.w6(32'h3b0603a6),
	.w7(32'hbad2daaf),
	.w8(32'h3ba06d69),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8ac0),
	.w1(32'h3b1ebd2f),
	.w2(32'h3ab90b70),
	.w3(32'h3b565de4),
	.w4(32'h3a6174b7),
	.w5(32'h3af03f33),
	.w6(32'h3c50e9d0),
	.w7(32'h3c12b860),
	.w8(32'h3a779991),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39842db7),
	.w1(32'hbb34bb9a),
	.w2(32'h39ac5e38),
	.w3(32'hba23e81f),
	.w4(32'h39c83903),
	.w5(32'h3b3d9d83),
	.w6(32'h3a791a42),
	.w7(32'h3b2bd594),
	.w8(32'h3b102c7c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389de9af),
	.w1(32'h3a7d2288),
	.w2(32'h3b1f2a07),
	.w3(32'h3a6f4207),
	.w4(32'h39aacfdf),
	.w5(32'hbadca64c),
	.w6(32'h3a25848e),
	.w7(32'h3a8aac38),
	.w8(32'hbac87cc3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec384d),
	.w1(32'hbac15100),
	.w2(32'hb8fe518b),
	.w3(32'hba53dbe0),
	.w4(32'hba900229),
	.w5(32'hbb4827fd),
	.w6(32'h3b2a8157),
	.w7(32'h3a13c25d),
	.w8(32'h3c2abd3d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d34b0),
	.w1(32'h3a301961),
	.w2(32'h3b32ccbb),
	.w3(32'h3b3e0239),
	.w4(32'hbb604e85),
	.w5(32'hba4ee55a),
	.w6(32'h3c5b2722),
	.w7(32'h3c038b12),
	.w8(32'hbb3084a3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba922245),
	.w1(32'hb9bb7614),
	.w2(32'h3a2fa091),
	.w3(32'hba2ea284),
	.w4(32'h38d35a2d),
	.w5(32'hba15f878),
	.w6(32'hbb86a57c),
	.w7(32'hbb4412ee),
	.w8(32'h3b2a66e1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0d5c8),
	.w1(32'hba1f4d42),
	.w2(32'h367aca41),
	.w3(32'h395f4afa),
	.w4(32'hba558918),
	.w5(32'h3b117a52),
	.w6(32'h3b0f41b5),
	.w7(32'h3b063ab7),
	.w8(32'h3b283358),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3798a11b),
	.w1(32'h3ac5c94e),
	.w2(32'h3b65d141),
	.w3(32'h3b0b8f3b),
	.w4(32'h3b487621),
	.w5(32'h398c6224),
	.w6(32'h3b914af8),
	.w7(32'h3bacac0d),
	.w8(32'h3a1f50b9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59987e),
	.w1(32'hba83126d),
	.w2(32'hba4d2a2d),
	.w3(32'hba5e4fda),
	.w4(32'hba8310e3),
	.w5(32'h39a3a644),
	.w6(32'hbb4a66ac),
	.w7(32'hb769b740),
	.w8(32'h3a009eab),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafc358),
	.w1(32'h3ae6a1e3),
	.w2(32'h3b588da2),
	.w3(32'hb9dd613c),
	.w4(32'h3a930614),
	.w5(32'h3abbcf8a),
	.w6(32'h3a5f01a7),
	.w7(32'h3acb1c3a),
	.w8(32'hbb1e0cbd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f6ecd),
	.w1(32'h3b0afa6e),
	.w2(32'h3a1e9a58),
	.w3(32'h3b1da977),
	.w4(32'hba40f7c5),
	.w5(32'h3a7f89a0),
	.w6(32'hbb157257),
	.w7(32'hbb840699),
	.w8(32'hbb414c24),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8357e5),
	.w1(32'h38bd8e97),
	.w2(32'h3b0a30c2),
	.w3(32'h39541e00),
	.w4(32'hbb14a248),
	.w5(32'hba2baac4),
	.w6(32'hbc0d79cd),
	.w7(32'hbc1d1c7d),
	.w8(32'h3aeb7563),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4b8a2),
	.w1(32'h3b91a278),
	.w2(32'h3b8b05af),
	.w3(32'h3b646ace),
	.w4(32'h3b33e4c3),
	.w5(32'hbb0330b9),
	.w6(32'h3bc9c983),
	.w7(32'h3b155eec),
	.w8(32'hba4ddf2a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac93779),
	.w1(32'hbab1b65f),
	.w2(32'hbaf81506),
	.w3(32'hba7415c0),
	.w4(32'hbab0be01),
	.w5(32'hba2f6323),
	.w6(32'h3b3cf382),
	.w7(32'h39b1a3b0),
	.w8(32'hba4d55bd),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47c888),
	.w1(32'h3b370fe3),
	.w2(32'hba930473),
	.w3(32'h39863e04),
	.w4(32'hb922025f),
	.w5(32'hb9423f6e),
	.w6(32'h3b0418bd),
	.w7(32'h3a2a0213),
	.w8(32'hba85bc4f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9586166),
	.w1(32'hba0f36fd),
	.w2(32'hba036804),
	.w3(32'hba887174),
	.w4(32'hba867279),
	.w5(32'h3acf66da),
	.w6(32'hbb66fc64),
	.w7(32'hbaaa520d),
	.w8(32'h3ac65157),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395113ce),
	.w1(32'hb95f8a1b),
	.w2(32'h39026008),
	.w3(32'h3a802ad6),
	.w4(32'h3aae3b23),
	.w5(32'h3aa8bbd2),
	.w6(32'h3b0401a0),
	.w7(32'h3ae5248c),
	.w8(32'h3a697dc8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dfe55),
	.w1(32'h39c7bfca),
	.w2(32'h3ad0845c),
	.w3(32'h3a7cfd61),
	.w4(32'h3a565ec0),
	.w5(32'h3b5224e8),
	.w6(32'hba377be9),
	.w7(32'h3a855ed4),
	.w8(32'h3b37a481),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa64165),
	.w1(32'hb916cc90),
	.w2(32'h3aff004f),
	.w3(32'hb91d4312),
	.w4(32'h3b808153),
	.w5(32'hba78daaa),
	.w6(32'h3b4520ba),
	.w7(32'h3bb10dcf),
	.w8(32'hbaec7c41),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0580ae),
	.w1(32'h3b16da33),
	.w2(32'h3b65ff29),
	.w3(32'h39d89e7d),
	.w4(32'hba292666),
	.w5(32'h3b6c0b3f),
	.w6(32'h3b63b966),
	.w7(32'hbb03fae9),
	.w8(32'h3afd9351),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac06101),
	.w1(32'hba5da8ef),
	.w2(32'h39d076ea),
	.w3(32'h3b1831cf),
	.w4(32'h3aedb8b5),
	.w5(32'h3b2ba01e),
	.w6(32'hbb11ba23),
	.w7(32'hb95239b3),
	.w8(32'h3a70b68a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39874a9b),
	.w1(32'hba30b637),
	.w2(32'h3aecfa3e),
	.w3(32'h3b3dd501),
	.w4(32'h3b4d93f4),
	.w5(32'hbac1ecc7),
	.w6(32'hbb21bdcb),
	.w7(32'h3bcc53f2),
	.w8(32'hbb68e646),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74ba51),
	.w1(32'hbb123c4d),
	.w2(32'h3a9736cb),
	.w3(32'hbac212ff),
	.w4(32'hbacdcd86),
	.w5(32'h3b236ccb),
	.w6(32'hbb014b0c),
	.w7(32'hbb206cf2),
	.w8(32'h3aa8b9c6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc1f93),
	.w1(32'hb9fa6205),
	.w2(32'h3affc270),
	.w3(32'hbac4c864),
	.w4(32'h3a46652e),
	.w5(32'hb9642a73),
	.w6(32'hbb256b26),
	.w7(32'hb883c9a1),
	.w8(32'h3af1c63c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f104fe),
	.w1(32'hba1fb920),
	.w2(32'h397a41a8),
	.w3(32'hb9f02887),
	.w4(32'hba4b30d9),
	.w5(32'h3b6f6c66),
	.w6(32'hba151cc0),
	.w7(32'h3a4e85d3),
	.w8(32'h3a0b2f61),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f225e),
	.w1(32'h3921e37e),
	.w2(32'h3a749a90),
	.w3(32'h39867129),
	.w4(32'h39b0ca60),
	.w5(32'h3ac15c05),
	.w6(32'hba0dc1d5),
	.w7(32'h3b816e22),
	.w8(32'h390643b7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ac341),
	.w1(32'h3952845b),
	.w2(32'h3acc34bf),
	.w3(32'h3a99c3e6),
	.w4(32'h3a8070ca),
	.w5(32'hbaf42af8),
	.w6(32'hbabbc233),
	.w7(32'h39b02a91),
	.w8(32'h3aeb40d7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3dbc9),
	.w1(32'h3b3e1a74),
	.w2(32'h3a0e62c8),
	.w3(32'h3a1b79f1),
	.w4(32'h3a132050),
	.w5(32'h3a83095a),
	.w6(32'h3be685ea),
	.w7(32'h3b3adbe5),
	.w8(32'h3a1cafb3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81d04a),
	.w1(32'h39538f12),
	.w2(32'h397f9e10),
	.w3(32'hb8556a70),
	.w4(32'hba9413f0),
	.w5(32'hb9f1a183),
	.w6(32'h3ac6a293),
	.w7(32'h39e7e9cc),
	.w8(32'h3a07f15f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19a49b),
	.w1(32'h3af103d7),
	.w2(32'h3afe9c80),
	.w3(32'hba57a4ae),
	.w4(32'hbaa7228c),
	.w5(32'h3ab29e8b),
	.w6(32'h3b2bc247),
	.w7(32'h3a735f7d),
	.w8(32'hba9b6899),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd9266),
	.w1(32'hbb084d36),
	.w2(32'h3a0ab173),
	.w3(32'hb9989ec6),
	.w4(32'h3a677827),
	.w5(32'h3a65ca38),
	.w6(32'hbb1a7f08),
	.w7(32'hba2d7e8f),
	.w8(32'h3b804a71),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a385191),
	.w1(32'hb9798b3b),
	.w2(32'h3b1539fd),
	.w3(32'hbac3af12),
	.w4(32'hba768910),
	.w5(32'h388f6d53),
	.w6(32'h3917c852),
	.w7(32'h3b469a3c),
	.w8(32'hba0937c3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe9014),
	.w1(32'hbb48deb3),
	.w2(32'h3a33c2f3),
	.w3(32'hbb233d38),
	.w4(32'hbac9a722),
	.w5(32'h3ad1caa5),
	.w6(32'hbb274c51),
	.w7(32'hbab36bde),
	.w8(32'hbb6519ac),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79b58a),
	.w1(32'hbb3734e5),
	.w2(32'hb89522cb),
	.w3(32'hba17be96),
	.w4(32'h39e85fe5),
	.w5(32'hb8955e13),
	.w6(32'hbb4afa35),
	.w7(32'hbb7d0fbe),
	.w8(32'hb9fb8382),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cbc317),
	.w1(32'h39fe4d01),
	.w2(32'h38ce2990),
	.w3(32'hb98d63de),
	.w4(32'hb863a924),
	.w5(32'h3b23285b),
	.w6(32'h3a2d2213),
	.w7(32'h3920596a),
	.w8(32'h3ab922b2),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e2272),
	.w1(32'h3abadbbc),
	.w2(32'h3a260b28),
	.w3(32'h3a8b5844),
	.w4(32'h39f409c2),
	.w5(32'h3a8b95a7),
	.w6(32'hbad49b9e),
	.w7(32'hba398bc9),
	.w8(32'h3aef0d7b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0522d7),
	.w1(32'h3967aeb3),
	.w2(32'h3b0163d8),
	.w3(32'h3a84523a),
	.w4(32'h3a8838d1),
	.w5(32'hbb2fd0e1),
	.w6(32'h37ddccba),
	.w7(32'hba25360e),
	.w8(32'hbb09e541),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04eaca),
	.w1(32'h3b96298b),
	.w2(32'h3b3be5ff),
	.w3(32'h3adea216),
	.w4(32'hba9a8794),
	.w5(32'hbab4dd8c),
	.w6(32'h3b95943f),
	.w7(32'hbb298fd4),
	.w8(32'h3af75499),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64509f),
	.w1(32'h3a3387bb),
	.w2(32'h3a24a5d3),
	.w3(32'h3a984547),
	.w4(32'hbad42ec5),
	.w5(32'hb9664e3a),
	.w6(32'h3b62ab67),
	.w7(32'hb9d82a7b),
	.w8(32'hba2ac5d1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62af44),
	.w1(32'hba4ab0c2),
	.w2(32'h39e1e235),
	.w3(32'hb9b560ea),
	.w4(32'hba0357d2),
	.w5(32'hbaa25131),
	.w6(32'hba35739b),
	.w7(32'hbab3cde5),
	.w8(32'hbaad7bca),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93bdc81),
	.w1(32'h3a189df9),
	.w2(32'h3af0520e),
	.w3(32'hb883d8fa),
	.w4(32'hba7178d9),
	.w5(32'hbadcd309),
	.w6(32'hba80be6e),
	.w7(32'hb9d2f7a7),
	.w8(32'h38a3ab39),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91d876),
	.w1(32'hbb2c9320),
	.w2(32'hb97884e5),
	.w3(32'hbac60514),
	.w4(32'hbb073612),
	.w5(32'hb97f9c1a),
	.w6(32'h3ab8dcf4),
	.w7(32'h3acb46ff),
	.w8(32'hbab81efd),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c0f3f),
	.w1(32'h3a206205),
	.w2(32'h3af848af),
	.w3(32'h39a8908b),
	.w4(32'hba0f3cc8),
	.w5(32'hba80434e),
	.w6(32'hba605d0c),
	.w7(32'hba6ad367),
	.w8(32'hba97a13e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb244e1b),
	.w1(32'hbb769ea5),
	.w2(32'hbb6d269a),
	.w3(32'hbb63e220),
	.w4(32'hbb0f24da),
	.w5(32'h3a2f3f18),
	.w6(32'h3a82e027),
	.w7(32'hba787c1f),
	.w8(32'hb8248bc3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b3478),
	.w1(32'hba20e912),
	.w2(32'h39fc2094),
	.w3(32'hba8a5f12),
	.w4(32'h3a54fa7c),
	.w5(32'hba08185a),
	.w6(32'hbaadb5bb),
	.w7(32'hb951e27c),
	.w8(32'hbadc46c2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd2320),
	.w1(32'h3b3ab3e9),
	.w2(32'h3b1015cd),
	.w3(32'h3ae8f669),
	.w4(32'h3af3280f),
	.w5(32'hb99f39d6),
	.w6(32'h3bd696c3),
	.w7(32'h3aba828b),
	.w8(32'hbb4112b1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa25e97),
	.w1(32'hba63b98b),
	.w2(32'hbad1dedb),
	.w3(32'hbaea83c9),
	.w4(32'h3908491a),
	.w5(32'hba8d41b5),
	.w6(32'h3b112654),
	.w7(32'h3a5c8aa2),
	.w8(32'hba9b85af),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a869607),
	.w1(32'h3a19dd3b),
	.w2(32'h3a869f44),
	.w3(32'hba94fc4c),
	.w4(32'hba06b0dc),
	.w5(32'h3a910cd2),
	.w6(32'hba10d256),
	.w7(32'hb905358d),
	.w8(32'h3986f515),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac255a2),
	.w1(32'hbac1ab2e),
	.w2(32'hbabd9841),
	.w3(32'hbb43764a),
	.w4(32'hba26da7a),
	.w5(32'hbabcc577),
	.w6(32'hbb1dddc5),
	.w7(32'hbb1a3b5c),
	.w8(32'hba66b50f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175487),
	.w1(32'hbb685b4d),
	.w2(32'hbb209426),
	.w3(32'hbb1d9c43),
	.w4(32'hbb28922d),
	.w5(32'hba767795),
	.w6(32'h3b348417),
	.w7(32'h3ab5f3b9),
	.w8(32'h39ba9bd4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0906bd),
	.w1(32'hbac4e3ab),
	.w2(32'h3af21a4e),
	.w3(32'h38f5c397),
	.w4(32'h3b6038d2),
	.w5(32'h3a97f948),
	.w6(32'h39a6146c),
	.w7(32'h3af11c68),
	.w8(32'h3a15929c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c3ec0),
	.w1(32'hbaa8ef36),
	.w2(32'hbab84073),
	.w3(32'hb961d7bd),
	.w4(32'hba2b6204),
	.w5(32'hbb4d004c),
	.w6(32'hba7552c8),
	.w7(32'hba58b5bc),
	.w8(32'hbb133f19),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad12241),
	.w1(32'hbb33fdcf),
	.w2(32'hba6fc2e5),
	.w3(32'hbb1be020),
	.w4(32'hba1633c5),
	.w5(32'h3aaa210e),
	.w6(32'hbaf8cd2d),
	.w7(32'hba994b72),
	.w8(32'h3adbf1e9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378c839d),
	.w1(32'h3a38cfd4),
	.w2(32'h39fe33c2),
	.w3(32'hb8de59a7),
	.w4(32'h39e3bc32),
	.w5(32'h3b386592),
	.w6(32'h3b2728ca),
	.w7(32'h3808c0e4),
	.w8(32'h3b351c05),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b691ca6),
	.w1(32'h3b0bafa1),
	.w2(32'h3b4b2c67),
	.w3(32'h3b8aaf88),
	.w4(32'h3b820bc7),
	.w5(32'hb85f2961),
	.w6(32'h3732ba81),
	.w7(32'h3b5d47f8),
	.w8(32'hbacfce84),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13db62),
	.w1(32'hbb00f270),
	.w2(32'h3a8c30d1),
	.w3(32'hbab3a1b4),
	.w4(32'hba03f5bb),
	.w5(32'hbac2371d),
	.w6(32'hbadaac51),
	.w7(32'h38965ff0),
	.w8(32'hbaa7c0f0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f276f),
	.w1(32'hb961032f),
	.w2(32'h3a0f1990),
	.w3(32'hbabdec6d),
	.w4(32'hba7389e4),
	.w5(32'h39e63ee7),
	.w6(32'hba45932b),
	.w7(32'hba050936),
	.w8(32'hb7ee3548),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a506cf9),
	.w1(32'h3abaa22f),
	.w2(32'hb9e635e4),
	.w3(32'h3a6e0135),
	.w4(32'h3b0489dd),
	.w5(32'h3a9720b5),
	.w6(32'hba276cef),
	.w7(32'hba33c52d),
	.w8(32'h3a47ce10),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf794b),
	.w1(32'h3ae4a4a2),
	.w2(32'h3b39e828),
	.w3(32'hb754840d),
	.w4(32'h3a4d299f),
	.w5(32'h3b37d211),
	.w6(32'hb9622e6a),
	.w7(32'h3a43e175),
	.w8(32'h3b3fd313),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840eb0),
	.w1(32'h3b3440c6),
	.w2(32'h3b517a4c),
	.w3(32'h3afb7902),
	.w4(32'h3b59e138),
	.w5(32'h3b9035c7),
	.w6(32'h3ac8fe68),
	.w7(32'h3a848695),
	.w8(32'h3b57a2a3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91882b),
	.w1(32'h3b5d67ab),
	.w2(32'h3b5d3c89),
	.w3(32'h3ba25562),
	.w4(32'h3ba1fee4),
	.w5(32'hb9926178),
	.w6(32'hbace86d8),
	.w7(32'hb88c7461),
	.w8(32'hbab73436),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba043710),
	.w1(32'hbab35771),
	.w2(32'hbb12ceff),
	.w3(32'hb910077c),
	.w4(32'hbb3657a1),
	.w5(32'hba90781c),
	.w6(32'hbad8ea94),
	.w7(32'hbb426d79),
	.w8(32'hba8bdba6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39146b0a),
	.w1(32'h3a8ad442),
	.w2(32'h3ae8b37b),
	.w3(32'h3a98f8d4),
	.w4(32'h3a8b2063),
	.w5(32'h3b1b9330),
	.w6(32'hba54e0a3),
	.w7(32'hb9a9ed01),
	.w8(32'hbb089c0a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babb81a),
	.w1(32'h3c5116bd),
	.w2(32'h3c191218),
	.w3(32'h3b9c3491),
	.w4(32'h3b40b7db),
	.w5(32'hbaf51756),
	.w6(32'hb9706716),
	.w7(32'hbb3f9a71),
	.w8(32'h39a71eb0),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c36e3),
	.w1(32'hb9139304),
	.w2(32'hbaa8ca6a),
	.w3(32'hbb405444),
	.w4(32'hba9afcd2),
	.w5(32'hba377d12),
	.w6(32'h3bcbadd0),
	.w7(32'h3b534bf8),
	.w8(32'h3b82e07d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432531),
	.w1(32'hbabc67b0),
	.w2(32'h3ae511e7),
	.w3(32'hba5d931c),
	.w4(32'h3a9d4911),
	.w5(32'h3a614123),
	.w6(32'hb9100a12),
	.w7(32'h3b49b625),
	.w8(32'h399000c5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399486c1),
	.w1(32'h3a00320a),
	.w2(32'hbb7f29f4),
	.w3(32'h3aacfe96),
	.w4(32'hbb37b2f5),
	.w5(32'h3a214f7a),
	.w6(32'h3a6e7f0d),
	.w7(32'hbb4fd416),
	.w8(32'h3b0e3840),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e748),
	.w1(32'h3aa37f2d),
	.w2(32'hbb31b59f),
	.w3(32'h3a008e2d),
	.w4(32'hbad44545),
	.w5(32'hbb1fbd4f),
	.w6(32'h3ac3e73d),
	.w7(32'hbb525dac),
	.w8(32'h3a84f9c4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbc529),
	.w1(32'h3b3c590d),
	.w2(32'hbab0da79),
	.w3(32'h3a6ab80f),
	.w4(32'hb94a362e),
	.w5(32'hbb27f009),
	.w6(32'h3ba47fb1),
	.w7(32'h3b82a27e),
	.w8(32'hbbb472bb),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1dad7),
	.w1(32'h3b7e6582),
	.w2(32'h3b5c5ffe),
	.w3(32'hbb376d83),
	.w4(32'hbb40e47b),
	.w5(32'h3a241c78),
	.w6(32'hbb833fad),
	.w7(32'hbb5cdc3c),
	.w8(32'h3a306005),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9db47),
	.w1(32'hbb833a96),
	.w2(32'hbb421b7f),
	.w3(32'hbb39a6fc),
	.w4(32'hbb79d6b4),
	.w5(32'hba54db06),
	.w6(32'hbb610272),
	.w7(32'hbb91bd12),
	.w8(32'h3ab771c1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95607fb),
	.w1(32'h3ad68283),
	.w2(32'hb9dff7d9),
	.w3(32'h3a6bceb4),
	.w4(32'hb9702574),
	.w5(32'hbb668fa7),
	.w6(32'h3a574929),
	.w7(32'h3a62295d),
	.w8(32'hbb8d0984),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0603f3),
	.w1(32'hba99b3d0),
	.w2(32'hbabdce1f),
	.w3(32'hbb90e635),
	.w4(32'hbb93c983),
	.w5(32'h39b145f8),
	.w6(32'hbb94cbcf),
	.w7(32'hbb89222f),
	.w8(32'h3a65ad80),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b047fe3),
	.w1(32'hb934f73e),
	.w2(32'h3ae7fee2),
	.w3(32'h3aef5f98),
	.w4(32'hba78fc82),
	.w5(32'h3a4f73a7),
	.w6(32'h3b0cca93),
	.w7(32'h3af9c3da),
	.w8(32'h3aa6f16a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15f58f),
	.w1(32'h3abd0b50),
	.w2(32'h3913b19f),
	.w3(32'h3abe7705),
	.w4(32'hbb27774e),
	.w5(32'hbb8bf515),
	.w6(32'h3a0b2be1),
	.w7(32'hbb4938d4),
	.w8(32'hbb1eb7cf),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f3360),
	.w1(32'hbb802931),
	.w2(32'hbb795e3c),
	.w3(32'hbc034f10),
	.w4(32'hbb884c2b),
	.w5(32'hbb8a7051),
	.w6(32'hbac4d319),
	.w7(32'hbafc5fa6),
	.w8(32'hbbbab439),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba62c17),
	.w1(32'hbb963aea),
	.w2(32'hbc3aaee8),
	.w3(32'hbb5e36e0),
	.w4(32'hbc2bd7c4),
	.w5(32'h3a99f1c5),
	.w6(32'hbb9c444b),
	.w7(32'hbc3145fa),
	.w8(32'h3b49762c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b1e8c),
	.w1(32'h3be1cc00),
	.w2(32'h3bb80387),
	.w3(32'h3b850a23),
	.w4(32'h39920a52),
	.w5(32'h3b5bfa47),
	.w6(32'h3c0f95b2),
	.w7(32'h3bc34c55),
	.w8(32'h3bd82683),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07a62f),
	.w1(32'h3bc54e56),
	.w2(32'h3b4fd0b2),
	.w3(32'h3b36447a),
	.w4(32'h3b5e8bad),
	.w5(32'hbb453cc8),
	.w6(32'h3ba95225),
	.w7(32'h3a738b5c),
	.w8(32'hbb0fffff),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb716728),
	.w1(32'hbb0b2a7a),
	.w2(32'h3913f6fa),
	.w3(32'hbaec2ffa),
	.w4(32'hb96d7fc6),
	.w5(32'h3be0652a),
	.w6(32'hbae475b6),
	.w7(32'hba884067),
	.w8(32'h3b84a349),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08ad55),
	.w1(32'h3b6394d4),
	.w2(32'h3ba40583),
	.w3(32'h3bbbb870),
	.w4(32'h3b306ac4),
	.w5(32'h392219ca),
	.w6(32'h3ab237c4),
	.w7(32'hba340040),
	.w8(32'hba2cf94a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2bf9),
	.w1(32'hb9b812b3),
	.w2(32'hbaf8de40),
	.w3(32'hb9376626),
	.w4(32'hb9e54d31),
	.w5(32'h3a960b45),
	.w6(32'hbabf055c),
	.w7(32'hbb720a7e),
	.w8(32'hbb17f605),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb202950),
	.w1(32'h38c935ee),
	.w2(32'h3b3e61f7),
	.w3(32'hbb3e1b91),
	.w4(32'h3b0c4191),
	.w5(32'hbaa5d9e0),
	.w6(32'hbafacd8c),
	.w7(32'hba375e72),
	.w8(32'hbabb7a7c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86386e),
	.w1(32'hba374fbc),
	.w2(32'h399a06f1),
	.w3(32'hbadade71),
	.w4(32'hbab3b3ca),
	.w5(32'h3a653f41),
	.w6(32'hbb1dd48b),
	.w7(32'hbb203a60),
	.w8(32'h3a387348),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedafdd),
	.w1(32'h3b9a8824),
	.w2(32'h3ba30b48),
	.w3(32'h3b7289c8),
	.w4(32'h3bbce4e9),
	.w5(32'hbb334d30),
	.w6(32'h3bada196),
	.w7(32'h3be7a1e0),
	.w8(32'hbb6fc920),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e467e0),
	.w1(32'hbaf90cf4),
	.w2(32'hb8a29f62),
	.w3(32'hba3036a8),
	.w4(32'hbb0dcf29),
	.w5(32'h3bcc9f63),
	.w6(32'h3a32175e),
	.w7(32'hb959fd13),
	.w8(32'h3ba63354),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d554f),
	.w1(32'h3b073b39),
	.w2(32'hb9721b57),
	.w3(32'h3b886a41),
	.w4(32'h3aac4ce4),
	.w5(32'hbc0b46a6),
	.w6(32'h3b0c7282),
	.w7(32'h3970bc7c),
	.w8(32'hbc00b70d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09b840),
	.w1(32'hbba72662),
	.w2(32'hbc350f70),
	.w3(32'hbb833751),
	.w4(32'hbc2818ee),
	.w5(32'hbb392170),
	.w6(32'hbae41d60),
	.w7(32'hbc062d3c),
	.w8(32'hbba1ea68),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba60ac1),
	.w1(32'hbad8a85f),
	.w2(32'hbb2460a3),
	.w3(32'hb99d3bba),
	.w4(32'hb990e721),
	.w5(32'h3aeedc00),
	.w6(32'hbb393e54),
	.w7(32'hbb05c4cb),
	.w8(32'h3b7ef61b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91577e),
	.w1(32'h3b894f23),
	.w2(32'h3b1c63f1),
	.w3(32'h3b6d7a05),
	.w4(32'h3b3ba6c9),
	.w5(32'h39a49f87),
	.w6(32'h3b3e3571),
	.w7(32'h3a8ae188),
	.w8(32'hbba48d42),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b828b07),
	.w1(32'h3b9375a3),
	.w2(32'h3bd5da23),
	.w3(32'h3b3b0f9b),
	.w4(32'h3b128179),
	.w5(32'hbb830684),
	.w6(32'h3a2e0dd2),
	.w7(32'h3b230339),
	.w8(32'hbbad53c4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23648a),
	.w1(32'hba9fa404),
	.w2(32'h3b8e8dfb),
	.w3(32'h3a0d6451),
	.w4(32'h3b9de66b),
	.w5(32'h3aeea91c),
	.w6(32'hbab6b401),
	.w7(32'h3b634210),
	.w8(32'hbadea273),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fa40a),
	.w1(32'h3ba4f566),
	.w2(32'h3b94a16c),
	.w3(32'h3b1a6c37),
	.w4(32'h3ba11bea),
	.w5(32'h3aed88bf),
	.w6(32'h3b7bdd6a),
	.w7(32'h3b6b0143),
	.w8(32'h3ac202cb),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a4c0b),
	.w1(32'h3bc3457f),
	.w2(32'h3ba14a26),
	.w3(32'hb8e26387),
	.w4(32'hbae6eac8),
	.w5(32'h3b7f7908),
	.w6(32'h3b538c92),
	.w7(32'hb9e1631e),
	.w8(32'h3ad5dd09),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b356d47),
	.w1(32'h3b3c2e9a),
	.w2(32'h3bc9ba56),
	.w3(32'h3b54c44a),
	.w4(32'h3bb4dbb4),
	.w5(32'hbb4abf58),
	.w6(32'h3bd99671),
	.w7(32'h3c01b69b),
	.w8(32'hbb094c72),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2504c),
	.w1(32'hbb1acb84),
	.w2(32'hbb67b46a),
	.w3(32'hbb81a7aa),
	.w4(32'hbaf8fbca),
	.w5(32'h3c53b246),
	.w6(32'hbb470494),
	.w7(32'hbb20b7d0),
	.w8(32'h3c52344c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule