module layer_10_featuremap_149(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39318fc3),
	.w1(32'hb8e134b5),
	.w2(32'h390a1679),
	.w3(32'h3946c200),
	.w4(32'hb7df29c3),
	.w5(32'h37b4e686),
	.w6(32'hb98b6975),
	.w7(32'hb9c426f8),
	.w8(32'h38ea1421),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb750f428),
	.w1(32'h3a405efa),
	.w2(32'h39e08a49),
	.w3(32'hb9f96cc6),
	.w4(32'h3940a7cc),
	.w5(32'hb9067519),
	.w6(32'h3b4502a0),
	.w7(32'h3b9b0455),
	.w8(32'h3b6f917c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378ac620),
	.w1(32'hb94edcab),
	.w2(32'hb8d424e0),
	.w3(32'h389d3520),
	.w4(32'hb8803550),
	.w5(32'hb864de0a),
	.w6(32'hb9335399),
	.w7(32'hb91ba8c3),
	.w8(32'hb9470af6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90af29c),
	.w1(32'hba9add30),
	.w2(32'hba9d6013),
	.w3(32'hb9220b0b),
	.w4(32'hba2c6c14),
	.w5(32'hba1d63ce),
	.w6(32'hb941afaa),
	.w7(32'hb834d456),
	.w8(32'hb996477c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92cc005),
	.w1(32'hb79a5fed),
	.w2(32'h36bde71f),
	.w3(32'hb936d278),
	.w4(32'hb8130871),
	.w5(32'h39077ad4),
	.w6(32'hb9331c04),
	.w7(32'h38a1c68a),
	.w8(32'h38d7a84b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7638536),
	.w1(32'h39ac85ba),
	.w2(32'h39c0c259),
	.w3(32'h38a79e5a),
	.w4(32'h39a15e6c),
	.w5(32'h39b4c8b7),
	.w6(32'h39aca7e3),
	.w7(32'h39bffcdc),
	.w8(32'h39baebf7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b934e0f),
	.w1(32'h389fcfb1),
	.w2(32'hbb45a735),
	.w3(32'hbad1d0e8),
	.w4(32'hbb2e9a32),
	.w5(32'h3b68ae63),
	.w6(32'hbba952c7),
	.w7(32'h3a4a3cd0),
	.w8(32'h3ba42e55),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91ba31),
	.w1(32'h3bf0ca48),
	.w2(32'h3b7504ab),
	.w3(32'h3c1da154),
	.w4(32'h3c055f86),
	.w5(32'h39f62b93),
	.w6(32'hbc0a288f),
	.w7(32'hbc0fc900),
	.w8(32'hbc1f4dbe),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b4b7d),
	.w1(32'hb63ed3fa),
	.w2(32'hb96047dc),
	.w3(32'h39de16fc),
	.w4(32'h37d16dfd),
	.w5(32'hb9451b00),
	.w6(32'h390d2ba6),
	.w7(32'hb9380d76),
	.w8(32'hb9560a76),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37556c3e),
	.w1(32'hba5fb243),
	.w2(32'hbb6e6c17),
	.w3(32'h3bc4ba9b),
	.w4(32'h3b884d83),
	.w5(32'h3b03a522),
	.w6(32'h39fb3f5c),
	.w7(32'h3aaa2ca5),
	.w8(32'h3ad86a91),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91657d9),
	.w1(32'hb998379d),
	.w2(32'hb98f28a3),
	.w3(32'hb80933ad),
	.w4(32'h38ca596e),
	.w5(32'hb8e61921),
	.w6(32'hb97d4760),
	.w7(32'hb989ee9b),
	.w8(32'hb9b4a247),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4631e6),
	.w1(32'hbbe7b335),
	.w2(32'hbb05f86d),
	.w3(32'h3afe6dbc),
	.w4(32'hbb89eebb),
	.w5(32'h3a07159b),
	.w6(32'hbc0f6ee2),
	.w7(32'hbbf6e661),
	.w8(32'hb98b66b0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a87a9),
	.w1(32'h3a43c35f),
	.w2(32'hba28e25a),
	.w3(32'h3b873539),
	.w4(32'h3b25dc22),
	.w5(32'h3b5bd0c5),
	.w6(32'hbb815548),
	.w7(32'hbb3864e9),
	.w8(32'hba6b8c46),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ef331),
	.w1(32'h3b8aced1),
	.w2(32'h3b3ba789),
	.w3(32'h3bd28250),
	.w4(32'h3beccf6f),
	.w5(32'h3bec49a2),
	.w6(32'h3abe4c24),
	.w7(32'h3b8ff6ae),
	.w8(32'h3bec566a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fe85c),
	.w1(32'hb9cfff35),
	.w2(32'hba8330a5),
	.w3(32'h3a98afee),
	.w4(32'hb78b0e53),
	.w5(32'hba297321),
	.w6(32'h3b3737bc),
	.w7(32'h3b3c4542),
	.w8(32'h3b0abb9c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f0702),
	.w1(32'h3b898974),
	.w2(32'hb995d4ce),
	.w3(32'h3b89f2e7),
	.w4(32'h3c033ea3),
	.w5(32'h3b2ec71a),
	.w6(32'h3aca7204),
	.w7(32'h3bf5acc3),
	.w8(32'h3aac32cb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85bfd4f),
	.w1(32'h3975b344),
	.w2(32'h393fa23b),
	.w3(32'h38d15256),
	.w4(32'h388eb6b1),
	.w5(32'hb869a4bf),
	.w6(32'h39e2ddc5),
	.w7(32'h39e4fad1),
	.w8(32'h3957aefa),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25c3e9),
	.w1(32'h3b0ff10c),
	.w2(32'h3b384a26),
	.w3(32'h3bac97dd),
	.w4(32'h3bb50d49),
	.w5(32'h3b8d887c),
	.w6(32'hbc56ca1b),
	.w7(32'hbc016a4a),
	.w8(32'hbb1f2b12),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73c6e6),
	.w1(32'h3ac1a5c2),
	.w2(32'h3ab96d0c),
	.w3(32'h3a9624f7),
	.w4(32'h3ae60435),
	.w5(32'h3b2ea3af),
	.w6(32'hbbc32486),
	.w7(32'hbba13e03),
	.w8(32'hbac8ebcc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7af8ad7),
	.w1(32'hb8a8d18e),
	.w2(32'hb88c8827),
	.w3(32'h38369944),
	.w4(32'hb915aa2d),
	.w5(32'hb8993f08),
	.w6(32'hb8973165),
	.w7(32'hb7f31c26),
	.w8(32'hb92f2b70),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ec012),
	.w1(32'h39a187f3),
	.w2(32'h39fec203),
	.w3(32'hb96d7ee2),
	.w4(32'h39a66492),
	.w5(32'h39e9ba93),
	.w6(32'h38fa6f14),
	.w7(32'h3923c0c3),
	.w8(32'h38ac4318),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a192ac),
	.w1(32'hba915cf2),
	.w2(32'hb9c6200f),
	.w3(32'h3a1a3a4b),
	.w4(32'hba2ef190),
	.w5(32'hb9ae6048),
	.w6(32'h3add0f08),
	.w7(32'h3a9957f9),
	.w8(32'h3a54e013),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64bec4),
	.w1(32'hbaeaabae),
	.w2(32'hbb1a5535),
	.w3(32'h3b26d645),
	.w4(32'h3adc021d),
	.w5(32'h391bf96d),
	.w6(32'hbbe4da88),
	.w7(32'hba4bf793),
	.w8(32'hbb69f07e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a481a17),
	.w1(32'h3a3692b2),
	.w2(32'h39aed619),
	.w3(32'h3b18cf92),
	.w4(32'h3aeb19d2),
	.w5(32'h3aa1f909),
	.w6(32'h3a31c69e),
	.w7(32'hb9577228),
	.w8(32'hba12e750),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b6c5e),
	.w1(32'h3ad89324),
	.w2(32'h3a519dde),
	.w3(32'h3b35a4ab),
	.w4(32'h3a925544),
	.w5(32'hbb187951),
	.w6(32'h3c2a28c2),
	.w7(32'h3be51ce9),
	.w8(32'h3b7d93a0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9ab1b),
	.w1(32'h39dcc518),
	.w2(32'hb83ffc92),
	.w3(32'h3a34d6b2),
	.w4(32'h3a369887),
	.w5(32'h39da9335),
	.w6(32'h39f41ce7),
	.w7(32'h3a416e4d),
	.w8(32'h3982ea53),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ac8f0),
	.w1(32'hb8999a00),
	.w2(32'hb8141a2e),
	.w3(32'hb989df09),
	.w4(32'hb828fb24),
	.w5(32'hb8976f98),
	.w6(32'hb87e7ea5),
	.w7(32'hb8a22373),
	.w8(32'hb97f9374),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd1cc1),
	.w1(32'h3add4c30),
	.w2(32'hbac9b1af),
	.w3(32'hbb4d976e),
	.w4(32'hbb9f7690),
	.w5(32'hbc1c5848),
	.w6(32'h3c7a59e7),
	.w7(32'h3bfb1125),
	.w8(32'h3af7af28),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962a55d),
	.w1(32'h398b3f5e),
	.w2(32'hb9a9d931),
	.w3(32'h38e1bbbe),
	.w4(32'h397d3a31),
	.w5(32'hb98d9a48),
	.w6(32'h3a238332),
	.w7(32'h38939fae),
	.w8(32'hb98bde74),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad26589),
	.w1(32'hb99f679a),
	.w2(32'hbaf503a5),
	.w3(32'h39346280),
	.w4(32'h3a8ad41f),
	.w5(32'hb9ae3072),
	.w6(32'h3c3dcb03),
	.w7(32'h3c0ee6a9),
	.w8(32'h3c02400d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d1b73),
	.w1(32'h390806bf),
	.w2(32'h394df8dd),
	.w3(32'h39056299),
	.w4(32'h395625a6),
	.w5(32'h397d7032),
	.w6(32'h38cfdfcd),
	.w7(32'h390e7c42),
	.w8(32'h38ea8c48),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938706b),
	.w1(32'h380fe0ef),
	.w2(32'h38b5266e),
	.w3(32'h394bbd67),
	.w4(32'h3863f257),
	.w5(32'h380a39b8),
	.w6(32'h3880c331),
	.w7(32'h38b32436),
	.w8(32'hb8889434),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac9321),
	.w1(32'h3a2c79ee),
	.w2(32'h39eb7ee6),
	.w3(32'h3b0b0551),
	.w4(32'h3afd0f8f),
	.w5(32'h3afcf27a),
	.w6(32'hbb8a7408),
	.w7(32'hbb3a4f99),
	.w8(32'hbac6afe8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ca0fa),
	.w1(32'h3a4ea3cc),
	.w2(32'h399d354c),
	.w3(32'h3ac4eec8),
	.w4(32'h3a436e03),
	.w5(32'hba9eb553),
	.w6(32'h3b37e44e),
	.w7(32'h3b1d479a),
	.w8(32'h3a6394de),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3703d47f),
	.w1(32'hba386094),
	.w2(32'hba448486),
	.w3(32'hb7f1fe78),
	.w4(32'hb9099076),
	.w5(32'hba1a5d63),
	.w6(32'hba815bc6),
	.w7(32'hba689b3a),
	.w8(32'h39b7a8e5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f4e1c),
	.w1(32'h3b1dfaa3),
	.w2(32'h3b8b3eb9),
	.w3(32'h3a9df70d),
	.w4(32'h3b0b3d95),
	.w5(32'h3b55bd43),
	.w6(32'hbc17b61d),
	.w7(32'hbb9f4256),
	.w8(32'hbae98eff),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9730ac),
	.w1(32'h3bd5338e),
	.w2(32'h3ac243fc),
	.w3(32'h3bf87f42),
	.w4(32'hbc1d600b),
	.w5(32'h3bb78d7e),
	.w6(32'h3a282ef5),
	.w7(32'h3b095576),
	.w8(32'h3c4a01c1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cfaef),
	.w1(32'hb8826378),
	.w2(32'h3a3c7488),
	.w3(32'hba45dc16),
	.w4(32'hbb784508),
	.w5(32'hbbba27fd),
	.w6(32'h3c45b708),
	.w7(32'h3be1a7b0),
	.w8(32'h3b469b59),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47ed9e),
	.w1(32'hbb210698),
	.w2(32'hba6b2900),
	.w3(32'hbb1863fe),
	.w4(32'hbbaea54f),
	.w5(32'hbbafe502),
	.w6(32'h3c51876c),
	.w7(32'h3b90ca36),
	.w8(32'hba382c3c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fcbd0b),
	.w1(32'hb9beab40),
	.w2(32'h390bd56e),
	.w3(32'h3962dddf),
	.w4(32'hb8be135c),
	.w5(32'h39f59b64),
	.w6(32'h3afb5577),
	.w7(32'h3b0825d4),
	.w8(32'h3ad27644),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78374b9),
	.w1(32'hb8d93887),
	.w2(32'h38f0ef66),
	.w3(32'h38c7d679),
	.w4(32'h367e1d3d),
	.w5(32'h3928bcce),
	.w6(32'hb7a03d01),
	.w7(32'h3887db35),
	.w8(32'h3898c054),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e358a),
	.w1(32'hb950fbd4),
	.w2(32'h3877d4e8),
	.w3(32'hb839c3d8),
	.w4(32'hb931bbb7),
	.w5(32'hb820db99),
	.w6(32'hb93b2f81),
	.w7(32'h3702d224),
	.w8(32'h39018625),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989ea7a),
	.w1(32'h3a32e670),
	.w2(32'h389015f3),
	.w3(32'h39987970),
	.w4(32'h39aa74dc),
	.w5(32'h389cc78e),
	.w6(32'h3a0f747f),
	.w7(32'h388d97fb),
	.w8(32'hba7e3749),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cd38f),
	.w1(32'h3be1714a),
	.w2(32'h3b1f4fef),
	.w3(32'h3b05c1a3),
	.w4(32'h3bfb9cd6),
	.w5(32'h3b70fb2b),
	.w6(32'h3be23254),
	.w7(32'h3af5a7ca),
	.w8(32'hbbc70bee),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e2d85),
	.w1(32'h39b10edd),
	.w2(32'hb9b25c6d),
	.w3(32'h3a1a85b8),
	.w4(32'hb8b53a4e),
	.w5(32'hbadc2e83),
	.w6(32'h3ba66c93),
	.w7(32'h3ada282e),
	.w8(32'hb99d7c85),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84efac),
	.w1(32'h3a7a0105),
	.w2(32'h3aa7502a),
	.w3(32'hba847a01),
	.w4(32'hba33e615),
	.w5(32'hbb00e642),
	.w6(32'hbaf2800e),
	.w7(32'hbb068d56),
	.w8(32'hbb3c6333),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3be56),
	.w1(32'hba712c89),
	.w2(32'hbb0094f5),
	.w3(32'h39a220ab),
	.w4(32'hb9108a0e),
	.w5(32'hbb030c69),
	.w6(32'h3b2fa083),
	.w7(32'h3a6a79c2),
	.w8(32'hb9ee2a3a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4ce9e),
	.w1(32'hb952a7ba),
	.w2(32'h3ae04862),
	.w3(32'h3bc2b29e),
	.w4(32'h3ba41402),
	.w5(32'h3be6565c),
	.w6(32'hbc74f5ee),
	.w7(32'hbc28b1fb),
	.w8(32'hbb85ab5a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ac351),
	.w1(32'hb8a38836),
	.w2(32'h388388df),
	.w3(32'hb989a919),
	.w4(32'hb9141dd6),
	.w5(32'hb88612b2),
	.w6(32'hb82f8f80),
	.w7(32'h38c6cacc),
	.w8(32'hb9322823),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc63f4),
	.w1(32'h38987b5c),
	.w2(32'h36553806),
	.w3(32'hb925c107),
	.w4(32'h39c74906),
	.w5(32'h39bd31a6),
	.w6(32'h39d6cfc3),
	.w7(32'h39c73c6c),
	.w8(32'h39504630),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfa9e8),
	.w1(32'h392e2925),
	.w2(32'h382d6623),
	.w3(32'h3a08ded6),
	.w4(32'h39c1a6b8),
	.w5(32'h37dd24bd),
	.w6(32'h399b73ed),
	.w7(32'h398ac4fc),
	.w8(32'h37f96eb6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08ce88),
	.w1(32'h3ac22034),
	.w2(32'hbacf30a2),
	.w3(32'hba0329e7),
	.w4(32'h392cf54b),
	.w5(32'hba0ea0b8),
	.w6(32'h39e666e3),
	.w7(32'h3aa9b8b7),
	.w8(32'hbac0513a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af1cc8),
	.w1(32'h3a8f8ee7),
	.w2(32'hba82624a),
	.w3(32'h3a6922d3),
	.w4(32'h3aa18ee5),
	.w5(32'h3a0a2be1),
	.w6(32'hba33c641),
	.w7(32'hb8cf838a),
	.w8(32'h37ce89ee),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a119a57),
	.w1(32'h3a1dfdae),
	.w2(32'h3a2f076c),
	.w3(32'h3c205924),
	.w4(32'h3bf1f48d),
	.w5(32'h3bea64aa),
	.w6(32'hbc012a70),
	.w7(32'hbbae3a0d),
	.w8(32'hba52b24c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad10164),
	.w1(32'h3a873bdc),
	.w2(32'hb9f1f0d6),
	.w3(32'h3b021972),
	.w4(32'h3a57e68e),
	.w5(32'hba3364d0),
	.w6(32'h3ad50e8f),
	.w7(32'hb9c7eca1),
	.w8(32'hbb14b5d0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912d734),
	.w1(32'h389766d7),
	.w2(32'h390e1638),
	.w3(32'h388ba786),
	.w4(32'h39822dd7),
	.w5(32'h39948912),
	.w6(32'h3a4c9752),
	.w7(32'h3a5cdbe1),
	.w8(32'h3a5579b7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38afc53a),
	.w1(32'h39a5ef4a),
	.w2(32'h394c47ce),
	.w3(32'h38d0196a),
	.w4(32'h39c69cbc),
	.w5(32'h39983eae),
	.w6(32'h39abd76d),
	.w7(32'h3906e9a5),
	.w8(32'hb68548bb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385c8511),
	.w1(32'hb9563f0d),
	.w2(32'hba04cacf),
	.w3(32'h396d2a29),
	.w4(32'hb9dbe397),
	.w5(32'hba1f3178),
	.w6(32'h39e4a716),
	.w7(32'h3a230ec8),
	.w8(32'h37e1d6b0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988ef5e),
	.w1(32'hb9865a32),
	.w2(32'hb9cadbd0),
	.w3(32'hb6e8af9a),
	.w4(32'hb87c6ab4),
	.w5(32'hb8bbb357),
	.w6(32'h397a8374),
	.w7(32'h38599e07),
	.w8(32'h38cbd34a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e2e83e),
	.w1(32'h39e1de82),
	.w2(32'h37dae53d),
	.w3(32'h39f72437),
	.w4(32'h3a416297),
	.w5(32'h39bff771),
	.w6(32'hb9ce4339),
	.w7(32'hb8bb3050),
	.w8(32'h37078cb8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10f445),
	.w1(32'h3a95d3cb),
	.w2(32'h396429c9),
	.w3(32'h3a7b2f00),
	.w4(32'h3afd03ee),
	.w5(32'h3a89d4c3),
	.w6(32'hbb3d926a),
	.w7(32'hbaccee66),
	.w8(32'hbadbfb0c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4be01a),
	.w1(32'h3b78cfaa),
	.w2(32'h3ab6ab10),
	.w3(32'h3b45b633),
	.w4(32'h3bb17982),
	.w5(32'h3b06b0dc),
	.w6(32'h3c1e8918),
	.w7(32'h3b9b187a),
	.w8(32'h3affbcc2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976671b),
	.w1(32'hb8be6bbd),
	.w2(32'hb9e79ea1),
	.w3(32'h39650c03),
	.w4(32'hb95da7dc),
	.w5(32'hb988f2d3),
	.w6(32'hb9df0fd3),
	.w7(32'hba16049b),
	.w8(32'hb9afbd28),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f52b72),
	.w1(32'hb95def92),
	.w2(32'hb93f6840),
	.w3(32'hb9ea3b66),
	.w4(32'hb8a6b8ad),
	.w5(32'hb8f450e2),
	.w6(32'hb8ce8a72),
	.w7(32'hb8b9a988),
	.w8(32'h38450998),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d5584),
	.w1(32'hb92efb58),
	.w2(32'hb9482c72),
	.w3(32'h38785a88),
	.w4(32'hb9139fac),
	.w5(32'hb940d426),
	.w6(32'hb94271e3),
	.w7(32'hb9976d47),
	.w8(32'hb9103993),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9475941),
	.w1(32'hb9691692),
	.w2(32'hb9dcd0df),
	.w3(32'hb90a7719),
	.w4(32'hb9b59cc6),
	.w5(32'hb9f87867),
	.w6(32'hb8da4abf),
	.w7(32'hb9ad8b5b),
	.w8(32'hb99778e4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc742653),
	.w1(32'h39513725),
	.w2(32'hbc0314b2),
	.w3(32'h3b53f935),
	.w4(32'h3b889f94),
	.w5(32'hbbbb4b3a),
	.w6(32'h3bb4750c),
	.w7(32'h3c001dab),
	.w8(32'h3b968c82),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81cebd),
	.w1(32'h3b64b4a7),
	.w2(32'h3b8191d4),
	.w3(32'hbbae2566),
	.w4(32'h39da0291),
	.w5(32'hba7699d4),
	.w6(32'hbca29f85),
	.w7(32'hbc1edfa9),
	.w8(32'hbc18457d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e2b87),
	.w1(32'h3b3e7a3b),
	.w2(32'hbb5e23c8),
	.w3(32'h3a218098),
	.w4(32'h3ae4c995),
	.w5(32'hbb3492fc),
	.w6(32'hbb1513e6),
	.w7(32'hbac75872),
	.w8(32'hbbb92831),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc50daf),
	.w1(32'h3964b688),
	.w2(32'hba907dde),
	.w3(32'hba0f7996),
	.w4(32'hbb3172df),
	.w5(32'hbba6ed78),
	.w6(32'h3c1ef62d),
	.w7(32'h3b88d3db),
	.w8(32'h3a9ff156),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ffff0),
	.w1(32'hb8cb7809),
	.w2(32'h33e4b585),
	.w3(32'hb99b73b5),
	.w4(32'hb8a66daf),
	.w5(32'hb8385574),
	.w6(32'hb972dc0f),
	.w7(32'hb91eed07),
	.w8(32'hb83b6cf6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9d2a9),
	.w1(32'h38f742fa),
	.w2(32'h3958ea93),
	.w3(32'hb825ab3e),
	.w4(32'h3913d76c),
	.w5(32'h3933f729),
	.w6(32'h38d17ee2),
	.w7(32'h39157b6f),
	.w8(32'h38b175a7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c1c45),
	.w1(32'h3927d08d),
	.w2(32'h396de9c1),
	.w3(32'h3805cd05),
	.w4(32'h38de7dc5),
	.w5(32'h3926d89a),
	.w6(32'h39003988),
	.w7(32'h38fccbc7),
	.w8(32'h38df5a68),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f9b5b),
	.w1(32'h3ae9fd32),
	.w2(32'h39411bd5),
	.w3(32'h3ab852a7),
	.w4(32'h3ac2c2c2),
	.w5(32'h37ddfe21),
	.w6(32'hbae44428),
	.w7(32'hbae63442),
	.w8(32'hbaf93b99),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9496869),
	.w1(32'hb9133a85),
	.w2(32'hb8993f24),
	.w3(32'hb9267435),
	.w4(32'hb8398d26),
	.w5(32'hb8113bda),
	.w6(32'hb8d9d519),
	.w7(32'hb8a34d46),
	.w8(32'h37c2abbe),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa32dec),
	.w1(32'hb99d8882),
	.w2(32'hba9731a3),
	.w3(32'h3b29aabd),
	.w4(32'h388b3bd3),
	.w5(32'h39646748),
	.w6(32'hbb170682),
	.w7(32'hbb1ff49b),
	.w8(32'h3a4c5398),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b715),
	.w1(32'h3b205ce5),
	.w2(32'h3b501500),
	.w3(32'h3b81de5d),
	.w4(32'h3b2fb04d),
	.w5(32'h3c0a3a15),
	.w6(32'hbc4caf9e),
	.w7(32'hbc09bf54),
	.w8(32'hbba00cb6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9975fd),
	.w1(32'h3aa7cae3),
	.w2(32'h3a88a2d4),
	.w3(32'h3a04478b),
	.w4(32'hb81db8c2),
	.w5(32'hba46e95a),
	.w6(32'h3bb6053a),
	.w7(32'h3b8834a9),
	.w8(32'h3b18d9ef),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc57ba),
	.w1(32'h3a5dce33),
	.w2(32'hba4f50b2),
	.w3(32'h3b5e8686),
	.w4(32'h3b1fd53f),
	.w5(32'h3883cdfc),
	.w6(32'hbaaba384),
	.w7(32'hb916fb35),
	.w8(32'hba38bd45),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82e351),
	.w1(32'hbb72d2bd),
	.w2(32'hba9373b9),
	.w3(32'h3b837bc8),
	.w4(32'h3a88d0bc),
	.w5(32'h39a03c52),
	.w6(32'hba2fb85c),
	.w7(32'h3a7cc8e9),
	.w8(32'h3b80b43d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab100b2),
	.w1(32'h3aeb3634),
	.w2(32'h3a56bb01),
	.w3(32'h3a4d26d1),
	.w4(32'h3a4df1a8),
	.w5(32'hba466c1a),
	.w6(32'h3b9d034f),
	.w7(32'h3ac91c51),
	.w8(32'h39869be9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39381d69),
	.w1(32'hba2bc08b),
	.w2(32'hb8b18d9d),
	.w3(32'h3b1da024),
	.w4(32'h3ac65e70),
	.w5(32'h3af1300d),
	.w6(32'hbb852acd),
	.w7(32'hbb30a2f8),
	.w8(32'hba2e14a9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397683c8),
	.w1(32'h36a8f838),
	.w2(32'h389409b2),
	.w3(32'h397ca66d),
	.w4(32'h383fffff),
	.w5(32'h3874069a),
	.w6(32'h38049078),
	.w7(32'h37bfe465),
	.w8(32'hb7f282f3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71552d7),
	.w1(32'h388fb2de),
	.w2(32'h38b4fcb5),
	.w3(32'h3883aaf5),
	.w4(32'h392a925f),
	.w5(32'h390226fe),
	.w6(32'h385fc2dc),
	.w7(32'h383173fa),
	.w8(32'h38b96825),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388bdb61),
	.w1(32'hb5c45e18),
	.w2(32'h3818e992),
	.w3(32'h38c0b4b3),
	.w4(32'hb8e8ff8e),
	.w5(32'hb998fe1b),
	.w6(32'h393c0ff3),
	.w7(32'hb8c56290),
	.w8(32'h393eafc9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a766e),
	.w1(32'h396bf971),
	.w2(32'hb91150ac),
	.w3(32'hb8234200),
	.w4(32'h399e7d9e),
	.w5(32'h38afdc80),
	.w6(32'h3a9d2279),
	.w7(32'h3a8a1ac7),
	.w8(32'h39a50a14),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b516b7a),
	.w1(32'h383acfdb),
	.w2(32'hbaaa940f),
	.w3(32'h3ab3c64f),
	.w4(32'hba33dfcc),
	.w5(32'hbae717d8),
	.w6(32'h3bc66f2b),
	.w7(32'h3b61b53d),
	.w8(32'h39091d74),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba130768),
	.w1(32'h387b4f6d),
	.w2(32'h37a78e07),
	.w3(32'hba1d4b23),
	.w4(32'h392a1f8b),
	.w5(32'h397f2bfe),
	.w6(32'hb7c34e2f),
	.w7(32'h399e9a11),
	.w8(32'h395f24ce),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af50769),
	.w1(32'h3ac87a8d),
	.w2(32'h3b0d8c9a),
	.w3(32'hbaa77963),
	.w4(32'h3a4990aa),
	.w5(32'hba6ec219),
	.w6(32'hb9c7cb88),
	.w7(32'h37121517),
	.w8(32'hbb823892),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3d37e),
	.w1(32'h3b3fee23),
	.w2(32'h3b0a63e4),
	.w3(32'h3af7425c),
	.w4(32'h3b4f4a88),
	.w5(32'h3b951649),
	.w6(32'hbc151550),
	.w7(32'hbbd9c91e),
	.w8(32'hbb3bcfaa),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b466cad),
	.w1(32'h3ad09837),
	.w2(32'hbb00e047),
	.w3(32'hba91a43a),
	.w4(32'hbb78e27b),
	.w5(32'hbb892d4c),
	.w6(32'h3bddb834),
	.w7(32'h3ad81590),
	.w8(32'hb9c4fd2e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd71cdd),
	.w1(32'hbc0ea76b),
	.w2(32'hbbae90eb),
	.w3(32'h3b4d6818),
	.w4(32'hbbd68456),
	.w5(32'hbb4da9c6),
	.w6(32'hbc3f106f),
	.w7(32'hba850148),
	.w8(32'h3b9debeb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58e250),
	.w1(32'h3a177e7f),
	.w2(32'h3b5e3e5f),
	.w3(32'h3ab69c40),
	.w4(32'hbb0c0a8d),
	.w5(32'hbb3f1746),
	.w6(32'h3b3b15bb),
	.w7(32'hbb0a1e7c),
	.w8(32'hbb815d23),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb806c5b),
	.w1(32'h3b2aa567),
	.w2(32'hbb16adf6),
	.w3(32'h3bae3573),
	.w4(32'h3c0ba9b3),
	.w5(32'h3b343ed5),
	.w6(32'hbba07d25),
	.w7(32'h3b3bf2b1),
	.w8(32'h3a78d310),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c693c7),
	.w1(32'h39da97c9),
	.w2(32'h3a869869),
	.w3(32'h3a997827),
	.w4(32'hba4e4333),
	.w5(32'hbb2f1784),
	.w6(32'h3b4f62f8),
	.w7(32'h3b41f525),
	.w8(32'h3b9d94ec),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67b026),
	.w1(32'h39994f52),
	.w2(32'hba4e9007),
	.w3(32'hba9d3728),
	.w4(32'hbad648b0),
	.w5(32'hbaf17bc1),
	.w6(32'h3c1139df),
	.w7(32'h3c0357e4),
	.w8(32'h3bea018b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa5301),
	.w1(32'h38dc138c),
	.w2(32'h385f09ce),
	.w3(32'hb895d8a8),
	.w4(32'h383ca8fa),
	.w5(32'hb831de7b),
	.w6(32'hb938acdc),
	.w7(32'hb8b2ad81),
	.w8(32'h395ac733),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8968a2),
	.w1(32'h3a7eb6e1),
	.w2(32'h3a2f67ed),
	.w3(32'h3b66040f),
	.w4(32'h3b80d568),
	.w5(32'h3b3df45e),
	.w6(32'hbbc90b87),
	.w7(32'hbb9f14bd),
	.w8(32'hbb03ae02),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11586a),
	.w1(32'hbbbecadf),
	.w2(32'hbc16c7b9),
	.w3(32'hba893e15),
	.w4(32'hbc1e602d),
	.w5(32'hbbfb6375),
	.w6(32'hb9bf5097),
	.w7(32'hbba21ea8),
	.w8(32'hbab01e89),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d06f1),
	.w1(32'h3c4b328d),
	.w2(32'h3b83a975),
	.w3(32'h3c691a4c),
	.w4(32'h3c26c13f),
	.w5(32'h3c4e5ba3),
	.w6(32'hbc988c08),
	.w7(32'hbbb2e7d2),
	.w8(32'hbb4d1ceb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f22c2),
	.w1(32'h3ac7ecc9),
	.w2(32'hbb28b43f),
	.w3(32'h3af7dfdc),
	.w4(32'h3ac0d56e),
	.w5(32'hbac242d2),
	.w6(32'h3c1bae68),
	.w7(32'h3bcca29e),
	.w8(32'h3a233bd5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b538044),
	.w1(32'h3ae7cb7c),
	.w2(32'h3b211fe6),
	.w3(32'h3b257637),
	.w4(32'h3a92e0a0),
	.w5(32'h3a1612c0),
	.w6(32'h3be1144d),
	.w7(32'h3b801003),
	.w8(32'h3b4bbe73),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399962c2),
	.w1(32'hbbdf072f),
	.w2(32'hbba5d238),
	.w3(32'h3c177047),
	.w4(32'hbae65e94),
	.w5(32'h3b3a0cd2),
	.w6(32'hbbc7f44a),
	.w7(32'h3ad53c82),
	.w8(32'h3c1f2f23),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33a22c),
	.w1(32'h39910030),
	.w2(32'h39968457),
	.w3(32'h3a55e36a),
	.w4(32'h3a4305a4),
	.w5(32'h3a06add5),
	.w6(32'h39d6d997),
	.w7(32'h3a5964cf),
	.w8(32'h3a15eac4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8ddb3),
	.w1(32'h3bccd097),
	.w2(32'hbb6da15c),
	.w3(32'h3c732baa),
	.w4(32'h3b65eda8),
	.w5(32'h3c07f498),
	.w6(32'hbb1cdcc0),
	.w7(32'hbbdaa118),
	.w8(32'hbacccc1b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8636ab),
	.w1(32'hbb3722ab),
	.w2(32'hbb8a43ac),
	.w3(32'h3b71d0b1),
	.w4(32'hbaa847ec),
	.w5(32'hba9eb008),
	.w6(32'hba35591d),
	.w7(32'hbb0e81b6),
	.w8(32'hbb8a3405),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9823314),
	.w1(32'hb977e3f3),
	.w2(32'hb928ae86),
	.w3(32'hb983b948),
	.w4(32'hb918d33a),
	.w5(32'hb8e7662a),
	.w6(32'h391d447f),
	.w7(32'h3921c9ca),
	.w8(32'h390ed8d2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaba2f6),
	.w1(32'h3b0db669),
	.w2(32'h3b21a1d2),
	.w3(32'hba47878c),
	.w4(32'h3b143ffd),
	.w5(32'h3ae4d47f),
	.w6(32'h3a8622d5),
	.w7(32'h3b503c8b),
	.w8(32'hba63d763),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfa30c),
	.w1(32'h3aad8bb2),
	.w2(32'h3a174e9a),
	.w3(32'h3b3d2c14),
	.w4(32'h3b70c239),
	.w5(32'h3b2fe75b),
	.w6(32'hbaf2eaee),
	.w7(32'h39dc8990),
	.w8(32'hba017af7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09045b),
	.w1(32'h3a990e1f),
	.w2(32'h3abd7dc7),
	.w3(32'h3ad100b9),
	.w4(32'h3a120586),
	.w5(32'hb9f3ffde),
	.w6(32'h3bca8d24),
	.w7(32'h3b6e900b),
	.w8(32'h3ae9f43b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7eb35),
	.w1(32'h39ef59f3),
	.w2(32'hb8e3d669),
	.w3(32'hba34d671),
	.w4(32'hbac862e0),
	.w5(32'hbb492d5b),
	.w6(32'h3bb5d5f7),
	.w7(32'h3a8a87ca),
	.w8(32'hbb099845),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8633d),
	.w1(32'h395a9ddf),
	.w2(32'hb9ff1a15),
	.w3(32'h38995840),
	.w4(32'hba352e33),
	.w5(32'hba555e88),
	.w6(32'h3b44748f),
	.w7(32'h3b2370b0),
	.w8(32'h3aad312e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a371b6a),
	.w1(32'hb9b3fde7),
	.w2(32'h3b7945f2),
	.w3(32'hbc054a64),
	.w4(32'hbabfa3f4),
	.w5(32'hba9237f3),
	.w6(32'hbc790c0a),
	.w7(32'hbc5761e1),
	.w8(32'hbc13b1b5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb969359),
	.w1(32'h3b93dc76),
	.w2(32'h3af08f8d),
	.w3(32'h3ba7c953),
	.w4(32'h3c1864c3),
	.w5(32'h3bd02523),
	.w6(32'h3b0ef261),
	.w7(32'h3c05acb2),
	.w8(32'h3bc1d1e8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49cdc4),
	.w1(32'h3a17f930),
	.w2(32'h3a13fbb6),
	.w3(32'h3ab4176c),
	.w4(32'h3a9875bf),
	.w5(32'h39ad27f1),
	.w6(32'h3add5080),
	.w7(32'h396e99de),
	.w8(32'hb9a162e4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3876693f),
	.w1(32'h39beaee8),
	.w2(32'h39701204),
	.w3(32'h39188f72),
	.w4(32'h39b2fe34),
	.w5(32'h3983aa64),
	.w6(32'h3a189ded),
	.w7(32'h39f98dfe),
	.w8(32'h39d30d39),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec914e),
	.w1(32'h3aba416c),
	.w2(32'h3a8b5296),
	.w3(32'h3a7273dd),
	.w4(32'h3ab3e84b),
	.w5(32'h3a46340c),
	.w6(32'h39fa3a6e),
	.w7(32'h3aa4fd49),
	.w8(32'h3a89369f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933b7b7),
	.w1(32'h39499aa3),
	.w2(32'h394e006d),
	.w3(32'h393468b3),
	.w4(32'h392c4d18),
	.w5(32'h39435c35),
	.w6(32'h39736bc5),
	.w7(32'h3941bcc3),
	.w8(32'h395c040d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39356e30),
	.w1(32'h37697b16),
	.w2(32'h39338579),
	.w3(32'h393af5a7),
	.w4(32'hb8cc701b),
	.w5(32'hb713de15),
	.w6(32'h37a313ab),
	.w7(32'hb59e1b1c),
	.w8(32'h38b3b5c4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e431b),
	.w1(32'h392d7cc7),
	.w2(32'h39861e7d),
	.w3(32'h3aa26770),
	.w4(32'h39b0e434),
	.w5(32'hba5908f9),
	.w6(32'h3abd7e92),
	.w7(32'hb9a89a12),
	.w8(32'hba0fd17a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9847010),
	.w1(32'hb96ac7e2),
	.w2(32'hb9791c54),
	.w3(32'hb8950862),
	.w4(32'hb7c8462d),
	.w5(32'hb84087bf),
	.w6(32'hb945a263),
	.w7(32'hb99c857c),
	.w8(32'hb9914eed),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf19a),
	.w1(32'hbb713072),
	.w2(32'hb99ff82e),
	.w3(32'h3b06b20b),
	.w4(32'h3a603e13),
	.w5(32'h3aca84bf),
	.w6(32'hbb9a5041),
	.w7(32'hbb742160),
	.w8(32'hbaaa1c26),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a511e04),
	.w1(32'h3a5bf4f9),
	.w2(32'hba9ce4ec),
	.w3(32'hb9a98d47),
	.w4(32'hb8e977a8),
	.w5(32'hbb07f39b),
	.w6(32'h3be9afee),
	.w7(32'h3bcb3b39),
	.w8(32'h3bb1ebbb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39534a70),
	.w1(32'hb99cabb2),
	.w2(32'hb9027339),
	.w3(32'h396a0c8b),
	.w4(32'hb9f5043f),
	.w5(32'hb9a2613a),
	.w6(32'hb9441cd5),
	.w7(32'hb952c367),
	.w8(32'h37ef1406),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37526661),
	.w1(32'hb7f6b946),
	.w2(32'h3932a70e),
	.w3(32'hb9957038),
	.w4(32'h395e018b),
	.w5(32'h3940f224),
	.w6(32'hb9097871),
	.w7(32'h3886c8ac),
	.w8(32'h390be8c5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916d229),
	.w1(32'hb7e016c8),
	.w2(32'h38e9c12b),
	.w3(32'h38bcc893),
	.w4(32'h38c337ea),
	.w5(32'h391b0ec1),
	.w6(32'hb8580b49),
	.w7(32'h37874d8f),
	.w8(32'hb7ce009f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e04fe),
	.w1(32'h3bfce057),
	.w2(32'h3b0b11cf),
	.w3(32'h398273cc),
	.w4(32'h3b956193),
	.w5(32'h3bc0981b),
	.w6(32'hbb4ca3b6),
	.w7(32'hbc52deda),
	.w8(32'hbb912bd1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bee8a),
	.w1(32'h3a3c51bb),
	.w2(32'h3c8ec11b),
	.w3(32'h3b8ea7a0),
	.w4(32'h3c8f8a07),
	.w5(32'h3d1ee175),
	.w6(32'hbd42ddf7),
	.w7(32'hbd42f162),
	.w8(32'hbcca0798),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3cf84),
	.w1(32'hbafe4f43),
	.w2(32'hbc251e03),
	.w3(32'h3cb6415e),
	.w4(32'h3c176d6d),
	.w5(32'h3c0a4b76),
	.w6(32'hbc2fbac1),
	.w7(32'hbc041b5e),
	.w8(32'hbc13f76a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc037b47),
	.w1(32'hbae46396),
	.w2(32'hba4d5196),
	.w3(32'hbbf73ddd),
	.w4(32'h3bc7cf6e),
	.w5(32'h3b2bf4ed),
	.w6(32'hbbc9c5e5),
	.w7(32'hbb99ef37),
	.w8(32'hbc08388e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1af0c6),
	.w1(32'hbbfc0891),
	.w2(32'hbc280d1a),
	.w3(32'h3ba8a303),
	.w4(32'hb9ae6775),
	.w5(32'hbb867009),
	.w6(32'hbc254102),
	.w7(32'hba43250f),
	.w8(32'hbbd726f5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc189fdd),
	.w1(32'hbc914b0a),
	.w2(32'hbc9b6ea6),
	.w3(32'hbb22a7ae),
	.w4(32'h3bd9f116),
	.w5(32'h3c7ac2b7),
	.w6(32'h3a78c0bd),
	.w7(32'hbadd8e8c),
	.w8(32'h3bc3ca29),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50e2e0),
	.w1(32'h3a4038c7),
	.w2(32'h3b21ccbe),
	.w3(32'h3caab29b),
	.w4(32'h3a0a31bf),
	.w5(32'h3a18baf4),
	.w6(32'hbb26109d),
	.w7(32'hbbba72c1),
	.w8(32'h3b00d5e0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3302e1),
	.w1(32'hbc03f043),
	.w2(32'h3af61128),
	.w3(32'h3c059fc5),
	.w4(32'h3c949278),
	.w5(32'h3d2ab647),
	.w6(32'hbd122f95),
	.w7(32'hbd459a1f),
	.w8(32'hbd061657),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c258b),
	.w1(32'hbc0b0e0b),
	.w2(32'hbbc85650),
	.w3(32'h3d254a42),
	.w4(32'h3bc70f83),
	.w5(32'hbaac8bfe),
	.w6(32'hbc5012ce),
	.w7(32'hbbb550a9),
	.w8(32'hbc0e4fb1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00c05f),
	.w1(32'h3b6ef68c),
	.w2(32'h3bf30c77),
	.w3(32'h3b38884c),
	.w4(32'h3b9373fc),
	.w5(32'h3c87a9ea),
	.w6(32'hbbb18314),
	.w7(32'hbc7014b9),
	.w8(32'hbb0b367d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba646bb),
	.w1(32'h3bfe074a),
	.w2(32'h3b9c8d22),
	.w3(32'h3c13aaf3),
	.w4(32'h3c7f50dd),
	.w5(32'h3c78bf49),
	.w6(32'hbc436537),
	.w7(32'hbc7e85b5),
	.w8(32'hbb9cb712),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a539),
	.w1(32'hbc3692d3),
	.w2(32'hbc4d2ec6),
	.w3(32'h3bee6a67),
	.w4(32'hbc0bd102),
	.w5(32'hbc9b69cc),
	.w6(32'h3ae12367),
	.w7(32'h3c5cd101),
	.w8(32'hba76de37),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e73de),
	.w1(32'hbc998bbe),
	.w2(32'hbc91ef22),
	.w3(32'hbc4b4c15),
	.w4(32'h3b280e1e),
	.w5(32'hbaa7de56),
	.w6(32'h3bf44a98),
	.w7(32'h3b97bd8f),
	.w8(32'h3b868a7a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc733a9c),
	.w1(32'h3b74dffd),
	.w2(32'h3a2c3e5c),
	.w3(32'h3c28c65b),
	.w4(32'h3bff1bfa),
	.w5(32'h3c5cc481),
	.w6(32'h39b491d6),
	.w7(32'h3bc60755),
	.w8(32'h3b971d26),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2884ff),
	.w1(32'h399bc5a2),
	.w2(32'hbaf5b917),
	.w3(32'h3bdbad97),
	.w4(32'hba4be99f),
	.w5(32'h3b0d0244),
	.w6(32'h3b08046b),
	.w7(32'hbb5043a7),
	.w8(32'hba99862f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b689ae),
	.w1(32'h3c8fc862),
	.w2(32'h3c53bd5d),
	.w3(32'h399c0012),
	.w4(32'hbbbfc0df),
	.w5(32'hb801f82a),
	.w6(32'h3cebdb81),
	.w7(32'h3cdb6f2b),
	.w8(32'h3cdb50d2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b4fa4),
	.w1(32'h3b81c595),
	.w2(32'hbb50a641),
	.w3(32'hbc108da0),
	.w4(32'h3c1bdcf3),
	.w5(32'h3ba02f80),
	.w6(32'h3c0b02c6),
	.w7(32'h3c180b47),
	.w8(32'h3b4dfe23),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1aeab),
	.w1(32'h3bd2d79e),
	.w2(32'h3c30be09),
	.w3(32'hbc1c0a30),
	.w4(32'h3c3a8098),
	.w5(32'h3ca8192a),
	.w6(32'hbc6fe973),
	.w7(32'hbcaa88e5),
	.w8(32'hbc011349),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c024371),
	.w1(32'hbb2e4344),
	.w2(32'hb9a3194f),
	.w3(32'h3c0c15a8),
	.w4(32'hba5accab),
	.w5(32'h3b23b636),
	.w6(32'hbb86986c),
	.w7(32'hbb819917),
	.w8(32'hbb02a912),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fc015),
	.w1(32'hba7a40c5),
	.w2(32'hbb50a367),
	.w3(32'h3b76d2bf),
	.w4(32'hba06b2e0),
	.w5(32'hbc58a472),
	.w6(32'h3c84a426),
	.w7(32'h3ca7a0f1),
	.w8(32'h3b5b376f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43bb3),
	.w1(32'hbb696c90),
	.w2(32'hbb33d746),
	.w3(32'hbb44548c),
	.w4(32'hbab5a34b),
	.w5(32'hbb9431c0),
	.w6(32'hbaecd2af),
	.w7(32'h3a1b4b1d),
	.w8(32'hbbea603f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad21bb),
	.w1(32'h3abc627a),
	.w2(32'h3b055116),
	.w3(32'h3b9fe92b),
	.w4(32'h3c215814),
	.w5(32'h3c5ed535),
	.w6(32'hbc64ea0a),
	.w7(32'hbc82ba8e),
	.w8(32'hbc1e0893),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0b03b),
	.w1(32'h3c03feda),
	.w2(32'h3c1c2d59),
	.w3(32'h3b014048),
	.w4(32'h3bc8ad26),
	.w5(32'h3c87f34a),
	.w6(32'hba1cd94e),
	.w7(32'hbc6e8d6b),
	.w8(32'h3b37a934),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36eec1),
	.w1(32'h3bce7a1c),
	.w2(32'hbc1d265f),
	.w3(32'h3c5c4fe8),
	.w4(32'hbc157d4b),
	.w5(32'hbc65d734),
	.w6(32'h3c41d17d),
	.w7(32'h3c05c733),
	.w8(32'h3b0ddde0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31794f),
	.w1(32'h3a354d44),
	.w2(32'hbb903e8c),
	.w3(32'hbc45e219),
	.w4(32'h3a98cdb8),
	.w5(32'h3bbc283d),
	.w6(32'h3b9d0524),
	.w7(32'hbae3c770),
	.w8(32'hbb575fa3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16c737),
	.w1(32'hba32c411),
	.w2(32'h3c0c1c9a),
	.w3(32'h3ba30e3c),
	.w4(32'h3befeee4),
	.w5(32'h3cacd9bc),
	.w6(32'hbc971c76),
	.w7(32'hbcc2f812),
	.w8(32'hbb97d152),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6799a3),
	.w1(32'h3b564033),
	.w2(32'hba8bdd0d),
	.w3(32'h3c00c1dd),
	.w4(32'hba99eb1f),
	.w5(32'hbc3bb7c5),
	.w6(32'h3c81b56c),
	.w7(32'h3b3d1617),
	.w8(32'h39d38cae),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad5a88),
	.w1(32'hbab8e3e8),
	.w2(32'hbbe9d7a2),
	.w3(32'hbaaff302),
	.w4(32'h3c392617),
	.w5(32'h3c618be2),
	.w6(32'h3bbb0bc0),
	.w7(32'h3b5b55d5),
	.w8(32'h3bb3d215),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac00018),
	.w1(32'h3b24c91b),
	.w2(32'h3baff37b),
	.w3(32'h3ba118f8),
	.w4(32'h3b86fc7f),
	.w5(32'h3c42bb1d),
	.w6(32'hbbd3404c),
	.w7(32'hbc336586),
	.w8(32'hbc06e9a6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a200c81),
	.w1(32'h3b74358d),
	.w2(32'hbb55785b),
	.w3(32'h3b3bae85),
	.w4(32'h3be97d5b),
	.w5(32'h3b298a66),
	.w6(32'h3b16263f),
	.w7(32'hbb792de6),
	.w8(32'hbbcfa6aa),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6218f5),
	.w1(32'h3bd56a98),
	.w2(32'hbba50cea),
	.w3(32'h3b265be0),
	.w4(32'h3c14f7a7),
	.w5(32'h3a960055),
	.w6(32'h3c912598),
	.w7(32'hbadc07c5),
	.w8(32'h3b18b23e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dc902),
	.w1(32'h3b348d0c),
	.w2(32'hbb68f98c),
	.w3(32'h39b9a282),
	.w4(32'hb8688bb2),
	.w5(32'hbba81057),
	.w6(32'h3c211a35),
	.w7(32'h3bcd389c),
	.w8(32'h3ba55f17),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3186e8),
	.w1(32'h3b0d641a),
	.w2(32'h3bcf75b8),
	.w3(32'h3a29232b),
	.w4(32'h3b1232b2),
	.w5(32'h3c07cd19),
	.w6(32'hbb9175a1),
	.w7(32'hbc2e5dc2),
	.w8(32'hbb3c908b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a8ccb),
	.w1(32'hba516deb),
	.w2(32'h3af29290),
	.w3(32'h3ad63dde),
	.w4(32'h3a264656),
	.w5(32'h3c18c47c),
	.w6(32'hbbbf73b0),
	.w7(32'hbc5defc8),
	.w8(32'hbbabe775),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa55718),
	.w1(32'hbc00b688),
	.w2(32'hbb5fedad),
	.w3(32'h3bed584c),
	.w4(32'hbbb58dc9),
	.w5(32'h3b315f60),
	.w6(32'hbc5d6310),
	.w7(32'hb9eede3d),
	.w8(32'hbbca95d3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0aebb),
	.w1(32'hbb6fabf5),
	.w2(32'hbaa37133),
	.w3(32'h3ab68bb0),
	.w4(32'hba243e32),
	.w5(32'h3a66f349),
	.w6(32'hbbdea119),
	.w7(32'hbb962152),
	.w8(32'hbbc33ced),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b706a18),
	.w1(32'h3b850a31),
	.w2(32'h3b59b6c1),
	.w3(32'h3bb7ad64),
	.w4(32'h3bd8746a),
	.w5(32'hb9c04ca9),
	.w6(32'h3c0cbd68),
	.w7(32'h3c20cc7d),
	.w8(32'h3b2efcde),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6d660),
	.w1(32'h3bb09349),
	.w2(32'h3bfaaac3),
	.w3(32'h3b892508),
	.w4(32'h3b9ff3ca),
	.w5(32'h3c19734c),
	.w6(32'hbb009535),
	.w7(32'hbc176d62),
	.w8(32'hbb9d4798),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1fd0e),
	.w1(32'hba07bc36),
	.w2(32'h3b3549e6),
	.w3(32'h3b21c359),
	.w4(32'h3c112e0a),
	.w5(32'h3bd2a1de),
	.w6(32'hbbe6b117),
	.w7(32'hbb84af57),
	.w8(32'hbad23027),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b220c2a),
	.w1(32'hbb731a00),
	.w2(32'hbbc7b94e),
	.w3(32'h3c1d2300),
	.w4(32'hb9b1c9b8),
	.w5(32'hbbee3a7a),
	.w6(32'hba45ea1a),
	.w7(32'h3a9387d9),
	.w8(32'hbbd2a8bd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec301),
	.w1(32'h3add1d1c),
	.w2(32'h3bf56220),
	.w3(32'hba0496e5),
	.w4(32'h3c0213d6),
	.w5(32'h3ca93a04),
	.w6(32'hbc79fa60),
	.w7(32'hbcd025ac),
	.w8(32'hbc293143),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf74a49),
	.w1(32'h3a10b821),
	.w2(32'hba3e5b2f),
	.w3(32'h3c3d5567),
	.w4(32'h3b9254f4),
	.w5(32'hbb7a7f53),
	.w6(32'h3a6507e1),
	.w7(32'h3b2621ed),
	.w8(32'hbbbd70e4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b203000),
	.w1(32'h3b40df7d),
	.w2(32'h3bf387e2),
	.w3(32'hbb49a985),
	.w4(32'hbbb9d962),
	.w5(32'h3aecdd0f),
	.w6(32'hbc1c9037),
	.w7(32'hbb8c40ed),
	.w8(32'hbb620a9d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cb857),
	.w1(32'hbc391e7b),
	.w2(32'hbc7885ad),
	.w3(32'hb9c37550),
	.w4(32'hbb02b243),
	.w5(32'hbbba12d8),
	.w6(32'hbbab0e5d),
	.w7(32'hbb7acf85),
	.w8(32'hbbdcd094),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f7130),
	.w1(32'hbab764c8),
	.w2(32'hbab4095b),
	.w3(32'h3b5dbbee),
	.w4(32'h3a4a0813),
	.w5(32'h3bdcb85f),
	.w6(32'hbb081fad),
	.w7(32'hbbe0d632),
	.w8(32'hbad6e41c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac17d0),
	.w1(32'hbc262b51),
	.w2(32'hbc8933cc),
	.w3(32'h3aced91e),
	.w4(32'hbc9e7067),
	.w5(32'hbd0659ef),
	.w6(32'h3ce5c9f8),
	.w7(32'h3d1cc42d),
	.w8(32'h3c36b346),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefe9d2),
	.w1(32'h3c3332dc),
	.w2(32'hbb03c706),
	.w3(32'hbc143ea5),
	.w4(32'hbc962bc1),
	.w5(32'hbd2701a2),
	.w6(32'h3d21a5ad),
	.w7(32'h3d3d54e7),
	.w8(32'h3c8c09da),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4094fe),
	.w1(32'h3badadbc),
	.w2(32'hbc09dd91),
	.w3(32'hbcec91c6),
	.w4(32'hbc5f0ad4),
	.w5(32'hbcf1b4ce),
	.w6(32'h3c98e9d0),
	.w7(32'h3ccbab51),
	.w8(32'h3b055038),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc365e74),
	.w1(32'hbb6ac05c),
	.w2(32'h3ba78b8e),
	.w3(32'hbcbfe766),
	.w4(32'h3b1244df),
	.w5(32'h3ba5aee5),
	.w6(32'hbbf7636c),
	.w7(32'h3af0949e),
	.w8(32'h3afe962b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb370b8),
	.w1(32'h3bb13031),
	.w2(32'hbba46b51),
	.w3(32'h3b4c85cd),
	.w4(32'h3bdb8b92),
	.w5(32'hbb1f9a2d),
	.w6(32'h3b97c060),
	.w7(32'hbb60cf6b),
	.w8(32'h3b193ebf),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06666c),
	.w1(32'hbb71a2c4),
	.w2(32'hbb910dc4),
	.w3(32'h3b9f5cda),
	.w4(32'h3bb03276),
	.w5(32'h3c31d49e),
	.w6(32'hbbede30b),
	.w7(32'hbc212c28),
	.w8(32'hbbdb7933),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5942c),
	.w1(32'h3c26971a),
	.w2(32'h3c275780),
	.w3(32'h3b723476),
	.w4(32'h3b378966),
	.w5(32'h3c2769a7),
	.w6(32'h3b6edccc),
	.w7(32'hbb7f8715),
	.w8(32'h3b8af5af),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6ad8e),
	.w1(32'h3b965e20),
	.w2(32'hbbe93a33),
	.w3(32'h3b4df702),
	.w4(32'hbc64f8a8),
	.w5(32'hbd12c407),
	.w6(32'h3ce34880),
	.w7(32'h3d174817),
	.w8(32'h3c40d1b7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ae1d7),
	.w1(32'h3c7645bd),
	.w2(32'h3c1c59a1),
	.w3(32'hbcf36f50),
	.w4(32'hba8e821c),
	.w5(32'h3bf1b65a),
	.w6(32'hbb18a97e),
	.w7(32'h3b42999a),
	.w8(32'h3b49c630),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25006c),
	.w1(32'hbb57aadd),
	.w2(32'h3c3053a2),
	.w3(32'h3c587c57),
	.w4(32'h3caacc67),
	.w5(32'h3d268a82),
	.w6(32'hbd02c708),
	.w7(32'hbd0d8c43),
	.w8(32'hbca8fb2d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be29590),
	.w1(32'hbbcde7b6),
	.w2(32'hbb13b11a),
	.w3(32'h3cd0ca9c),
	.w4(32'h3bb64138),
	.w5(32'h3b7b4c00),
	.w6(32'hbc14c90d),
	.w7(32'hbc82d444),
	.w8(32'hbc21fb38),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1f109),
	.w1(32'hbb84d05c),
	.w2(32'hbafa2cc4),
	.w3(32'h3bd190c3),
	.w4(32'h39be4a0c),
	.w5(32'hbb3b9ae6),
	.w6(32'hbb53c582),
	.w7(32'hbb1025be),
	.w8(32'hbb24971c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09a4a4),
	.w1(32'h3a856128),
	.w2(32'h3bfa6195),
	.w3(32'h38e40f6c),
	.w4(32'hbbbbaf97),
	.w5(32'h3b8ffa35),
	.w6(32'hb9a01547),
	.w7(32'h3bb30fe3),
	.w8(32'hbbbece25),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b049c52),
	.w1(32'h3c18fea5),
	.w2(32'hbb8d2ea1),
	.w3(32'h3b18bbbe),
	.w4(32'hbba024cd),
	.w5(32'hbca4a1c0),
	.w6(32'h3c225586),
	.w7(32'h3c61d386),
	.w8(32'h3b89eac5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0c6b7),
	.w1(32'h3b449f70),
	.w2(32'hbbafcafb),
	.w3(32'hba185f53),
	.w4(32'hbc077af8),
	.w5(32'hbc1ff23c),
	.w6(32'h3bc574ca),
	.w7(32'h3b7ddf10),
	.w8(32'hbc7170fc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc696e69),
	.w1(32'hbaaad0af),
	.w2(32'hbaed2672),
	.w3(32'hbbbc2596),
	.w4(32'h3b625533),
	.w5(32'h3a723923),
	.w6(32'hbb1f6470),
	.w7(32'hbaac5447),
	.w8(32'hbbc4fe29),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2ffd),
	.w1(32'h3bb67dde),
	.w2(32'h3be3f230),
	.w3(32'h3b726879),
	.w4(32'h3c316728),
	.w5(32'h3cb5c6fb),
	.w6(32'hbcd06d6d),
	.w7(32'hbd021257),
	.w8(32'hbc804446),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b319431),
	.w1(32'h3ad5123a),
	.w2(32'hba045dce),
	.w3(32'h3ba1b051),
	.w4(32'h3ade6214),
	.w5(32'hbc3b9c37),
	.w6(32'h3be6a117),
	.w7(32'h3a15a724),
	.w8(32'hbbf2bcc5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79fd78),
	.w1(32'hbb694d66),
	.w2(32'hbbf57d1c),
	.w3(32'h3ae103eb),
	.w4(32'h39be8092),
	.w5(32'h3a51a080),
	.w6(32'hbafbfa6b),
	.w7(32'hbbec9fd3),
	.w8(32'h3b15d884),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d00d3),
	.w1(32'hbafebbe9),
	.w2(32'hbb7ddcb6),
	.w3(32'hbbd30f6c),
	.w4(32'h3ae4b5e9),
	.w5(32'hbc3598ad),
	.w6(32'hbbaaa310),
	.w7(32'h3be78d6f),
	.w8(32'hbb8706d1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b391926),
	.w1(32'hbbfae51a),
	.w2(32'hbc328d31),
	.w3(32'hbbe29ba5),
	.w4(32'hbc238958),
	.w5(32'hbc9b09fd),
	.w6(32'h3c2acc80),
	.w7(32'h3ca40ff9),
	.w8(32'h3b83a8b8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8c7b),
	.w1(32'h3a6c5cb9),
	.w2(32'hb9e0e1ec),
	.w3(32'hbb7a9df8),
	.w4(32'h3b298265),
	.w5(32'hba198674),
	.w6(32'h3b2c7998),
	.w7(32'h3b633cb3),
	.w8(32'hba04eed1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2300f),
	.w1(32'h3b8a2276),
	.w2(32'hbbc030c0),
	.w3(32'h3b070f4e),
	.w4(32'hbb34729e),
	.w5(32'hbc314b19),
	.w6(32'h3b3173ee),
	.w7(32'h3b888081),
	.w8(32'hbb1ce5c7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb829c97),
	.w1(32'hbb96ce13),
	.w2(32'hbba7118e),
	.w3(32'hbb64d2ad),
	.w4(32'hbc02817f),
	.w5(32'hbbd88c50),
	.w6(32'hbbaa5b92),
	.w7(32'h3a403202),
	.w8(32'h3aa04c31),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4e7c7),
	.w1(32'h3b47c565),
	.w2(32'hb940677c),
	.w3(32'h3bbd856d),
	.w4(32'hba1bdb14),
	.w5(32'h3b2d9e63),
	.w6(32'h3bf8f599),
	.w7(32'h3b8bcbd9),
	.w8(32'h3b2610a3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803fde),
	.w1(32'h3b345ec5),
	.w2(32'h3c69b414),
	.w3(32'h3b125a12),
	.w4(32'h39f33b04),
	.w5(32'h3c9db016),
	.w6(32'hbc323f64),
	.w7(32'hbca542ae),
	.w8(32'hbc1034d8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d262),
	.w1(32'h3c9d974d),
	.w2(32'hbafdbe9c),
	.w3(32'h3bbfa0d0),
	.w4(32'hbc45029d),
	.w5(32'hbd3ff87d),
	.w6(32'h3d39daa5),
	.w7(32'h3d528722),
	.w8(32'h3c9b45df),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ad94),
	.w1(32'h3aecf062),
	.w2(32'hb9ad93a6),
	.w3(32'hbd1dabef),
	.w4(32'h3b859ee6),
	.w5(32'hbb4cd5a4),
	.w6(32'h3c118786),
	.w7(32'h3bcc3e52),
	.w8(32'hbb50e2c7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72ab64),
	.w1(32'h3b16e2f3),
	.w2(32'h3bf99b2c),
	.w3(32'h3b2fc6e7),
	.w4(32'h3b981375),
	.w5(32'h3c86063f),
	.w6(32'hbbd6033d),
	.w7(32'hbc8dd6e6),
	.w8(32'hbbfdb15f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7e95f),
	.w1(32'h3c212464),
	.w2(32'h3bed85c6),
	.w3(32'h3c460211),
	.w4(32'h3c43011e),
	.w5(32'h3c9eafd6),
	.w6(32'hbc8283ac),
	.w7(32'hbcbfa7f1),
	.w8(32'hbc0f3637),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b997f71),
	.w1(32'h3ac000dd),
	.w2(32'h3c00e9b8),
	.w3(32'h3c089776),
	.w4(32'h3b465036),
	.w5(32'h3c622d6d),
	.w6(32'hbb65498e),
	.w7(32'hbc58e4de),
	.w8(32'hbb2b1695),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba07027),
	.w1(32'h3b3f9863),
	.w2(32'h3a06202c),
	.w3(32'h3ba5d2f0),
	.w4(32'h3bc5a607),
	.w5(32'h3a7eaa1c),
	.w6(32'hbb6a60d3),
	.w7(32'hbb37e452),
	.w8(32'hbbaa07f9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedd13d),
	.w1(32'hbc035656),
	.w2(32'hbc9bd737),
	.w3(32'h3af98de5),
	.w4(32'hbc53b469),
	.w5(32'hbc671b65),
	.w6(32'h3caa869d),
	.w7(32'h3c9796a9),
	.w8(32'hb9bfd813),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc947799),
	.w1(32'h3b6d0a39),
	.w2(32'h3b4786e7),
	.w3(32'h3b6a173b),
	.w4(32'hb93c833b),
	.w5(32'h3c288ded),
	.w6(32'h3a3e3f41),
	.w7(32'hbc39e42f),
	.w8(32'h3a5914ca),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baffbed),
	.w1(32'hbb515d49),
	.w2(32'hbbc84336),
	.w3(32'h3ba022c0),
	.w4(32'hbad097c7),
	.w5(32'hbc45fe61),
	.w6(32'hbc29cace),
	.w7(32'h39746a7a),
	.w8(32'hbbbb79d7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a38fe),
	.w1(32'hb99ca491),
	.w2(32'hba2fe7b6),
	.w3(32'h3a87a52a),
	.w4(32'h3c6933a5),
	.w5(32'h3c593c9a),
	.w6(32'hbbb71d2d),
	.w7(32'hbba88d2e),
	.w8(32'hbb584f86),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd105cd),
	.w1(32'h3c408711),
	.w2(32'h3c47846d),
	.w3(32'h3c8a0878),
	.w4(32'h3c72bc92),
	.w5(32'h3c96a7ef),
	.w6(32'hba9a093d),
	.w7(32'hbc60a1b9),
	.w8(32'hba16e6d3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a088b),
	.w1(32'h3b0b34cc),
	.w2(32'h3bd3056b),
	.w3(32'h3bbd769f),
	.w4(32'hbb6cac02),
	.w5(32'h3b86a13d),
	.w6(32'hbb28405e),
	.w7(32'hbb0ba192),
	.w8(32'hbb1bf1c7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5af614),
	.w1(32'hba6e37de),
	.w2(32'h3b92c231),
	.w3(32'h3b221a79),
	.w4(32'h3b92f8fb),
	.w5(32'h3b85cbcd),
	.w6(32'hbc02678f),
	.w7(32'hbaeaaf01),
	.w8(32'hbb9fd0f9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b292872),
	.w1(32'h3a3a6e68),
	.w2(32'hba644d13),
	.w3(32'h3b88110f),
	.w4(32'h3a85968f),
	.w5(32'hbad6729b),
	.w6(32'h3b94d5c6),
	.w7(32'h3a9dfbaa),
	.w8(32'h3a8e5388),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67ca7b),
	.w1(32'h3b0050a5),
	.w2(32'h3bba3e5a),
	.w3(32'hbc1ce185),
	.w4(32'h39b02e3b),
	.w5(32'hbb7b8bbb),
	.w6(32'hbc940857),
	.w7(32'hbc64f3a9),
	.w8(32'hbc576da8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79238e),
	.w1(32'h3b89aedd),
	.w2(32'h3b8f279d),
	.w3(32'h390e2781),
	.w4(32'h3a6c4c71),
	.w5(32'hbb2e2aaf),
	.w6(32'hbbcb349c),
	.w7(32'hba174fff),
	.w8(32'hbb5cce58),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b410d7c),
	.w1(32'hbb38ad10),
	.w2(32'hbb927a0f),
	.w3(32'h3ac60a20),
	.w4(32'hb9d2bfe2),
	.w5(32'hbb7362a0),
	.w6(32'hbae3f299),
	.w7(32'hbac15310),
	.w8(32'hbbe7f6e8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44ea9f),
	.w1(32'hbc16b492),
	.w2(32'hbb95b4e9),
	.w3(32'h3b5a68dd),
	.w4(32'hbca3746f),
	.w5(32'hbc9d8666),
	.w6(32'h3cb1650f),
	.w7(32'h3cb11904),
	.w8(32'h3c5e83b7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95b02b),
	.w1(32'h3b8c72d4),
	.w2(32'h3c070fcb),
	.w3(32'hbba64ba9),
	.w4(32'h3b4f3837),
	.w5(32'h3c1f2f39),
	.w6(32'hba934d04),
	.w7(32'hbbd4ac08),
	.w8(32'h3af815ab),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6bea0),
	.w1(32'h3b02efc1),
	.w2(32'h3b9d8358),
	.w3(32'h3b559d0b),
	.w4(32'h3b7d5459),
	.w5(32'h3b8b3943),
	.w6(32'hbbc5efbb),
	.w7(32'hbb5c1719),
	.w8(32'hb9e7526e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1adee4),
	.w1(32'h3c52e229),
	.w2(32'h3cb72406),
	.w3(32'h3bca52db),
	.w4(32'h3b39067d),
	.w5(32'h3cc5b082),
	.w6(32'hbc3324fe),
	.w7(32'hbcbdd93a),
	.w8(32'h3aafd80e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35200d),
	.w1(32'hba975f56),
	.w2(32'h3b14e21f),
	.w3(32'h3ba92958),
	.w4(32'hb85f1f25),
	.w5(32'h3c40f3ad),
	.w6(32'hbc847bcd),
	.w7(32'hbc9f3321),
	.w8(32'hbbdef031),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb3f56),
	.w1(32'hbbcd3158),
	.w2(32'hbc337e05),
	.w3(32'h3bc5675d),
	.w4(32'hbc4ccff9),
	.w5(32'hbccdf5d5),
	.w6(32'h3b9abe37),
	.w7(32'h3c9c2bc1),
	.w8(32'h3b2699d4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11f75a),
	.w1(32'h3ba35988),
	.w2(32'h3bddd0f9),
	.w3(32'hbc891e1c),
	.w4(32'h3c495267),
	.w5(32'h3c5cca4b),
	.w6(32'h3b177b30),
	.w7(32'hbb8aa8f1),
	.w8(32'hba9ad067),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33c2e1),
	.w1(32'h3c01f11a),
	.w2(32'h3c28bba4),
	.w3(32'h3c5f6810),
	.w4(32'h3a043363),
	.w5(32'h3b788f69),
	.w6(32'h3c5e2e37),
	.w7(32'h3c0af170),
	.w8(32'h3acde2b2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81c5ed),
	.w1(32'hbc014ee2),
	.w2(32'hbc1e1b43),
	.w3(32'h3a739530),
	.w4(32'hb99d436a),
	.w5(32'hbb0fe67a),
	.w6(32'hbc103988),
	.w7(32'hbb7bdfc7),
	.w8(32'hbbfad71e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1474a2),
	.w1(32'hbc3fd1eb),
	.w2(32'hbc36f626),
	.w3(32'hb97f12b0),
	.w4(32'h3be2cb02),
	.w5(32'h3ca7714f),
	.w6(32'hbcde05e1),
	.w7(32'hbd089992),
	.w8(32'hbcd870e6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb57bd),
	.w1(32'hbae6dbed),
	.w2(32'hbba58faa),
	.w3(32'h3c6bdf3c),
	.w4(32'hbb468dd0),
	.w5(32'hbb7f0389),
	.w6(32'hbbb6ced7),
	.w7(32'hbbdf4eb5),
	.w8(32'hba8454a3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad68dc),
	.w1(32'h3b812c41),
	.w2(32'hbc8a3d24),
	.w3(32'hbb423868),
	.w4(32'h3c7194f0),
	.w5(32'h3c23a7fc),
	.w6(32'hbbd4028b),
	.w7(32'hbcdd364b),
	.w8(32'hbc543cff),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b528c6),
	.w1(32'hb9ef7b99),
	.w2(32'h3add93f1),
	.w3(32'h3c8384cb),
	.w4(32'h3bf2ddd3),
	.w5(32'h3b9009d6),
	.w6(32'hbc019463),
	.w7(32'hbb46368d),
	.w8(32'hbc185966),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7b09e),
	.w1(32'h3bd72c67),
	.w2(32'h3c5e6cf0),
	.w3(32'h3a666a86),
	.w4(32'h3c45e3dc),
	.w5(32'h3ca0d064),
	.w6(32'hbc833f17),
	.w7(32'hbc4f0c98),
	.w8(32'hbba30443),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf26bf3),
	.w1(32'h3bc4c124),
	.w2(32'hbb45a123),
	.w3(32'h3c4a1f7d),
	.w4(32'h3c098be6),
	.w5(32'hbc3a5d9b),
	.w6(32'h3bd44329),
	.w7(32'h3cb459bf),
	.w8(32'h39b695f0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea4dd7),
	.w1(32'h3a793f7d),
	.w2(32'hbbf29258),
	.w3(32'hbbf6bca6),
	.w4(32'hbb8e2558),
	.w5(32'hba909a91),
	.w6(32'hba9d457d),
	.w7(32'h3b88d4d7),
	.w8(32'hb9fe4feb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6ca4c),
	.w1(32'h3bb517d4),
	.w2(32'h3c172037),
	.w3(32'h3bf4aa0c),
	.w4(32'h3bf8fe81),
	.w5(32'h3cbc3acf),
	.w6(32'hbcb3bcf3),
	.w7(32'hbcf20e15),
	.w8(32'h3acd29db),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc9309),
	.w1(32'h3b6efb5d),
	.w2(32'h3c1dce8d),
	.w3(32'h3bde07d0),
	.w4(32'h3b442330),
	.w5(32'h3c9432f7),
	.w6(32'hbc5fd975),
	.w7(32'hbcc428f2),
	.w8(32'hbc49679b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7639),
	.w1(32'h3b362603),
	.w2(32'h3b36201b),
	.w3(32'h3c09f59a),
	.w4(32'h3aa0d0eb),
	.w5(32'h3c23aeeb),
	.w6(32'hbb1a3400),
	.w7(32'hbc2c2565),
	.w8(32'h39050a5c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba07d53),
	.w1(32'h3ba1a8af),
	.w2(32'h3ba66c96),
	.w3(32'h3bcc81a7),
	.w4(32'h3beeaefe),
	.w5(32'h3c4a2156),
	.w6(32'hbc424151),
	.w7(32'hbc76a395),
	.w8(32'hbc109ad4),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79481d),
	.w1(32'hbbb1aeae),
	.w2(32'hbbf3f78f),
	.w3(32'h3b8c1ca6),
	.w4(32'h3b2e0c97),
	.w5(32'hbac329c0),
	.w6(32'hbc039f01),
	.w7(32'hbb742a87),
	.w8(32'hbc33612b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd292db),
	.w1(32'hba1f289c),
	.w2(32'h3ba16dde),
	.w3(32'hb9f38c0c),
	.w4(32'hbad7f7f9),
	.w5(32'h3c365765),
	.w6(32'hbb64777b),
	.w7(32'hbc5793b2),
	.w8(32'hba4cb29e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea3177),
	.w1(32'h3b285272),
	.w2(32'h3af34743),
	.w3(32'h3ba4dfc5),
	.w4(32'hbadf59de),
	.w5(32'h3be87c4b),
	.w6(32'hba9a92cd),
	.w7(32'hbc15beee),
	.w8(32'h3a62c7e2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6927cc),
	.w1(32'hbb93dda4),
	.w2(32'hbc24b3c6),
	.w3(32'h3b3050c8),
	.w4(32'hbc964594),
	.w5(32'hbd0309c2),
	.w6(32'h3c3156c2),
	.w7(32'h3cc39b0f),
	.w8(32'h3b99470e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50dcbb),
	.w1(32'h3bb944d6),
	.w2(32'h3c69d740),
	.w3(32'hbce7c986),
	.w4(32'h3c1d42e8),
	.w5(32'h3cc92542),
	.w6(32'hbc6b00b9),
	.w7(32'hbca0425a),
	.w8(32'hbbb17b6e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc82c6),
	.w1(32'h3baac46a),
	.w2(32'hbc008417),
	.w3(32'h3c922325),
	.w4(32'h3afde457),
	.w5(32'hbc2d9184),
	.w6(32'h3c2845d9),
	.w7(32'h3cb57a3d),
	.w8(32'h3c45b8c9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac74c7a),
	.w1(32'h3bf4f5c9),
	.w2(32'h3c9aae97),
	.w3(32'hbc988dd3),
	.w4(32'h3c65af04),
	.w5(32'h3cfe7ca5),
	.w6(32'hbcb1a7d4),
	.w7(32'hbce6135b),
	.w8(32'hbc265328),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2488f9),
	.w1(32'hbc335481),
	.w2(32'hbca6aecf),
	.w3(32'h3c9d3179),
	.w4(32'hbb2d8028),
	.w5(32'hbbd94399),
	.w6(32'hbb87a611),
	.w7(32'hba126a4d),
	.w8(32'hbc22fc51),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6f842),
	.w1(32'h3c64d314),
	.w2(32'h3be469cd),
	.w3(32'hbbb498e4),
	.w4(32'h3ac4982f),
	.w5(32'h3b15bfea),
	.w6(32'h3c888d6c),
	.w7(32'h3c5248c5),
	.w8(32'h3c93583e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33ae16),
	.w1(32'h3b91eb73),
	.w2(32'h3b5e1186),
	.w3(32'hb94c35f1),
	.w4(32'h39edec0e),
	.w5(32'h3c5ab2f9),
	.w6(32'hbb479f4f),
	.w7(32'hbc5d62be),
	.w8(32'h3b161f4e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc1b88),
	.w1(32'hbb263544),
	.w2(32'h3b5678e7),
	.w3(32'h3bad7c8e),
	.w4(32'h3b882123),
	.w5(32'h3c892349),
	.w6(32'hbc711726),
	.w7(32'hbcb82673),
	.w8(32'hbc35075d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ba1fd),
	.w1(32'hbb21ff86),
	.w2(32'h3b87ad2a),
	.w3(32'h3c293ccb),
	.w4(32'h3beb572b),
	.w5(32'h3cba1815),
	.w6(32'hbc93fc57),
	.w7(32'hbcdf5c85),
	.w8(32'hbc4d638f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78ba44),
	.w1(32'h39c305d9),
	.w2(32'hbc3a4f75),
	.w3(32'h3c99cbeb),
	.w4(32'hbb90ad15),
	.w5(32'hbc6fe330),
	.w6(32'hbb4f9f76),
	.w7(32'hbbbd488f),
	.w8(32'hbc0a650e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48bdaa),
	.w1(32'hbb0bc981),
	.w2(32'hbb9dd6c5),
	.w3(32'hbc8169c8),
	.w4(32'hbc12aed0),
	.w5(32'hbc75ca64),
	.w6(32'h3b819183),
	.w7(32'h3c678be8),
	.w8(32'hba831e87),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb538db3),
	.w1(32'hb9fea769),
	.w2(32'h3c137785),
	.w3(32'hbb3989f9),
	.w4(32'h3c062880),
	.w5(32'h3cc81914),
	.w6(32'hbc823119),
	.w7(32'hbca73808),
	.w8(32'hbc9b0ef3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce7002),
	.w1(32'hbacb398b),
	.w2(32'h3b666650),
	.w3(32'h3caf4142),
	.w4(32'h3c849942),
	.w5(32'h3cbd252e),
	.w6(32'hbcb6d48e),
	.w7(32'hbcb41ccb),
	.w8(32'hbc9dd402),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae72a9f),
	.w1(32'h3b129c05),
	.w2(32'h3bb6bb91),
	.w3(32'h3c6eccc9),
	.w4(32'h3bec5d5d),
	.w5(32'h3c95b08b),
	.w6(32'hbc7159d5),
	.w7(32'hbcc72527),
	.w8(32'hbc272e48),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c1766),
	.w1(32'hba73f850),
	.w2(32'hbc41aae3),
	.w3(32'h3c0b549b),
	.w4(32'hbc178aad),
	.w5(32'hbc7615f9),
	.w6(32'hbc0c919d),
	.w7(32'hbc475c45),
	.w8(32'hbc80455f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8326db),
	.w1(32'hbc6617a9),
	.w2(32'h3b1af20f),
	.w3(32'hbcb4cac7),
	.w4(32'h3c9285e3),
	.w5(32'h3d5296d4),
	.w6(32'hbd2f4270),
	.w7(32'hbd5dab03),
	.w8(32'hbd0bb113),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f04d4f),
	.w1(32'h3c617a6c),
	.w2(32'h3c511234),
	.w3(32'h3d1f5a4e),
	.w4(32'h3caea515),
	.w5(32'h3caf1559),
	.w6(32'h3c0def1c),
	.w7(32'hbbaecbc6),
	.w8(32'hbb42df0e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0005fc),
	.w1(32'hb91d5f7d),
	.w2(32'hb83fe6a9),
	.w3(32'h3be9df71),
	.w4(32'h377819d6),
	.w5(32'h3782d5b6),
	.w6(32'hb8e5eec0),
	.w7(32'h38d3eddc),
	.w8(32'h392c6432),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe2cdb),
	.w1(32'h3b4bf785),
	.w2(32'h3bc7a0fe),
	.w3(32'hbb3c4221),
	.w4(32'hbaeacfc9),
	.w5(32'hbb71505c),
	.w6(32'hbb39d2b7),
	.w7(32'hbb8b3db8),
	.w8(32'hbbab2996),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule