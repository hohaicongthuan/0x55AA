module layer_10_featuremap_449(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b099bf1),
	.w1(32'hbaace86c),
	.w2(32'h3b544991),
	.w3(32'hbbe2cce8),
	.w4(32'h3b3e06fe),
	.w5(32'h3afa96ad),
	.w6(32'hba9c1a2b),
	.w7(32'h39fe8422),
	.w8(32'hbb942f73),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4f1e2),
	.w1(32'h3b0ecb9a),
	.w2(32'h3bcaaa7b),
	.w3(32'h3c14d665),
	.w4(32'hba6ad63f),
	.w5(32'h3c88c543),
	.w6(32'h3c1f333e),
	.w7(32'h3a86aead),
	.w8(32'h3c38760e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01071c),
	.w1(32'h3a0d199b),
	.w2(32'hbc4ce62a),
	.w3(32'hbbca4f59),
	.w4(32'hbbbd2fee),
	.w5(32'hbcd5507c),
	.w6(32'h3aecc70b),
	.w7(32'hbb83cf68),
	.w8(32'hbc26128c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a9400),
	.w1(32'hbb575a3f),
	.w2(32'h3c81197a),
	.w3(32'hbc470d4d),
	.w4(32'h3c42b9fb),
	.w5(32'h3d27d24a),
	.w6(32'hbc49e694),
	.w7(32'h3b9dfd68),
	.w8(32'hb9a3714d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb660c5c),
	.w1(32'hbb97b7b1),
	.w2(32'hbbd88678),
	.w3(32'hbc0993ac),
	.w4(32'hbbe0615c),
	.w5(32'hbb9a834c),
	.w6(32'h3991fcf2),
	.w7(32'hbc24dbbe),
	.w8(32'hbbbdb6a8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba929a5f),
	.w1(32'hbb333eb4),
	.w2(32'h38aa258d),
	.w3(32'h3bd426b2),
	.w4(32'hbbb1f2f4),
	.w5(32'h3b45749e),
	.w6(32'h3ac9c9ad),
	.w7(32'hbab67b40),
	.w8(32'h3ba7630f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe90a3),
	.w1(32'h3b8069b7),
	.w2(32'hbbd6c8f9),
	.w3(32'h3bb527a4),
	.w4(32'hbaa36aa7),
	.w5(32'hbc276e7c),
	.w6(32'h3afe5bda),
	.w7(32'hbb23e082),
	.w8(32'h3b9e9955),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac706ac),
	.w1(32'hbad7e107),
	.w2(32'hbad3493f),
	.w3(32'h3b16a256),
	.w4(32'h3aff7c2c),
	.w5(32'hbb11a028),
	.w6(32'hbacd28ba),
	.w7(32'h3b739690),
	.w8(32'hb78b4c8a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c6bdf),
	.w1(32'hbbbdfa32),
	.w2(32'hbbb5daa1),
	.w3(32'h3ba2eaca),
	.w4(32'h3b8d4ffa),
	.w5(32'h3c4c0944),
	.w6(32'h3b8962fc),
	.w7(32'h3b978bdb),
	.w8(32'h3b14d063),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07e002),
	.w1(32'hbbb6af3b),
	.w2(32'h3bbd8aea),
	.w3(32'hba93e666),
	.w4(32'hbb260cbd),
	.w5(32'h3c9657f4),
	.w6(32'h3a43bd5c),
	.w7(32'h3b758245),
	.w8(32'hb9b9578a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e953e),
	.w1(32'hbb8224f6),
	.w2(32'h3ab6aa4b),
	.w3(32'h3ab7470d),
	.w4(32'h3c51bde3),
	.w5(32'hbc26f311),
	.w6(32'hbb9f45ad),
	.w7(32'hbac7b942),
	.w8(32'hbc3b0b40),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8bd9c),
	.w1(32'hbbd667ad),
	.w2(32'hbb589563),
	.w3(32'hba965fce),
	.w4(32'hbc10a5f7),
	.w5(32'h3b2aa1f1),
	.w6(32'hbb0057f2),
	.w7(32'h3b9f5dbf),
	.w8(32'h3b802c5c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb294e0b),
	.w1(32'hbbd1e6a3),
	.w2(32'h3b865573),
	.w3(32'h3bab7b91),
	.w4(32'h3ae45ed8),
	.w5(32'h3d330521),
	.w6(32'hbaa98d6b),
	.w7(32'hba9f033a),
	.w8(32'h3b16bc0b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11e89d),
	.w1(32'hbb9aa161),
	.w2(32'hbc2f4f36),
	.w3(32'hbc4a0e7a),
	.w4(32'hbbca4c90),
	.w5(32'hbc827c82),
	.w6(32'hbc7f0f49),
	.w7(32'h39a154da),
	.w8(32'hbc387f27),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc5061),
	.w1(32'h3bb9c76f),
	.w2(32'h3bc4704e),
	.w3(32'hbb335e72),
	.w4(32'h3b67907a),
	.w5(32'hbb20a80f),
	.w6(32'hbbcf61fc),
	.w7(32'h3bcd50c7),
	.w8(32'h3bc97003),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4833cb),
	.w1(32'h3b0755a1),
	.w2(32'h3963dc52),
	.w3(32'hbb0b949b),
	.w4(32'h3c256ac9),
	.w5(32'hba73c968),
	.w6(32'h3afa8f13),
	.w7(32'h3bcc875e),
	.w8(32'hbb532ab6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18ef9e),
	.w1(32'hbad912a7),
	.w2(32'hbbd341ab),
	.w3(32'h3b8b91a2),
	.w4(32'hbb0ca858),
	.w5(32'hbc023ea8),
	.w6(32'hba2ea1bb),
	.w7(32'hbb43c196),
	.w8(32'hbb7a5bbb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cde3e9),
	.w1(32'h3be0b857),
	.w2(32'h3a7e0131),
	.w3(32'hb99d345d),
	.w4(32'h3bf77a19),
	.w5(32'hbc2a8369),
	.w6(32'hbb92297b),
	.w7(32'hb9da2510),
	.w8(32'hbc1e3655),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd36282),
	.w1(32'hbb6a61ce),
	.w2(32'hbb692a4a),
	.w3(32'hbbe25ebd),
	.w4(32'hbaf1d169),
	.w5(32'h3b0588d0),
	.w6(32'hbb6dee09),
	.w7(32'h3ac1f4f7),
	.w8(32'h3b5eeceb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab20d6e),
	.w1(32'hbba11625),
	.w2(32'hbba5e8c8),
	.w3(32'h3b27f5b8),
	.w4(32'hbc5a5f37),
	.w5(32'hbc9142ba),
	.w6(32'h3acbc595),
	.w7(32'hbc25c12d),
	.w8(32'hbb2b08fd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc83d3d),
	.w1(32'h3b0d0b8c),
	.w2(32'hbaaf46d9),
	.w3(32'hbc2b0175),
	.w4(32'h3b0eb9e3),
	.w5(32'hbadf30e3),
	.w6(32'hbbb0b4ff),
	.w7(32'h3ac7c007),
	.w8(32'h3bad000f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad89893),
	.w1(32'h3b953b06),
	.w2(32'h3b2c8623),
	.w3(32'h3b0bb9d9),
	.w4(32'h3b96f09a),
	.w5(32'hbc158d60),
	.w6(32'hbb29a95d),
	.w7(32'h3a522ad2),
	.w8(32'h3ba76120),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6548c),
	.w1(32'hbb21ea48),
	.w2(32'hbc0efc99),
	.w3(32'hbb898965),
	.w4(32'hbc08d2a5),
	.w5(32'h3ba643ac),
	.w6(32'hbb892d82),
	.w7(32'h3a2355fc),
	.w8(32'hbb56a0d6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aa280),
	.w1(32'hbba03e59),
	.w2(32'hbc03549b),
	.w3(32'hbb338e94),
	.w4(32'hbb903414),
	.w5(32'hbb126778),
	.w6(32'hbb4833b5),
	.w7(32'hbb84042c),
	.w8(32'hbbd1eed7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c907a),
	.w1(32'hbb03dba3),
	.w2(32'hbc0c6a88),
	.w3(32'h3b85ca64),
	.w4(32'hbb24dab3),
	.w5(32'hbb4ec2ef),
	.w6(32'hba8c8b3f),
	.w7(32'h3b513f46),
	.w8(32'hbb081c3f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa932c4),
	.w1(32'hbc0a0cc6),
	.w2(32'hbb1b2b28),
	.w3(32'hbb33799d),
	.w4(32'hbc0d6c26),
	.w5(32'h3a11c9b8),
	.w6(32'hbb639ab2),
	.w7(32'hbb33df68),
	.w8(32'h3aeb3b33),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bb798),
	.w1(32'h3af71376),
	.w2(32'hba858ec0),
	.w3(32'h3ba0784d),
	.w4(32'h3b50323f),
	.w5(32'h3bc0cb04),
	.w6(32'hba44968d),
	.w7(32'h3b98ff9c),
	.w8(32'h3ae3b2f4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8e8e),
	.w1(32'hba680332),
	.w2(32'h3b39f9fa),
	.w3(32'hbb53d9a4),
	.w4(32'hbb8d81bc),
	.w5(32'h3c0ddfc1),
	.w6(32'hbac8202d),
	.w7(32'hba8527b9),
	.w8(32'h3bb66f4f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d17c2),
	.w1(32'hbb29f70f),
	.w2(32'hbc5d2702),
	.w3(32'h3b535d9e),
	.w4(32'hbb8483ff),
	.w5(32'h39dbf134),
	.w6(32'h3b9df2bf),
	.w7(32'h3beae1ea),
	.w8(32'hbbc721da),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e8f71),
	.w1(32'hbbb17d30),
	.w2(32'hbb9afc71),
	.w3(32'h3a4f5c85),
	.w4(32'hbb4b3db0),
	.w5(32'hb9b38fa3),
	.w6(32'hbba2d9f4),
	.w7(32'h3ad6e570),
	.w8(32'hbb0e40e4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6a79b),
	.w1(32'hbbe78ae1),
	.w2(32'hbb3bf771),
	.w3(32'h3ac3f156),
	.w4(32'hbc01b364),
	.w5(32'hbb903c14),
	.w6(32'hbae676a4),
	.w7(32'hbb848cde),
	.w8(32'hbac3dfcd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6f847),
	.w1(32'h3b43ac8a),
	.w2(32'h3b4930d0),
	.w3(32'hba0fc0de),
	.w4(32'h3b160364),
	.w5(32'h3b377c49),
	.w6(32'hbc13725b),
	.w7(32'h3bc23f48),
	.w8(32'h3b047730),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd520d8),
	.w1(32'h3be62f1b),
	.w2(32'hbbc15dcc),
	.w3(32'hbc551144),
	.w4(32'h3acbbe07),
	.w5(32'hbc49bf41),
	.w6(32'hbc407a17),
	.w7(32'h3916215b),
	.w8(32'hbb8d551a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06fa22),
	.w1(32'hbbab6dc6),
	.w2(32'hbc3faf0f),
	.w3(32'hba348eac),
	.w4(32'hbb97cfa1),
	.w5(32'hbc078598),
	.w6(32'hb9b4282c),
	.w7(32'hbb93cf81),
	.w8(32'hba7157a1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2567a),
	.w1(32'h3c75f528),
	.w2(32'h3b49f689),
	.w3(32'h39b37793),
	.w4(32'h3b8c9726),
	.w5(32'h3b174900),
	.w6(32'h3a38fd66),
	.w7(32'h3c1429e7),
	.w8(32'hbacfae9a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb6ef),
	.w1(32'h39851ea0),
	.w2(32'h3b8fc790),
	.w3(32'hbab3c570),
	.w4(32'h3891ff46),
	.w5(32'h3c1a013f),
	.w6(32'hbc3aeaaa),
	.w7(32'h3b179b0c),
	.w8(32'hba80a3e8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bcf87),
	.w1(32'h3b91ad62),
	.w2(32'h3c24b6e8),
	.w3(32'hbb738ca6),
	.w4(32'h3c1971a3),
	.w5(32'h3c3191db),
	.w6(32'hbb9fdaa4),
	.w7(32'h3c00227b),
	.w8(32'h3b905ad1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd14982),
	.w1(32'h3b473e9f),
	.w2(32'h3bb285cc),
	.w3(32'hba9d37d6),
	.w4(32'h3bc044a2),
	.w5(32'h3c6c1154),
	.w6(32'hbbe64553),
	.w7(32'h3bf277e7),
	.w8(32'h3bb70abb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d5b9d),
	.w1(32'h3a9eaec4),
	.w2(32'hbc2ba700),
	.w3(32'hbc586afb),
	.w4(32'h39d7ebfa),
	.w5(32'hbc71d588),
	.w6(32'hbc4cf6d9),
	.w7(32'hbb1afec5),
	.w8(32'hbc014ab8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b9d17),
	.w1(32'h38ca159e),
	.w2(32'h3c3504f3),
	.w3(32'h3b84cd52),
	.w4(32'hbba2b3ff),
	.w5(32'h3ca2f6c0),
	.w6(32'h3b979d96),
	.w7(32'h3b085dea),
	.w8(32'h3bc6b379),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baab030),
	.w1(32'hbc76d9eb),
	.w2(32'h3b11a184),
	.w3(32'h3b22cffa),
	.w4(32'hbcd2f9c2),
	.w5(32'h3cf65550),
	.w6(32'h3a9b20e7),
	.w7(32'hbc5d221c),
	.w8(32'h3ae80512),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc507fe7),
	.w1(32'hb7a53b18),
	.w2(32'h3bbbdec1),
	.w3(32'hbb8d51ea),
	.w4(32'hbbac0878),
	.w5(32'h3c9d2ba9),
	.w6(32'hbb7745df),
	.w7(32'hbb7aba28),
	.w8(32'h3b39f880),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16feaa),
	.w1(32'hbbab9ff8),
	.w2(32'h3bdb920a),
	.w3(32'hbb75df50),
	.w4(32'h3b5523ba),
	.w5(32'h3d0a0ad3),
	.w6(32'hbbc445bd),
	.w7(32'h3bf44f50),
	.w8(32'hbbb2ee4e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099caf),
	.w1(32'h3a803d6c),
	.w2(32'h3bd7a3cf),
	.w3(32'hbc55842e),
	.w4(32'h3b36cf55),
	.w5(32'hba535a50),
	.w6(32'hbbecdd91),
	.w7(32'h3b5d06cd),
	.w8(32'hb9a6db0c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e2307),
	.w1(32'hb9047ae4),
	.w2(32'h3b9ebb66),
	.w3(32'hbb6a3be5),
	.w4(32'h3b81c2f4),
	.w5(32'h3c7370a4),
	.w6(32'h3a84456a),
	.w7(32'h3b1e05d0),
	.w8(32'h3bbcf1b0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9347d87),
	.w1(32'hbb4027ae),
	.w2(32'h3a06fae6),
	.w3(32'hba00825a),
	.w4(32'h3c22759d),
	.w5(32'h3ab49d3a),
	.w6(32'h3ade2366),
	.w7(32'h3bafc958),
	.w8(32'h3a389b5f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b7bab),
	.w1(32'hbc1d59bb),
	.w2(32'hbadd846c),
	.w3(32'hba3f2ecc),
	.w4(32'h3a9e4cd5),
	.w5(32'h3bf40546),
	.w6(32'h3a25238f),
	.w7(32'h3bc6490c),
	.w8(32'hbbf122fa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb2442),
	.w1(32'hbb554335),
	.w2(32'h3b55fa00),
	.w3(32'hbbf0cc52),
	.w4(32'h3b32f31b),
	.w5(32'h3bca0c1a),
	.w6(32'hbc3edeb1),
	.w7(32'h3b4282ca),
	.w8(32'h3ba797a9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ad864),
	.w1(32'hbb413840),
	.w2(32'hbc0dac3c),
	.w3(32'hbb2ae04d),
	.w4(32'hbc00a7c6),
	.w5(32'hbc872b5f),
	.w6(32'hbbc0acdf),
	.w7(32'hba78c7ab),
	.w8(32'hbb879fed),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd07ee),
	.w1(32'h3aa0012a),
	.w2(32'h3ae3b190),
	.w3(32'h3c35d060),
	.w4(32'hbb35a358),
	.w5(32'h3b70e2ee),
	.w6(32'h3c2c1455),
	.w7(32'h3beb13c0),
	.w8(32'h3b1b6558),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22dd65),
	.w1(32'h394adb8f),
	.w2(32'hbb82b3c1),
	.w3(32'h3b8244b9),
	.w4(32'hbba32cb9),
	.w5(32'hb9ca97b6),
	.w6(32'hbc1e9aa6),
	.w7(32'hbb165f04),
	.w8(32'hbbc79db7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d9dbd),
	.w1(32'h3b977e61),
	.w2(32'hbc05f020),
	.w3(32'h3b8458fa),
	.w4(32'h3b1da051),
	.w5(32'hbbc694ae),
	.w6(32'h3a4beb7e),
	.w7(32'h3b150b3d),
	.w8(32'hba9ee537),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4466ec),
	.w1(32'hbb2e1ace),
	.w2(32'hbbaffa27),
	.w3(32'hbb0bdeb8),
	.w4(32'hbbe69582),
	.w5(32'hbbd6e637),
	.w6(32'hbb3981ff),
	.w7(32'h3ae76ba2),
	.w8(32'hba719d37),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2520d7),
	.w1(32'h3a3eb296),
	.w2(32'hbadac763),
	.w3(32'h3b89d7c1),
	.w4(32'hbb602655),
	.w5(32'hbc4e6cd8),
	.w6(32'h3b4ade5b),
	.w7(32'h3ba43176),
	.w8(32'hbaf2ecd0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f7770),
	.w1(32'h3bacc9a2),
	.w2(32'h3b79682b),
	.w3(32'h3ac8b6b7),
	.w4(32'hba1e8e63),
	.w5(32'h3b3b0dcd),
	.w6(32'hbb3556f0),
	.w7(32'h3c07e419),
	.w8(32'hbb996f3f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6eae5),
	.w1(32'h3a95cbdf),
	.w2(32'hb92a1137),
	.w3(32'hbb9954b7),
	.w4(32'hbb4b517e),
	.w5(32'hbb81b10e),
	.w6(32'hbb934af4),
	.w7(32'h3b98bfa5),
	.w8(32'h3b797bb4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a3485),
	.w1(32'hba63bcda),
	.w2(32'hbb9016b2),
	.w3(32'hbc13ce16),
	.w4(32'h3a6aa812),
	.w5(32'h3a84aca0),
	.w6(32'hbb9337e6),
	.w7(32'hbc03742d),
	.w8(32'h3a7e3dc5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b730fef),
	.w1(32'h3bc1c02a),
	.w2(32'h3ab055df),
	.w3(32'h3bc11a1f),
	.w4(32'hbbf9e6ce),
	.w5(32'hbc2f9b90),
	.w6(32'h3b8664a5),
	.w7(32'hbc270b5e),
	.w8(32'hbab4b941),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9ef1),
	.w1(32'hbb773702),
	.w2(32'hbc0e17b9),
	.w3(32'h3ab138d2),
	.w4(32'hbc23a985),
	.w5(32'hbbd2babb),
	.w6(32'hbbfc4276),
	.w7(32'hbb4027a6),
	.w8(32'hbc0bf25f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aead2e),
	.w1(32'hbb910126),
	.w2(32'hbb95a4f4),
	.w3(32'hb9844e87),
	.w4(32'hbbfb495a),
	.w5(32'hbb655eb1),
	.w6(32'hbac5ae0b),
	.w7(32'hbc08c300),
	.w8(32'hbadb2d99),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc328478),
	.w1(32'h3b21c749),
	.w2(32'hbc77ee95),
	.w3(32'h3bb8728c),
	.w4(32'h3be49bdf),
	.w5(32'hbc283530),
	.w6(32'h3bbe73cb),
	.w7(32'h38fbf891),
	.w8(32'hbc0efeed),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085abd),
	.w1(32'h3af29da5),
	.w2(32'h3b1be0dc),
	.w3(32'h3aa303fc),
	.w4(32'hbb088c96),
	.w5(32'hbb5b665a),
	.w6(32'hbbb0e1d3),
	.w7(32'h3a2b9d89),
	.w8(32'h3ba9bd37),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23635a),
	.w1(32'h3a62ef5e),
	.w2(32'h3b884f75),
	.w3(32'hbb35960c),
	.w4(32'h3b21b154),
	.w5(32'h3c4aa7dd),
	.w6(32'h3bdc0aa1),
	.w7(32'hbac6b7c4),
	.w8(32'hbc85ee90),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13e209),
	.w1(32'hbb8103b5),
	.w2(32'hbbcd39c3),
	.w3(32'hbc473a9f),
	.w4(32'hbbfe9ba5),
	.w5(32'h3aa8bd7d),
	.w6(32'hbc22fecb),
	.w7(32'hbbcac475),
	.w8(32'hbbe9d1fd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba205b52),
	.w1(32'h3b9d72d1),
	.w2(32'h3b9c7476),
	.w3(32'h3bb1b333),
	.w4(32'h3bf81113),
	.w5(32'h3b5232e7),
	.w6(32'h3b6e3e92),
	.w7(32'hba20f130),
	.w8(32'hbb563556),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30ff64),
	.w1(32'hbb4f048b),
	.w2(32'hbc6430a6),
	.w3(32'h394bc805),
	.w4(32'hbc34cef1),
	.w5(32'hbc46fe5f),
	.w6(32'hb884e1f6),
	.w7(32'hbbab18c8),
	.w8(32'hbba8400c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf32e08),
	.w1(32'hbbe19c4d),
	.w2(32'h38ffe9aa),
	.w3(32'h3b437ac2),
	.w4(32'hbae2faf7),
	.w5(32'h3aa91f1d),
	.w6(32'h3b82de57),
	.w7(32'h3b154987),
	.w8(32'h3ba69910),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37fead),
	.w1(32'hb967a57c),
	.w2(32'hbc5229bb),
	.w3(32'h3b37bc27),
	.w4(32'hbbb4ad54),
	.w5(32'hbc49884b),
	.w6(32'hbbabc34a),
	.w7(32'hbbb45037),
	.w8(32'hbbbac622),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2f7b2),
	.w1(32'hbb81e074),
	.w2(32'h3b41b1f3),
	.w3(32'hbbca391e),
	.w4(32'hbc424028),
	.w5(32'h3c5194c5),
	.w6(32'hbbef62a5),
	.w7(32'hbbafcd3e),
	.w8(32'h3b3dc3f7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa58da9),
	.w1(32'hbb0b402e),
	.w2(32'h3b319173),
	.w3(32'hbb7e2ef4),
	.w4(32'h3b4d8a93),
	.w5(32'h3ab47485),
	.w6(32'hbb5e2a87),
	.w7(32'h3bf11359),
	.w8(32'h3b14e5eb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4076e),
	.w1(32'h3b8f99c1),
	.w2(32'h3b02e8f9),
	.w3(32'h3b851c94),
	.w4(32'h3a334e23),
	.w5(32'h3bebc464),
	.w6(32'h3bda854c),
	.w7(32'hbaaed85e),
	.w8(32'h39caef95),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b451966),
	.w1(32'hbb34b918),
	.w2(32'h3b6234a2),
	.w3(32'h3a94bb11),
	.w4(32'h3b5f3652),
	.w5(32'h3b961f66),
	.w6(32'hba857829),
	.w7(32'hbbadfb16),
	.w8(32'hbb050aa0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6724d6),
	.w1(32'h3ac59c04),
	.w2(32'h3b9a7223),
	.w3(32'hbc2d60ca),
	.w4(32'hbb9360ce),
	.w5(32'hbc015d51),
	.w6(32'hbb507486),
	.w7(32'hbb8c09c6),
	.w8(32'hba8efe2f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba22108),
	.w1(32'hb9c470f2),
	.w2(32'h37b6bba4),
	.w3(32'hba6da6a9),
	.w4(32'h3ac9573f),
	.w5(32'h3b8f8d8f),
	.w6(32'h3b3fe986),
	.w7(32'h3a2e2479),
	.w8(32'hbbb12df0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a096896),
	.w1(32'h3a052c61),
	.w2(32'hbbe14c18),
	.w3(32'hbb130e32),
	.w4(32'hbbb70299),
	.w5(32'hbbff7f5d),
	.w6(32'hbb1d0796),
	.w7(32'hbb391743),
	.w8(32'h3b811a01),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39456d6c),
	.w1(32'h38e0c963),
	.w2(32'h3840c771),
	.w3(32'hbc24976c),
	.w4(32'h3c25f081),
	.w5(32'h3c9e1137),
	.w6(32'hbba8efdb),
	.w7(32'hbb9e5e06),
	.w8(32'hbc15d458),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9fe87),
	.w1(32'h3a9ecba7),
	.w2(32'hb9fb3f82),
	.w3(32'h3b5f691e),
	.w4(32'h3bb1d691),
	.w5(32'hb9a56bff),
	.w6(32'hbb9035db),
	.w7(32'h3bc8d216),
	.w8(32'h3bd31f47),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26604e),
	.w1(32'hbb780e24),
	.w2(32'hbb8794bd),
	.w3(32'h39830ec7),
	.w4(32'hbac7ec29),
	.w5(32'hbc28ba0d),
	.w6(32'h3be758a5),
	.w7(32'h3bbad651),
	.w8(32'h3c0186a4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae454f3),
	.w1(32'h398e31d5),
	.w2(32'h3ba1c202),
	.w3(32'hbc29081b),
	.w4(32'h3a5c0d48),
	.w5(32'h3b4bc921),
	.w6(32'h3c004af0),
	.w7(32'hbaf38e40),
	.w8(32'hbb6ea23f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c243db5),
	.w1(32'hbb6fde72),
	.w2(32'hbba7f808),
	.w3(32'h3b726aa4),
	.w4(32'h3bbbaac6),
	.w5(32'h3badf5c4),
	.w6(32'h3b6640ab),
	.w7(32'h3b9c0b63),
	.w8(32'hba7adf0b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d845f),
	.w1(32'h3b29d88f),
	.w2(32'hba0b70b1),
	.w3(32'hbac1f141),
	.w4(32'hbb699157),
	.w5(32'hbac135bd),
	.w6(32'h3a3b0031),
	.w7(32'h3c1ae55a),
	.w8(32'h3b8c8b67),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c7054),
	.w1(32'hbafe27ab),
	.w2(32'h38129b64),
	.w3(32'h3bd52ae0),
	.w4(32'hba9ff2f1),
	.w5(32'hb90b180f),
	.w6(32'h3c1b03ca),
	.w7(32'hbb808aff),
	.w8(32'hbb200ff2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba450873),
	.w1(32'hbb2c1d63),
	.w2(32'hbb881b48),
	.w3(32'hbad36dff),
	.w4(32'h3be76b15),
	.w5(32'h3b9c1c33),
	.w6(32'h394e68d1),
	.w7(32'hbb086868),
	.w8(32'hbbbc91c3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba158076),
	.w1(32'hbabe21e5),
	.w2(32'hb9a52611),
	.w3(32'h3a67c4d1),
	.w4(32'h3bc43cf5),
	.w5(32'h3c05480c),
	.w6(32'hbb15056d),
	.w7(32'hbae09d9f),
	.w8(32'hbb50ea9d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d71df),
	.w1(32'h3a9bfd95),
	.w2(32'h3b40f04f),
	.w3(32'hbb772f76),
	.w4(32'hbc2b8086),
	.w5(32'hbc19939e),
	.w6(32'hbbdc61fc),
	.w7(32'hbb2af0fa),
	.w8(32'hbb3deafd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994b56f),
	.w1(32'hba9211f7),
	.w2(32'h3a3d1a74),
	.w3(32'hb9d73ac9),
	.w4(32'hba53a88f),
	.w5(32'hbb97b306),
	.w6(32'h3a74690f),
	.w7(32'hba73c3ec),
	.w8(32'hbadbcb2b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f4345),
	.w1(32'h3b0cbae4),
	.w2(32'h39e39b17),
	.w3(32'h3ac9a7b2),
	.w4(32'hba661831),
	.w5(32'hbb3a0366),
	.w6(32'hbb549989),
	.w7(32'h3a6e2023),
	.w8(32'hbb1ed22a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e2e1b),
	.w1(32'h3a10e73f),
	.w2(32'hbaff30bb),
	.w3(32'h39e9677b),
	.w4(32'hbb831e00),
	.w5(32'hbb160461),
	.w6(32'h39e73669),
	.w7(32'hbaefd3d4),
	.w8(32'hbb164955),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1ddfa),
	.w1(32'hbb3e4509),
	.w2(32'hbc298c8a),
	.w3(32'hbb6b979d),
	.w4(32'h3bcab835),
	.w5(32'h3c37721e),
	.w6(32'h3bb767fb),
	.w7(32'h39cf8cc3),
	.w8(32'hb9c79d22),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb304d32),
	.w1(32'hbb3c6503),
	.w2(32'hba0ef8f1),
	.w3(32'hbb50e873),
	.w4(32'hbbe74784),
	.w5(32'hbb828c6d),
	.w6(32'hbb677c6a),
	.w7(32'h3aeb0c69),
	.w8(32'hbb4c6632),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb5b46),
	.w1(32'hbb588b06),
	.w2(32'hbbae29c2),
	.w3(32'hbb3639eb),
	.w4(32'hbb4aac98),
	.w5(32'hbbba6b6b),
	.w6(32'hbc054f7a),
	.w7(32'hbb747106),
	.w8(32'hbb759164),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde0308),
	.w1(32'h3afa56f5),
	.w2(32'h3b9c8f89),
	.w3(32'hba1f7264),
	.w4(32'h3b892027),
	.w5(32'h3a649221),
	.w6(32'h3b53fe86),
	.w7(32'hbae5b977),
	.w8(32'h3b91ae4d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f55b4),
	.w1(32'h3ad64b6b),
	.w2(32'h3c354755),
	.w3(32'h3c07683b),
	.w4(32'h3be76395),
	.w5(32'h3c004f4d),
	.w6(32'h3b97c0b3),
	.w7(32'hba3f4965),
	.w8(32'hbbbe8d87),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ddf8),
	.w1(32'h3ba93b28),
	.w2(32'h3c02e50d),
	.w3(32'hbb7de821),
	.w4(32'h3af63d20),
	.w5(32'h3b463a0d),
	.w6(32'hbc34a168),
	.w7(32'h3ab11f9f),
	.w8(32'hbb025bc4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a16b3),
	.w1(32'hbb879cde),
	.w2(32'hbc07556d),
	.w3(32'h3ac056cf),
	.w4(32'h3c4a8105),
	.w5(32'h3c8079fb),
	.w6(32'hbabc75f4),
	.w7(32'h389b5899),
	.w8(32'h3b57cf62),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab34cfb),
	.w1(32'h3bd60809),
	.w2(32'hbb979aff),
	.w3(32'h3b5cec71),
	.w4(32'hbbeaae8d),
	.w5(32'hbbe7fb9a),
	.w6(32'h3b43deaf),
	.w7(32'hbb104906),
	.w8(32'h3a081c93),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd43176),
	.w1(32'h3b531f9d),
	.w2(32'hbb01e36e),
	.w3(32'h3bdb5b97),
	.w4(32'hbb81c803),
	.w5(32'h3b18c1a0),
	.w6(32'h3bf69680),
	.w7(32'hb912ac4f),
	.w8(32'h3b884644),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21676a),
	.w1(32'h39406bff),
	.w2(32'hbbaa6eef),
	.w3(32'h3b85a4ad),
	.w4(32'h397ef5fd),
	.w5(32'hbb6469b1),
	.w6(32'hbb4c29b3),
	.w7(32'hbaa0d54c),
	.w8(32'hbb80e15f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc121f5),
	.w1(32'h3a239505),
	.w2(32'hbb304a32),
	.w3(32'hbaec717a),
	.w4(32'hbab0b14c),
	.w5(32'h3b0af0a9),
	.w6(32'hbbf5a2d4),
	.w7(32'hb98f6878),
	.w8(32'hbb0ff4c0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c759f),
	.w1(32'hbb313061),
	.w2(32'hbc3210f3),
	.w3(32'hba8099aa),
	.w4(32'h3b305e6e),
	.w5(32'h3ba144df),
	.w6(32'hba2a2392),
	.w7(32'h3c27aad3),
	.w8(32'h3c065dd3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc186b9e),
	.w1(32'hbb6fa650),
	.w2(32'hbb598c57),
	.w3(32'h3b5e5c67),
	.w4(32'h3ae1cb30),
	.w5(32'h3c1211a7),
	.w6(32'h3bbb9343),
	.w7(32'h3af7832c),
	.w8(32'hbaac9b01),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6488d),
	.w1(32'hbb1a29fa),
	.w2(32'hbb5c37d6),
	.w3(32'hbb5337a7),
	.w4(32'hbb98549c),
	.w5(32'hbb211843),
	.w6(32'hbaa9dadd),
	.w7(32'hbc031ba1),
	.w8(32'hbb903471),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4d1f),
	.w1(32'h3b033988),
	.w2(32'hbbf739c3),
	.w3(32'h3bcaf049),
	.w4(32'hbb5d2bcc),
	.w5(32'hb7f58842),
	.w6(32'hbc161dfc),
	.w7(32'hbba532ff),
	.w8(32'h3ad11ee2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38178),
	.w1(32'hbc03cfef),
	.w2(32'h3b20d395),
	.w3(32'hb81cd2f4),
	.w4(32'hbb3487cd),
	.w5(32'hbc2bf6b4),
	.w6(32'h3c01109d),
	.w7(32'hb9968e1b),
	.w8(32'hbbce6f30),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5295d5),
	.w1(32'hbbdaf7ed),
	.w2(32'h3acc1847),
	.w3(32'hba3bd7bf),
	.w4(32'h3b7dc45e),
	.w5(32'h3c0253ba),
	.w6(32'hbb860375),
	.w7(32'hba96bf7f),
	.w8(32'hbbeb6836),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10a368),
	.w1(32'hbb093037),
	.w2(32'hba92c18d),
	.w3(32'hbbe76178),
	.w4(32'hba391232),
	.w5(32'hb9f5d014),
	.w6(32'hbb683e33),
	.w7(32'hb9dc30ed),
	.w8(32'hba837719),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf43130),
	.w1(32'h3b6c9b75),
	.w2(32'h3b9580b7),
	.w3(32'h3aa874aa),
	.w4(32'hba0da737),
	.w5(32'hbb268c56),
	.w6(32'hbb6b7600),
	.w7(32'hba6d9b18),
	.w8(32'hbb2e2c89),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1ebf8),
	.w1(32'h3a9a8b5b),
	.w2(32'h3a0753f4),
	.w3(32'hbbbe7853),
	.w4(32'hbac5d5d7),
	.w5(32'hbbec2bd5),
	.w6(32'hb9c54f74),
	.w7(32'hbb2c285d),
	.w8(32'hbaa3fe3e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2cbe6),
	.w1(32'hbb71d99e),
	.w2(32'h3a4b087d),
	.w3(32'hbb285227),
	.w4(32'h3b62a424),
	.w5(32'h3c09c9ca),
	.w6(32'hbb862347),
	.w7(32'hbb5b494c),
	.w8(32'hbbb94164),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d1be4),
	.w1(32'hba05a8a4),
	.w2(32'h380c15ef),
	.w3(32'h3b65efe6),
	.w4(32'h3b9844d2),
	.w5(32'h3bec93a9),
	.w6(32'hbae2ae87),
	.w7(32'hbaa8fdfb),
	.w8(32'hbbde2d3f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b782579),
	.w1(32'h39ee75d2),
	.w2(32'h3bb80a8e),
	.w3(32'h3c35c8b5),
	.w4(32'hbb8c8b22),
	.w5(32'h3a94fa92),
	.w6(32'hbc080fc3),
	.w7(32'hbbd78fda),
	.w8(32'hba9a309f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4e75a),
	.w1(32'h3b1f7c2c),
	.w2(32'hba82e537),
	.w3(32'hbb59b697),
	.w4(32'hbb214a07),
	.w5(32'hbb744256),
	.w6(32'hba735f36),
	.w7(32'h3bb8e882),
	.w8(32'h3b89f87e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48b92b),
	.w1(32'h3beb22f4),
	.w2(32'hbb3957d8),
	.w3(32'hbb7ce12c),
	.w4(32'hbbb0d2f7),
	.w5(32'hbbb5e683),
	.w6(32'h3a251f5f),
	.w7(32'h3ba30d2d),
	.w8(32'h3c05ba71),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1bc6),
	.w1(32'hbc2c5d6c),
	.w2(32'hbc7bc5df),
	.w3(32'h3bb02b3b),
	.w4(32'h3c2c97f2),
	.w5(32'h3d09af22),
	.w6(32'h3bceec5b),
	.w7(32'hbbda349f),
	.w8(32'hbc468670),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d3571),
	.w1(32'hbc141767),
	.w2(32'hbb2e4028),
	.w3(32'hbbade94e),
	.w4(32'h3aba9e90),
	.w5(32'h3b0c52d0),
	.w6(32'hbbc373e9),
	.w7(32'h3b114b7a),
	.w8(32'hbb3734fa),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a3de0),
	.w1(32'h3b6e80e5),
	.w2(32'hbb4fc19a),
	.w3(32'h3b154f1c),
	.w4(32'h3b77f3bb),
	.w5(32'h3aa06b6b),
	.w6(32'h3a2ba390),
	.w7(32'hba99ce67),
	.w8(32'h3abad2b4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39952164),
	.w1(32'h3bcc28a2),
	.w2(32'hba17b234),
	.w3(32'hbaaa6737),
	.w4(32'hbb17e592),
	.w5(32'hbbc59931),
	.w6(32'h3b1203ea),
	.w7(32'h3a87eda7),
	.w8(32'h3ad1f831),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78954aa),
	.w1(32'h3c195f97),
	.w2(32'h3c2fd89b),
	.w3(32'h3c17cd22),
	.w4(32'h3c4e046c),
	.w5(32'h3b687760),
	.w6(32'hbacd538e),
	.w7(32'hbb9a00cc),
	.w8(32'hbc52120c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c212ed6),
	.w1(32'hbb9601dd),
	.w2(32'hbbaba1de),
	.w3(32'hbb62c642),
	.w4(32'hbc152bb1),
	.w5(32'hbb820c97),
	.w6(32'hbc388525),
	.w7(32'hbb736985),
	.w8(32'hbaaf44f9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2761),
	.w1(32'h3ba9b84c),
	.w2(32'hbc00ddd1),
	.w3(32'hbc1857e8),
	.w4(32'hbadc0a32),
	.w5(32'hbc28919b),
	.w6(32'h3a5d7896),
	.w7(32'hb953c90a),
	.w8(32'h3abf27c8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb22a1),
	.w1(32'h3ac4cbb2),
	.w2(32'h3a046046),
	.w3(32'hba8b8126),
	.w4(32'h3b9f80e7),
	.w5(32'h3c139bbb),
	.w6(32'h3afaf0b9),
	.w7(32'h3afaecae),
	.w8(32'h3ac1a127),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3481a6),
	.w1(32'hbbf09e24),
	.w2(32'hbbdfb194),
	.w3(32'h3b5baa4d),
	.w4(32'hba7c5d40),
	.w5(32'hb85c5373),
	.w6(32'h3b875391),
	.w7(32'h3b2384f5),
	.w8(32'h3b53b7e3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9784d8),
	.w1(32'h3b86ba01),
	.w2(32'hbb21312b),
	.w3(32'h3ad49104),
	.w4(32'hbb6bbefe),
	.w5(32'hba121611),
	.w6(32'h3bb17105),
	.w7(32'h38c6965c),
	.w8(32'h3b88b1f8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ae01d),
	.w1(32'h3bb78b7e),
	.w2(32'hb6aa16e6),
	.w3(32'h3bb23832),
	.w4(32'h3b0e2d33),
	.w5(32'h3a7edd9b),
	.w6(32'h3bab7630),
	.w7(32'h3c0b08a3),
	.w8(32'h3bbf1407),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba184f6),
	.w1(32'h3b12d090),
	.w2(32'h3ba8712e),
	.w3(32'h3b93da51),
	.w4(32'h3c131367),
	.w5(32'h3c80e4fe),
	.w6(32'hbacf7afc),
	.w7(32'hbb8069b2),
	.w8(32'hbbaaadb4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b832baf),
	.w1(32'hbb95ed38),
	.w2(32'h3b892045),
	.w3(32'hb9ac8fe0),
	.w4(32'h3c3b3ac8),
	.w5(32'h3ca40737),
	.w6(32'hbbb331e8),
	.w7(32'hbc3803d1),
	.w8(32'hbbf546ae),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32aac8),
	.w1(32'hbc005559),
	.w2(32'hbb999769),
	.w3(32'hbc04c055),
	.w4(32'hbbee5605),
	.w5(32'hba7d0cc6),
	.w6(32'hbc027ffa),
	.w7(32'hbb8ec1bb),
	.w8(32'hbbcacc2c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15d124),
	.w1(32'hba74d4cb),
	.w2(32'h3aa2ab8a),
	.w3(32'hbbbea79a),
	.w4(32'hbb84d3b8),
	.w5(32'hbbb6f9e2),
	.w6(32'hbb8e9347),
	.w7(32'hbb19ab1e),
	.w8(32'h3bcff36c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea8387),
	.w1(32'hbb8fdfef),
	.w2(32'hbb3b8bb3),
	.w3(32'hbc12d039),
	.w4(32'h3b929e43),
	.w5(32'h3b4b5ede),
	.w6(32'hbaeee6c0),
	.w7(32'hbb0ad9c2),
	.w8(32'hba477e86),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad3938),
	.w1(32'hbba704d9),
	.w2(32'hba123edd),
	.w3(32'h3b562c8e),
	.w4(32'h3b6412b1),
	.w5(32'h3af459ae),
	.w6(32'hbaab0002),
	.w7(32'h3b55b82d),
	.w8(32'hb984eff7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01da4e),
	.w1(32'hbadedfbf),
	.w2(32'hbbf039d9),
	.w3(32'hbb660d9c),
	.w4(32'hbb51e997),
	.w5(32'h3c70fae8),
	.w6(32'hbad2ed09),
	.w7(32'hbb85c4c9),
	.w8(32'hbc4d391a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69bec2),
	.w1(32'hbb4e7b49),
	.w2(32'h3b77056c),
	.w3(32'h3b575463),
	.w4(32'h3c7ba99c),
	.w5(32'h3c59beb9),
	.w6(32'hbc3203ef),
	.w7(32'hbbf643a1),
	.w8(32'hbba071bc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c287bfb),
	.w1(32'h3a50dbce),
	.w2(32'hbabeff29),
	.w3(32'h3acd5927),
	.w4(32'h3bb5223f),
	.w5(32'h3baab4bc),
	.w6(32'hbb5f2e7c),
	.w7(32'hb99bd437),
	.w8(32'h3a1e1068),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad9bf9),
	.w1(32'hbb95b85f),
	.w2(32'hbb47d482),
	.w3(32'h3b6b03ca),
	.w4(32'h3afb5163),
	.w5(32'hb8e9a519),
	.w6(32'hbb325ec0),
	.w7(32'h3b9b0a9e),
	.w8(32'h3b822edd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc3258),
	.w1(32'h3bee4959),
	.w2(32'h39e7b303),
	.w3(32'hbaaf96cf),
	.w4(32'hba26a8c5),
	.w5(32'h3abe70b6),
	.w6(32'hbad8e671),
	.w7(32'h3b32f5f8),
	.w8(32'h3b32f994),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b094694),
	.w1(32'h3be31071),
	.w2(32'h3bdbdb96),
	.w3(32'hbb147388),
	.w4(32'hbaf3ab28),
	.w5(32'hbb838b17),
	.w6(32'h3afe2267),
	.w7(32'h3b00eebc),
	.w8(32'h3a2920fb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbddd66),
	.w1(32'h3aa790ec),
	.w2(32'h3b799841),
	.w3(32'hba44fc25),
	.w4(32'h3c0573a6),
	.w5(32'hbb819d3a),
	.w6(32'h3b1b2a29),
	.w7(32'hbac05f2f),
	.w8(32'hbbd96faa),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03e35d),
	.w1(32'hbb0da717),
	.w2(32'h3a30ea35),
	.w3(32'hbbfd9029),
	.w4(32'h3bd995b3),
	.w5(32'h3c05e6d5),
	.w6(32'hbc07c907),
	.w7(32'hbb585731),
	.w8(32'hbb705e73),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854eec),
	.w1(32'h3c440113),
	.w2(32'h3ca231ef),
	.w3(32'h3b57bb81),
	.w4(32'hbb62207a),
	.w5(32'hbba464f0),
	.w6(32'h3b60466a),
	.w7(32'h3b06870c),
	.w8(32'h3a007eea),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e4695),
	.w1(32'h3ac1ab30),
	.w2(32'hbb86e109),
	.w3(32'hba8d6fce),
	.w4(32'h3a8d5431),
	.w5(32'hba477111),
	.w6(32'hb8c67303),
	.w7(32'h39812903),
	.w8(32'hbb61ad27),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7316a4),
	.w1(32'hbb683954),
	.w2(32'hbb74f64a),
	.w3(32'h3af06783),
	.w4(32'h3c42c05b),
	.w5(32'h3c10b684),
	.w6(32'h3a952988),
	.w7(32'hbbd494d8),
	.w8(32'hbc0cdbdb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb8170),
	.w1(32'hbb0c4823),
	.w2(32'hbae86926),
	.w3(32'hbbf348e3),
	.w4(32'hbb930ab6),
	.w5(32'hbb4b0ce5),
	.w6(32'h3aa32a94),
	.w7(32'h3b10023c),
	.w8(32'hbabea011),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba227b6),
	.w1(32'h3bb2aa7b),
	.w2(32'h3b1ab1b7),
	.w3(32'hbb2ad686),
	.w4(32'hbb97e933),
	.w5(32'hbacb55b4),
	.w6(32'hbb7b3a7a),
	.w7(32'hbb54ee26),
	.w8(32'h3a8248e7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b247be9),
	.w1(32'h3a84c966),
	.w2(32'hbb57ecfa),
	.w3(32'h3bcc99eb),
	.w4(32'h39de62ef),
	.w5(32'h3af29249),
	.w6(32'h3a6d72f1),
	.w7(32'h3a94e085),
	.w8(32'h3bc42ef4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989ae26),
	.w1(32'h39df5dc6),
	.w2(32'h3b00ede4),
	.w3(32'h3b82a5b4),
	.w4(32'h3a25520d),
	.w5(32'hb7cf32cd),
	.w6(32'h3bbaf71b),
	.w7(32'h39623bb6),
	.w8(32'h3b08a2df),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2d07c),
	.w1(32'hbacce17f),
	.w2(32'h3acb736a),
	.w3(32'hba07ace1),
	.w4(32'hbb3e4228),
	.w5(32'hbbab1ff3),
	.w6(32'h3b050c0c),
	.w7(32'hbb161dca),
	.w8(32'hbb2b5bb4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa240f1),
	.w1(32'h3b27f20e),
	.w2(32'hbb2da386),
	.w3(32'hbba1ed48),
	.w4(32'hbabbb9d6),
	.w5(32'hbb658583),
	.w6(32'hba82c8ad),
	.w7(32'h3a9367f3),
	.w8(32'hba93e0ee),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0284c9),
	.w1(32'h3ac79a56),
	.w2(32'h3b0862d7),
	.w3(32'hba0419e9),
	.w4(32'h3bbeca44),
	.w5(32'hbb6af09c),
	.w6(32'hbb7b7b9b),
	.w7(32'h3b2417fb),
	.w8(32'h3b5a36dd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19a52f),
	.w1(32'h3a7440bc),
	.w2(32'hb9b580e5),
	.w3(32'hbb320b40),
	.w4(32'hbb16c609),
	.w5(32'hbb3b1d3c),
	.w6(32'h3ae8d145),
	.w7(32'hba3fd4fd),
	.w8(32'hbbc9954b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8d397),
	.w1(32'hb93b49e2),
	.w2(32'hbb471168),
	.w3(32'hbb8290ce),
	.w4(32'hba80ec6c),
	.w5(32'hbc03cebb),
	.w6(32'hbbb7e999),
	.w7(32'hbb018b82),
	.w8(32'hbb115c67),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24069b),
	.w1(32'hbb92ff6d),
	.w2(32'hbc31c68a),
	.w3(32'h3a352a3f),
	.w4(32'h3b91a25a),
	.w5(32'h3b4d3449),
	.w6(32'hbb0681e0),
	.w7(32'h3b67149f),
	.w8(32'h3adc338c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab031a),
	.w1(32'hbb87b20e),
	.w2(32'hbb3bd912),
	.w3(32'h3b698b49),
	.w4(32'hbc2910ce),
	.w5(32'hbb8db7b8),
	.w6(32'h3b4656af),
	.w7(32'hbb6e5be5),
	.w8(32'hbb2b78cd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1f4f),
	.w1(32'hbaa92f04),
	.w2(32'h3acda79f),
	.w3(32'hbc0e29bd),
	.w4(32'h3b8b4332),
	.w5(32'hbba5da27),
	.w6(32'hba829601),
	.w7(32'h3a516496),
	.w8(32'hbba25119),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb4edf),
	.w1(32'h3a8be7d3),
	.w2(32'hbb61fdca),
	.w3(32'hba829eb4),
	.w4(32'h3b9ce0b9),
	.w5(32'h3a448c92),
	.w6(32'h3b5a3907),
	.w7(32'h3bbadad3),
	.w8(32'hbb188fbe),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995c015),
	.w1(32'h3b5d0e35),
	.w2(32'h3b0d0dd8),
	.w3(32'h3bde0e92),
	.w4(32'h397b4260),
	.w5(32'h3b5b0522),
	.w6(32'h3b5ef3b7),
	.w7(32'hba9db7e2),
	.w8(32'h3b8851c1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaec8dc),
	.w1(32'hba9724a6),
	.w2(32'hbb3cee36),
	.w3(32'hbb74e957),
	.w4(32'hbba7b47f),
	.w5(32'hbbae979e),
	.w6(32'hbb064e41),
	.w7(32'hbb744d06),
	.w8(32'hbb5f16f1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0310f7),
	.w1(32'hbb2331bd),
	.w2(32'hbbd6f850),
	.w3(32'hb9f51586),
	.w4(32'h3aea3f2b),
	.w5(32'hbbd5a636),
	.w6(32'hb94252fb),
	.w7(32'h3b1c58f3),
	.w8(32'h3a88744f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a5432),
	.w1(32'hbae3436d),
	.w2(32'h3a7a6aad),
	.w3(32'hbc16a3b0),
	.w4(32'hbb0fe146),
	.w5(32'hba200e34),
	.w6(32'hbbd8abdf),
	.w7(32'hbaf70204),
	.w8(32'hbbd243a0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e4750),
	.w1(32'hbb2b463c),
	.w2(32'hbb8023f1),
	.w3(32'hbb6cde2e),
	.w4(32'hbb9372db),
	.w5(32'hbb5bb72d),
	.w6(32'hbb207e62),
	.w7(32'h3b8f5476),
	.w8(32'h3baa0412),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910ba51),
	.w1(32'h3a8ab712),
	.w2(32'hbb3cfafa),
	.w3(32'hbbb2e009),
	.w4(32'hbbc48f37),
	.w5(32'hbc491470),
	.w6(32'h3c0f2575),
	.w7(32'hbb46debd),
	.w8(32'hbb990024),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aa7bd),
	.w1(32'hba01e5d0),
	.w2(32'hbb4122df),
	.w3(32'hbb8d8858),
	.w4(32'h3b3fa4f6),
	.w5(32'h3b96f890),
	.w6(32'hbba322a8),
	.w7(32'h3be1e705),
	.w8(32'h38ce93ec),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbd727),
	.w1(32'hb89f4664),
	.w2(32'hba123fed),
	.w3(32'hbaa79211),
	.w4(32'h3abe4f36),
	.w5(32'h3992fcd8),
	.w6(32'h3a829e20),
	.w7(32'h3b513d38),
	.w8(32'h3b12cba8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab728d0),
	.w1(32'hbbbdba38),
	.w2(32'hbc480b07),
	.w3(32'hba22b5cc),
	.w4(32'hbb488ac6),
	.w5(32'hbc399199),
	.w6(32'h3b830093),
	.w7(32'hba7ee120),
	.w8(32'hbb584755),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2287a2),
	.w1(32'hbbd5da9f),
	.w2(32'h3ad4c90a),
	.w3(32'hb7113c26),
	.w4(32'h3ba71419),
	.w5(32'h3bcf7352),
	.w6(32'hba800a4b),
	.w7(32'hbad41b2e),
	.w8(32'hbb4cb4f4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0474c3),
	.w1(32'h3b214b1b),
	.w2(32'hbaac7a39),
	.w3(32'h3b9ec825),
	.w4(32'h3bb71bfb),
	.w5(32'h3a2f5889),
	.w6(32'hba97f6a8),
	.w7(32'h3b9dd7ac),
	.w8(32'h3b024fd4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999672b),
	.w1(32'hbb272e7f),
	.w2(32'hb9bdec93),
	.w3(32'h3ac8354f),
	.w4(32'hbaa15b77),
	.w5(32'hbb911d7c),
	.w6(32'h3b9b5ea2),
	.w7(32'h3a4f05df),
	.w8(32'hbb028a41),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e2473),
	.w1(32'h3ba5a5b4),
	.w2(32'hbb7ae2d8),
	.w3(32'hbb7e07cb),
	.w4(32'hbc295a18),
	.w5(32'hbc7e0467),
	.w6(32'h3abf677c),
	.w7(32'hbaa9606b),
	.w8(32'hb9a2119f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbde7a8),
	.w1(32'h3b27da43),
	.w2(32'hb9c81ad5),
	.w3(32'h3a136060),
	.w4(32'hb9baccdc),
	.w5(32'h3b6a424f),
	.w6(32'hbb3f54c0),
	.w7(32'hbb71ff3f),
	.w8(32'hba5963d8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b924ab8),
	.w1(32'h3c260e68),
	.w2(32'h3a7ff624),
	.w3(32'h3b48db25),
	.w4(32'hb9905b4f),
	.w5(32'h3b941a4b),
	.w6(32'h3b1dc383),
	.w7(32'hbbd491a8),
	.w8(32'hbb93ca99),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0271e1),
	.w1(32'h3a5e2a6c),
	.w2(32'hbb850c0c),
	.w3(32'hbb39a840),
	.w4(32'hbbcb9db3),
	.w5(32'hbc1b4f8c),
	.w6(32'h3a63066c),
	.w7(32'hbbde7447),
	.w8(32'h3a34694b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fae7),
	.w1(32'hbb7f48a4),
	.w2(32'hbb698d67),
	.w3(32'hb93a7db1),
	.w4(32'h3909ea2e),
	.w5(32'h38c4f682),
	.w6(32'h386c2c7f),
	.w7(32'hbbd75dfe),
	.w8(32'hbb8e0536),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a3324),
	.w1(32'h3b7d50fe),
	.w2(32'hbab20b20),
	.w3(32'hbb9ef4d7),
	.w4(32'h3a2c432e),
	.w5(32'hbbaaf80b),
	.w6(32'hbad45d79),
	.w7(32'hbb00cc84),
	.w8(32'hba85c6db),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71280b),
	.w1(32'h3ad61184),
	.w2(32'hbadb1222),
	.w3(32'hba2835e7),
	.w4(32'hba056a08),
	.w5(32'h3b29a7dd),
	.w6(32'hbb96bedf),
	.w7(32'hbb090adb),
	.w8(32'hbb6e8623),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917fafc),
	.w1(32'hbb93cc73),
	.w2(32'hbbb64d9b),
	.w3(32'h39757643),
	.w4(32'hbaddf325),
	.w5(32'hbb0ac41a),
	.w6(32'hbb6b6ab5),
	.w7(32'h3a5c63d6),
	.w8(32'h3b0348d8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec56c0),
	.w1(32'h3b48e19a),
	.w2(32'h3c618cd3),
	.w3(32'hb82b89b4),
	.w4(32'h3abcd536),
	.w5(32'h3a9967ac),
	.w6(32'h3b7604c5),
	.w7(32'hba315d95),
	.w8(32'hbb8a6173),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf598fd),
	.w1(32'hbac2e9c1),
	.w2(32'hbb013250),
	.w3(32'hbb6203b5),
	.w4(32'hbb560809),
	.w5(32'hbc0489c9),
	.w6(32'hbb7440d9),
	.w7(32'h3b000b64),
	.w8(32'hbb5d0640),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd83b78),
	.w1(32'h3b875360),
	.w2(32'h3b7467e1),
	.w3(32'hbbaaa0b2),
	.w4(32'hba9fda9b),
	.w5(32'h3aabd7e7),
	.w6(32'hbb728c76),
	.w7(32'h392f8cf8),
	.w8(32'hbb632f51),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dd8b9),
	.w1(32'h3bd7bc91),
	.w2(32'hba5288c1),
	.w3(32'h3b85d172),
	.w4(32'h394deec5),
	.w5(32'hbb71acb1),
	.w6(32'hbbd52dd5),
	.w7(32'hbaaef5e2),
	.w8(32'hbb88006f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab790eb),
	.w1(32'hbab73488),
	.w2(32'hbaf44be5),
	.w3(32'h3b9c9726),
	.w4(32'hbaf38333),
	.w5(32'hb8a96dee),
	.w6(32'hbb027bd1),
	.w7(32'h3ac058fd),
	.w8(32'h388096b7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e9968),
	.w1(32'h3accf220),
	.w2(32'h3a94a2af),
	.w3(32'hbba24049),
	.w4(32'hbb2ad72d),
	.w5(32'hbb81ff60),
	.w6(32'hbb6da250),
	.w7(32'hbb1d1c01),
	.w8(32'hba919cde),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4def17),
	.w1(32'hbb6ac27a),
	.w2(32'hbb4162a4),
	.w3(32'hbadf5796),
	.w4(32'hbbb62d13),
	.w5(32'hbbe6b185),
	.w6(32'h3aa55279),
	.w7(32'h3b61ba6b),
	.w8(32'h3aff84d1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1bdfc),
	.w1(32'hba957bbc),
	.w2(32'hbbdb5749),
	.w3(32'hbaf917d8),
	.w4(32'hbb673f5f),
	.w5(32'hbc388d03),
	.w6(32'h3bce13d0),
	.w7(32'h3bce2545),
	.w8(32'h3a93c698),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb3a24),
	.w1(32'hba278311),
	.w2(32'hbb9590a7),
	.w3(32'hbba38949),
	.w4(32'h3aa78888),
	.w5(32'hbb645aa3),
	.w6(32'h3b60ccd7),
	.w7(32'hbb9a3740),
	.w8(32'h3a1b59c3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b246254),
	.w1(32'hbbe2bab8),
	.w2(32'hbb6c60a0),
	.w3(32'hba9734eb),
	.w4(32'h3b78dd31),
	.w5(32'hbba0cc27),
	.w6(32'h3ae15dad),
	.w7(32'h3b945951),
	.w8(32'h3ad57f13),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa959e),
	.w1(32'hba7fafb9),
	.w2(32'hbb0514eb),
	.w3(32'hbb54deff),
	.w4(32'h3935ad9f),
	.w5(32'h39f87cd7),
	.w6(32'hbaa050f6),
	.w7(32'hbad07d7e),
	.w8(32'hba6d933b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fbcd6),
	.w1(32'hbab3363d),
	.w2(32'h3a62718d),
	.w3(32'hbb7d2454),
	.w4(32'hbab103b2),
	.w5(32'h3a878d9c),
	.w6(32'hbb5edc6f),
	.w7(32'h3aafd463),
	.w8(32'h3af98f79),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50e904),
	.w1(32'hbbb96140),
	.w2(32'hbbc416ea),
	.w3(32'hba3fa865),
	.w4(32'hbac2943d),
	.w5(32'hba712e52),
	.w6(32'hb8dc6ec4),
	.w7(32'hbb924a48),
	.w8(32'h3a8cb385),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d8ee8),
	.w1(32'h3b1c53a2),
	.w2(32'hba5535ba),
	.w3(32'hbab7eb1d),
	.w4(32'h3b6babb7),
	.w5(32'hbb462eef),
	.w6(32'hbba94334),
	.w7(32'h3b64e13c),
	.w8(32'h3ba59ccf),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2bcf),
	.w1(32'h3b8b33be),
	.w2(32'h3be9b2ed),
	.w3(32'h3b3bffdd),
	.w4(32'hbb0f9f5d),
	.w5(32'hbb68eabe),
	.w6(32'h3add1bee),
	.w7(32'h3a13e956),
	.w8(32'h3bc16cd0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2a0ac),
	.w1(32'h3b9c1175),
	.w2(32'hbb11c119),
	.w3(32'hba971bf4),
	.w4(32'hbb4898d4),
	.w5(32'hbc1d7f0e),
	.w6(32'h3a5e5be4),
	.w7(32'hba2d7f3e),
	.w8(32'h3a42d737),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ea0eb),
	.w1(32'hba822b53),
	.w2(32'hba5010e4),
	.w3(32'h3ba1417e),
	.w4(32'h3a894433),
	.w5(32'hbb836045),
	.w6(32'h3a3acae3),
	.w7(32'hbc19cdc4),
	.w8(32'hbc01f896),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c353a),
	.w1(32'h3b8e68ac),
	.w2(32'hbb7d4999),
	.w3(32'hbbc67dbf),
	.w4(32'h3b03c51f),
	.w5(32'h39ece7f8),
	.w6(32'hbba84f32),
	.w7(32'h3a2a08c2),
	.w8(32'h3a173c97),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7504),
	.w1(32'h3b827588),
	.w2(32'h3b9603ad),
	.w3(32'h3a8c9989),
	.w4(32'h3bbbc0d4),
	.w5(32'h3a650b70),
	.w6(32'h3a2d82d6),
	.w7(32'h3bdcd823),
	.w8(32'h3b9da6e6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cafe4),
	.w1(32'h3bd84a45),
	.w2(32'hbbcc928a),
	.w3(32'hba165482),
	.w4(32'hbb9583ac),
	.w5(32'hbbbb42e7),
	.w6(32'h3b10042f),
	.w7(32'h3ab069ea),
	.w8(32'h3af8d36c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb478ddb),
	.w1(32'hbb554684),
	.w2(32'h3abade7c),
	.w3(32'h3a93a85e),
	.w4(32'h3a6da640),
	.w5(32'h3bb9e04f),
	.w6(32'hbb0f6584),
	.w7(32'hba1d31de),
	.w8(32'hbb4eb517),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fcc61),
	.w1(32'hbb36add0),
	.w2(32'hbbb1738c),
	.w3(32'h3baca2ed),
	.w4(32'hbab25de0),
	.w5(32'hbb4659e7),
	.w6(32'hbb96d904),
	.w7(32'h36f680e4),
	.w8(32'h3afad71c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd2aff),
	.w1(32'hb869e463),
	.w2(32'h3a2023e7),
	.w3(32'hbbfc6d7f),
	.w4(32'h3b811a33),
	.w5(32'hba69d582),
	.w6(32'h3a2561dc),
	.w7(32'hbb59ab9a),
	.w8(32'h3a1cb3c3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb43465),
	.w1(32'h3bb9f736),
	.w2(32'h3c1a9d3c),
	.w3(32'hbb98c158),
	.w4(32'hbbaa56a2),
	.w5(32'hbb8f18e0),
	.w6(32'hba9d0819),
	.w7(32'hbc11dc6d),
	.w8(32'hbbdcaa41),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dedc6),
	.w1(32'h3c47beb4),
	.w2(32'h3c31bf7b),
	.w3(32'hbb3b9f08),
	.w4(32'h3bef88c8),
	.w5(32'h3c76d53a),
	.w6(32'hbadfceb7),
	.w7(32'h3b118c33),
	.w8(32'h3ba8715b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4af91),
	.w1(32'h385f627a),
	.w2(32'h3be4b840),
	.w3(32'h3bafabbc),
	.w4(32'hba8a1432),
	.w5(32'h3cff6608),
	.w6(32'hbb87b394),
	.w7(32'h3bc8cca1),
	.w8(32'h3c70dae4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab23b25),
	.w1(32'hbb85c201),
	.w2(32'hbbe03788),
	.w3(32'h3c2da7f4),
	.w4(32'hbb5c763f),
	.w5(32'hbb8e24d7),
	.w6(32'h3b2c7082),
	.w7(32'h3ad65852),
	.w8(32'hbb5c5ec2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b994d03),
	.w1(32'hbc34cf30),
	.w2(32'hbc9a7a45),
	.w3(32'hbbd41185),
	.w4(32'hbc732008),
	.w5(32'hbc9095b5),
	.w6(32'hbbcd808f),
	.w7(32'hbc66ed68),
	.w8(32'hbcabe1cf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8356d3),
	.w1(32'hbbfc8872),
	.w2(32'hbc4c76e1),
	.w3(32'hbc6125f0),
	.w4(32'hbd0c891d),
	.w5(32'hbd2aac03),
	.w6(32'hbc2a76f0),
	.w7(32'hbc5c1905),
	.w8(32'hbc66e2f9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25c5bb),
	.w1(32'h39fcf953),
	.w2(32'h3af4aff0),
	.w3(32'hbcfa2e9c),
	.w4(32'hbc0c56b2),
	.w5(32'hbb02199c),
	.w6(32'hbc4cae21),
	.w7(32'hbbe0b1a9),
	.w8(32'hbc0bbfc0),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b656fe7),
	.w1(32'h3b336e3d),
	.w2(32'hbb80caf1),
	.w3(32'hbaa7ed08),
	.w4(32'h3b006b2e),
	.w5(32'hbc09bcf0),
	.w6(32'hbbaca49a),
	.w7(32'hbb7cc59a),
	.w8(32'h3bbd8f14),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39950c3e),
	.w1(32'hbca67e35),
	.w2(32'hbcbd5377),
	.w3(32'h3aa8ca69),
	.w4(32'hbc9f8bb3),
	.w5(32'hbc355b7e),
	.w6(32'h3be41ece),
	.w7(32'hbc0ba6b4),
	.w8(32'hbce32bf2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2264eb),
	.w1(32'h3baa2c70),
	.w2(32'h3b29379b),
	.w3(32'hbc81b408),
	.w4(32'hbb5b2d4e),
	.w5(32'hbb98922d),
	.w6(32'hbcb3901b),
	.w7(32'h39405a3d),
	.w8(32'hbbe3e83b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a3ec),
	.w1(32'h3be0d61c),
	.w2(32'hbb85fb4a),
	.w3(32'hba38ac38),
	.w4(32'h3bd8146f),
	.w5(32'h3c706f39),
	.w6(32'hbc4c0672),
	.w7(32'hbc0d2eeb),
	.w8(32'h3c01db4d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43db90),
	.w1(32'h3c272885),
	.w2(32'h3c1e5e07),
	.w3(32'h3be9e048),
	.w4(32'h3c0a362d),
	.w5(32'h3bbed6af),
	.w6(32'h3ae07b51),
	.w7(32'h3c8856d6),
	.w8(32'h3c8c07a7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa0d40),
	.w1(32'hba709bcc),
	.w2(32'hb8213798),
	.w3(32'h3c7cbee6),
	.w4(32'h3b4d2fe0),
	.w5(32'h3baeec81),
	.w6(32'h3c93bec4),
	.w7(32'h3afc1a3a),
	.w8(32'h3b152648),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9078261),
	.w1(32'h3afc09bf),
	.w2(32'h3bf1987d),
	.w3(32'h3ba4151e),
	.w4(32'h3c3c3549),
	.w5(32'h3cd90106),
	.w6(32'hbac526bd),
	.w7(32'h3b0a0963),
	.w8(32'h3c8e8042),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ca39d),
	.w1(32'hba653d1c),
	.w2(32'h3a36ac2a),
	.w3(32'h3c542091),
	.w4(32'h3b37ae00),
	.w5(32'h3c2c1653),
	.w6(32'hb8cc99a4),
	.w7(32'h3aa1d040),
	.w8(32'h3c9e4d2d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6b63c),
	.w1(32'h3ba0ce5c),
	.w2(32'hbb4244d8),
	.w3(32'h3a1c0675),
	.w4(32'h399d5708),
	.w5(32'h3b889ca3),
	.w6(32'hbb395c92),
	.w7(32'hbb89a1c2),
	.w8(32'h3b29093f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15de57),
	.w1(32'h3aa63222),
	.w2(32'hbb37f55b),
	.w3(32'h3b0b96cd),
	.w4(32'hbab69bf8),
	.w5(32'h39f62621),
	.w6(32'h39256824),
	.w7(32'h3a8d4d07),
	.w8(32'hbb5838b5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1c2be),
	.w1(32'hbb9167ce),
	.w2(32'hbc3563d6),
	.w3(32'hbb3d7f02),
	.w4(32'hbbde6b44),
	.w5(32'hbbcf7779),
	.w6(32'hbbe0a8f4),
	.w7(32'hbb5439b7),
	.w8(32'hbc08ee31),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebe96e),
	.w1(32'hbc10ce4b),
	.w2(32'hbcad46a6),
	.w3(32'hbb928a5d),
	.w4(32'hbc42f901),
	.w5(32'hbc330354),
	.w6(32'hbc217715),
	.w7(32'hbc04d431),
	.w8(32'hbce1ffc8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ec35b),
	.w1(32'h3b1d5fb0),
	.w2(32'hbb652c48),
	.w3(32'hbc67b766),
	.w4(32'hba932ad0),
	.w5(32'hbb4822a7),
	.w6(32'hbc2b558a),
	.w7(32'hbb9e4ffc),
	.w8(32'h3c333a03),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae32311),
	.w1(32'h3a9e0c2f),
	.w2(32'h3b9a9621),
	.w3(32'h3b9270cd),
	.w4(32'h3bc40147),
	.w5(32'h3b3291f1),
	.w6(32'hba7082ef),
	.w7(32'h3932a8ee),
	.w8(32'hbc16b349),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399357d7),
	.w1(32'h3b95bdab),
	.w2(32'h3b18468b),
	.w3(32'hbaea4ce8),
	.w4(32'hbb0da72d),
	.w5(32'hbc0fbf3d),
	.w6(32'hbbab2cbc),
	.w7(32'h3b4e27b8),
	.w8(32'hbbd52541),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c605),
	.w1(32'h3bae13cf),
	.w2(32'h3c1cf52a),
	.w3(32'h397e0554),
	.w4(32'h3c18948b),
	.w5(32'h3c7af88c),
	.w6(32'h3bc991ad),
	.w7(32'h3adcc95d),
	.w8(32'hbb3480ab),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36d970),
	.w1(32'h3b8d6a1f),
	.w2(32'h3c6ddae9),
	.w3(32'h39af546b),
	.w4(32'h3c8e6ef9),
	.w5(32'h3d082fe6),
	.w6(32'hbb2351a9),
	.w7(32'h3c0b3ba9),
	.w8(32'h3ca7d389),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e8f59),
	.w1(32'hbaa1255d),
	.w2(32'hbb3fa5cf),
	.w3(32'h3c8d97c3),
	.w4(32'h3b51d05b),
	.w5(32'hbb2f8fac),
	.w6(32'h3c0943ba),
	.w7(32'h3b2effe4),
	.w8(32'h3b9841bd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a642e7b),
	.w1(32'hbb367e23),
	.w2(32'hbbb46883),
	.w3(32'h3b046a98),
	.w4(32'h3c3a6b52),
	.w5(32'h3cfdfdcf),
	.w6(32'h3bdc7a52),
	.w7(32'h3c27c8bd),
	.w8(32'h3c9697cc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedd87b),
	.w1(32'h3c2a8c1d),
	.w2(32'hbc11f041),
	.w3(32'h3c01b395),
	.w4(32'hbba39c93),
	.w5(32'hbc2a037d),
	.w6(32'h3ad850ca),
	.w7(32'hbc84f56b),
	.w8(32'hbcf3ed6d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a5bc8),
	.w1(32'hbbb10cb4),
	.w2(32'hbc052632),
	.w3(32'hbc562150),
	.w4(32'hbc3be79a),
	.w5(32'hbbd5f36e),
	.w6(32'hbc3736cd),
	.w7(32'hbc0fa919),
	.w8(32'hbc618509),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc766204),
	.w1(32'h3a4aa90f),
	.w2(32'h3acc65f8),
	.w3(32'hbbb3a62b),
	.w4(32'h3aa3892c),
	.w5(32'hbae9d6f0),
	.w6(32'hb8883e3f),
	.w7(32'hba91c3ea),
	.w8(32'h3b56a780),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beac227),
	.w1(32'hbb95f8b6),
	.w2(32'h3bb9836b),
	.w3(32'h3b819f48),
	.w4(32'h39a7fc3a),
	.w5(32'hbc098976),
	.w6(32'hba843e41),
	.w7(32'h3b8acf59),
	.w8(32'h3b2b1e41),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea69ea),
	.w1(32'h3b9fa913),
	.w2(32'hbb42a2e7),
	.w3(32'hba27dc54),
	.w4(32'h3b0b8fae),
	.w5(32'h3a5ceac0),
	.w6(32'h392a721c),
	.w7(32'hbba8ba52),
	.w8(32'hbc1d0c08),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1039),
	.w1(32'hb985a0a0),
	.w2(32'hbb8377f4),
	.w3(32'hbb9f7bc4),
	.w4(32'hbb36a9a3),
	.w5(32'hbae31276),
	.w6(32'hbac14595),
	.w7(32'hba6a82b7),
	.w8(32'h3bd37801),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4344a7),
	.w1(32'hbafdb0bd),
	.w2(32'hbc53fdcd),
	.w3(32'hbbb53884),
	.w4(32'h3ab2becd),
	.w5(32'hbb157686),
	.w6(32'h3bbe8b80),
	.w7(32'hbc1b43bd),
	.w8(32'hbb40407d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ff204),
	.w1(32'h3baccf3c),
	.w2(32'h398db68b),
	.w3(32'h3b9e2073),
	.w4(32'hbb27a8be),
	.w5(32'hb9888308),
	.w6(32'h3b98afeb),
	.w7(32'hbb6d6fb9),
	.w8(32'hbc1bfe2e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab50f15),
	.w1(32'hbb2b033f),
	.w2(32'hbb9e64fe),
	.w3(32'hbb42132f),
	.w4(32'hbb3b4eac),
	.w5(32'h3b8b9d2f),
	.w6(32'h39196b61),
	.w7(32'h3b9687cf),
	.w8(32'h3bd1cc27),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33c32f),
	.w1(32'h3bcedb4b),
	.w2(32'h3c5386f3),
	.w3(32'h3aaeb5d4),
	.w4(32'h3bbe34ae),
	.w5(32'h3d04afda),
	.w6(32'h3be30c98),
	.w7(32'hbc4b17a6),
	.w8(32'h3bde88c1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1606de),
	.w1(32'hba1bf954),
	.w2(32'hbb32799e),
	.w3(32'h3c079f24),
	.w4(32'h3878bf76),
	.w5(32'h3a1090d4),
	.w6(32'hbc358a7a),
	.w7(32'h3bb5213b),
	.w8(32'h3c08ee2a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45f213),
	.w1(32'h3b70cb59),
	.w2(32'h3c98c5b7),
	.w3(32'h3c1b145e),
	.w4(32'h3aad940f),
	.w5(32'h3a1e3c26),
	.w6(32'hbac415a3),
	.w7(32'hba94787b),
	.w8(32'hbc39d31c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27d4c7),
	.w1(32'h38a3927c),
	.w2(32'h3c41c209),
	.w3(32'hbb7eebea),
	.w4(32'h3bf291a3),
	.w5(32'h3be708fb),
	.w6(32'hbc39a5b2),
	.w7(32'h3be0e5b7),
	.w8(32'h3b1fd148),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccaad7),
	.w1(32'h3b10ab04),
	.w2(32'h3a6cea65),
	.w3(32'hbb554447),
	.w4(32'h3b9f8aa9),
	.w5(32'h3d0234cf),
	.w6(32'h3b94e20d),
	.w7(32'hbb5c94a4),
	.w8(32'h3b83d60e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f5885),
	.w1(32'h3b802e2f),
	.w2(32'h3b4ea301),
	.w3(32'h3c4c939a),
	.w4(32'h3c02ee15),
	.w5(32'h3d078b16),
	.w6(32'h3bb86aaf),
	.w7(32'hbb762efc),
	.w8(32'h3b2bca78),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfabe6),
	.w1(32'h3b689e15),
	.w2(32'h3c0313b9),
	.w3(32'h3c6eea91),
	.w4(32'h398d10ce),
	.w5(32'h3c1e47e9),
	.w6(32'h3be9d193),
	.w7(32'h3b931a80),
	.w8(32'h39e304ce),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd9ef6),
	.w1(32'hbb0d1e0b),
	.w2(32'h37621f24),
	.w3(32'h3b4fb1a2),
	.w4(32'hbc09e6a1),
	.w5(32'h3b7b373b),
	.w6(32'hb87f9f5d),
	.w7(32'h3b01b265),
	.w8(32'hba05286f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a5e9c),
	.w1(32'hbb74c870),
	.w2(32'hbc9c090e),
	.w3(32'h3b3cfd77),
	.w4(32'hbc3cccdb),
	.w5(32'hbccf4b50),
	.w6(32'hbbcb5f6f),
	.w7(32'hbc26018b),
	.w8(32'hbc21552e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bebcc),
	.w1(32'h3ad75fad),
	.w2(32'h3a71dd75),
	.w3(32'hbc4854b5),
	.w4(32'h3a29dfde),
	.w5(32'hbbd6b20b),
	.w6(32'h392c8cf3),
	.w7(32'hbbc32371),
	.w8(32'hbc3aaf12),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9688),
	.w1(32'hba3d9d11),
	.w2(32'h3b44fb4b),
	.w3(32'hbab87bf9),
	.w4(32'h3acbf16c),
	.w5(32'h3b9ece85),
	.w6(32'hbb11183b),
	.w7(32'h3ad162a6),
	.w8(32'h3bcd654f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f953b),
	.w1(32'hbb63f0a5),
	.w2(32'hbc30ebca),
	.w3(32'h3bca556c),
	.w4(32'hbb3e5246),
	.w5(32'hbb2d7cde),
	.w6(32'hb96020fc),
	.w7(32'h3a66b148),
	.w8(32'h3b2eb978),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1338b),
	.w1(32'h3c29cf59),
	.w2(32'h3c5ac8a3),
	.w3(32'hba35bd3e),
	.w4(32'h3beb4bc1),
	.w5(32'h3a6f1d6d),
	.w6(32'hba9374d3),
	.w7(32'hbbf92e3f),
	.w8(32'hbc4cdfc7),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80c3a4),
	.w1(32'h3c162263),
	.w2(32'h3c418fd4),
	.w3(32'h3b80b165),
	.w4(32'h3c31840f),
	.w5(32'h3c186c6f),
	.w6(32'h3ad2f993),
	.w7(32'hba951c77),
	.w8(32'h3c192e8b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e6ca7),
	.w1(32'hbc57d4db),
	.w2(32'hbcfa6224),
	.w3(32'h3c457414),
	.w4(32'hbc90d68b),
	.w5(32'hbc0369f5),
	.w6(32'hbb3736cf),
	.w7(32'hbcc94fda),
	.w8(32'hbd34138d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc993d95),
	.w1(32'hbb9129a9),
	.w2(32'hbb61d80a),
	.w3(32'hbc9497d5),
	.w4(32'hba9b01d5),
	.w5(32'h3b38fe87),
	.w6(32'hbcf96f71),
	.w7(32'h3b82ed9c),
	.w8(32'h3c2f112f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77f475),
	.w1(32'h3b3452b3),
	.w2(32'hb9eafc37),
	.w3(32'h3adf0d6b),
	.w4(32'h3c3ad076),
	.w5(32'h3b08c21d),
	.w6(32'hbb0f7f86),
	.w7(32'h3baf1ae8),
	.w8(32'h3c696221),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82dbc1),
	.w1(32'h3bf437f4),
	.w2(32'h3bd124c0),
	.w3(32'h3c1740c4),
	.w4(32'h3aea41c2),
	.w5(32'h3a1b54a4),
	.w6(32'hb9612b9d),
	.w7(32'h3b7b722a),
	.w8(32'h3b855005),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88ea8),
	.w1(32'h390e9c1f),
	.w2(32'h3ad38d94),
	.w3(32'h3b13ecb3),
	.w4(32'h3a7fb51f),
	.w5(32'h3b2c7e61),
	.w6(32'h3a302145),
	.w7(32'h3b3d58fc),
	.w8(32'hbb052135),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62ed80),
	.w1(32'h3b85ce78),
	.w2(32'h3b180cf8),
	.w3(32'hbb0a05ae),
	.w4(32'h3b8b5504),
	.w5(32'h3a31acc8),
	.w6(32'h3bc7bf32),
	.w7(32'h3ab69de1),
	.w8(32'h3b80dd3c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad65f51),
	.w1(32'h3b4512d7),
	.w2(32'h3c3d3157),
	.w3(32'h3b3785c7),
	.w4(32'h3bd9523e),
	.w5(32'h3d06f8d8),
	.w6(32'h3bc23db5),
	.w7(32'h3bb6e2b2),
	.w8(32'h3c86fb52),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8148b7),
	.w1(32'hbacaf472),
	.w2(32'h3abc9c0e),
	.w3(32'h3c02781d),
	.w4(32'h3ba6b7cb),
	.w5(32'h3c959a51),
	.w6(32'h3ba98f25),
	.w7(32'hbaaa097f),
	.w8(32'h3b412125),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c078e27),
	.w1(32'h3aa7f450),
	.w2(32'h3b9234c4),
	.w3(32'h3bf1ec86),
	.w4(32'h3a7a1ce7),
	.w5(32'h3bd05333),
	.w6(32'hbc22ee85),
	.w7(32'hbbadef05),
	.w8(32'hbc06f405),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4719dc),
	.w1(32'h3bdae4dc),
	.w2(32'h3bd7964d),
	.w3(32'h3c10f1c6),
	.w4(32'hbb954466),
	.w5(32'hbb01b6ba),
	.w6(32'hba0692fc),
	.w7(32'hbb8659c3),
	.w8(32'h3b8e5b1a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule