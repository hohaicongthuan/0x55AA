module layer_8_featuremap_70(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a782fb1),
	.w1(32'hba476f1a),
	.w2(32'hbb9a005c),
	.w3(32'hbab92735),
	.w4(32'hbb6a8106),
	.w5(32'hbbbf6dc9),
	.w6(32'h3ac4b1cf),
	.w7(32'hbafc0764),
	.w8(32'h3b8b28f2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e5459),
	.w1(32'hb9cb8649),
	.w2(32'hbb53b4ed),
	.w3(32'h3a91c348),
	.w4(32'hbb516a2d),
	.w5(32'hbb87b359),
	.w6(32'h3b36d72c),
	.w7(32'h39bfaafc),
	.w8(32'h3b51c5a7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b029b83),
	.w1(32'hba466c95),
	.w2(32'hbb69ed73),
	.w3(32'h3850729e),
	.w4(32'hbb36dc3b),
	.w5(32'hbb89c676),
	.w6(32'h3ab41682),
	.w7(32'hba8d7122),
	.w8(32'hbbb32aa2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb7d07),
	.w1(32'h3b4770c1),
	.w2(32'hbb37a7a8),
	.w3(32'h3bcc8cc9),
	.w4(32'h3bbeeda3),
	.w5(32'h3b1de1d4),
	.w6(32'hba1a7a5d),
	.w7(32'h3a8cf2bd),
	.w8(32'h3b571af2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefe218),
	.w1(32'hbb122cfa),
	.w2(32'hbbd42eb8),
	.w3(32'hb98f1cee),
	.w4(32'hbb87de75),
	.w5(32'hbc196fed),
	.w6(32'h3aad2057),
	.w7(32'hbad517c3),
	.w8(32'h3d372a14),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce81a3e),
	.w1(32'h3a6ec542),
	.w2(32'hbd01996e),
	.w3(32'h3c2851bc),
	.w4(32'hbcaeb68f),
	.w5(32'hbd33ee26),
	.w6(32'h3cca6b48),
	.w7(32'hbb03933d),
	.w8(32'h3b65d544),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1e53b),
	.w1(32'hbaacb2ce),
	.w2(32'hbb9fa1fb),
	.w3(32'h3a835b37),
	.w4(32'hbb56bfa5),
	.w5(32'hbba0af37),
	.w6(32'h3ad15ec9),
	.w7(32'hbadc06e4),
	.w8(32'h3b46ab0b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae03b0),
	.w1(32'hbb273f3d),
	.w2(32'hbbcfbc7f),
	.w3(32'hba53eb3d),
	.w4(32'hbb8faee6),
	.w5(32'hbc227523),
	.w6(32'h3abb0d58),
	.w7(32'hbab02bb7),
	.w8(32'h3b9a4cae),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b317305),
	.w1(32'hbb0b88b7),
	.w2(32'hbbbf154d),
	.w3(32'h3a773742),
	.w4(32'hbba5cb1e),
	.w5(32'hbbdfccda),
	.w6(32'h3b196b6b),
	.w7(32'hba178613),
	.w8(32'hbbffba5a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa49c1d),
	.w1(32'hb9df563e),
	.w2(32'h3c4d961c),
	.w3(32'h3bdd671b),
	.w4(32'h3c1dd44e),
	.w5(32'h3b79a51c),
	.w6(32'hbb0de826),
	.w7(32'h3b8eeaf5),
	.w8(32'h3b02d28b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a493d6b),
	.w1(32'hbb7f9d51),
	.w2(32'hbbf008a9),
	.w3(32'hba9cca2f),
	.w4(32'hbb83bbed),
	.w5(32'hbbee9499),
	.w6(32'hb9a77cfb),
	.w7(32'hbb642709),
	.w8(32'h3b843e33),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b307c40),
	.w1(32'hba376d48),
	.w2(32'hbb9f64f0),
	.w3(32'h39fcb5af),
	.w4(32'hbb7d2338),
	.w5(32'hbbbcb4aa),
	.w6(32'h3b093582),
	.w7(32'hbaa4d905),
	.w8(32'h3abfd651),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5713c2),
	.w1(32'hbb412854),
	.w2(32'hbbc74224),
	.w3(32'h3a595b02),
	.w4(32'hbb6e4c1f),
	.w5(32'hbba49134),
	.w6(32'h38bff65d),
	.w7(32'hbadf64d0),
	.w8(32'h3d4dd221),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d014d3f),
	.w1(32'h3a8210ac),
	.w2(32'hbd113915),
	.w3(32'h3c445eea),
	.w4(32'hbcc09adc),
	.w5(32'hbd461ecf),
	.w6(32'h3ce40e42),
	.w7(32'hbaf9a093),
	.w8(32'h3cca9aea),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81d2c0),
	.w1(32'h3aa17063),
	.w2(32'hbc954a59),
	.w3(32'h3b985186),
	.w4(32'hbc4b05f9),
	.w5(32'hbcdebfbc),
	.w6(32'h3c71c59f),
	.w7(32'hbb0d47dc),
	.w8(32'h3a8327ac),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28d466),
	.w1(32'hbb0d9050),
	.w2(32'hbae115ce),
	.w3(32'hba5e454a),
	.w4(32'hbb22afa2),
	.w5(32'hba8788b0),
	.w6(32'h3aa79bb2),
	.w7(32'h3a9a7348),
	.w8(32'h3b0a247b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5df34),
	.w1(32'h3b96ec0a),
	.w2(32'h3ab1d26c),
	.w3(32'hba1bfa60),
	.w4(32'h3a1b7df1),
	.w5(32'hbb983bd7),
	.w6(32'h3b529c50),
	.w7(32'hb9473ad6),
	.w8(32'hba3ddea9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c53dac),
	.w1(32'hbb08a9e1),
	.w2(32'hbb93262c),
	.w3(32'h3a8df97f),
	.w4(32'hbb162e7a),
	.w5(32'hbb162f09),
	.w6(32'hbabf7762),
	.w7(32'hbaa4b615),
	.w8(32'hbb03e549),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb458e74),
	.w1(32'hbbbbd481),
	.w2(32'hbb9f7828),
	.w3(32'hbab045c2),
	.w4(32'hbbd23f4e),
	.w5(32'hbbfc3ea2),
	.w6(32'h3985f2c3),
	.w7(32'h3b87d099),
	.w8(32'hbcc103e7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1fba2),
	.w1(32'hbbb640ad),
	.w2(32'hbcb993f4),
	.w3(32'hbbb997b0),
	.w4(32'hbc8e6fdc),
	.w5(32'hbc93a30a),
	.w6(32'hbb9fc6d3),
	.w7(32'hbc202eff),
	.w8(32'hbca275d6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b1009),
	.w1(32'hb8b22889),
	.w2(32'h3c37928f),
	.w3(32'hbb927367),
	.w4(32'h3c1a58ba),
	.w5(32'h3c8e62c4),
	.w6(32'hbc1b4527),
	.w7(32'h39ba00ea),
	.w8(32'h3bd2aec6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85803c),
	.w1(32'hbade8b20),
	.w2(32'hbc13e9fb),
	.w3(32'h3a5905f0),
	.w4(32'hbbba3441),
	.w5(32'hbc46ecde),
	.w6(32'h3b492076),
	.w7(32'hbb34825b),
	.w8(32'hbd17caa1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7340b),
	.w1(32'hba913d39),
	.w2(32'h3ce05ad6),
	.w3(32'hbb93b3c8),
	.w4(32'h3cb73731),
	.w5(32'h3d3c3cf8),
	.w6(32'hbca367b9),
	.w7(32'h3b98ed2a),
	.w8(32'hbb09a9d2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb907972),
	.w1(32'hbaa0d1d3),
	.w2(32'hbafd14e2),
	.w3(32'hbb864a31),
	.w4(32'hbb89db7c),
	.w5(32'hbb2d4037),
	.w6(32'hba0b9830),
	.w7(32'h3a8289c8),
	.w8(32'hbc4995cd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156650),
	.w1(32'hbc22542b),
	.w2(32'h3bb567c4),
	.w3(32'h39da2510),
	.w4(32'h3b18200e),
	.w5(32'h3c3e5a4f),
	.w6(32'hbc268f00),
	.w7(32'h3b15c3f3),
	.w8(32'hbd0e42f8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca7833),
	.w1(32'hba95ab67),
	.w2(32'h3cd22cf1),
	.w3(32'hbb8daba0),
	.w4(32'h3caa4dd6),
	.w5(32'h3d304824),
	.w6(32'hbc9a13af),
	.w7(32'h3b8ccd6b),
	.w8(32'hbcf36228),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad638f),
	.w1(32'hba8b15c3),
	.w2(32'h3cb367af),
	.w3(32'hbb78922b),
	.w4(32'h3c912d5e),
	.w5(32'h3d168cbc),
	.w6(32'hbc84c74c),
	.w7(32'h3b6a5fbd),
	.w8(32'hbc990253),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fa9bc),
	.w1(32'h385746d8),
	.w2(32'h3c79e53a),
	.w3(32'hbb1a483a),
	.w4(32'h3c4069e3),
	.w5(32'h3ca30a24),
	.w6(32'hbc00a7b5),
	.w7(32'h3b87f27d),
	.w8(32'hbc4dd9fc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bb7ef),
	.w1(32'hbc0dfa43),
	.w2(32'hba86548f),
	.w3(32'hbc14797a),
	.w4(32'hbc14d121),
	.w5(32'h3a8b67a9),
	.w6(32'hbc513b80),
	.w7(32'hbbe2ef29),
	.w8(32'h3b57245f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20ec93),
	.w1(32'hb974a481),
	.w2(32'hbb5c1b9e),
	.w3(32'h3a2c7511),
	.w4(32'hbb2291fe),
	.w5(32'hbb86ff6c),
	.w6(32'h3af717af),
	.w7(32'hba3494c5),
	.w8(32'hbc335315),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc070000),
	.w1(32'hbbb0575a),
	.w2(32'hbc1b6e41),
	.w3(32'hbc3d43c4),
	.w4(32'hbb30bd12),
	.w5(32'h3b720f24),
	.w6(32'hbc0525ec),
	.w7(32'hbc44cc33),
	.w8(32'hbd0b5b0b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6b400),
	.w1(32'hbba5999f),
	.w2(32'h3c95350b),
	.w3(32'hbc002dc4),
	.w4(32'h3c4ea065),
	.w5(32'h3cfc0a18),
	.w6(32'hbc94faea),
	.w7(32'h3aa9ec54),
	.w8(32'hbc1c0cb4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc337fe5),
	.w1(32'hbb42f69c),
	.w2(32'hbc004db0),
	.w3(32'hbbe75c4d),
	.w4(32'hbb7d15bc),
	.w5(32'hbb4e572e),
	.w6(32'hbc252745),
	.w7(32'hbbfd982a),
	.w8(32'hbb49e2f9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f14d8),
	.w1(32'h3ae3a654),
	.w2(32'hbbe0b8fd),
	.w3(32'hbaa949a4),
	.w4(32'hbb57f4c3),
	.w5(32'hba6eac25),
	.w6(32'hbb4cdd67),
	.w7(32'hbbae45c5),
	.w8(32'h3d348c98),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce2e70d),
	.w1(32'h3a5f7259),
	.w2(32'hbcfedba5),
	.w3(32'h3c2b4e89),
	.w4(32'hbca9733a),
	.w5(32'hbd2e12c4),
	.w6(32'h3cc7dfe5),
	.w7(32'hbaded373),
	.w8(32'hba25e4f1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e4e1b),
	.w1(32'hbb4db5ed),
	.w2(32'hbba3d601),
	.w3(32'hbaf89e71),
	.w4(32'hbbae6149),
	.w5(32'hbbb036d4),
	.w6(32'h392b229f),
	.w7(32'h3a8baa38),
	.w8(32'hbc9e8a32),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59b7ca),
	.w1(32'hbbe84c93),
	.w2(32'h3c09b921),
	.w3(32'hbb589353),
	.w4(32'h3bcab6c0),
	.w5(32'h3c3e69a6),
	.w6(32'hbc2d92c0),
	.w7(32'h3b029077),
	.w8(32'h3ba93134),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62587b),
	.w1(32'hb9741e13),
	.w2(32'hbb8d03c9),
	.w3(32'h39e44c7b),
	.w4(32'hbb538731),
	.w5(32'hbbc0787f),
	.w6(32'h3b346286),
	.w7(32'hba908ded),
	.w8(32'h3d1e838e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc80648),
	.w1(32'h3b3a0a52),
	.w2(32'hbced04cc),
	.w3(32'h3be143ed),
	.w4(32'hbca18797),
	.w5(32'hbd3ad996),
	.w6(32'h3cc63705),
	.w7(32'hbb7f76d5),
	.w8(32'hbcb3116d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81482e),
	.w1(32'hbb649821),
	.w2(32'h3c4f4ba6),
	.w3(32'hbb8c4bfe),
	.w4(32'h3c1a5836),
	.w5(32'h3c9b9664),
	.w6(32'hbc335154),
	.w7(32'h3b209cc8),
	.w8(32'hbc70c31d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29ff58),
	.w1(32'hb9c29cf4),
	.w2(32'h3c32d3c5),
	.w3(32'hbaf2903b),
	.w4(32'h3c1051a5),
	.w5(32'h3c9385e5),
	.w6(32'hbc01ba17),
	.w7(32'h3ae9b583),
	.w8(32'hb931c478),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ed313),
	.w1(32'hb8ef27d7),
	.w2(32'hb9cd9ee1),
	.w3(32'h399f7c9e),
	.w4(32'hb82b360f),
	.w5(32'hb9f6a832),
	.w6(32'h38f588f5),
	.w7(32'h391cbcf0),
	.w8(32'h3935b9fc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c840d),
	.w1(32'hbb86e52f),
	.w2(32'hbaa5e40f),
	.w3(32'hba97ad6a),
	.w4(32'hbb95d32a),
	.w5(32'hb98b82e0),
	.w6(32'hbb446ae2),
	.w7(32'hbb3aa4c2),
	.w8(32'hb9ec1bc5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1d29d),
	.w1(32'hb805c8ba),
	.w2(32'hb98d06dc),
	.w3(32'h39972d55),
	.w4(32'hb91e6d1b),
	.w5(32'hba09bcd2),
	.w6(32'hb8b85cf8),
	.w7(32'h389d7b8a),
	.w8(32'h39967c56),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398eb557),
	.w1(32'h39a665cd),
	.w2(32'h38d5ebcf),
	.w3(32'h39cf629f),
	.w4(32'h3995f535),
	.w5(32'h38095e4d),
	.w6(32'h3a0e2b78),
	.w7(32'h39dcc884),
	.w8(32'hb85e032e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31d878),
	.w1(32'h3a788d39),
	.w2(32'hb9215325),
	.w3(32'h39f76af5),
	.w4(32'h399f1d4f),
	.w5(32'hb98038ed),
	.w6(32'h3a058fdc),
	.w7(32'h39c2e2e8),
	.w8(32'h3a41f549),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9ed00),
	.w1(32'h3a9050a4),
	.w2(32'h3ac5798c),
	.w3(32'hb842065d),
	.w4(32'hbad29b4d),
	.w5(32'h3aebb437),
	.w6(32'hbb044e34),
	.w7(32'hba6efb58),
	.w8(32'hb97f97ae),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ca9ae),
	.w1(32'hba561dee),
	.w2(32'hb94e7dbe),
	.w3(32'hba662f4c),
	.w4(32'hb9b71395),
	.w5(32'hb8295b4a),
	.w6(32'hba2bd347),
	.w7(32'hb9a2e1fc),
	.w8(32'h38c90ca3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c458d0),
	.w1(32'h38d2e6dd),
	.w2(32'h3940d098),
	.w3(32'h3a6f4704),
	.w4(32'h3a95e7f6),
	.w5(32'h3aa59adc),
	.w6(32'h39831dea),
	.w7(32'h391da6a0),
	.w8(32'h39843545),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fb846),
	.w1(32'h3a06cec7),
	.w2(32'h390e567f),
	.w3(32'h39ee2bc5),
	.w4(32'h39e5dbe5),
	.w5(32'h393e3775),
	.w6(32'h3a0de1fb),
	.w7(32'h39c766f4),
	.w8(32'hb99fb086),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96161d1),
	.w1(32'hb9ac81c2),
	.w2(32'hb9b25f13),
	.w3(32'h38d46688),
	.w4(32'hb9182b36),
	.w5(32'hb9eba91e),
	.w6(32'hb9171419),
	.w7(32'hb747ac6d),
	.w8(32'hba6cb901),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0a221),
	.w1(32'hba2c9a7c),
	.w2(32'hba7268e6),
	.w3(32'h38013a37),
	.w4(32'hb9be1f59),
	.w5(32'hba6f358f),
	.w6(32'hb9c53b81),
	.w7(32'hb8bfd597),
	.w8(32'hbb235384),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8483a),
	.w1(32'h3a6398ca),
	.w2(32'h3a411ad4),
	.w3(32'hbb86f5ef),
	.w4(32'hb8bf7388),
	.w5(32'hb8f1e6cc),
	.w6(32'h3a897d3e),
	.w7(32'hb96e51e0),
	.w8(32'hba0c38f0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38652a),
	.w1(32'hba249ed9),
	.w2(32'h397a4e48),
	.w3(32'hb9940432),
	.w4(32'hb98046d8),
	.w5(32'h39fa34ce),
	.w6(32'hb9bdd04a),
	.w7(32'h39cdec93),
	.w8(32'h3a361750),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e965c),
	.w1(32'hbab3fd1f),
	.w2(32'hba54590e),
	.w3(32'hba9a66e2),
	.w4(32'hbab16f3b),
	.w5(32'h394afd50),
	.w6(32'hbb3ef482),
	.w7(32'hbafaac8e),
	.w8(32'hba2c2a22),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82ffcc),
	.w1(32'h3aa0e875),
	.w2(32'hbb51a0f7),
	.w3(32'hb9f9e72c),
	.w4(32'hbab22a1e),
	.w5(32'hbb2a7961),
	.w6(32'hba3e9b48),
	.w7(32'hbb1b153a),
	.w8(32'hba427e9b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89968f5),
	.w1(32'h3af5913d),
	.w2(32'h38d15e66),
	.w3(32'h39bc7d25),
	.w4(32'hba0eefa3),
	.w5(32'h379e177d),
	.w6(32'hba344799),
	.w7(32'hb9b9b608),
	.w8(32'h3a0b117c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad84109),
	.w1(32'hbb1c460e),
	.w2(32'hb99eeb4e),
	.w3(32'hba72104d),
	.w4(32'hba828f8f),
	.w5(32'hba8b35de),
	.w6(32'hbb4f9438),
	.w7(32'hb9bf3895),
	.w8(32'h3a5ea389),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a81c06),
	.w1(32'hb865ff6c),
	.w2(32'h39f1facb),
	.w3(32'h3aaad493),
	.w4(32'h3a88c8d3),
	.w5(32'h3ab2463b),
	.w6(32'h3a16f990),
	.w7(32'h3a4c96fb),
	.w8(32'hbb37b5c8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e4261),
	.w1(32'hbab51b08),
	.w2(32'hba962596),
	.w3(32'hbb1eecbe),
	.w4(32'hba96d297),
	.w5(32'hbb13411d),
	.w6(32'hbb095217),
	.w7(32'hbb0f1184),
	.w8(32'h39bf78dc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add72fa),
	.w1(32'h39ff6579),
	.w2(32'h3a15953f),
	.w3(32'hba98ff8a),
	.w4(32'hbaa0d039),
	.w5(32'hbb065369),
	.w6(32'hb990aef6),
	.w7(32'hba5be646),
	.w8(32'hba8104f8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bf9df),
	.w1(32'h39b86bc3),
	.w2(32'h3815ed13),
	.w3(32'hba82e0cd),
	.w4(32'hb9fb25a8),
	.w5(32'hb9951b81),
	.w6(32'hb9493ee7),
	.w7(32'hb893876e),
	.w8(32'h3846a931),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e451b1),
	.w1(32'hb919c918),
	.w2(32'hb971a8ea),
	.w3(32'h3a714460),
	.w4(32'h3941f69b),
	.w5(32'hb9895226),
	.w6(32'h3962664a),
	.w7(32'h3a005258),
	.w8(32'hbb27c4bc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba169c54),
	.w1(32'hbb250fcb),
	.w2(32'hba4c3708),
	.w3(32'hbb509011),
	.w4(32'hbb890105),
	.w5(32'hbb2c4b83),
	.w6(32'hbb3a67fa),
	.w7(32'hbb0e7a56),
	.w8(32'hb8f3d416),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861edf0),
	.w1(32'hb936d982),
	.w2(32'hba0aba9b),
	.w3(32'h39f8ebe8),
	.w4(32'hb9488270),
	.w5(32'hba3a655c),
	.w6(32'hb7087827),
	.w7(32'hb941ca91),
	.w8(32'hb9b9a204),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ba465),
	.w1(32'hb946640f),
	.w2(32'hb9bc4291),
	.w3(32'hb8a91914),
	.w4(32'hb9a5eb18),
	.w5(32'hb9fb2e84),
	.w6(32'hb984f08f),
	.w7(32'hb94218b7),
	.w8(32'hba04376d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986d457),
	.w1(32'hb9b005eb),
	.w2(32'hb9c29d25),
	.w3(32'hb6a975d4),
	.w4(32'hb956feed),
	.w5(32'hb9f148df),
	.w6(32'hb979bd8e),
	.w7(32'hb90ae7b4),
	.w8(32'hb8f80b38),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2a470),
	.w1(32'hbb09a5c3),
	.w2(32'hbacd9ebc),
	.w3(32'hbae42c74),
	.w4(32'hbac1af11),
	.w5(32'hba7fc5cc),
	.w6(32'hba2bb271),
	.w7(32'hbac3a0df),
	.w8(32'h3921f6c2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6b635),
	.w1(32'h39cd223d),
	.w2(32'h395f85af),
	.w3(32'h39a2779e),
	.w4(32'h39873d3c),
	.w5(32'h3901e6a4),
	.w6(32'h39f5454d),
	.w7(32'h39ad65b6),
	.w8(32'h3a993497),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e40936),
	.w1(32'hb8b615e7),
	.w2(32'h39fb57e1),
	.w3(32'h3a8ca10e),
	.w4(32'h3a006eb4),
	.w5(32'h3a6dcd8f),
	.w6(32'h3a407b82),
	.w7(32'h3aa17cdb),
	.w8(32'hba0deb15),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9579780),
	.w1(32'hb978ffa0),
	.w2(32'hb9d89cbd),
	.w3(32'h39c5b19e),
	.w4(32'hb881ae8c),
	.w5(32'hba10b988),
	.w6(32'hb9322066),
	.w7(32'h37b72966),
	.w8(32'h39be712c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a143d88),
	.w1(32'h3a277596),
	.w2(32'h3998340e),
	.w3(32'h39dc6baf),
	.w4(32'h3a0c0eb0),
	.w5(32'h3974a59c),
	.w6(32'h3a2613d5),
	.w7(32'h39ec7c80),
	.w8(32'hba2dc6e3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be633a),
	.w1(32'hb9ad92f9),
	.w2(32'hba2141f7),
	.w3(32'h394fdbf7),
	.w4(32'hb9153787),
	.w5(32'hba55728f),
	.w6(32'hb990b825),
	.w7(32'hb8db3a97),
	.w8(32'hba59e1b5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20ee97),
	.w1(32'hbafd002b),
	.w2(32'hba44a447),
	.w3(32'hbb54e625),
	.w4(32'hba2b4642),
	.w5(32'hb9120a4b),
	.w6(32'h3a76b3da),
	.w7(32'hbaa1ea0e),
	.w8(32'hba1fb9b5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cbf51),
	.w1(32'hb8bb874e),
	.w2(32'hb9a4aaa3),
	.w3(32'hb9f3e7a4),
	.w4(32'hb8d1c6b2),
	.w5(32'hba023139),
	.w6(32'h398780d0),
	.w7(32'h3868a802),
	.w8(32'hb9da7b7e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf0941),
	.w1(32'hb9103611),
	.w2(32'hb99312bb),
	.w3(32'h396454a6),
	.w4(32'hb8e08cfd),
	.w5(32'hb9f76343),
	.w6(32'hb94537fb),
	.w7(32'h3790f71c),
	.w8(32'hb9b46ea7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa68c9),
	.w1(32'hb8bc47da),
	.w2(32'hb9ad831a),
	.w3(32'h38f34739),
	.w4(32'hb881e712),
	.w5(32'hb9ab7022),
	.w6(32'h38081e45),
	.w7(32'h36a29aaa),
	.w8(32'h3abeb262),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed9a85),
	.w1(32'hb92d6c0b),
	.w2(32'h3a1e6d9d),
	.w3(32'h3ac12b01),
	.w4(32'h3a3ef0ff),
	.w5(32'h3a96aca4),
	.w6(32'h3a577224),
	.w7(32'h3ab46556),
	.w8(32'h3a3ef250),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39888607),
	.w1(32'hb850aa46),
	.w2(32'h3972d5ad),
	.w3(32'h3a515413),
	.w4(32'h3923b4f6),
	.w5(32'h39982a69),
	.w6(32'h39a5c86e),
	.w7(32'h3a66a3a9),
	.w8(32'hb84e3b4c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6417a),
	.w1(32'h390ab32a),
	.w2(32'hb9217052),
	.w3(32'h373ff48d),
	.w4(32'hb9cf0da3),
	.w5(32'hb9576928),
	.w6(32'h37a6cfba),
	.w7(32'hb9b2611a),
	.w8(32'hbb0559d7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadacb7f),
	.w1(32'hbb57f765),
	.w2(32'hbb4c6e79),
	.w3(32'hbb85e709),
	.w4(32'hbae0869f),
	.w5(32'hb9cff766),
	.w6(32'hbb80fce6),
	.w7(32'hbba92aef),
	.w8(32'hb9b875ad),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b5e8c),
	.w1(32'h38e1f735),
	.w2(32'hb91e74de),
	.w3(32'h391658a7),
	.w4(32'hb8e708e5),
	.w5(32'hb9189314),
	.w6(32'h38fdd5c1),
	.w7(32'h3915d8ac),
	.w8(32'h39c335cd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02ed02),
	.w1(32'h3aacf318),
	.w2(32'h3a06f78b),
	.w3(32'h39a10765),
	.w4(32'h3a66d621),
	.w5(32'h3a0e905c),
	.w6(32'h3a133a5b),
	.w7(32'h39b8250f),
	.w8(32'hbaf03ded),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93e83b),
	.w1(32'h3bd0c386),
	.w2(32'h3b97915e),
	.w3(32'hb9b74450),
	.w4(32'h3b21761c),
	.w5(32'h3b0f34ab),
	.w6(32'h3b3df77f),
	.w7(32'h3affe37a),
	.w8(32'hb90b2c0f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d719b6),
	.w1(32'h392bcdab),
	.w2(32'h3997cc14),
	.w3(32'h3a074737),
	.w4(32'h399a7aaf),
	.w5(32'h3985ac17),
	.w6(32'h39a9a207),
	.w7(32'h3a5dd22f),
	.w8(32'h387bfdc3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9496a),
	.w1(32'h38d2e66b),
	.w2(32'hb89945a2),
	.w3(32'h398e4e2b),
	.w4(32'h393d855e),
	.w5(32'hb723359a),
	.w6(32'h39c69a1e),
	.w7(32'h39b33a50),
	.w8(32'h39856e00),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38284c31),
	.w1(32'h39101727),
	.w2(32'h39869b89),
	.w3(32'h3a9cfdfb),
	.w4(32'h3ac6014e),
	.w5(32'h3adcbdec),
	.w6(32'h39a56cdd),
	.w7(32'h39516e35),
	.w8(32'h3a426254),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a089432),
	.w1(32'h39a099e3),
	.w2(32'h394a568f),
	.w3(32'h39bc230d),
	.w4(32'h39ba1ace),
	.w5(32'h38bcb679),
	.w6(32'h39b1df86),
	.w7(32'h38efd65b),
	.w8(32'hbb33f9f9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43b809),
	.w1(32'hbb02c20f),
	.w2(32'hbae32d9c),
	.w3(32'hbb6cf8f2),
	.w4(32'hbb510c64),
	.w5(32'hbb006a9d),
	.w6(32'hbb4a66ba),
	.w7(32'hbb593e16),
	.w8(32'h397f21a8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387144b7),
	.w1(32'h392f0835),
	.w2(32'h398d85c8),
	.w3(32'h3a977598),
	.w4(32'h3abee2e2),
	.w5(32'h3ad32a2f),
	.w6(32'h39af2dfb),
	.w7(32'h3960bc0c),
	.w8(32'h396404ea),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f0942),
	.w1(32'h38e7ff37),
	.w2(32'h394cc2ef),
	.w3(32'h3a82a2cb),
	.w4(32'h3a9ee20b),
	.w5(32'h3ab0d948),
	.w6(32'h3984eab2),
	.w7(32'h39274c21),
	.w8(32'hba7241c9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ddaa3),
	.w1(32'hba505f95),
	.w2(32'hb83cd19d),
	.w3(32'hb9b9a1b7),
	.w4(32'hba2fa6a2),
	.w5(32'hb925c763),
	.w6(32'hba4be520),
	.w7(32'h3858bb63),
	.w8(32'h37f4a77d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba949690),
	.w1(32'h3a1e9066),
	.w2(32'h3aad126e),
	.w3(32'hbaae1805),
	.w4(32'hba7934ff),
	.w5(32'h3a8a2d2e),
	.w6(32'h3a869c1c),
	.w7(32'h39b3919b),
	.w8(32'hb93bb92c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9251cb9),
	.w1(32'hb951f516),
	.w2(32'hb97739c3),
	.w3(32'h382dd536),
	.w4(32'hb8a271f9),
	.w5(32'hb990e256),
	.w6(32'hb8ec7669),
	.w7(32'hb7106aa4),
	.w8(32'hbaaf25a8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c0878),
	.w1(32'h3a458d8a),
	.w2(32'hb96c806b),
	.w3(32'hbac6b134),
	.w4(32'hbabf8501),
	.w5(32'hbaa25025),
	.w6(32'hbaaa5bcc),
	.w7(32'hba857c48),
	.w8(32'hbaceb5db),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2fc6f),
	.w1(32'hba197dce),
	.w2(32'hb9cfbf7e),
	.w3(32'hb8a9e2cf),
	.w4(32'hba5f38ef),
	.w5(32'hba9ce9fb),
	.w6(32'hba0f6c72),
	.w7(32'h3947c8a6),
	.w8(32'h39ba3648),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb009b9a),
	.w1(32'hbb5e2fe3),
	.w2(32'hbb107b19),
	.w3(32'hba9be275),
	.w4(32'hbb0ae7c5),
	.w5(32'hbae43aae),
	.w6(32'hba4e5540),
	.w7(32'hba29bbbb),
	.w8(32'hb9fa12d4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac59d1),
	.w1(32'h3b8174fa),
	.w2(32'h3b10c4c8),
	.w3(32'hbaf1d767),
	.w4(32'hbaaa11de),
	.w5(32'hba14e7d8),
	.w6(32'h3afb262e),
	.w7(32'hba8ec098),
	.w8(32'h3aa6a8c9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2a3ec),
	.w1(32'hb96d52b7),
	.w2(32'h3a083fdd),
	.w3(32'h3a9cd2b3),
	.w4(32'h3a136178),
	.w5(32'h3a80977f),
	.w6(32'h3a229d42),
	.w7(32'h3a9727ce),
	.w8(32'h3a4597d5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a568f59),
	.w1(32'h3a4ad2a5),
	.w2(32'h391e7227),
	.w3(32'h3a50662b),
	.w4(32'h39b8e4b4),
	.w5(32'hb648cc39),
	.w6(32'h3a1b03ae),
	.w7(32'h398ddea7),
	.w8(32'hbad12116),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d3b5c),
	.w1(32'hba910d6e),
	.w2(32'hb9975dc7),
	.w3(32'hbab86c17),
	.w4(32'hba5b9c36),
	.w5(32'hba4cc4b1),
	.w6(32'hbaefeeda),
	.w7(32'hba612c7d),
	.w8(32'hb9e4f553),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c91ce),
	.w1(32'hb9c9d380),
	.w2(32'hb9e4dc81),
	.w3(32'h393c924f),
	.w4(32'hb9099b51),
	.w5(32'hba08bb9a),
	.w6(32'hb92061db),
	.w7(32'h37633894),
	.w8(32'h3af8258a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34adc5),
	.w1(32'h3867f7eb),
	.w2(32'h3a37c7ba),
	.w3(32'h3afe509c),
	.w4(32'h3a12929b),
	.w5(32'h3a894ea7),
	.w6(32'h3a25922b),
	.w7(32'h3b04afae),
	.w8(32'hbae751d5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbd09b),
	.w1(32'hba8c4340),
	.w2(32'hb9dc7766),
	.w3(32'hba81acf7),
	.w4(32'hbaa3cf6c),
	.w5(32'hba417494),
	.w6(32'hbabd0d23),
	.w7(32'hb9d9aaa6),
	.w8(32'h38e780fc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b215c2),
	.w1(32'h38628296),
	.w2(32'h38a5b2f7),
	.w3(32'h39c916c9),
	.w4(32'h3a067459),
	.w5(32'h3a1645d7),
	.w6(32'h38b108ae),
	.w7(32'h37ebcf38),
	.w8(32'h36f25ccb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882396d),
	.w1(32'h388ea648),
	.w2(32'hb77fb493),
	.w3(32'h37d5f0e6),
	.w4(32'h383d3d4d),
	.w5(32'h3803f228),
	.w6(32'h38c37d9a),
	.w7(32'h38bb5ab2),
	.w8(32'hb81e21f2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865a580),
	.w1(32'h38998b77),
	.w2(32'h3840e017),
	.w3(32'h38b20c76),
	.w4(32'h3891a008),
	.w5(32'h380a83f4),
	.w6(32'h38966c27),
	.w7(32'h3880b0f5),
	.w8(32'h37d84318),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5995345),
	.w1(32'h37353129),
	.w2(32'h37547291),
	.w3(32'h3734601e),
	.w4(32'h379e9f3d),
	.w5(32'h37c57633),
	.w6(32'h37851b15),
	.w7(32'h37d964a2),
	.w8(32'h37fdf01d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5fb2395),
	.w1(32'hb6e06896),
	.w2(32'hb72b1f99),
	.w3(32'hb7210954),
	.w4(32'hb74f014e),
	.w5(32'hb72fe445),
	.w6(32'hb77eee12),
	.w7(32'hb7328e5c),
	.w8(32'hb6cbb9d1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a4ba1c),
	.w1(32'h37444359),
	.w2(32'h36670c1c),
	.w3(32'h38620827),
	.w4(32'h37f588fb),
	.w5(32'h3771f565),
	.w6(32'h37fb9512),
	.w7(32'h37c02d4b),
	.w8(32'h37797494),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8048e3e),
	.w1(32'hb7e29700),
	.w2(32'hb6cedf6d),
	.w3(32'hb706a971),
	.w4(32'hb687f722),
	.w5(32'hb64ee5e7),
	.w6(32'hb8189486),
	.w7(32'hb82d63b3),
	.w8(32'hb8192c5b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aa7216),
	.w1(32'hb7fa27d0),
	.w2(32'hb7d12051),
	.w3(32'hb7666017),
	.w4(32'hb734d465),
	.w5(32'hb6a1d2b7),
	.w6(32'hb7eb002c),
	.w7(32'hb8058fba),
	.w8(32'hb7afe62d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37844bc6),
	.w1(32'h36a40e24),
	.w2(32'h37870ab1),
	.w3(32'hb72c4b34),
	.w4(32'hb741235a),
	.w5(32'h37b59aed),
	.w6(32'hb739e454),
	.w7(32'hb5fe2de5),
	.w8(32'h3798f9c1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d45ba7),
	.w1(32'h36347318),
	.w2(32'hb43056e6),
	.w3(32'hb606d3c2),
	.w4(32'hb251b4a2),
	.w5(32'hb61b5c37),
	.w6(32'h34ca2561),
	.w7(32'h33c3891d),
	.w8(32'hb5b227af),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h353ec556),
	.w1(32'h370f6edb),
	.w2(32'h372c8973),
	.w3(32'h377364d0),
	.w4(32'h379c3c5b),
	.w5(32'h370a1dd2),
	.w6(32'h377909bf),
	.w7(32'h373afb73),
	.w8(32'hb7104335),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366a9179),
	.w1(32'h36e1c60e),
	.w2(32'h360ac98a),
	.w3(32'h37cd31d5),
	.w4(32'h37f6d1b3),
	.w5(32'h369d6b4a),
	.w6(32'h376eb785),
	.w7(32'h376da7ac),
	.w8(32'h355ee886),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63cef59),
	.w1(32'hb7282960),
	.w2(32'hb6ca43d1),
	.w3(32'h36b2bc6c),
	.w4(32'h36ac0b32),
	.w5(32'h37192bad),
	.w6(32'hb7cbd6be),
	.w7(32'hb7994b17),
	.w8(32'hb751eafa),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373d05a7),
	.w1(32'h382dca1c),
	.w2(32'h3773ff87),
	.w3(32'h37e510cc),
	.w4(32'h38536485),
	.w5(32'h382ed413),
	.w6(32'h38269d0b),
	.w7(32'h37e8f97e),
	.w8(32'hb7aa0fe7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb351c0a1),
	.w1(32'hb44fedf8),
	.w2(32'hb460f675),
	.w3(32'hb49561d7),
	.w4(32'hb50e9a72),
	.w5(32'h34aa31e6),
	.w6(32'h351a4f35),
	.w7(32'h34bdd5a2),
	.w8(32'h356c1783),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34d58c5d),
	.w1(32'hb5e99a86),
	.w2(32'hb50e21a6),
	.w3(32'h35a0ba58),
	.w4(32'h349cac0f),
	.w5(32'hb6298edf),
	.w6(32'h357a0e6c),
	.w7(32'hb56ef4d9),
	.w8(32'hb75d4948),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c45c68),
	.w1(32'hb70c3f2f),
	.w2(32'hb81c5a04),
	.w3(32'h3867d8c4),
	.w4(32'h385b1ae5),
	.w5(32'h3797b204),
	.w6(32'h380aa5f7),
	.w7(32'h380254a5),
	.w8(32'h374dcf93),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c66927),
	.w1(32'hb7bbddd4),
	.w2(32'hb81dfc6c),
	.w3(32'h36e37204),
	.w4(32'hb7fe1c85),
	.w5(32'hb853b7e0),
	.w6(32'hb6c1144a),
	.w7(32'hb833fdf6),
	.w8(32'hb844d370),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71c5baa),
	.w1(32'hb71a0b24),
	.w2(32'hb718f166),
	.w3(32'hb78803a5),
	.w4(32'hb76f166c),
	.w5(32'hb73eceae),
	.w6(32'hb761efca),
	.w7(32'hb7b15cb2),
	.w8(32'hb75cd86c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65426eb),
	.w1(32'hb74c1b54),
	.w2(32'hb79d45b6),
	.w3(32'hb783f5b9),
	.w4(32'hb7b25137),
	.w5(32'hb7891cb5),
	.w6(32'hb7a73345),
	.w7(32'hb7b84715),
	.w8(32'hb78e6edb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d7df2c),
	.w1(32'hb6fa0c10),
	.w2(32'hb709055c),
	.w3(32'h3694aef9),
	.w4(32'hb5863361),
	.w5(32'h3606809f),
	.w6(32'h3641ec4e),
	.w7(32'h364f3fbe),
	.w8(32'h368292f3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6be6282),
	.w1(32'h37864f68),
	.w2(32'h3584b22a),
	.w3(32'h374e8ccb),
	.w4(32'h371a6e34),
	.w5(32'h380c6278),
	.w6(32'h37d2e2eb),
	.w7(32'h380a78d1),
	.w8(32'h38171253),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75ac07a),
	.w1(32'h364d99ba),
	.w2(32'hb714640d),
	.w3(32'h361fe8b1),
	.w4(32'hb72eb315),
	.w5(32'hb80c6cb4),
	.w6(32'hb706e9fc),
	.w7(32'hb78519f2),
	.w8(32'hb82e07a6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368d03ff),
	.w1(32'hb73a914c),
	.w2(32'hb842cf25),
	.w3(32'hb77e1c1b),
	.w4(32'hb76ea738),
	.w5(32'hb7605554),
	.w6(32'hb64b09dc),
	.w7(32'hb750b4fc),
	.w8(32'hb84ce30f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule