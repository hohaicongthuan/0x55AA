module layer_10_featuremap_171(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10927d),
	.w1(32'h3b940a92),
	.w2(32'h3c71d672),
	.w3(32'hba0a1455),
	.w4(32'h39039d89),
	.w5(32'h3a030a86),
	.w6(32'h3b6a2ea1),
	.w7(32'h3b31c32d),
	.w8(32'h3abbc8e1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16bd69),
	.w1(32'h3ac3598b),
	.w2(32'h39e68d5a),
	.w3(32'h3abdb193),
	.w4(32'h39bcfa20),
	.w5(32'hb93d5bed),
	.w6(32'h3aac5434),
	.w7(32'h3a1e9796),
	.w8(32'hb9fdbc4d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de0eef),
	.w1(32'h3aa0394d),
	.w2(32'h3ad5fd15),
	.w3(32'hbab1f5aa),
	.w4(32'hbaced9f4),
	.w5(32'hbb060f40),
	.w6(32'h39dd70ac),
	.w7(32'hbaa45e44),
	.w8(32'hba5a9ed5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb0150),
	.w1(32'hbb75def7),
	.w2(32'hbbd7e560),
	.w3(32'hbb199089),
	.w4(32'h3aae4aa4),
	.w5(32'hb932c0ed),
	.w6(32'hbac706e9),
	.w7(32'hbb1fc572),
	.w8(32'hba800723),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89c4fe),
	.w1(32'h3b1411ad),
	.w2(32'hba5e87d3),
	.w3(32'hbb4db3c5),
	.w4(32'h3b74ff63),
	.w5(32'h3b323e5b),
	.w6(32'h3a5abb2d),
	.w7(32'h3a90c859),
	.w8(32'h3b2ee2cb),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f2a8),
	.w1(32'hbaf41a9f),
	.w2(32'hbb61faab),
	.w3(32'h3ae97246),
	.w4(32'hba29b6c1),
	.w5(32'hbb251d29),
	.w6(32'hbac74971),
	.w7(32'hbb033bd9),
	.w8(32'hba3aad74),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0493c),
	.w1(32'h3b328782),
	.w2(32'h39936818),
	.w3(32'hbaa5cf49),
	.w4(32'hb9c69402),
	.w5(32'hb9754da7),
	.w6(32'h3a91c2e2),
	.w7(32'hb96c317e),
	.w8(32'hbac77bbf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba690aeb),
	.w1(32'h39abffa4),
	.w2(32'hb9d492e6),
	.w3(32'hbafb6931),
	.w4(32'h3a5c57c4),
	.w5(32'h3a11332d),
	.w6(32'hb8add111),
	.w7(32'hba7a85d3),
	.w8(32'hb8b8b5c1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d8f24),
	.w1(32'hbacda7ef),
	.w2(32'h3954cd8c),
	.w3(32'h39b304ff),
	.w4(32'hbaa42263),
	.w5(32'hb97cf299),
	.w6(32'hbac23d50),
	.w7(32'hba8726ea),
	.w8(32'hba58a157),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95bbdc0),
	.w1(32'h3b2ac89d),
	.w2(32'h3b45b5c9),
	.w3(32'hb83d74c0),
	.w4(32'h3a60ed8d),
	.w5(32'h3adfee81),
	.w6(32'h3abd30ef),
	.w7(32'h39e4df37),
	.w8(32'h3ac692eb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca16c8),
	.w1(32'hbaa3d6f2),
	.w2(32'h3a275f04),
	.w3(32'hbaa06a71),
	.w4(32'h3af2e74a),
	.w5(32'h3b06a449),
	.w6(32'h3a4b640a),
	.w7(32'hb93cb366),
	.w8(32'h3a2cc6ff),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c26a4),
	.w1(32'hba9707a8),
	.w2(32'hbb17d253),
	.w3(32'h395f748a),
	.w4(32'h3b1da615),
	.w5(32'h3a962c88),
	.w6(32'hba906661),
	.w7(32'hbad193b3),
	.w8(32'hba610101),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ff6e),
	.w1(32'h38cd291f),
	.w2(32'h3a45e26d),
	.w3(32'hba4206c6),
	.w4(32'hb920f894),
	.w5(32'h3a561060),
	.w6(32'hba28d1ed),
	.w7(32'hbaafd499),
	.w8(32'h3949ae29),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd68ff),
	.w1(32'hb9dedd98),
	.w2(32'hbb000c12),
	.w3(32'h3a198820),
	.w4(32'h3aa6721b),
	.w5(32'h385e46a0),
	.w6(32'hba125905),
	.w7(32'hbb39fc1d),
	.w8(32'hbb42d3ba),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0df27d),
	.w1(32'h3b2212aa),
	.w2(32'hbb09c497),
	.w3(32'h3a78e6e1),
	.w4(32'h3c2aef18),
	.w5(32'h3c08db49),
	.w6(32'h3a147ec1),
	.w7(32'h3a04ecb0),
	.w8(32'h3b8adf08),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02507c),
	.w1(32'hba8bda09),
	.w2(32'hba043dc9),
	.w3(32'hbabe504d),
	.w4(32'hba4df4ac),
	.w5(32'h399118ea),
	.w6(32'hbaa4e856),
	.w7(32'hbaba4670),
	.w8(32'hb91eb7bd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67d397),
	.w1(32'h3a0baf4b),
	.w2(32'hba89fe0e),
	.w3(32'hb9f5339c),
	.w4(32'h39db0e48),
	.w5(32'hba894343),
	.w6(32'hba2776e1),
	.w7(32'hba9cca05),
	.w8(32'hbabeac03),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadb665),
	.w1(32'h3af935e8),
	.w2(32'h3b1eac37),
	.w3(32'h37e8c946),
	.w4(32'hba69ac5a),
	.w5(32'h3a6ac0cf),
	.w6(32'hb6bdf93d),
	.w7(32'h396e2892),
	.w8(32'hb9af4a3a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba551628),
	.w1(32'h3a853817),
	.w2(32'h39365e99),
	.w3(32'hbb23eb50),
	.w4(32'h3a81c940),
	.w5(32'h3a32262c),
	.w6(32'hba3886a5),
	.w7(32'hba962759),
	.w8(32'hba81859d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f4d84),
	.w1(32'hbad7cf4e),
	.w2(32'h39b59db9),
	.w3(32'hba8291bc),
	.w4(32'hba8ffd9c),
	.w5(32'hb99b58e2),
	.w6(32'hbad199be),
	.w7(32'hba164c11),
	.w8(32'hba715669),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba304949),
	.w1(32'hbaef8506),
	.w2(32'hbaa280fa),
	.w3(32'hb884471e),
	.w4(32'h38ae378f),
	.w5(32'h38a86bc1),
	.w6(32'hba9f158a),
	.w7(32'hba8390f9),
	.w8(32'hbac6a6b1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9212be),
	.w1(32'h3b90aca0),
	.w2(32'h3c37f9be),
	.w3(32'hb93f871c),
	.w4(32'h3926dc75),
	.w5(32'hba038a9b),
	.w6(32'h3b32028f),
	.w7(32'hbb9d66ba),
	.w8(32'h372b9d66),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf2a80),
	.w1(32'hb9d4e333),
	.w2(32'h3a8acfc0),
	.w3(32'h3bbf9b1e),
	.w4(32'hbaaa4ff9),
	.w5(32'h3a87ce1a),
	.w6(32'h3afba916),
	.w7(32'h3984daa8),
	.w8(32'h3b0fb354),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dea21),
	.w1(32'h39b60e66),
	.w2(32'h3a3116b4),
	.w3(32'h368ca9fb),
	.w4(32'h3a088c1b),
	.w5(32'h3acbb6be),
	.w6(32'h394d2058),
	.w7(32'hba6922ca),
	.w8(32'h3a0eaf6b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4f188),
	.w1(32'hbaa0837a),
	.w2(32'hb9b30b2a),
	.w3(32'h3a471d78),
	.w4(32'h3a6af61c),
	.w5(32'h3a35de16),
	.w6(32'h38edf061),
	.w7(32'h3a30af57),
	.w8(32'hb9bcadfe),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd4305),
	.w1(32'h3abec44c),
	.w2(32'h3adcd107),
	.w3(32'hb9bed63c),
	.w4(32'h3b10b2d1),
	.w5(32'h3b15ec48),
	.w6(32'hba63091d),
	.w7(32'hb9bad9f7),
	.w8(32'h3917366f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45c4bd),
	.w1(32'hba79d4a8),
	.w2(32'hb9a269df),
	.w3(32'hb9f7b1a2),
	.w4(32'hb9d7c6d8),
	.w5(32'hb913ac9b),
	.w6(32'hba8642d0),
	.w7(32'hba481ff2),
	.w8(32'hba3aac4f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93eac23),
	.w1(32'hbafc875f),
	.w2(32'hba8346fd),
	.w3(32'h398d095c),
	.w4(32'h39220c9d),
	.w5(32'hb983ee13),
	.w6(32'hba92f777),
	.w7(32'hba83d34f),
	.w8(32'hba78bdb0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb3ca8),
	.w1(32'h3aa50b40),
	.w2(32'hba5dc65c),
	.w3(32'hb9877107),
	.w4(32'h3a955235),
	.w5(32'hbae3c35b),
	.w6(32'h3b1f2dce),
	.w7(32'hba9e47ac),
	.w8(32'h390dc209),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90275f),
	.w1(32'h39c48d3d),
	.w2(32'h3ad1290f),
	.w3(32'hb9064843),
	.w4(32'h39e24b76),
	.w5(32'h3a95ce9e),
	.w6(32'h3a420c56),
	.w7(32'h39fcd658),
	.w8(32'h3acd3bc6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab45ed3),
	.w1(32'hba935305),
	.w2(32'hba7ddd78),
	.w3(32'h3a75a184),
	.w4(32'hb9b2f0e8),
	.w5(32'hba12f34d),
	.w6(32'hba4b63f6),
	.w7(32'hba440fdc),
	.w8(32'hba2e51e4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9ab12),
	.w1(32'hba5cd53d),
	.w2(32'hba41c9b0),
	.w3(32'hb9ca0be5),
	.w4(32'hb98c1e70),
	.w5(32'hb9a8f879),
	.w6(32'hba878db3),
	.w7(32'hba91e964),
	.w8(32'hba825a69),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba232a48),
	.w1(32'h39c1b466),
	.w2(32'h3b87f485),
	.w3(32'hba5393fb),
	.w4(32'h3aae53ef),
	.w5(32'hb8bafcdd),
	.w6(32'h38308922),
	.w7(32'hba702a09),
	.w8(32'hb9658aa8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95842a),
	.w1(32'h3abaa202),
	.w2(32'h3b7a6d99),
	.w3(32'h3ad19870),
	.w4(32'hb91abf19),
	.w5(32'h3b94ad70),
	.w6(32'hba2cc473),
	.w7(32'h3ae3e2c7),
	.w8(32'h394908df),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d77be1),
	.w1(32'hb9c08bef),
	.w2(32'h3ab0715a),
	.w3(32'h3a8fef02),
	.w4(32'hba879a45),
	.w5(32'hba59799b),
	.w6(32'hba6076b6),
	.w7(32'h39b1d3ce),
	.w8(32'hba9c9267),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99f183),
	.w1(32'hbabbd119),
	.w2(32'hba8b7422),
	.w3(32'hbb159b2e),
	.w4(32'hb96695bf),
	.w5(32'hba4e98e4),
	.w6(32'hba841b04),
	.w7(32'hba7a8ab9),
	.w8(32'hba6621c0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8e912),
	.w1(32'hb927402d),
	.w2(32'hbad4fe01),
	.w3(32'hb9cac974),
	.w4(32'h3a3aaf2b),
	.w5(32'h3ab41cb6),
	.w6(32'h3a5ad3a9),
	.w7(32'hb9e65d11),
	.w8(32'h394a3599),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a343e37),
	.w1(32'h3b19a8a0),
	.w2(32'h3ac35dea),
	.w3(32'h39b538ca),
	.w4(32'hba09b528),
	.w5(32'hbb158c2d),
	.w6(32'h3b88ff7f),
	.w7(32'h3a93a5f7),
	.w8(32'hbaa4a696),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d861af),
	.w1(32'hbae88ce5),
	.w2(32'hbaf1ed4e),
	.w3(32'hba76a63d),
	.w4(32'hba977d76),
	.w5(32'hbb43654f),
	.w6(32'h3a0775b1),
	.w7(32'hba3dcd38),
	.w8(32'hbb06382c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba053763),
	.w1(32'h39279215),
	.w2(32'hba133727),
	.w3(32'hb982d823),
	.w4(32'hb8719b39),
	.w5(32'h3a630053),
	.w6(32'hb9e2f167),
	.w7(32'hb8c6a6a3),
	.w8(32'hba19b363),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d79c4),
	.w1(32'h39d31c35),
	.w2(32'h3aba3b64),
	.w3(32'hba9354ca),
	.w4(32'h3a8d9a66),
	.w5(32'h3aba9fcd),
	.w6(32'h3a93614a),
	.w7(32'h3a9c6aca),
	.w8(32'h3af16fd8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9774af),
	.w1(32'hb9eee567),
	.w2(32'hb98373b1),
	.w3(32'h3ab2414e),
	.w4(32'h3a61e807),
	.w5(32'h3abc7b43),
	.w6(32'hbac29bfe),
	.w7(32'hb99fc2e9),
	.w8(32'hbb0c6b26),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa56066),
	.w1(32'hb88eab11),
	.w2(32'h39f989b7),
	.w3(32'hbaa0fad1),
	.w4(32'hba44f6a0),
	.w5(32'hb9775419),
	.w6(32'h37f9c6a8),
	.w7(32'hba6cb825),
	.w8(32'hb99a2099),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd3bf3),
	.w1(32'h3b9f53bc),
	.w2(32'h3b58d699),
	.w3(32'hba384a36),
	.w4(32'h3adabcc6),
	.w5(32'h3b0b6bf7),
	.w6(32'h3b14413e),
	.w7(32'h3ae1cfd3),
	.w8(32'h3b21cc6d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad34931),
	.w1(32'h3b728a95),
	.w2(32'h3bfd0ae5),
	.w3(32'h3a70b38d),
	.w4(32'h3a59ef31),
	.w5(32'h3a9d5391),
	.w6(32'h3b65bd5d),
	.w7(32'hb78336ad),
	.w8(32'hbabacf45),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38909d2f),
	.w1(32'h3b84bca1),
	.w2(32'h3b3c7ddd),
	.w3(32'h3aae052a),
	.w4(32'hb9a8e55c),
	.w5(32'h3aa9aa11),
	.w6(32'h3ac71810),
	.w7(32'hbae26fe2),
	.w8(32'hba24e5c5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395362c0),
	.w1(32'h383c40dd),
	.w2(32'hbb3e864f),
	.w3(32'hb951f7ed),
	.w4(32'h3bb1e74f),
	.w5(32'h3c05e3b1),
	.w6(32'h3a8a8a56),
	.w7(32'h3abc3d00),
	.w8(32'h3b278a0e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba811516),
	.w1(32'hb91f74f5),
	.w2(32'h3ad7c875),
	.w3(32'h3ac7074c),
	.w4(32'hba8be2ee),
	.w5(32'h39d07450),
	.w6(32'hba937e2a),
	.w7(32'hbad1f3c8),
	.w8(32'hba97e5ca),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa24f8),
	.w1(32'hba7a69b0),
	.w2(32'h3a1772cf),
	.w3(32'hb96591ea),
	.w4(32'hba311141),
	.w5(32'hb9b1a2b0),
	.w6(32'hba65e274),
	.w7(32'hba010a98),
	.w8(32'hba10215d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ec026d),
	.w1(32'h39f6dc2f),
	.w2(32'hba92694d),
	.w3(32'hb9322049),
	.w4(32'h3ab1513e),
	.w5(32'h3a075a6b),
	.w6(32'h3a44975d),
	.w7(32'hba0febc8),
	.w8(32'h38a29d14),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b3af5),
	.w1(32'h3b5d052a),
	.w2(32'hbaa39ca1),
	.w3(32'h3a76875a),
	.w4(32'h3a93140e),
	.w5(32'h3a3f12cf),
	.w6(32'h3a449e7f),
	.w7(32'hba6ec703),
	.w8(32'hbabdc4ca),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba488f5f),
	.w1(32'hbb5af0ca),
	.w2(32'h3a7d8e5b),
	.w3(32'hba209c17),
	.w4(32'h3a8e40b6),
	.w5(32'h3b0ac321),
	.w6(32'hbafcafee),
	.w7(32'h3b2692c6),
	.w8(32'hbb008e43),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb918885),
	.w1(32'hbaa4c420),
	.w2(32'hbb1a1091),
	.w3(32'h3aea4205),
	.w4(32'hb7f7c2ab),
	.w5(32'hba858d79),
	.w6(32'hba3c658d),
	.w7(32'hbae775b4),
	.w8(32'hba033b75),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ef0ee),
	.w1(32'h3b1e1813),
	.w2(32'hb8b61b19),
	.w3(32'hb7c61fd8),
	.w4(32'h3b0cb09c),
	.w5(32'h3b56126c),
	.w6(32'hb93cdb09),
	.w7(32'h3a7106ff),
	.w8(32'h3ad502de),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade709d),
	.w1(32'h3a12f63c),
	.w2(32'hb843dc2b),
	.w3(32'h39dec709),
	.w4(32'h3983669c),
	.w5(32'hba1bad1a),
	.w6(32'h3805683f),
	.w7(32'hb9c6557e),
	.w8(32'hba2d471a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f02d68),
	.w1(32'h3997a427),
	.w2(32'h3b347ed1),
	.w3(32'hba805b17),
	.w4(32'h3b2680f5),
	.w5(32'h3b32dced),
	.w6(32'h3b37e2b8),
	.w7(32'h3b22f3b4),
	.w8(32'h3b474951),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b083a90),
	.w1(32'h3af6bc0c),
	.w2(32'hba1ef79f),
	.w3(32'h3b0cedde),
	.w4(32'hba1dcd38),
	.w5(32'h38168058),
	.w6(32'h3a009dbc),
	.w7(32'hba24de8f),
	.w8(32'hba89134f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25fabb),
	.w1(32'h3b73938e),
	.w2(32'hbb0f0f04),
	.w3(32'hb81b21cc),
	.w4(32'h3b46efb5),
	.w5(32'h3b27a48e),
	.w6(32'hba4243f3),
	.w7(32'hbb1bd86c),
	.w8(32'hb9bcaae9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace4643),
	.w1(32'h3a7bf109),
	.w2(32'h3ae6139c),
	.w3(32'h3a81e2c9),
	.w4(32'hba39f291),
	.w5(32'hba91612a),
	.w6(32'h3a280f43),
	.w7(32'h39a858d4),
	.w8(32'hbad3e958),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c8820),
	.w1(32'hb9c1a363),
	.w2(32'hb9a1bd03),
	.w3(32'hbae20e72),
	.w4(32'h3954f960),
	.w5(32'h37b2f958),
	.w6(32'hb8993bce),
	.w7(32'hb9eee35e),
	.w8(32'hb9d9ba20),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9840d8a),
	.w1(32'h3aa51159),
	.w2(32'h3b0788f6),
	.w3(32'h3843bdd3),
	.w4(32'hb8756554),
	.w5(32'h3aae0fee),
	.w6(32'hb8be3dab),
	.w7(32'h397eaf16),
	.w8(32'hb9eeb867),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e744b8),
	.w1(32'h39382551),
	.w2(32'h3a118ae4),
	.w3(32'hb9b4e92d),
	.w4(32'h38a40e8a),
	.w5(32'hb8afd130),
	.w6(32'h3a534603),
	.w7(32'hba27de0f),
	.w8(32'hba4ccb34),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44514b),
	.w1(32'h3a05956c),
	.w2(32'h3c78644d),
	.w3(32'h39f089f8),
	.w4(32'h3ae9316b),
	.w5(32'h3b68103c),
	.w6(32'h3b2980e9),
	.w7(32'h3a4d0a4a),
	.w8(32'hbb600e02),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb538993),
	.w1(32'h3b162801),
	.w2(32'h3ac33189),
	.w3(32'h3b2026dd),
	.w4(32'h3a690e74),
	.w5(32'h39c76f08),
	.w6(32'h3ae925f5),
	.w7(32'h3abf39a6),
	.w8(32'h3a3e6b37),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e722f5),
	.w1(32'h39ded151),
	.w2(32'hba748d66),
	.w3(32'h39244a02),
	.w4(32'hba14e5e5),
	.w5(32'hba7adab8),
	.w6(32'h39014f3b),
	.w7(32'hbac1369f),
	.w8(32'hba94d591),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7bf2b),
	.w1(32'h3b3b8411),
	.w2(32'hbacd1862),
	.w3(32'hbae68c76),
	.w4(32'h3a69fe80),
	.w5(32'h398e7807),
	.w6(32'hb9973e70),
	.w7(32'hbb1529ed),
	.w8(32'hbaeac4c3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02d380),
	.w1(32'h398e81b2),
	.w2(32'h3b081699),
	.w3(32'h3a9e6bc6),
	.w4(32'h3a6ed4dc),
	.w5(32'h3aeaf461),
	.w6(32'h3a01e1c2),
	.w7(32'h3ac6d064),
	.w8(32'h3b064db0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac62ce6),
	.w1(32'hb9bf6322),
	.w2(32'h3680b257),
	.w3(32'h3a42afe2),
	.w4(32'hb9922409),
	.w5(32'h3969be2f),
	.w6(32'h3a7f9591),
	.w7(32'h3a3416d7),
	.w8(32'h3adaff0e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa75fa1),
	.w1(32'hba9d80c3),
	.w2(32'hbaa76415),
	.w3(32'h39f71609),
	.w4(32'hba250eee),
	.w5(32'hba66561a),
	.w6(32'hb9a15a69),
	.w7(32'hba340430),
	.w8(32'hba44e5c3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c79e5),
	.w1(32'h3b734414),
	.w2(32'hbad5a4d2),
	.w3(32'hba05ea92),
	.w4(32'h3a7d76da),
	.w5(32'h3b3511b5),
	.w6(32'h3a77bc98),
	.w7(32'hbad75fa2),
	.w8(32'h3a0a7981),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9268ba),
	.w1(32'h3a323bca),
	.w2(32'h3b00e395),
	.w3(32'h3a89929b),
	.w4(32'hba862eaf),
	.w5(32'hba49ab04),
	.w6(32'h39ace6be),
	.w7(32'h3a2651b8),
	.w8(32'hbaa9433f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801163),
	.w1(32'hba5420a0),
	.w2(32'hba93d11c),
	.w3(32'hbaea09e2),
	.w4(32'hba03299f),
	.w5(32'hba69372b),
	.w6(32'hba4c0336),
	.w7(32'hba813e9a),
	.w8(32'hba358670),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b55382),
	.w1(32'hba56622f),
	.w2(32'hba265d5f),
	.w3(32'hb874fc12),
	.w4(32'hb93d854f),
	.w5(32'hb9cdc212),
	.w6(32'hb998d7b1),
	.w7(32'hba1c5e35),
	.w8(32'hba2d0e48),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8dd75),
	.w1(32'hbabe88ad),
	.w2(32'hba8da8e5),
	.w3(32'hb98bb762),
	.w4(32'hba1cc135),
	.w5(32'hba420b42),
	.w6(32'hbadb50df),
	.w7(32'hba920fd6),
	.w8(32'hba93c1c0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4eabb9),
	.w1(32'hba7c56bb),
	.w2(32'hba32dcec),
	.w3(32'hba74039c),
	.w4(32'h3830b87a),
	.w5(32'hb9d50695),
	.w6(32'h386b0039),
	.w7(32'h38b1e263),
	.w8(32'hbaaeeb01),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab23710),
	.w1(32'h3a1186f3),
	.w2(32'hb8b5d190),
	.w3(32'hbad54a78),
	.w4(32'h3c01b914),
	.w5(32'h3c192282),
	.w6(32'hbb176757),
	.w7(32'h3a6fed16),
	.w8(32'hba1f6fc8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4025b3),
	.w1(32'h3a81a5e0),
	.w2(32'hba40d04f),
	.w3(32'h3b27ca8c),
	.w4(32'h3b08014b),
	.w5(32'h3a04eb6d),
	.w6(32'h3a917bae),
	.w7(32'hba42adf7),
	.w8(32'h3ab19e07),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b7fd4),
	.w1(32'hb93e44f4),
	.w2(32'h3beb03c6),
	.w3(32'h3ab6f33c),
	.w4(32'hba253da5),
	.w5(32'h3ae13bf9),
	.w6(32'hba88b420),
	.w7(32'h39369451),
	.w8(32'hbb00ccb3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8909d4),
	.w1(32'h3a7f046d),
	.w2(32'hb9ec6038),
	.w3(32'h37d39574),
	.w4(32'hb9d79fc2),
	.w5(32'hba4074b1),
	.w6(32'hbac0ccfa),
	.w7(32'hbb2720ff),
	.w8(32'hba64481d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33542a),
	.w1(32'hba6c4909),
	.w2(32'hba82664e),
	.w3(32'hbac3dec3),
	.w4(32'h390fca3a),
	.w5(32'h39473196),
	.w6(32'hba64ac50),
	.w7(32'hba976ce7),
	.w8(32'hb985b7f3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a8e6c),
	.w1(32'hb9eee64b),
	.w2(32'hb8b05f44),
	.w3(32'hb98586a1),
	.w4(32'h39879191),
	.w5(32'h3a47aeb0),
	.w6(32'h3a5b35c4),
	.w7(32'h3a0bfe59),
	.w8(32'h3ae38783),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ed09c),
	.w1(32'hba01c3bd),
	.w2(32'hbb1b3a46),
	.w3(32'h39dc27e0),
	.w4(32'hbaea197d),
	.w5(32'hbb039cd3),
	.w6(32'hbb0ebd0a),
	.w7(32'hbb29afc2),
	.w8(32'hbb49fea7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07d46d),
	.w1(32'hba5f53d2),
	.w2(32'h3a1dafa1),
	.w3(32'hbb201850),
	.w4(32'hb7be9448),
	.w5(32'hb747d193),
	.w6(32'hb999f798),
	.w7(32'h39c83ded),
	.w8(32'hb920f06b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9366cf7),
	.w1(32'h3a858efb),
	.w2(32'h3b20fd1d),
	.w3(32'hb99e388b),
	.w4(32'hba2a3293),
	.w5(32'hba678a3c),
	.w6(32'h3a8d4f63),
	.w7(32'h38ae00d6),
	.w8(32'hba34f168),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921ec72),
	.w1(32'hbab14d1d),
	.w2(32'h3a588974),
	.w3(32'hba572792),
	.w4(32'hba23ca79),
	.w5(32'hb9a52c04),
	.w6(32'hbaba17c6),
	.w7(32'hbac8d4e2),
	.w8(32'hbabf132f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f96546),
	.w1(32'h3a26533d),
	.w2(32'hba17a027),
	.w3(32'hba4577cc),
	.w4(32'h39035935),
	.w5(32'hba03342a),
	.w6(32'h39b4a988),
	.w7(32'hba2bec29),
	.w8(32'hba3c43d1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ea7529),
	.w1(32'hbabc55cb),
	.w2(32'h3a9c7335),
	.w3(32'hb90a775c),
	.w4(32'hb9a50ba8),
	.w5(32'h3a8ff4b0),
	.w6(32'hbb1a207a),
	.w7(32'h3aa56838),
	.w8(32'hba9f6614),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22cdaf),
	.w1(32'hba7aefce),
	.w2(32'hba495d7f),
	.w3(32'hb9c181cb),
	.w4(32'hb89d8acb),
	.w5(32'hb97b9335),
	.w6(32'hba046af8),
	.w7(32'hb9fa6a28),
	.w8(32'hba39b3e3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be16fb),
	.w1(32'h3a207d56),
	.w2(32'h3a2fb8f9),
	.w3(32'hb93fc1b1),
	.w4(32'h39ae2a89),
	.w5(32'h3a1db429),
	.w6(32'hb90c48dd),
	.w7(32'hb91417e2),
	.w8(32'h390eea76),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b13519),
	.w1(32'hb9cb0c05),
	.w2(32'hb9e8de5d),
	.w3(32'hb93a49cc),
	.w4(32'h3a5e9400),
	.w5(32'h3a381de7),
	.w6(32'hb9cb4b70),
	.w7(32'hba268f0e),
	.w8(32'hb9ba17fa),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2823a),
	.w1(32'hbab564f7),
	.w2(32'hba7f754e),
	.w3(32'h39dd6e83),
	.w4(32'hba6d7a4d),
	.w5(32'hbac10b39),
	.w6(32'hb8a63865),
	.w7(32'hba4ffac0),
	.w8(32'hba978614),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f4dac),
	.w1(32'h3a716b06),
	.w2(32'h3ad29f18),
	.w3(32'hbabaa700),
	.w4(32'hbaca0cc7),
	.w5(32'h399b9d83),
	.w6(32'h3a06ba84),
	.w7(32'hb93b6196),
	.w8(32'hb9b1b220),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996e65f),
	.w1(32'hb8be9890),
	.w2(32'h3a0d1900),
	.w3(32'hb9630eb2),
	.w4(32'hba87560b),
	.w5(32'hbab45f2a),
	.w6(32'h3abe7739),
	.w7(32'h3a08c61a),
	.w8(32'h3a63bcd1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1babc4),
	.w1(32'h3a5696ad),
	.w2(32'h3a64dc2e),
	.w3(32'hbac099bb),
	.w4(32'h3a4bc448),
	.w5(32'h3a8ce552),
	.w6(32'h3ac84cc1),
	.w7(32'h3a900002),
	.w8(32'h3b536424),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a922a83),
	.w1(32'h3a97c671),
	.w2(32'h3b2f9994),
	.w3(32'h3993d2e9),
	.w4(32'hbaa6c83f),
	.w5(32'hb9593c48),
	.w6(32'hb9fcc4f2),
	.w7(32'hba989f80),
	.w8(32'h385acb57),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e00a0f),
	.w1(32'h3b3f9f85),
	.w2(32'h3abaf14f),
	.w3(32'hbaa55a63),
	.w4(32'hba94aeda),
	.w5(32'hbaba657a),
	.w6(32'h3a8b7560),
	.w7(32'hba792e07),
	.w8(32'h3a2db7d3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b195076),
	.w1(32'h393bc86d),
	.w2(32'h3a2e8b86),
	.w3(32'h3a6d6144),
	.w4(32'hb9fe2fee),
	.w5(32'h3a3ffef2),
	.w6(32'h37e8fbdd),
	.w7(32'h38e078fc),
	.w8(32'h3a71e66d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb899b),
	.w1(32'h39d569fb),
	.w2(32'h3babb448),
	.w3(32'h3a72327d),
	.w4(32'h39e7f019),
	.w5(32'h3a6df268),
	.w6(32'h3a8c825d),
	.w7(32'h38f7202c),
	.w8(32'hba2b1b2e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a4f7d),
	.w1(32'h39a632cf),
	.w2(32'hba0ca17f),
	.w3(32'h3ab7c437),
	.w4(32'hbab3a9b1),
	.w5(32'hba10bd53),
	.w6(32'hba3e23c0),
	.w7(32'hba90f756),
	.w8(32'hbb094159),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad02db8),
	.w1(32'hba953be0),
	.w2(32'hbb0cf43d),
	.w3(32'hbaa14333),
	.w4(32'h3a11f56d),
	.w5(32'hba5543f9),
	.w6(32'h39ad9460),
	.w7(32'hba307c98),
	.w8(32'hb98aa32c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c6483),
	.w1(32'h3be73b51),
	.w2(32'hba46ea70),
	.w3(32'h3a5d94cd),
	.w4(32'h3ace555d),
	.w5(32'h3b3a9ae4),
	.w6(32'h3b5183fc),
	.w7(32'hbae5e261),
	.w8(32'hba8408ac),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b680d4d),
	.w1(32'h3bb2bd10),
	.w2(32'hbb37042e),
	.w3(32'h3a9eb3cf),
	.w4(32'h3b021cd3),
	.w5(32'h3b154394),
	.w6(32'h3a24ae9c),
	.w7(32'hba71d324),
	.w8(32'h3aa915fa),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf9bea),
	.w1(32'h37bba26e),
	.w2(32'hbb27905a),
	.w3(32'h3bf42bf2),
	.w4(32'h3ac7c790),
	.w5(32'h3aa005d1),
	.w6(32'h3a2332dc),
	.w7(32'hbb3871f8),
	.w8(32'h3a979c93),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d6d45),
	.w1(32'hba367920),
	.w2(32'hbaed16a3),
	.w3(32'h3b0c0567),
	.w4(32'hb95fa827),
	.w5(32'hba793578),
	.w6(32'hba6b49a5),
	.w7(32'hbaa6a285),
	.w8(32'hba4929cd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9816a77),
	.w1(32'h38cc5b1f),
	.w2(32'hba33f2dc),
	.w3(32'hb9462676),
	.w4(32'h3a67506b),
	.w5(32'h3a83e542),
	.w6(32'h39baf0f9),
	.w7(32'hba931e6e),
	.w8(32'h3a714551),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea42fe),
	.w1(32'hba706bc1),
	.w2(32'h3a83e8ec),
	.w3(32'h3a97639b),
	.w4(32'hba2b9e26),
	.w5(32'hb989b2b3),
	.w6(32'hba3d0719),
	.w7(32'hb9c9f586),
	.w8(32'hba38928e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9b592),
	.w1(32'h373b4b70),
	.w2(32'h3b6e81ca),
	.w3(32'h3848eb58),
	.w4(32'hbb0cb172),
	.w5(32'hbb0b3bd7),
	.w6(32'h3a616cda),
	.w7(32'hba9bdcff),
	.w8(32'hbac348d3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e0419),
	.w1(32'hbad35df4),
	.w2(32'hba43e99a),
	.w3(32'hbaa416c2),
	.w4(32'hba004a80),
	.w5(32'hb9a78688),
	.w6(32'hba9db6c1),
	.w7(32'hba801fb3),
	.w8(32'hbaad743a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20e262),
	.w1(32'h3a1f87e6),
	.w2(32'hba662667),
	.w3(32'hba709105),
	.w4(32'h3a8476ce),
	.w5(32'h3a90f648),
	.w6(32'hb9aa958b),
	.w7(32'hbb02cdb2),
	.w8(32'h39f3142f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39dda2),
	.w1(32'h3ac6425c),
	.w2(32'h3b569685),
	.w3(32'h3a8bc8ed),
	.w4(32'hba26d4ea),
	.w5(32'hb986bafc),
	.w6(32'h398a1895),
	.w7(32'hbaf795ca),
	.w8(32'hbb48dd2f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5c189),
	.w1(32'hbafa2b16),
	.w2(32'hb99d1203),
	.w3(32'hb81cb3de),
	.w4(32'hba77975f),
	.w5(32'hb9a629f5),
	.w6(32'hba7c6cde),
	.w7(32'hba2b638a),
	.w8(32'hbaa596a1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63f0c8),
	.w1(32'h3a2f57db),
	.w2(32'h3c6ff5b2),
	.w3(32'h394fd4c9),
	.w4(32'h3b25628c),
	.w5(32'h3bce209c),
	.w6(32'h3a938a11),
	.w7(32'h3b905c96),
	.w8(32'hbb084b6d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb495a5e),
	.w1(32'hbae9c584),
	.w2(32'hbae2cb58),
	.w3(32'h3afbba26),
	.w4(32'hba246089),
	.w5(32'hba943009),
	.w6(32'hba609124),
	.w7(32'hbab0b151),
	.w8(32'hbaaa1a96),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad61432),
	.w1(32'hba4feb01),
	.w2(32'h3a283eec),
	.w3(32'hbaa1dc4d),
	.w4(32'hba883e91),
	.w5(32'hb97cd4a0),
	.w6(32'hbab6366a),
	.w7(32'hb9f7d7aa),
	.w8(32'hba955126),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccd47f),
	.w1(32'h39bcf74f),
	.w2(32'h3b2a9899),
	.w3(32'hbac06747),
	.w4(32'h39f4962e),
	.w5(32'h3a914c3b),
	.w6(32'h3a4d7a5e),
	.w7(32'h38b6b244),
	.w8(32'hb5dd1214),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b70b8),
	.w1(32'h3910166f),
	.w2(32'hbb10481c),
	.w3(32'h3ac1d3f1),
	.w4(32'h3acf6ac5),
	.w5(32'h390b7349),
	.w6(32'h3a153885),
	.w7(32'hbaec2f5e),
	.w8(32'h392f7697),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd45ff),
	.w1(32'hba3317c3),
	.w2(32'hba8e2439),
	.w3(32'h3ad4b3d9),
	.w4(32'h390d2b12),
	.w5(32'hb9d4b46a),
	.w6(32'hb9f45707),
	.w7(32'hba8f5397),
	.w8(32'hba06ea9f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9ebac),
	.w1(32'hbaa4f221),
	.w2(32'hbae3f29c),
	.w3(32'h3995a0ad),
	.w4(32'h39042949),
	.w5(32'hba6cda1a),
	.w6(32'hba540fab),
	.w7(32'hbad9d86b),
	.w8(32'hba03ccb7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9342a32),
	.w1(32'h3b3e605d),
	.w2(32'h3b7c0ec3),
	.w3(32'hb85bc42d),
	.w4(32'hb9172086),
	.w5(32'hba89c3a0),
	.w6(32'h3a28c760),
	.w7(32'hbb86f41c),
	.w8(32'hbb04499f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbe1cc),
	.w1(32'h3b6a4696),
	.w2(32'hba133773),
	.w3(32'h3b692f3d),
	.w4(32'h3a7f7364),
	.w5(32'h39921f78),
	.w6(32'h3a20a554),
	.w7(32'hbac46f6a),
	.w8(32'hbae55aa0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f1bce),
	.w1(32'hbb168126),
	.w2(32'hbaf77a25),
	.w3(32'hba905c80),
	.w4(32'hbab2c7f3),
	.w5(32'hbae093ff),
	.w6(32'hbb0297a5),
	.w7(32'hbb191466),
	.w8(32'hbb23ba70),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfc485),
	.w1(32'hbb167016),
	.w2(32'hba969a46),
	.w3(32'hbaf21b01),
	.w4(32'hbab7cf89),
	.w5(32'hbabc0b64),
	.w6(32'hbb10b1e0),
	.w7(32'hbaf055c7),
	.w8(32'hbac2c6ca),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c10496),
	.w1(32'h398e697e),
	.w2(32'hb8ea0d26),
	.w3(32'hb80b7c80),
	.w4(32'h3a8d8c3e),
	.w5(32'h39d47b7c),
	.w6(32'h3a83c2c4),
	.w7(32'h399212eb),
	.w8(32'h39b63744),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c507ec),
	.w1(32'h3c025f61),
	.w2(32'h3bf86da4),
	.w3(32'h3a28f4dd),
	.w4(32'h3a501b83),
	.w5(32'hba102e00),
	.w6(32'h3b09b551),
	.w7(32'hbb49d45c),
	.w8(32'hbb0e0dad),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acff913),
	.w1(32'hbad47e8a),
	.w2(32'hbb8a7beb),
	.w3(32'h3ba8cb17),
	.w4(32'hbab0a340),
	.w5(32'hbb3f3205),
	.w6(32'hba80ff9c),
	.w7(32'hbb168c97),
	.w8(32'hba431876),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba767ea7),
	.w1(32'hbb08d7a0),
	.w2(32'hbab5c3f0),
	.w3(32'hba7e2e94),
	.w4(32'hba4caa0c),
	.w5(32'hba66475c),
	.w6(32'hba9fac26),
	.w7(32'hba8b04e1),
	.w8(32'hba9869f1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cabd8),
	.w1(32'h39f7d1ff),
	.w2(32'h39e21b16),
	.w3(32'hb9f2a1e9),
	.w4(32'h39e21128),
	.w5(32'h39d1a2c3),
	.w6(32'h399320e2),
	.w7(32'h3889cd4e),
	.w8(32'h39b6b52b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a007dd7),
	.w1(32'h39ef0131),
	.w2(32'h39cf20b0),
	.w3(32'h3a2b07ef),
	.w4(32'h3a574170),
	.w5(32'h3a77dbc9),
	.w6(32'h3a5f21ae),
	.w7(32'h3a0f7fd7),
	.w8(32'h3a81da11),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a890519),
	.w1(32'h39825e99),
	.w2(32'h3ac81490),
	.w3(32'h3a326dcc),
	.w4(32'hb97cc0a2),
	.w5(32'h3a883c16),
	.w6(32'hba81d431),
	.w7(32'hb99fa988),
	.w8(32'h39baf671),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d39ac9),
	.w1(32'hb96a8b3d),
	.w2(32'hb9d81f59),
	.w3(32'h39ae1e53),
	.w4(32'hb98d778b),
	.w5(32'hb9cc0aa7),
	.w6(32'hb944365b),
	.w7(32'hb92af812),
	.w8(32'hb984998b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb9f2f),
	.w1(32'h39d11ed0),
	.w2(32'h3802681e),
	.w3(32'hb8ad4600),
	.w4(32'h38d1880a),
	.w5(32'h38eb6669),
	.w6(32'h3a477080),
	.w7(32'h39ee16a9),
	.w8(32'h39399d8e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af32d8),
	.w1(32'hba3c6cbb),
	.w2(32'hba27fc42),
	.w3(32'h3905c9e3),
	.w4(32'hb9824e34),
	.w5(32'hb94dcf50),
	.w6(32'h387e09b7),
	.w7(32'h384f39b7),
	.w8(32'h398b2f8e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b27b5),
	.w1(32'hb986be68),
	.w2(32'hb786b84d),
	.w3(32'hba1e61e8),
	.w4(32'hb9bab4f1),
	.w5(32'h39575fb1),
	.w6(32'hb982657d),
	.w7(32'hba0a2b20),
	.w8(32'hb8c4387d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce4b98),
	.w1(32'h3a5f2967),
	.w2(32'h3a922015),
	.w3(32'hb9ac117b),
	.w4(32'h3a66f2df),
	.w5(32'h3ac69cd3),
	.w6(32'h3a13873f),
	.w7(32'h3a70edf0),
	.w8(32'h3ad4f280),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a978a73),
	.w1(32'hb99fcd8d),
	.w2(32'h362baaeb),
	.w3(32'h3a845a94),
	.w4(32'hb9ebd720),
	.w5(32'h398a414a),
	.w6(32'hb8b61c85),
	.w7(32'hb9b8d61d),
	.w8(32'h3a18f8c2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b05a67),
	.w1(32'h3a589c9a),
	.w2(32'h3a9f6b2e),
	.w3(32'hba5505c9),
	.w4(32'h3a1f95d4),
	.w5(32'h3aaf2587),
	.w6(32'h3a4566db),
	.w7(32'h3a36e4f1),
	.w8(32'h3ac39fea),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7d212),
	.w1(32'h39c11268),
	.w2(32'h3967dfc3),
	.w3(32'h3a9e5962),
	.w4(32'h391f2682),
	.w5(32'h3a6c2e2c),
	.w6(32'h39fd91c1),
	.w7(32'h39c28556),
	.w8(32'h3aba1abc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a851b74),
	.w1(32'hba1117b1),
	.w2(32'h396cc074),
	.w3(32'h39f204a5),
	.w4(32'hba7db645),
	.w5(32'h38bbd54f),
	.w6(32'hb9a3fd50),
	.w7(32'hba004caa),
	.w8(32'h386471ff),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a130d),
	.w1(32'h388bf29b),
	.w2(32'hb9bfce0f),
	.w3(32'hba6bf6d8),
	.w4(32'h393536b9),
	.w5(32'h393fba0f),
	.w6(32'h39b8ace0),
	.w7(32'h39c4c2b2),
	.w8(32'h3a1b0517),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39025578),
	.w1(32'h3a189984),
	.w2(32'h3ad926c1),
	.w3(32'hb99a24b5),
	.w4(32'h3a262082),
	.w5(32'h3b061c20),
	.w6(32'h3a89613c),
	.w7(32'h3a93438b),
	.w8(32'h3af85c91),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c6de4),
	.w1(32'h3a3639cd),
	.w2(32'h3a3f7aa3),
	.w3(32'h3a43beb3),
	.w4(32'h39f61606),
	.w5(32'h3a2209be),
	.w6(32'h39f95274),
	.w7(32'h39d155a8),
	.w8(32'h3a1dc5be),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6bb0b),
	.w1(32'h3a906407),
	.w2(32'h3ab2d7e5),
	.w3(32'h3a2e03e0),
	.w4(32'h3a9896fe),
	.w5(32'h3af219cf),
	.w6(32'h3aec1b80),
	.w7(32'h3af039ba),
	.w8(32'h3b3ee7f9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0743c5),
	.w1(32'hba56f590),
	.w2(32'hb99190b2),
	.w3(32'h3a66c6e5),
	.w4(32'hb98ebd5f),
	.w5(32'h3a3a7807),
	.w6(32'h3a31b6e8),
	.w7(32'h3a6588e1),
	.w8(32'h3a9da31a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d5481),
	.w1(32'h37a50ae7),
	.w2(32'h3946b14c),
	.w3(32'h394fb32b),
	.w4(32'h39988926),
	.w5(32'h39dd723d),
	.w6(32'h395d0054),
	.w7(32'h39b0d5ca),
	.w8(32'h39db0c93),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a259955),
	.w1(32'h3994411b),
	.w2(32'h3712e66f),
	.w3(32'h3a3106ec),
	.w4(32'h388b22bf),
	.w5(32'h39a214b1),
	.w6(32'hb9960436),
	.w7(32'hb8e4e8f1),
	.w8(32'hb9b7b72f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c043a2),
	.w1(32'h38939f10),
	.w2(32'hb9ed2ba0),
	.w3(32'h38f24cb0),
	.w4(32'hb8f687a5),
	.w5(32'hba08620e),
	.w6(32'h36b911ae),
	.w7(32'hb9271bb3),
	.w8(32'hb980e774),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ef85b),
	.w1(32'hba5777c4),
	.w2(32'h38fceccb),
	.w3(32'hba728d19),
	.w4(32'hb9796a21),
	.w5(32'h3a899cf1),
	.w6(32'h396d950b),
	.w7(32'h3a3ddcda),
	.w8(32'h3af76e83),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0df18e),
	.w1(32'h3a9d5c46),
	.w2(32'h3a2f999a),
	.w3(32'hb944ad1e),
	.w4(32'h3a3ee724),
	.w5(32'h3a8ad319),
	.w6(32'hb8e11e2c),
	.w7(32'h39dc5192),
	.w8(32'h3a4eb42a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d554f),
	.w1(32'h39cfc65a),
	.w2(32'h3a0bafdc),
	.w3(32'h3a1e10f0),
	.w4(32'h39ccede0),
	.w5(32'h3a03d815),
	.w6(32'h3979920e),
	.w7(32'h39c585a0),
	.w8(32'h3a2a0c7d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a77b4),
	.w1(32'h38c7090a),
	.w2(32'hb9323732),
	.w3(32'h39d00ea1),
	.w4(32'hb9ddfb13),
	.w5(32'h3abf19fd),
	.w6(32'hb9dcda8d),
	.w7(32'hb85de911),
	.w8(32'h3aade806),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929339b),
	.w1(32'h3931b6da),
	.w2(32'h3a040583),
	.w3(32'h39e2d917),
	.w4(32'h39a3b22b),
	.w5(32'h3a9903e0),
	.w6(32'h38f62644),
	.w7(32'h3990b5db),
	.w8(32'h3a51d828),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38308ade),
	.w1(32'h39f0e08d),
	.w2(32'h3a446359),
	.w3(32'hb9a9b6aa),
	.w4(32'h3a283433),
	.w5(32'h3a972254),
	.w6(32'h3a2d0bd2),
	.w7(32'h39c2c135),
	.w8(32'h3a9aae87),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e3418),
	.w1(32'hba269dee),
	.w2(32'h38102cde),
	.w3(32'h3a223e91),
	.w4(32'hb9d31050),
	.w5(32'h39b45c92),
	.w6(32'hb70ab220),
	.w7(32'hb91a0b99),
	.w8(32'h37e28abe),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb948e63c),
	.w1(32'hb8c69571),
	.w2(32'hba222591),
	.w3(32'h38acf5cd),
	.w4(32'hb99c9fa4),
	.w5(32'hb9d309d2),
	.w6(32'h39be9b95),
	.w7(32'h39939a51),
	.w8(32'h387fe5c3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d65131),
	.w1(32'h39e87996),
	.w2(32'h39ca9412),
	.w3(32'hb99bd964),
	.w4(32'h399bcbf5),
	.w5(32'h39c10555),
	.w6(32'h395da3cf),
	.w7(32'h39b906ba),
	.w8(32'h39e1a94a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ced361),
	.w1(32'hb78cbcde),
	.w2(32'h3a11d524),
	.w3(32'hb7d28bd8),
	.w4(32'hb8c940ba),
	.w5(32'h3a8ddbb6),
	.w6(32'hb9dc7f85),
	.w7(32'hb9a2939a),
	.w8(32'h3a16118e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af826ac),
	.w1(32'h3a3bc9f8),
	.w2(32'hb935b0d2),
	.w3(32'h3a857353),
	.w4(32'h3a7025b5),
	.w5(32'hb93e0746),
	.w6(32'h3a1ffe26),
	.w7(32'h3a807558),
	.w8(32'h3a58c673),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9460ec4),
	.w1(32'hba38023d),
	.w2(32'hba6e3381),
	.w3(32'hb8d64e14),
	.w4(32'hba47c5cf),
	.w5(32'hba6d5f0f),
	.w6(32'hba492772),
	.w7(32'hba515765),
	.w8(32'hba6af7d4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b05907),
	.w1(32'h3992f0f7),
	.w2(32'h39ef1cf1),
	.w3(32'hb98bd82f),
	.w4(32'h39870bb7),
	.w5(32'h39b6b337),
	.w6(32'h38aa77d7),
	.w7(32'h39784db7),
	.w8(32'h39b0f481),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14651e),
	.w1(32'h39a9b56a),
	.w2(32'h398a04ac),
	.w3(32'h39fd137b),
	.w4(32'h39c02b07),
	.w5(32'h3995b8bf),
	.w6(32'h399eafe5),
	.w7(32'h3996ed14),
	.w8(32'h3999a030),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a131d95),
	.w1(32'h3a4651bd),
	.w2(32'h3aae6d40),
	.w3(32'h39695090),
	.w4(32'h38be9ac0),
	.w5(32'h3ab90fb6),
	.w6(32'h39b69ca2),
	.w7(32'h393d45a2),
	.w8(32'h39dc002b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388adc13),
	.w1(32'hb9edcad2),
	.w2(32'h38fb607d),
	.w3(32'h3983ab0c),
	.w4(32'hb9135ba8),
	.w5(32'hb899c188),
	.w6(32'hba09ac62),
	.w7(32'h398b9e8b),
	.w8(32'h39e90fa7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b85068),
	.w1(32'h39ba4764),
	.w2(32'h3a3dd964),
	.w3(32'h38e69b30),
	.w4(32'hb804290f),
	.w5(32'h3a3d90d2),
	.w6(32'h39c4bd86),
	.w7(32'h384611f9),
	.w8(32'h3a06c6a3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959dc57),
	.w1(32'h398b24f3),
	.w2(32'h38f7dd03),
	.w3(32'hb8095da3),
	.w4(32'h39a8f932),
	.w5(32'h39aa41da),
	.w6(32'h398426f8),
	.w7(32'h39ae5641),
	.w8(32'h3994f02c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9deee08),
	.w1(32'h3919db38),
	.w2(32'hb99d1a69),
	.w3(32'hba1579ae),
	.w4(32'hb9b6b14e),
	.w5(32'hba5d2f60),
	.w6(32'hba2d1946),
	.w7(32'h3925290b),
	.w8(32'hb9a0cc44),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f8858f),
	.w1(32'hba1bebad),
	.w2(32'hba66e08e),
	.w3(32'hb84a44cf),
	.w4(32'hba263e24),
	.w5(32'hba346b56),
	.w6(32'hba108aaf),
	.w7(32'hba289788),
	.w8(32'hba1c9bb5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58ce00),
	.w1(32'h39e07262),
	.w2(32'h39a2427f),
	.w3(32'hba680c33),
	.w4(32'h3a1d87b7),
	.w5(32'h3a0c95e7),
	.w6(32'h39cf26e9),
	.w7(32'h3a0ae1a1),
	.w8(32'h3a38579b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88142f9),
	.w1(32'hba081a92),
	.w2(32'h3a09c4d3),
	.w3(32'hb9d10710),
	.w4(32'hba816f83),
	.w5(32'h39e36c7d),
	.w6(32'hb9fcbf9e),
	.w7(32'hba577a82),
	.w8(32'h38e13d87),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6db6d),
	.w1(32'hb9c75398),
	.w2(32'h39316297),
	.w3(32'hb9ddb2d6),
	.w4(32'hb98db8e6),
	.w5(32'h3a27836e),
	.w6(32'hb99c8bab),
	.w7(32'hb9098199),
	.w8(32'h3aa0ba65),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8b334),
	.w1(32'h38265aef),
	.w2(32'hb8bc8497),
	.w3(32'hba4116f1),
	.w4(32'hb920fd23),
	.w5(32'hb9304002),
	.w6(32'h397f4234),
	.w7(32'h3a2114dc),
	.w8(32'h399eb8b5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a267b65),
	.w1(32'h393ddfc5),
	.w2(32'h3a40c3ed),
	.w3(32'hb8db8a1d),
	.w4(32'h37ec6504),
	.w5(32'h3a64c580),
	.w6(32'h38f84de9),
	.w7(32'hb984606d),
	.w8(32'h3a9141ab),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be7f78),
	.w1(32'hba842763),
	.w2(32'hbaa2ec2d),
	.w3(32'h3972f0e0),
	.w4(32'hba8d5971),
	.w5(32'hba9b4ca5),
	.w6(32'hba54fc14),
	.w7(32'hba6cc673),
	.w8(32'hba2b21ad),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52a8f7),
	.w1(32'h3b0030d4),
	.w2(32'h3a9d0bde),
	.w3(32'h3a850379),
	.w4(32'h3b0dfeb8),
	.w5(32'h3b035ab9),
	.w6(32'h3aec33ad),
	.w7(32'h3b248daa),
	.w8(32'h3b33c434),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882b80e),
	.w1(32'h39d7e1f2),
	.w2(32'h3949b503),
	.w3(32'h395fd562),
	.w4(32'h386f50e0),
	.w5(32'h38b30679),
	.w6(32'h3a65994f),
	.w7(32'h39d661a3),
	.w8(32'h39f118c5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f6379),
	.w1(32'hba7d5416),
	.w2(32'hb90d592f),
	.w3(32'h3727a5bc),
	.w4(32'hba11c63f),
	.w5(32'h3a219f13),
	.w6(32'hba527db4),
	.w7(32'hb9c487df),
	.w8(32'h3a8bb4ff),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b194f),
	.w1(32'hb9ba130e),
	.w2(32'hb9b4df59),
	.w3(32'hba181378),
	.w4(32'hb97f1feb),
	.w5(32'hb6de916e),
	.w6(32'hb9bdf895),
	.w7(32'hb9993a8f),
	.w8(32'hb96f1c24),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b4af3),
	.w1(32'h39882caa),
	.w2(32'h3a2888a4),
	.w3(32'hba13de80),
	.w4(32'h39467dd4),
	.w5(32'h3a8e6148),
	.w6(32'hb8166d17),
	.w7(32'h39e13cd4),
	.w8(32'h3aab9372),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a091fee),
	.w1(32'h3a1db3a4),
	.w2(32'h3a114f98),
	.w3(32'h3a031019),
	.w4(32'h3a3d950e),
	.w5(32'h3a1e4068),
	.w6(32'h3a38055b),
	.w7(32'h3a39f076),
	.w8(32'h3a600942),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89265b),
	.w1(32'h39f9bf3c),
	.w2(32'hb69d0c7a),
	.w3(32'h3a6f96d2),
	.w4(32'h398510cd),
	.w5(32'h385bca87),
	.w6(32'h3a0d7f7a),
	.w7(32'h39b05c6a),
	.w8(32'h39b5d809),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3fea1),
	.w1(32'hba209225),
	.w2(32'h3a3ebe2c),
	.w3(32'h39a44363),
	.w4(32'hb82dc839),
	.w5(32'h3a78b634),
	.w6(32'h38f5a58b),
	.w7(32'h39567edc),
	.w8(32'h3a2574f9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4e7a9),
	.w1(32'h39710050),
	.w2(32'h3a45d86a),
	.w3(32'h3a8512a3),
	.w4(32'h39bf4aa5),
	.w5(32'h3aa2e3d9),
	.w6(32'h38b8354d),
	.w7(32'h3a7e51e3),
	.w8(32'h3ab7dd8d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebf2d6),
	.w1(32'hb9294607),
	.w2(32'h3931b0a5),
	.w3(32'h3a203c7d),
	.w4(32'hb92d8d64),
	.w5(32'h38de890e),
	.w6(32'hb9d4bda2),
	.w7(32'hb995b2f9),
	.w8(32'hb9876cbe),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1bdf0),
	.w1(32'hb72df06c),
	.w2(32'hb973657f),
	.w3(32'hb92eb00b),
	.w4(32'hb8bb7d9e),
	.w5(32'hb855029f),
	.w6(32'h371c4d85),
	.w7(32'hb789fc0c),
	.w8(32'h38cd9afe),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90fdd6f),
	.w1(32'hba58f435),
	.w2(32'hba8e458a),
	.w3(32'hb8c3a782),
	.w4(32'hba5e6f45),
	.w5(32'hba7dc01c),
	.w6(32'hba730d0e),
	.w7(32'hba7d4a8d),
	.w8(32'hba8d9ca5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea16ab),
	.w1(32'h3a075f08),
	.w2(32'h3a444460),
	.w3(32'hb9e76b4f),
	.w4(32'h398b9fb1),
	.w5(32'h3a1f3a22),
	.w6(32'h3a17bb09),
	.w7(32'h3a1ebb50),
	.w8(32'h3a5209a4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c57ebe),
	.w1(32'h39b84e2c),
	.w2(32'h3947058c),
	.w3(32'h38d6cc04),
	.w4(32'h39fd0c3a),
	.w5(32'h3937264a),
	.w6(32'h3a32e41d),
	.w7(32'h39c15d6d),
	.w8(32'h3a90bb51),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa309d7),
	.w1(32'hb78fe4a6),
	.w2(32'hb987720e),
	.w3(32'h3a5c5fe5),
	.w4(32'h38c46658),
	.w5(32'hb9643e06),
	.w6(32'hb977ac0d),
	.w7(32'hb92a4922),
	.w8(32'hb721681b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93194e),
	.w1(32'h3b23fca2),
	.w2(32'h3af21685),
	.w3(32'h387e8a99),
	.w4(32'h3adfcc96),
	.w5(32'h3b158eaf),
	.w6(32'h39a26aad),
	.w7(32'h3a2c4570),
	.w8(32'h3b0e5007),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04b4ab),
	.w1(32'h39182d4c),
	.w2(32'h39be394f),
	.w3(32'h397818f5),
	.w4(32'hb920cb0c),
	.w5(32'h3a15959b),
	.w6(32'hb9342b07),
	.w7(32'h387d5ad9),
	.w8(32'h3a21d2fa),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9949c0f),
	.w1(32'h39ba15a7),
	.w2(32'h3a0609bc),
	.w3(32'hb94458f1),
	.w4(32'h39b06029),
	.w5(32'h39f5c6d0),
	.w6(32'h398159ff),
	.w7(32'h39ce3b97),
	.w8(32'h3a007900),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ce73e),
	.w1(32'h3a1a073c),
	.w2(32'h3a10d9a9),
	.w3(32'h3a41b5ad),
	.w4(32'h391a890b),
	.w5(32'h39f54d0e),
	.w6(32'h38ba67aa),
	.w7(32'h3a09cb02),
	.w8(32'h3a126b3a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aefd14),
	.w1(32'hba149cb2),
	.w2(32'hba5152df),
	.w3(32'hb802f57d),
	.w4(32'hba3287cd),
	.w5(32'hba50de59),
	.w6(32'hb9da7f23),
	.w7(32'hba0aad39),
	.w8(32'hba069b7b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba701521),
	.w1(32'h39c26941),
	.w2(32'hb78f7df5),
	.w3(32'hba3f0844),
	.w4(32'h39ae8493),
	.w5(32'h390cc10e),
	.w6(32'h39b8fa09),
	.w7(32'h39b7065b),
	.w8(32'h392ff08e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89cb37a),
	.w1(32'hb93e0642),
	.w2(32'hb5b684c8),
	.w3(32'hb95807ef),
	.w4(32'hb8bbc5a5),
	.w5(32'hb76f6ab6),
	.w6(32'h3988ae29),
	.w7(32'hba1b2836),
	.w8(32'h39ebae01),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a996624),
	.w1(32'hba0468ac),
	.w2(32'hb9e80cbc),
	.w3(32'h3aa998c8),
	.w4(32'hba046496),
	.w5(32'hb9e38419),
	.w6(32'hb9ab0a29),
	.w7(32'h3982f9df),
	.w8(32'h3a50b911),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5b26d),
	.w1(32'h390ee23c),
	.w2(32'h3a20800d),
	.w3(32'hba8578dc),
	.w4(32'hb9fa998f),
	.w5(32'h399bc870),
	.w6(32'hba410afd),
	.w7(32'hb9a24648),
	.w8(32'h38ced7ad),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c963ce),
	.w1(32'h393f9cfc),
	.w2(32'h3a06dc60),
	.w3(32'hb90ea1bd),
	.w4(32'h397de844),
	.w5(32'h3a1ace9f),
	.w6(32'h398eeacb),
	.w7(32'h39ae0872),
	.w8(32'h3a1e02e6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab960da),
	.w1(32'h3800dfa4),
	.w2(32'hb7300418),
	.w3(32'h3a453123),
	.w4(32'hb9a0c8a3),
	.w5(32'h399168b7),
	.w6(32'h398565cb),
	.w7(32'hba3f26dc),
	.w8(32'h3a00c8ab),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a54ad6),
	.w1(32'h3832ddd4),
	.w2(32'hb9cbf1a4),
	.w3(32'hb8a532df),
	.w4(32'hb8dd2331),
	.w5(32'hb9bca4bf),
	.w6(32'h37706d1d),
	.w7(32'hb9268587),
	.w8(32'hb964d11b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec19d8),
	.w1(32'h3a03f1f3),
	.w2(32'h39bbbc4a),
	.w3(32'hba011b8a),
	.w4(32'h3a2fd9ef),
	.w5(32'h3a17ab98),
	.w6(32'h3a0dd597),
	.w7(32'h3a0a2f56),
	.w8(32'h3a169f24),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a220df6),
	.w1(32'h39ab9827),
	.w2(32'h3974e3d8),
	.w3(32'h3a30c549),
	.w4(32'h3a05c228),
	.w5(32'h3a07977b),
	.w6(32'h39cfaef4),
	.w7(32'h39f3bbe2),
	.w8(32'h3a1ade4b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a308e04),
	.w1(32'h39c4eab9),
	.w2(32'h398769c2),
	.w3(32'h3a3270e2),
	.w4(32'h39dd135c),
	.w5(32'h39ca2805),
	.w6(32'h398158ff),
	.w7(32'h39ca4e8e),
	.w8(32'h39cf98a1),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ec039),
	.w1(32'h391836ba),
	.w2(32'h3995405e),
	.w3(32'h39c83b52),
	.w4(32'hb94e20c4),
	.w5(32'h39b1778e),
	.w6(32'hb81fe834),
	.w7(32'hb98bcda1),
	.w8(32'h39171302),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d66b6a),
	.w1(32'hb9d29a43),
	.w2(32'h39c6ec13),
	.w3(32'h3983d04f),
	.w4(32'h38946b54),
	.w5(32'hb842937e),
	.w6(32'h3a695541),
	.w7(32'h3adad29f),
	.w8(32'h3a73d307),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b9e9c),
	.w1(32'h3a3232fd),
	.w2(32'h3aa3df88),
	.w3(32'hb81e964d),
	.w4(32'h3a239596),
	.w5(32'h3ab0bf0f),
	.w6(32'h3a67c3c2),
	.w7(32'h3a2a6a94),
	.w8(32'h3acbfe18),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64b4a2),
	.w1(32'h391b0a74),
	.w2(32'hb9060c88),
	.w3(32'h3a54b1f8),
	.w4(32'hb97a7865),
	.w5(32'hb95bdb6b),
	.w6(32'h390aef37),
	.w7(32'h3916dacd),
	.w8(32'hb9be412b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba088cef),
	.w1(32'hb60a98b1),
	.w2(32'h3a12c08b),
	.w3(32'hba157df6),
	.w4(32'hb9a5c54d),
	.w5(32'h3a345384),
	.w6(32'h3915655d),
	.w7(32'h394018d6),
	.w8(32'h3a4fda87),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0029be),
	.w1(32'h39d7e4ee),
	.w2(32'h3a53592e),
	.w3(32'h3962ece7),
	.w4(32'h390e0f7e),
	.w5(32'h3a80598c),
	.w6(32'hb8135c91),
	.w7(32'hb91cbaed),
	.w8(32'h3a619ff9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b97b3),
	.w1(32'h3a70fa3a),
	.w2(32'h3a8af340),
	.w3(32'h3ae7a4fa),
	.w4(32'h3a9a626c),
	.w5(32'h3a92f216),
	.w6(32'hb887c831),
	.w7(32'h3a53f450),
	.w8(32'h3ac77d27),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e4eff),
	.w1(32'h37aeba82),
	.w2(32'h389a2cf2),
	.w3(32'hb9aeec01),
	.w4(32'h3819675a),
	.w5(32'h392683d3),
	.w6(32'hb856209e),
	.w7(32'h385b1778),
	.w8(32'h38c26cf8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380d888c),
	.w1(32'hb9baad11),
	.w2(32'hb9897d3a),
	.w3(32'h393e9e93),
	.w4(32'hb962186e),
	.w5(32'h386df563),
	.w6(32'hb9c41765),
	.w7(32'hb8197a41),
	.w8(32'hb94825c6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983ffa4),
	.w1(32'h396a4cce),
	.w2(32'h381f490d),
	.w3(32'h39b985cb),
	.w4(32'hb7caa0d5),
	.w5(32'hb9540979),
	.w6(32'h3a8afc67),
	.w7(32'h3a79a191),
	.w8(32'h3a108594),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380904c5),
	.w1(32'hba50b972),
	.w2(32'h3a6fd6e0),
	.w3(32'hb95c3463),
	.w4(32'hba18c329),
	.w5(32'h3a89f92f),
	.w6(32'hb9d51fce),
	.w7(32'hb985054d),
	.w8(32'h3ac8a3ba),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c4abe),
	.w1(32'hb8c80a0b),
	.w2(32'h3999c6aa),
	.w3(32'hb9e3eadf),
	.w4(32'hba0862f9),
	.w5(32'h3a1072e2),
	.w6(32'hba001050),
	.w7(32'hb9a1d0df),
	.w8(32'h39c775ca),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f7369),
	.w1(32'h3a45e42e),
	.w2(32'h3a302bc9),
	.w3(32'hba1bc76a),
	.w4(32'h39b6cc5e),
	.w5(32'h39ebfea9),
	.w6(32'h3a16005a),
	.w7(32'h3a349426),
	.w8(32'h3a0a3560),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1569db),
	.w1(32'h395c7f3d),
	.w2(32'h399d3349),
	.w3(32'h39c011bf),
	.w4(32'h3951d569),
	.w5(32'h39823b77),
	.w6(32'h38c1d990),
	.w7(32'h3972a7b6),
	.w8(32'h39ae247d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ce243),
	.w1(32'hb8a75344),
	.w2(32'hb9ae57f5),
	.w3(32'h3a1c7bc3),
	.w4(32'hb6a21360),
	.w5(32'hb923f104),
	.w6(32'h3744a58f),
	.w7(32'hb816bb17),
	.w8(32'hb7c76327),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9976a20),
	.w1(32'h3a11be51),
	.w2(32'h3a272a50),
	.w3(32'hb99fce8d),
	.w4(32'h3a122cce),
	.w5(32'h39acc829),
	.w6(32'h39d95c06),
	.w7(32'h39df4c0e),
	.w8(32'h39a151d6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f03eb),
	.w1(32'h3b035a1c),
	.w2(32'h3ac20df5),
	.w3(32'h3b13a487),
	.w4(32'h3b2514d6),
	.w5(32'h3aa4feee),
	.w6(32'h3a80431b),
	.w7(32'h3a825848),
	.w8(32'h3a8434e8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90270a4),
	.w1(32'hba177ceb),
	.w2(32'hb8036f0a),
	.w3(32'hba44485d),
	.w4(32'hbaaf2058),
	.w5(32'h3902fc4c),
	.w6(32'hba7a0cbb),
	.w7(32'hba6297ef),
	.w8(32'h39ebd29d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c04b5),
	.w1(32'h382ae076),
	.w2(32'h39a48bcd),
	.w3(32'hb9f4a712),
	.w4(32'h38a4a52b),
	.w5(32'hb96f41a4),
	.w6(32'h3a8a9c6f),
	.w7(32'h3a62122b),
	.w8(32'hb893be9b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b1f68),
	.w1(32'hb8c0e5ea),
	.w2(32'h37f31c9f),
	.w3(32'h3941d9ea),
	.w4(32'hb9c9642c),
	.w5(32'hb9ca982f),
	.w6(32'hb99871af),
	.w7(32'hb9e5dbd2),
	.w8(32'hb9c94ac2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925c4ae),
	.w1(32'h39bfe0c3),
	.w2(32'h36e3b1d4),
	.w3(32'hb9852f39),
	.w4(32'h39794f39),
	.w5(32'h396fe469),
	.w6(32'h3a020d60),
	.w7(32'h39d786fa),
	.w8(32'h3986d111),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be1ceb),
	.w1(32'h398e32bb),
	.w2(32'h39c7f092),
	.w3(32'h38245055),
	.w4(32'h38e7914d),
	.w5(32'h383311c7),
	.w6(32'h3a01e1d2),
	.w7(32'h3a0bd711),
	.w8(32'h3987d3f6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f5a7b),
	.w1(32'hba1fab1e),
	.w2(32'hb951fad4),
	.w3(32'h396cc838),
	.w4(32'hba04d967),
	.w5(32'hba0f4baa),
	.w6(32'hb9beae7f),
	.w7(32'hb9a10a31),
	.w8(32'hba7ca660),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba617ecd),
	.w1(32'hb7abac02),
	.w2(32'h394b3429),
	.w3(32'hba83c5f5),
	.w4(32'h390d2149),
	.w5(32'h39a34978),
	.w6(32'hb7aec036),
	.w7(32'hb8570525),
	.w8(32'h37df7e71),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d7d1fd),
	.w1(32'h3728cdf1),
	.w2(32'hb9d12705),
	.w3(32'hb888e479),
	.w4(32'hb814b6da),
	.w5(32'hb98aa519),
	.w6(32'hb8b2fdcc),
	.w7(32'hb94a0c75),
	.w8(32'hb98f60cf),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93984f3),
	.w1(32'hb981df19),
	.w2(32'h3a95c554),
	.w3(32'hb98b2ec9),
	.w4(32'hba171b82),
	.w5(32'h3aa2923d),
	.w6(32'h3910ffa5),
	.w7(32'hb8ee442a),
	.w8(32'h3a2d2aa5),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7208837),
	.w1(32'h38fb59a4),
	.w2(32'h38f2a411),
	.w3(32'h38cc9664),
	.w4(32'h39c744b7),
	.w5(32'hb8971115),
	.w6(32'h3a05c7f9),
	.w7(32'hb8e25a2a),
	.w8(32'h3a5b20aa),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba085dee),
	.w1(32'h3a81c69b),
	.w2(32'h3a8d3ac9),
	.w3(32'hba0348e7),
	.w4(32'h38f14c98),
	.w5(32'h3a04f7f8),
	.w6(32'h39fbd2ce),
	.w7(32'h396ae7c1),
	.w8(32'h39ab5673),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eec86),
	.w1(32'h3a9f8952),
	.w2(32'h3ac0d4c7),
	.w3(32'h39ac8523),
	.w4(32'h3aa1f2fe),
	.w5(32'h3ad1c89f),
	.w6(32'h3aba1a2d),
	.w7(32'h3a8cf960),
	.w8(32'h3afc9a29),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2949b),
	.w1(32'h39eb89d0),
	.w2(32'h3a14be73),
	.w3(32'h3ab20025),
	.w4(32'h3a1e7296),
	.w5(32'h3a7b517b),
	.w6(32'h39ab74a1),
	.w7(32'h3a08bd45),
	.w8(32'h3a8ba6cc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef1b9d),
	.w1(32'h39bd1047),
	.w2(32'h39d0e62e),
	.w3(32'h3a0a55b3),
	.w4(32'h3a1ed0ab),
	.w5(32'h3a0e7f20),
	.w6(32'h3a16721d),
	.w7(32'h39fb725f),
	.w8(32'h3a34345e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bf1d2),
	.w1(32'h3a166783),
	.w2(32'h3a18b444),
	.w3(32'h3a6625d1),
	.w4(32'h3a18d86d),
	.w5(32'h3a696839),
	.w6(32'h39c12787),
	.w7(32'h3a0e6a6e),
	.w8(32'h3a60aada),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a278f27),
	.w1(32'h39d442e4),
	.w2(32'h38143ec4),
	.w3(32'h3a293eff),
	.w4(32'h39b3e3dd),
	.w5(32'h399ac07d),
	.w6(32'h3a2aaa79),
	.w7(32'h3a199b2b),
	.w8(32'h3a1294f3),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976a800),
	.w1(32'h39639c40),
	.w2(32'h3a025ab3),
	.w3(32'h397c04e4),
	.w4(32'h39a5b8e6),
	.w5(32'h3a08f06f),
	.w6(32'h39523391),
	.w7(32'h39cc5a14),
	.w8(32'h3a091d79),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a307ca2),
	.w1(32'h39f5101e),
	.w2(32'h39c325a7),
	.w3(32'h3a13a4c5),
	.w4(32'h3a298108),
	.w5(32'h3a05d6e6),
	.w6(32'h3a20afe8),
	.w7(32'h3a0fad78),
	.w8(32'h3a4ef486),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c3a29),
	.w1(32'h3a1fe038),
	.w2(32'h3a6ba74e),
	.w3(32'h3a4e5029),
	.w4(32'h3a2046c4),
	.w5(32'h3a6de718),
	.w6(32'h3a23439f),
	.w7(32'h3a71dfd2),
	.w8(32'h3a2d5733),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c152b),
	.w1(32'h39fa40ad),
	.w2(32'h3a451611),
	.w3(32'h3a934523),
	.w4(32'h3a0af068),
	.w5(32'h3a31257f),
	.w6(32'h3a9516b4),
	.w7(32'h3a7641c8),
	.w8(32'h3a5fffff),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b3d32),
	.w1(32'h3a449418),
	.w2(32'h3b07a8ec),
	.w3(32'h39d586eb),
	.w4(32'h3a1a4e82),
	.w5(32'h3b18f0da),
	.w6(32'h3893c632),
	.w7(32'h39c4b4df),
	.w8(32'h3ab34c21),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3962a3),
	.w1(32'h3a68661b),
	.w2(32'h3aa53a11),
	.w3(32'h39da73b7),
	.w4(32'h39bd6c9e),
	.w5(32'h3ac65194),
	.w6(32'hb9008dfd),
	.w7(32'h398493e4),
	.w8(32'h3a989747),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4223df),
	.w1(32'h3a5d29ea),
	.w2(32'h3a75dc4d),
	.w3(32'h39f537a0),
	.w4(32'h3a0de638),
	.w5(32'h3a8aa792),
	.w6(32'h3a373195),
	.w7(32'h3a1ce669),
	.w8(32'h3a97e5ad),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e12fa),
	.w1(32'h3aaecf98),
	.w2(32'h3ae211c8),
	.w3(32'h3a1c930a),
	.w4(32'h3ac46a6c),
	.w5(32'h3ad52a41),
	.w6(32'h3ab267f0),
	.w7(32'h3ad03980),
	.w8(32'h3ac92550),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae47945),
	.w1(32'h3a256c9a),
	.w2(32'h3a10cb0d),
	.w3(32'h3ad8a358),
	.w4(32'h3a7011a8),
	.w5(32'h3a49678c),
	.w6(32'h3a635f8e),
	.w7(32'h3a4d7524),
	.w8(32'h3a90b190),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87a8f3),
	.w1(32'h3a2150dd),
	.w2(32'h3a007e15),
	.w3(32'h3a9324a4),
	.w4(32'h3a518117),
	.w5(32'h3a387c61),
	.w6(32'h3a36432d),
	.w7(32'h3a289fdb),
	.w8(32'h3a36af36),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a558c65),
	.w1(32'h3a2119f5),
	.w2(32'h3a1fed29),
	.w3(32'h3a5ce2ac),
	.w4(32'h3a5054db),
	.w5(32'h3a54cc5d),
	.w6(32'h3a3262a4),
	.w7(32'h3a352a5a),
	.w8(32'h3a4435c4),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa07fc9),
	.w1(32'h3a5acc51),
	.w2(32'h3ab3db00),
	.w3(32'h3a8cbba0),
	.w4(32'h3a71ebd7),
	.w5(32'h3b1da078),
	.w6(32'h3a9aef59),
	.w7(32'h3ade85cf),
	.w8(32'h3b11e9a4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a8c14),
	.w1(32'hb92cc14a),
	.w2(32'hba1c7f7f),
	.w3(32'h3a86b3b7),
	.w4(32'hb94b0646),
	.w5(32'hba0bb423),
	.w6(32'hb9424332),
	.w7(32'hb9bafb15),
	.w8(32'hb9647cb6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de1255),
	.w1(32'h3818ca2a),
	.w2(32'hb7dc7662),
	.w3(32'hba680997),
	.w4(32'hb8fd5350),
	.w5(32'h39044194),
	.w6(32'h385a4926),
	.w7(32'h38b4c866),
	.w8(32'hb7f7aafe),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd17cc),
	.w1(32'hb697cf61),
	.w2(32'h39db53a9),
	.w3(32'h39c5d65f),
	.w4(32'h36e12473),
	.w5(32'h39c989d2),
	.w6(32'hb8db193a),
	.w7(32'h39b06174),
	.w8(32'h398d57df),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec082b),
	.w1(32'h3a054076),
	.w2(32'h39df3b4d),
	.w3(32'h39d0e40c),
	.w4(32'h3a309a5f),
	.w5(32'h3a1ed4bc),
	.w6(32'h3a1e276e),
	.w7(32'h3a24a0ab),
	.w8(32'h3a5319f6),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6daded),
	.w1(32'h39ab5772),
	.w2(32'h39ba18a8),
	.w3(32'h3a510740),
	.w4(32'hb77a1318),
	.w5(32'h3a8f60b4),
	.w6(32'h39f766f9),
	.w7(32'h3a010a8a),
	.w8(32'h3a726231),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f67ff),
	.w1(32'h392e3e3a),
	.w2(32'h3a3ebb55),
	.w3(32'h3a71571b),
	.w4(32'h39cc605e),
	.w5(32'h3a438680),
	.w6(32'h391b193f),
	.w7(32'h3a395c7a),
	.w8(32'h3a56fd89),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a851584),
	.w1(32'h39e7efa0),
	.w2(32'h3a163b5a),
	.w3(32'h3a7c0d3c),
	.w4(32'h39c85098),
	.w5(32'h3a229512),
	.w6(32'hb7454495),
	.w7(32'h39d26ecc),
	.w8(32'h3a2fdbc2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a69b9),
	.w1(32'hb860328a),
	.w2(32'hb8f673d5),
	.w3(32'h3a0bab52),
	.w4(32'hb838eab8),
	.w5(32'hb90ac8cf),
	.w6(32'hb82b42f9),
	.w7(32'hb8c0a6a9),
	.w8(32'hb88dff06),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe763b),
	.w1(32'h39bada05),
	.w2(32'h38b2ba41),
	.w3(32'h38a3a7cf),
	.w4(32'hb966bdf7),
	.w5(32'h390e4348),
	.w6(32'hb8fafaeb),
	.w7(32'h385d1bdf),
	.w8(32'h3974513f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule