module layer_8_featuremap_177(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe2a50),
	.w1(32'hba402511),
	.w2(32'hbba5b698),
	.w3(32'h3b91a8c8),
	.w4(32'hbc1b39d7),
	.w5(32'hbb79ede6),
	.w6(32'hbb65d195),
	.w7(32'h3c7145af),
	.w8(32'h3c90a0ad),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26847e),
	.w1(32'hbb30044a),
	.w2(32'hb93ed658),
	.w3(32'hbab72477),
	.w4(32'h3b14b9d7),
	.w5(32'h3bba3cff),
	.w6(32'hbb15b9c8),
	.w7(32'h39d13211),
	.w8(32'hba501c31),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb386a),
	.w1(32'hbaf2555e),
	.w2(32'hbbe5a88a),
	.w3(32'h39715fad),
	.w4(32'hbb7fbc98),
	.w5(32'hbb8d638f),
	.w6(32'h3b3fb399),
	.w7(32'h3bd5a707),
	.w8(32'h3c51b653),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bdeae),
	.w1(32'hbc9052fb),
	.w2(32'hbc72ed6f),
	.w3(32'hb979e7d4),
	.w4(32'hbc9fbd92),
	.w5(32'hbcb9833d),
	.w6(32'hbb86dbe4),
	.w7(32'h3c5ea266),
	.w8(32'h3c8a3334),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d711d),
	.w1(32'hbaf7280c),
	.w2(32'hba9b3113),
	.w3(32'hbc380575),
	.w4(32'h3acaa3e0),
	.w5(32'h3b9b5672),
	.w6(32'hbb388122),
	.w7(32'h3a9e0606),
	.w8(32'h3a012892),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d8b2f),
	.w1(32'hbc6518c9),
	.w2(32'hbcc5d524),
	.w3(32'h3b1b97ad),
	.w4(32'hbc438bce),
	.w5(32'hbc415b9a),
	.w6(32'h39a18e04),
	.w7(32'hbcc6df59),
	.w8(32'hbc46a640),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc412d0f),
	.w1(32'h3a225e59),
	.w2(32'h3a8d2064),
	.w3(32'hbb80e4b6),
	.w4(32'hbb69c0d5),
	.w5(32'hbb33c3c7),
	.w6(32'hbb7378a7),
	.w7(32'hbbb2e358),
	.w8(32'hbad90ee4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c95f2),
	.w1(32'hbb2e8bb7),
	.w2(32'h3bdc88b8),
	.w3(32'h3b07fdab),
	.w4(32'hbac06f57),
	.w5(32'h3b779a96),
	.w6(32'hbb466adb),
	.w7(32'hb9b4b3b6),
	.w8(32'h3bc82917),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ecf3c),
	.w1(32'h3b35e67b),
	.w2(32'h3aba21e6),
	.w3(32'hbbb17914),
	.w4(32'h3b86131d),
	.w5(32'h3b527ba1),
	.w6(32'hbad373a0),
	.w7(32'hbb66cf0f),
	.w8(32'hbb3358a5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaced807),
	.w1(32'hbbc58480),
	.w2(32'hbc4ada14),
	.w3(32'h3aa663b3),
	.w4(32'h3b08d24a),
	.w5(32'h38157011),
	.w6(32'hbb94cfc1),
	.w7(32'hbc3efa3e),
	.w8(32'hbb22f0d4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf0178),
	.w1(32'hbc2e8b25),
	.w2(32'h3c685204),
	.w3(32'hbbb1fd17),
	.w4(32'hbc987bc5),
	.w5(32'hbbcdce86),
	.w6(32'hba985883),
	.w7(32'h3ca2565d),
	.w8(32'h3b962794),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c900cfe),
	.w1(32'h3bbdeb0e),
	.w2(32'hbb18519f),
	.w3(32'hb96390cf),
	.w4(32'h3a1eb7eb),
	.w5(32'hbae18898),
	.w6(32'h3bac65bf),
	.w7(32'h3b09b6ef),
	.w8(32'hbb3bd644),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb7e57),
	.w1(32'h3c17177b),
	.w2(32'h3c1acf40),
	.w3(32'hb9868307),
	.w4(32'h3c0be666),
	.w5(32'h3c3fd00b),
	.w6(32'hbb93fae2),
	.w7(32'h39bb9580),
	.w8(32'h3b4c45c9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba2df2),
	.w1(32'hbd15b277),
	.w2(32'hbd485a46),
	.w3(32'hb9c6f51a),
	.w4(32'hbc9ffd0e),
	.w5(32'hbd02d7b2),
	.w6(32'hbc8f955f),
	.w7(32'hbc853b20),
	.w8(32'hbc38b15f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0691a5),
	.w1(32'h3afef6d3),
	.w2(32'h3ad631fa),
	.w3(32'hbcc9764e),
	.w4(32'hbb49ed5e),
	.w5(32'hbb0c63ee),
	.w6(32'hbb75c920),
	.w7(32'hbb0f42bd),
	.w8(32'hba7849f8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a07837),
	.w1(32'h3bce0372),
	.w2(32'h3bbe01fa),
	.w3(32'h384cae40),
	.w4(32'hbb88d7bd),
	.w5(32'hbc16cd13),
	.w6(32'hbbc63ee1),
	.w7(32'hbba9945e),
	.w8(32'hba75dc16),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb796b79),
	.w1(32'hbc7d01be),
	.w2(32'hbcda8371),
	.w3(32'hbb7c7637),
	.w4(32'hbc84122e),
	.w5(32'hbcadbd47),
	.w6(32'hbc84e40e),
	.w7(32'hbc696df9),
	.w8(32'hbcb2ae98),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7db953),
	.w1(32'h3c0236b0),
	.w2(32'h3b89b54c),
	.w3(32'hbca628f6),
	.w4(32'h3ba39b0a),
	.w5(32'h3c20b1d0),
	.w6(32'h3b7fbaa1),
	.w7(32'h3bbae3f6),
	.w8(32'h3c3f5282),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14ac23),
	.w1(32'hbc5ebdab),
	.w2(32'hbc902808),
	.w3(32'h3bc5246f),
	.w4(32'h3bccdcab),
	.w5(32'hbb9e0a2f),
	.w6(32'hbc498131),
	.w7(32'hbc2ebd8d),
	.w8(32'h3b4b4b9d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8902e2),
	.w1(32'h3b60de47),
	.w2(32'hba8f31a6),
	.w3(32'hbc027fb4),
	.w4(32'h3a9204ca),
	.w5(32'hba8c32d5),
	.w6(32'h3b39cd8b),
	.w7(32'hbb29cb94),
	.w8(32'hbabe5c0f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14e227),
	.w1(32'h3c2e9dff),
	.w2(32'h3bef1d55),
	.w3(32'h39d19ff9),
	.w4(32'h3be5f666),
	.w5(32'h3c6d11aa),
	.w6(32'h3bd885f1),
	.w7(32'h3bda1fce),
	.w8(32'hbb998276),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881e37),
	.w1(32'hbc23ea29),
	.w2(32'hbbba426e),
	.w3(32'h3ba768c2),
	.w4(32'hbc527d34),
	.w5(32'hbc2d26e5),
	.w6(32'h3b46dce1),
	.w7(32'hbbffd421),
	.w8(32'hbc3f4180),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fdef7),
	.w1(32'hbb685fb4),
	.w2(32'hbc945904),
	.w3(32'hbb48cdec),
	.w4(32'hbb46cdd6),
	.w5(32'hbbe36e03),
	.w6(32'h3b874d77),
	.w7(32'hbb82db8c),
	.w8(32'hbb768aa5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcad1e8),
	.w1(32'hbb9ed89d),
	.w2(32'hbba57f9d),
	.w3(32'hbacbe6bd),
	.w4(32'hbbd2b414),
	.w5(32'hbb3d6bd9),
	.w6(32'hbb53cfd7),
	.w7(32'hbc39d0a0),
	.w8(32'hbbacfdba),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d4c80),
	.w1(32'hbbf15871),
	.w2(32'hbad38fe4),
	.w3(32'h38473dd7),
	.w4(32'hbbad561d),
	.w5(32'h3bf4f231),
	.w6(32'hbb8a3086),
	.w7(32'hbacbda50),
	.w8(32'h3b38df15),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4eab19),
	.w1(32'h3c2be292),
	.w2(32'h3c1cdea9),
	.w3(32'h3bdd5e14),
	.w4(32'h3988c32b),
	.w5(32'h3bed02e5),
	.w6(32'h3b8e7b83),
	.w7(32'h3ac2d6b6),
	.w8(32'hbb5acf5c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc68a4c),
	.w1(32'h3b672380),
	.w2(32'h3c491da0),
	.w3(32'h3c1ac02d),
	.w4(32'h3be6fb4d),
	.w5(32'h3b320867),
	.w6(32'h3bb35930),
	.w7(32'h3c16653f),
	.w8(32'h3b637272),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9345ca9),
	.w1(32'hbbbc4ef6),
	.w2(32'h3c884410),
	.w3(32'hbbb8eecb),
	.w4(32'h3b6bbb5b),
	.w5(32'hbabbd06c),
	.w6(32'hbacb9238),
	.w7(32'h3c4f24d9),
	.w8(32'h3c5dc1a8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8642c7),
	.w1(32'h3b6741c0),
	.w2(32'h3b9c0b3c),
	.w3(32'h3be1339a),
	.w4(32'hbba0f77d),
	.w5(32'hbb4c0dd1),
	.w6(32'h3a41bef3),
	.w7(32'hbb0b77e8),
	.w8(32'h3aa273f1),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09a12d),
	.w1(32'h3aaa6bc5),
	.w2(32'h3c0094ca),
	.w3(32'hbb81d984),
	.w4(32'h3c3c998a),
	.w5(32'h3c87336b),
	.w6(32'hbb6657cf),
	.w7(32'h3b033d09),
	.w8(32'h3acc5644),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ea1c2),
	.w1(32'h3a61e4fb),
	.w2(32'h3abcab08),
	.w3(32'h3c4fe9d2),
	.w4(32'h3b341def),
	.w5(32'h3a8b2585),
	.w6(32'hbace4be7),
	.w7(32'hbb237c61),
	.w8(32'h3c1be6fd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05a08a),
	.w1(32'h3c13273e),
	.w2(32'h3c6d5ab7),
	.w3(32'hbae9e794),
	.w4(32'h3ba3c419),
	.w5(32'h3c442b27),
	.w6(32'h3b990d11),
	.w7(32'h3bc8b001),
	.w8(32'hbb5ae851),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d6901),
	.w1(32'hbc32bd03),
	.w2(32'hbc9d6b46),
	.w3(32'h3bd91407),
	.w4(32'hbc660dd4),
	.w5(32'hbcb682cf),
	.w6(32'hbc042ae4),
	.w7(32'hbbae5fee),
	.w8(32'hbb578149),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e8ae2),
	.w1(32'hbd086c5d),
	.w2(32'hbda6f95c),
	.w3(32'hbc3dcc8e),
	.w4(32'hbce546fb),
	.w5(32'hbd638365),
	.w6(32'hbcef1a98),
	.w7(32'hbd3992f1),
	.w8(32'hbca0a668),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd42429d),
	.w1(32'h3c05a66f),
	.w2(32'h3b85f352),
	.w3(32'hbd14c93b),
	.w4(32'h3b8813f2),
	.w5(32'h3be8b7c6),
	.w6(32'h3bd46ff0),
	.w7(32'h3b68014e),
	.w8(32'h3b900560),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb929d),
	.w1(32'h3c8bf829),
	.w2(32'h3cf53c27),
	.w3(32'h3ba5ec62),
	.w4(32'h3c8d3f70),
	.w5(32'h3ce3957f),
	.w6(32'h3aeb0b0c),
	.w7(32'h3b9b12a9),
	.w8(32'h3c0ca1bf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c855454),
	.w1(32'h3bcd3ef5),
	.w2(32'h3c0e379a),
	.w3(32'h3c39538d),
	.w4(32'h3993b827),
	.w5(32'h3b46bbed),
	.w6(32'h3be3a0b0),
	.w7(32'h3beb83f9),
	.w8(32'h3b8131dd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf31eaf),
	.w1(32'h3b6a6f82),
	.w2(32'h3bed0de2),
	.w3(32'h3b080f78),
	.w4(32'hbad850ba),
	.w5(32'h3b730e0f),
	.w6(32'hb8f38a7a),
	.w7(32'h3c001493),
	.w8(32'h3ba99a7d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb28c16),
	.w1(32'h3c8b9b9d),
	.w2(32'h3cdd9fcb),
	.w3(32'h3b95453e),
	.w4(32'h3c8adff1),
	.w5(32'h3c6891e0),
	.w6(32'hbb1fbd19),
	.w7(32'h3c400ae8),
	.w8(32'h3c130417),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6fe9c),
	.w1(32'h3b2bff71),
	.w2(32'h3c7ae0f1),
	.w3(32'h39d85818),
	.w4(32'h3b008eb9),
	.w5(32'h3c2bd741),
	.w6(32'hbb61907a),
	.w7(32'hbabb9b43),
	.w8(32'hbb8efd54),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f2f81),
	.w1(32'h3c43b2cf),
	.w2(32'h3c0154f5),
	.w3(32'h3bcad051),
	.w4(32'h3c358497),
	.w5(32'h3c19680e),
	.w6(32'h3c1dfc52),
	.w7(32'h3c059429),
	.w8(32'h3c2f2508),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b1f31),
	.w1(32'hbb4d92d4),
	.w2(32'hbbf4b418),
	.w3(32'h3c5058b2),
	.w4(32'h3b1f5e14),
	.w5(32'hbb94b2ff),
	.w6(32'hbb9b8ea2),
	.w7(32'hbbd39e01),
	.w8(32'h3a0964eb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abedc0d),
	.w1(32'hba3bcfb3),
	.w2(32'hbb085ec1),
	.w3(32'h3b09fe4c),
	.w4(32'hbb1df618),
	.w5(32'hbb694a16),
	.w6(32'h3b87e643),
	.w7(32'h3c08975b),
	.w8(32'hbb0889a8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa72469),
	.w1(32'h3c927451),
	.w2(32'h3d0f5fe7),
	.w3(32'hb9c50a02),
	.w4(32'h3c903c97),
	.w5(32'h3cba48a9),
	.w6(32'h3c2ff248),
	.w7(32'h3ca61a15),
	.w8(32'h3c933a9a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce11f6a),
	.w1(32'hbc90828d),
	.w2(32'hbd0ea3d4),
	.w3(32'h3c97c050),
	.w4(32'hbcd7cdd9),
	.w5(32'hbcfd7898),
	.w6(32'hbb8ddc65),
	.w7(32'hbcc2806b),
	.w8(32'hbcf1ae5a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a1072),
	.w1(32'h3ba03f31),
	.w2(32'h3af4bef4),
	.w3(32'hbcbf57c8),
	.w4(32'h3b98bdbe),
	.w5(32'h3bbac0b0),
	.w6(32'h3bc4fc39),
	.w7(32'hbaf9298a),
	.w8(32'h3a7721a4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22e866),
	.w1(32'hbc01b6a5),
	.w2(32'hbae9cbdb),
	.w3(32'h399f8072),
	.w4(32'hbba8f1f1),
	.w5(32'hbbbbfec0),
	.w6(32'hbc5e64e0),
	.w7(32'hbaf0ad99),
	.w8(32'h3b8027ca),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96f8ae),
	.w1(32'h3d0ca84c),
	.w2(32'h3d6b9239),
	.w3(32'hbbc9a55e),
	.w4(32'h3cd0bf46),
	.w5(32'h3d427060),
	.w6(32'h3c362323),
	.w7(32'h3cc91fdb),
	.w8(32'h3cc25903),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0b549a),
	.w1(32'h3d0b7177),
	.w2(32'h3d3f3056),
	.w3(32'h3d037a82),
	.w4(32'h3d0007a2),
	.w5(32'h3d2db274),
	.w6(32'h3c7211ab),
	.w7(32'h3ce95501),
	.w8(32'h3cdebcae),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdfc50b),
	.w1(32'hb8ff815b),
	.w2(32'h3b9aff82),
	.w3(32'h3ce6340a),
	.w4(32'h3be6ec98),
	.w5(32'hb8cf007b),
	.w6(32'h3b075a34),
	.w7(32'hba5bb6ea),
	.w8(32'h3c43964a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38bfc1),
	.w1(32'h3a95424e),
	.w2(32'hbc0e4ff0),
	.w3(32'h3b998257),
	.w4(32'h3a6f45ec),
	.w5(32'hbc1a6f3e),
	.w6(32'h3a9641bc),
	.w7(32'hbbf319cf),
	.w8(32'h399541c5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb051313),
	.w1(32'hbb6d1ff1),
	.w2(32'h3acbc8cc),
	.w3(32'hbab0ae95),
	.w4(32'h38a92114),
	.w5(32'h3bb09996),
	.w6(32'h3b273c36),
	.w7(32'hb7b3aa96),
	.w8(32'h3829d19d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ef85a),
	.w1(32'hbb65a6ba),
	.w2(32'h3b5f84b6),
	.w3(32'h3bbe382f),
	.w4(32'hbb71d9fe),
	.w5(32'h3b8a69d6),
	.w6(32'hbbcf5e56),
	.w7(32'h3bbaeb54),
	.w8(32'hba163e99),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4057d2),
	.w1(32'h3b259f6d),
	.w2(32'h3c91303b),
	.w3(32'hbb02ccf7),
	.w4(32'h3b20267c),
	.w5(32'h3c641772),
	.w6(32'h3bbd84fe),
	.w7(32'h3c84b72a),
	.w8(32'hbb1c64cc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3aff),
	.w1(32'h382f8b53),
	.w2(32'hbc0b0c1d),
	.w3(32'h3b9845d3),
	.w4(32'h3c5e0198),
	.w5(32'hbbf78a2b),
	.w6(32'h3a747b97),
	.w7(32'hbafe6e91),
	.w8(32'h3b0e9b39),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7385f1),
	.w1(32'h3ba14f8e),
	.w2(32'hbafc6a2e),
	.w3(32'hbc07bae4),
	.w4(32'h3bfb8aa6),
	.w5(32'hbbbd76b1),
	.w6(32'h3c4ba9c4),
	.w7(32'h3bec9b6a),
	.w8(32'h3b740a66),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7134c4),
	.w1(32'h3ba4868b),
	.w2(32'hbbeaf100),
	.w3(32'h3b9346c1),
	.w4(32'hb9a1824d),
	.w5(32'hbc31cd6a),
	.w6(32'h3ad251f1),
	.w7(32'h3b49918a),
	.w8(32'h39dba67a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9292b0),
	.w1(32'h3a908d0c),
	.w2(32'hbc19b43e),
	.w3(32'h3a7fab1c),
	.w4(32'hb9b98f0f),
	.w5(32'hbbcbaade),
	.w6(32'h386995d2),
	.w7(32'hbbbb51db),
	.w8(32'hbb5496e8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc064acc),
	.w1(32'hbb7a4bde),
	.w2(32'hbbd83b9c),
	.w3(32'hbc18bc70),
	.w4(32'hbbaf337d),
	.w5(32'hbc088f8d),
	.w6(32'hbb68da06),
	.w7(32'hbb30c15a),
	.w8(32'hbb4a7b71),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec19a5),
	.w1(32'hbc2a9d2f),
	.w2(32'hbc8d0b6b),
	.w3(32'hbc17e86c),
	.w4(32'hbc43d404),
	.w5(32'hbbf37f29),
	.w6(32'hbb328cba),
	.w7(32'hbbdae55a),
	.w8(32'hbc7e4484),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc685795),
	.w1(32'hbbff37f3),
	.w2(32'hbaa9288d),
	.w3(32'hbb8592f2),
	.w4(32'hbc024855),
	.w5(32'hbbef5d8d),
	.w6(32'hbc4c3cd2),
	.w7(32'hbac81949),
	.w8(32'h3b6fd715),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963b5b9),
	.w1(32'h3c4e3864),
	.w2(32'h3c12d8a2),
	.w3(32'hbbe3c571),
	.w4(32'h3b9e211c),
	.w5(32'h3be6b7ef),
	.w6(32'h3a50cc86),
	.w7(32'hba9dc3c0),
	.w8(32'hbb2c7473),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befea32),
	.w1(32'h3b999cfd),
	.w2(32'h3c7583c9),
	.w3(32'h3c30843c),
	.w4(32'h3b9b92af),
	.w5(32'h3c98606e),
	.w6(32'h3bad094c),
	.w7(32'h3b1f3c90),
	.w8(32'h3b681096),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2794ba),
	.w1(32'h3bb39607),
	.w2(32'h39238a57),
	.w3(32'h3c7fbe8b),
	.w4(32'h3b7d5bb3),
	.w5(32'h3a909a36),
	.w6(32'h3c156df8),
	.w7(32'h3a854c11),
	.w8(32'h3b8ffdf6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5c341),
	.w1(32'h3b89db5b),
	.w2(32'h3ba7cccc),
	.w3(32'hbb9e58be),
	.w4(32'h3a332c0d),
	.w5(32'h3b9a2742),
	.w6(32'h3a8862e4),
	.w7(32'hba56bb86),
	.w8(32'hbbc70079),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39904d8f),
	.w1(32'h3c4eaebd),
	.w2(32'h3c83f8d3),
	.w3(32'h3a1a0ad9),
	.w4(32'h3a78f375),
	.w5(32'h3cb88c7e),
	.w6(32'hba81d09e),
	.w7(32'h3a3552b1),
	.w8(32'h3ab5f671),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b00e7),
	.w1(32'h3c81622d),
	.w2(32'h3d0d3ada),
	.w3(32'h3c628b37),
	.w4(32'h3c0835e6),
	.w5(32'h3ca34bff),
	.w6(32'h3c0d39d8),
	.w7(32'h3cf235e6),
	.w8(32'h3c3e12d5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5f155),
	.w1(32'h3c8324a5),
	.w2(32'h3c177978),
	.w3(32'h3c4c14d0),
	.w4(32'h3b88ce9a),
	.w5(32'hbad7db49),
	.w6(32'h3c14f3e5),
	.w7(32'h3bb7d147),
	.w8(32'h3b412b9f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7de6a6),
	.w1(32'hbcb3393b),
	.w2(32'hbd2ab7ad),
	.w3(32'h3b6c704e),
	.w4(32'hbc16ae62),
	.w5(32'hbd0e7c1c),
	.w6(32'hbc2d7c72),
	.w7(32'hbc9cd765),
	.w8(32'hbba4bb15),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b9840),
	.w1(32'h3c0b26aa),
	.w2(32'h39a54403),
	.w3(32'hbc6b41a1),
	.w4(32'hb9d08e44),
	.w5(32'h3c032983),
	.w6(32'h3c28af56),
	.w7(32'h3b97aeef),
	.w8(32'h3c076feb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc15675),
	.w1(32'hba9ea1a4),
	.w2(32'h3c50cfda),
	.w3(32'h3b8078d2),
	.w4(32'hbace6ba3),
	.w5(32'h3baeef66),
	.w6(32'h3a17e7c7),
	.w7(32'h3c486768),
	.w8(32'hbb532e8d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfe882),
	.w1(32'hbcdb1670),
	.w2(32'hbd251bd6),
	.w3(32'h3b2cc313),
	.w4(32'hbc816ab1),
	.w5(32'hbd108a2c),
	.w6(32'hbc01f52f),
	.w7(32'hbc22edb7),
	.w8(32'hbc32231c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f7ee9),
	.w1(32'h3bbe32c7),
	.w2(32'hbb8a3628),
	.w3(32'hbbea984c),
	.w4(32'h3b17dfcc),
	.w5(32'hbac4e672),
	.w6(32'h3c153bb4),
	.w7(32'h3bddcb7b),
	.w8(32'h3b8a80a6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc190b2d),
	.w1(32'hbbba4bda),
	.w2(32'hbb7d24e9),
	.w3(32'hbb2f5b5c),
	.w4(32'hbb98dced),
	.w5(32'hbc02ce66),
	.w6(32'hbbaef086),
	.w7(32'hba3b9d44),
	.w8(32'h3b26cc85),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb538685),
	.w1(32'h3b341248),
	.w2(32'h3b7d4ead),
	.w3(32'hbc2c3862),
	.w4(32'hb9f32240),
	.w5(32'h3c04e8ee),
	.w6(32'h3a95497e),
	.w7(32'hb9ef77c2),
	.w8(32'hbc05513d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc98ccd),
	.w1(32'hbbbc167a),
	.w2(32'h3a693824),
	.w3(32'h3aee2932),
	.w4(32'hbb4b72a2),
	.w5(32'hbaddf2e2),
	.w6(32'h38fe8306),
	.w7(32'h3c1595e2),
	.w8(32'hba14d71c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd17864),
	.w1(32'h3b47c7d7),
	.w2(32'h3bad0900),
	.w3(32'hbc1699e0),
	.w4(32'hbb363162),
	.w5(32'h39e58049),
	.w6(32'hb99b232d),
	.w7(32'hbae89b87),
	.w8(32'h3af308c4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6561e7),
	.w1(32'hbbbd8d1e),
	.w2(32'h3a95895c),
	.w3(32'h3b805f24),
	.w4(32'hbbd180c3),
	.w5(32'hbab97d1c),
	.w6(32'hba77fc62),
	.w7(32'h3bb8c497),
	.w8(32'h3ba5e3de),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3889c5d7),
	.w1(32'hbb8f7ce0),
	.w2(32'hbbb5bd95),
	.w3(32'hbb4819bf),
	.w4(32'hbb7954ee),
	.w5(32'hbbec1a25),
	.w6(32'hbaf9273b),
	.w7(32'h3b2fad29),
	.w8(32'h3c487ecb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babd0dd),
	.w1(32'hbbf45e79),
	.w2(32'hbaf5abac),
	.w3(32'hbb83b95c),
	.w4(32'h39ec8bde),
	.w5(32'hbbc5a841),
	.w6(32'h3a8d9b55),
	.w7(32'h3bda6092),
	.w8(32'h3c55efaa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3adb8a),
	.w1(32'hbc595bb1),
	.w2(32'hbc8583cc),
	.w3(32'h3bef4e86),
	.w4(32'hbbc9a08e),
	.w5(32'hbc3bacf6),
	.w6(32'hbc054404),
	.w7(32'hbb4848fd),
	.w8(32'h3be20109),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8843a7),
	.w1(32'hbccd3919),
	.w2(32'hbd091c1c),
	.w3(32'h3abbb89a),
	.w4(32'hbbebd2d5),
	.w5(32'hbd00788b),
	.w6(32'hbcd50c5a),
	.w7(32'hbca5bf71),
	.w8(32'hbbccca31),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8036bd),
	.w1(32'hbc484ab7),
	.w2(32'hbc269cbe),
	.w3(32'hbc5ee34b),
	.w4(32'hbc2c4cc2),
	.w5(32'hbc38defc),
	.w6(32'h3b0b3b7a),
	.w7(32'h3aa83996),
	.w8(32'hbbbed128),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb837e41),
	.w1(32'hbbc262d0),
	.w2(32'hbc60183e),
	.w3(32'hbc2fcc0c),
	.w4(32'hbba0f620),
	.w5(32'hbc3364e8),
	.w6(32'h3a69f892),
	.w7(32'hbc32355a),
	.w8(32'hbb088726),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc95aa),
	.w1(32'hbcc1e6da),
	.w2(32'hbcffcb8f),
	.w3(32'hbc214b15),
	.w4(32'hbcb8cfe0),
	.w5(32'hbce60ba1),
	.w6(32'hbc553df7),
	.w7(32'hbbd2c556),
	.w8(32'h3c1344d2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f767c),
	.w1(32'h3b6380f3),
	.w2(32'hbbaa362d),
	.w3(32'hbc77400c),
	.w4(32'h3b266e1a),
	.w5(32'h3ae70800),
	.w6(32'h3a1c669a),
	.w7(32'h3aa31e4b),
	.w8(32'h3b6ce39b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa96266),
	.w1(32'h3b28a0b3),
	.w2(32'h3b5a02c9),
	.w3(32'h3a8e01a0),
	.w4(32'h3bbc99c3),
	.w5(32'h3bcc7d04),
	.w6(32'h3b21bf79),
	.w7(32'h3ba7dde7),
	.w8(32'h3b6ea4b5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09e82b),
	.w1(32'hbabd7e40),
	.w2(32'h3b8aaa56),
	.w3(32'h3bb026e6),
	.w4(32'hbc786058),
	.w5(32'hbbb0c97c),
	.w6(32'h3c3aca6c),
	.w7(32'h3ba4107b),
	.w8(32'hbabd56d5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba05736),
	.w1(32'hbb0cd3db),
	.w2(32'hbba8f5b7),
	.w3(32'h3a653828),
	.w4(32'hbbd85c72),
	.w5(32'hbc03f5a8),
	.w6(32'hba39f192),
	.w7(32'h3a8dd108),
	.w8(32'h3b824888),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03737b),
	.w1(32'h3c819fdc),
	.w2(32'h3c5b5482),
	.w3(32'hbbe95524),
	.w4(32'h3c4510cb),
	.w5(32'h3c27beab),
	.w6(32'h3c660b04),
	.w7(32'h3c9ba419),
	.w8(32'h3c28f38b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43affd),
	.w1(32'hbc0afbc3),
	.w2(32'hbc6b32f5),
	.w3(32'h3c5450f6),
	.w4(32'hbc06192e),
	.w5(32'hbcae0c49),
	.w6(32'h3b81d610),
	.w7(32'h3b9a6996),
	.w8(32'hba949500),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf24d3a),
	.w1(32'hbd155d39),
	.w2(32'hbd88a5dc),
	.w3(32'hbb98626d),
	.w4(32'hbcd1e094),
	.w5(32'hbd5a6ba2),
	.w6(32'hbcd3035a),
	.w7(32'hbd0df852),
	.w8(32'hbcfedf4e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3b3d6b),
	.w1(32'h3a922e94),
	.w2(32'hba0224e8),
	.w3(32'hbd159b8b),
	.w4(32'h3b05fe66),
	.w5(32'h3ad048d8),
	.w6(32'h3b955449),
	.w7(32'h3adb047a),
	.w8(32'hbb4393ee),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb827535),
	.w1(32'h39e94659),
	.w2(32'h3ba2a65a),
	.w3(32'hba35c607),
	.w4(32'h3af102c4),
	.w5(32'h3b84ec18),
	.w6(32'h3acc659d),
	.w7(32'h3b3b5fd7),
	.w8(32'h3b13c8f3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dbb54),
	.w1(32'h3bf95cf5),
	.w2(32'h3b0cd1ac),
	.w3(32'h3b67bee5),
	.w4(32'h3c2aa818),
	.w5(32'h3bfbcb09),
	.w6(32'hbb99301c),
	.w7(32'h3abd0349),
	.w8(32'hbac66237),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a1a5c),
	.w1(32'hbb689723),
	.w2(32'hbb921b61),
	.w3(32'hbb47dc52),
	.w4(32'hbba987e2),
	.w5(32'hbbc3f5ed),
	.w6(32'hbb728fc3),
	.w7(32'hbb603383),
	.w8(32'hbb1fc51b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc14e14),
	.w1(32'hbab1d744),
	.w2(32'hbb8f82bc),
	.w3(32'hbbef3cdb),
	.w4(32'h39c5c8fe),
	.w5(32'hbb8695a2),
	.w6(32'hba631f71),
	.w7(32'hbbf419ef),
	.w8(32'hbb77de9d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c820d),
	.w1(32'h3c57f23a),
	.w2(32'h3cbd7873),
	.w3(32'hbbd282af),
	.w4(32'h3c039698),
	.w5(32'h3c3abe67),
	.w6(32'h3c263cdd),
	.w7(32'h3c4448f8),
	.w8(32'h3c55a34e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59224b),
	.w1(32'h3cc690f7),
	.w2(32'h3d3b4c48),
	.w3(32'hb8c090c3),
	.w4(32'h3cc18aa5),
	.w5(32'h3d0fa2e5),
	.w6(32'h3bb4b905),
	.w7(32'h3cc07429),
	.w8(32'h3c88593d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8dcb5),
	.w1(32'hbc06bf7a),
	.w2(32'hbb4a6b4e),
	.w3(32'h3c72cdbf),
	.w4(32'hbbca8863),
	.w5(32'hbc2a0270),
	.w6(32'h3bd9dd19),
	.w7(32'h3c3bbcc0),
	.w8(32'h3bb1ce6e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb325d3b),
	.w1(32'h3c13ef24),
	.w2(32'h3bd331f3),
	.w3(32'hbb96ff5d),
	.w4(32'h3b3720fe),
	.w5(32'hbb05b3e6),
	.w6(32'h3a42f2a6),
	.w7(32'h3b6fe905),
	.w8(32'h3c30fdf4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14a0eb),
	.w1(32'hbc7d1152),
	.w2(32'hbcff2bce),
	.w3(32'hbb10594e),
	.w4(32'hbbd38b40),
	.w5(32'hbc14d191),
	.w6(32'hba932605),
	.w7(32'hbc8fbd88),
	.w8(32'hbbd815cf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d02d2),
	.w1(32'hbd05d129),
	.w2(32'hbd73a889),
	.w3(32'hbc790e8c),
	.w4(32'hbcc05853),
	.w5(32'hbd18472a),
	.w6(32'hbc9bc507),
	.w7(32'hbcc55fb3),
	.w8(32'hbc5df8d0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1861c5),
	.w1(32'h3c571b1e),
	.w2(32'h3c56706a),
	.w3(32'hbd0e0e3c),
	.w4(32'h3aedb003),
	.w5(32'h3c977642),
	.w6(32'h3bbd88f2),
	.w7(32'h3c484509),
	.w8(32'h3c1eae34),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e856c),
	.w1(32'h3cc1f2af),
	.w2(32'h3c86f7f0),
	.w3(32'h3c8f67c7),
	.w4(32'h3c83ce4a),
	.w5(32'h3b33adaa),
	.w6(32'h3bd7d211),
	.w7(32'h3bdb3b61),
	.w8(32'h3bb3a797),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfed860),
	.w1(32'hbb0cb8b9),
	.w2(32'hba303161),
	.w3(32'hbb98a700),
	.w4(32'hbb97f44d),
	.w5(32'hbb9409f3),
	.w6(32'hbb89539f),
	.w7(32'hbb9d9b34),
	.w8(32'hbc17d44b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc069fd1),
	.w1(32'h3aed0bef),
	.w2(32'h3bac6a19),
	.w3(32'hbc2632dd),
	.w4(32'h3b9147d6),
	.w5(32'h3bc9a68c),
	.w6(32'h3b85e54f),
	.w7(32'h3a3f9db7),
	.w8(32'h3b1c31ac),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c7ec8),
	.w1(32'h3b1b742f),
	.w2(32'hbba2e9ab),
	.w3(32'h3be5f28a),
	.w4(32'h3b74858b),
	.w5(32'h3b42edc3),
	.w6(32'hbb5eea5c),
	.w7(32'hbaa7402b),
	.w8(32'h3b327bad),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0059a),
	.w1(32'h3c4ba22d),
	.w2(32'h3c0e09ca),
	.w3(32'hbba5f4b4),
	.w4(32'h3b234b2d),
	.w5(32'h3b87fe69),
	.w6(32'h3b945fca),
	.w7(32'h3bb4e628),
	.w8(32'h3a92c181),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48ff98),
	.w1(32'hbaf7b5b5),
	.w2(32'h3a8333a1),
	.w3(32'hba964a98),
	.w4(32'h3afd4234),
	.w5(32'h3b934255),
	.w6(32'hbb0b5bc6),
	.w7(32'h3b160523),
	.w8(32'hbb009444),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db067a),
	.w1(32'hbcd494cb),
	.w2(32'hbd4be806),
	.w3(32'hb9e491e3),
	.w4(32'hbce5da93),
	.w5(32'hbd4f29dc),
	.w6(32'hbc1d4d4d),
	.w7(32'hbc2e8bb5),
	.w8(32'hbc97c71d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d054c),
	.w1(32'h3bc49829),
	.w2(32'h3b6a80a4),
	.w3(32'hbd15afb6),
	.w4(32'h3a445c88),
	.w5(32'h3b1e3586),
	.w6(32'h3c0d92b4),
	.w7(32'hba7cb2ef),
	.w8(32'hbb9909c9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57560c),
	.w1(32'hbc76a30f),
	.w2(32'hbd26f139),
	.w3(32'h3973802e),
	.w4(32'hbc946ee9),
	.w5(32'hbcb8ed7b),
	.w6(32'hbbaf698a),
	.w7(32'hbcbc4601),
	.w8(32'hbc8d0b8a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2db71),
	.w1(32'h3b647472),
	.w2(32'h3cab3914),
	.w3(32'hbabd5f91),
	.w4(32'h3c053f92),
	.w5(32'h3c6f5f05),
	.w6(32'h3bdc270e),
	.w7(32'h3c9b7030),
	.w8(32'h3c8b20f8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c788ef1),
	.w1(32'h3b8a439a),
	.w2(32'h3b197b0a),
	.w3(32'h3c320a3b),
	.w4(32'hba6aa133),
	.w5(32'hbaae77b5),
	.w6(32'h3b143517),
	.w7(32'h3bd5e6de),
	.w8(32'h3bc1131c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ad1e7),
	.w1(32'hbab9ae1b),
	.w2(32'h3ba8e250),
	.w3(32'hbb3f81a6),
	.w4(32'h3adafc1a),
	.w5(32'h3c04a06f),
	.w6(32'hbb5da66a),
	.w7(32'h3b7d53a3),
	.w8(32'hbb3bd71a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad93e33),
	.w1(32'hbbd90d81),
	.w2(32'hbb9e4f56),
	.w3(32'h3af9f0d4),
	.w4(32'hbb128278),
	.w5(32'h3aa93f93),
	.w6(32'hbc02e144),
	.w7(32'hbc081c0a),
	.w8(32'hbc2da805),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0aee03),
	.w1(32'hbc53c2cb),
	.w2(32'hbd1532bf),
	.w3(32'h3b509ec3),
	.w4(32'hbc451af0),
	.w5(32'hbd0f7634),
	.w6(32'hbc1cb098),
	.w7(32'hbcdf2acd),
	.w8(32'hbc6d0aff),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb212e4),
	.w1(32'hbcbbee75),
	.w2(32'hbd21e12d),
	.w3(32'hbc97ddfc),
	.w4(32'hb956da7a),
	.w5(32'hbd05b2c0),
	.w6(32'hbc2ba5d0),
	.w7(32'hbccbe09d),
	.w8(32'hbb904e4a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b49ff),
	.w1(32'hbbbad63b),
	.w2(32'hbc1131e8),
	.w3(32'hbcd9f5a1),
	.w4(32'hbc0974a2),
	.w5(32'hbc109bc8),
	.w6(32'hbad275f6),
	.w7(32'hbae6c884),
	.w8(32'hbb5854b2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98adc2),
	.w1(32'hbc8b551f),
	.w2(32'hbd43df51),
	.w3(32'hbc4c212f),
	.w4(32'hbc553e60),
	.w5(32'hbd23cb41),
	.w6(32'hbc34704a),
	.w7(32'hbc96bf14),
	.w8(32'hbb25d386),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc965342),
	.w1(32'hbba0d1ae),
	.w2(32'hbc027b76),
	.w3(32'hbc91f9d7),
	.w4(32'hbc33f17c),
	.w5(32'hbbfcbd5a),
	.w6(32'hbbb18711),
	.w7(32'h3c1fcc79),
	.w8(32'h3be27b5b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b57bf),
	.w1(32'hbb850adb),
	.w2(32'hbba055e1),
	.w3(32'hbbcad8cf),
	.w4(32'hb9557e71),
	.w5(32'h39eb2df0),
	.w6(32'hb9d42427),
	.w7(32'hbb3a3bc0),
	.w8(32'hbb9c0c48),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75bb6),
	.w1(32'hbb9efdc1),
	.w2(32'hbc79a5ee),
	.w3(32'hbb6bfc6b),
	.w4(32'hbbb23e4e),
	.w5(32'hbc21fea4),
	.w6(32'hbb38892a),
	.w7(32'hbc42d6d3),
	.w8(32'hbba3e7f5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4b0a3),
	.w1(32'hbcbe9367),
	.w2(32'hbd399f1e),
	.w3(32'h3acd76ef),
	.w4(32'h3b82dfeb),
	.w5(32'hbc6531c2),
	.w6(32'hbca41024),
	.w7(32'hbcf6a659),
	.w8(32'hbc1a3380),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6767a),
	.w1(32'h3ce83fd8),
	.w2(32'h3d5dec00),
	.w3(32'hbc713c74),
	.w4(32'h3cd7db60),
	.w5(32'h3d4861a9),
	.w6(32'h3c576ddf),
	.w7(32'h3cc356d9),
	.w8(32'h3cb3951d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08170d),
	.w1(32'h39ab2b89),
	.w2(32'hbb0bc1dc),
	.w3(32'h3cf6ebd8),
	.w4(32'h3a323a88),
	.w5(32'hbafb4551),
	.w6(32'h3a24ba14),
	.w7(32'hba5baf94),
	.w8(32'h3a9dae6d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2af616),
	.w1(32'h3a3be593),
	.w2(32'hbc0a813d),
	.w3(32'h38e75ebb),
	.w4(32'h3b3d02d8),
	.w5(32'hbc348f0a),
	.w6(32'h3b507a0c),
	.w7(32'hbc2ca2d0),
	.w8(32'hbb57378d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule