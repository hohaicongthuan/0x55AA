// This module converts an integer (0 - 255) of a colour value
// to a corresponding [0 - 1] single-precision floating-point scale

module Colour_Int_To_Float(data_i, data_o);
    input      [7:0] data_i;
    output reg [31:0] data_o;

    always @ (data_i) begin
        case (data_i)
        8'h00: data_o = 32'h00000000;
        8'h01: data_o = 32'h3b808081;
        8'h02: data_o = 32'h3c008081;
        8'h03: data_o = 32'h3c40c0c1;
        8'h04: data_o = 32'h3c808081;
        8'h05: data_o = 32'h3ca0a0a1;
        8'h06: data_o = 32'h3cc0c0c1;
        8'h07: data_o = 32'h3ce0e0e1;
        8'h08: data_o = 32'h3d008081;
        8'h09: data_o = 32'h3d109091;
        8'h0a: data_o = 32'h3d20a0a1;
        8'h0b: data_o = 32'h3d30b0b1;
        8'h0c: data_o = 32'h3d40c0c1;
        8'h0d: data_o = 32'h3d50d0d1;
        8'h0e: data_o = 32'h3d60e0e1;
        8'h0f: data_o = 32'h3d70f0f1;
        8'h10: data_o = 32'h3d808081;
        8'h11: data_o = 32'h3d888889;
        8'h12: data_o = 32'h3d909091;
        8'h13: data_o = 32'h3d989899;
        8'h14: data_o = 32'h3da0a0a1;
        8'h15: data_o = 32'h3da8a8a9;
        8'h16: data_o = 32'h3db0b0b1;
        8'h17: data_o = 32'h3db8b8b9;
        8'h18: data_o = 32'h3dc0c0c1;
        8'h19: data_o = 32'h3dc8c8c9;
        8'h1a: data_o = 32'h3dd0d0d1;
        8'h1b: data_o = 32'h3dd8d8d9;
        8'h1c: data_o = 32'h3de0e0e1;
        8'h1d: data_o = 32'h3de8e8e9;
        8'h1e: data_o = 32'h3df0f0f1;
        8'h1f: data_o = 32'h3df8f8f9;
        8'h20: data_o = 32'h3e008081;
        8'h21: data_o = 32'h3e048485;
        8'h22: data_o = 32'h3e088889;
        8'h23: data_o = 32'h3e0c8c8d;
        8'h24: data_o = 32'h3e109091;
        8'h25: data_o = 32'h3e149495;
        8'h26: data_o = 32'h3e189899;
        8'h27: data_o = 32'h3e1c9c9d;
        8'h28: data_o = 32'h3e20a0a1;
        8'h29: data_o = 32'h3e24a4a5;
        8'h2a: data_o = 32'h3e28a8a9;
        8'h2b: data_o = 32'h3e2cacad;
        8'h2c: data_o = 32'h3e30b0b1;
        8'h2d: data_o = 32'h3e34b4b5;
        8'h2e: data_o = 32'h3e38b8b9;
        8'h2f: data_o = 32'h3e3cbcbd;
        8'h30: data_o = 32'h3e40c0c1;
        8'h31: data_o = 32'h3e44c4c5;
        8'h32: data_o = 32'h3e48c8c9;
        8'h33: data_o = 32'h3e4ccccd;
        8'h34: data_o = 32'h3e50d0d1;
        8'h35: data_o = 32'h3e54d4d5;
        8'h36: data_o = 32'h3e58d8d9;
        8'h37: data_o = 32'h3e5cdcdd;
        8'h38: data_o = 32'h3e60e0e1;
        8'h39: data_o = 32'h3e64e4e5;
        8'h3a: data_o = 32'h3e68e8e9;
        8'h3b: data_o = 32'h3e6ceced;
        8'h3c: data_o = 32'h3e70f0f1;
        8'h3d: data_o = 32'h3e74f4f5;
        8'h3e: data_o = 32'h3e78f8f9;
        8'h3f: data_o = 32'h3e7cfcfd;
        8'h40: data_o = 32'h3e808081;
        8'h41: data_o = 32'h3e828283;
        8'h42: data_o = 32'h3e848485;
        8'h43: data_o = 32'h3e868687;
        8'h44: data_o = 32'h3e888889;
        8'h45: data_o = 32'h3e8a8a8b;
        8'h46: data_o = 32'h3e8c8c8d;
        8'h47: data_o = 32'h3e8e8e8f;
        8'h48: data_o = 32'h3e909091;
        8'h49: data_o = 32'h3e929293;
        8'h4a: data_o = 32'h3e949495;
        8'h4b: data_o = 32'h3e969697;
        8'h4c: data_o = 32'h3e989899;
        8'h4d: data_o = 32'h3e9a9a9b;
        8'h4e: data_o = 32'h3e9c9c9d;
        8'h4f: data_o = 32'h3e9e9e9f;
        8'h50: data_o = 32'h3ea0a0a1;
        8'h51: data_o = 32'h3ea2a2a3;
        8'h52: data_o = 32'h3ea4a4a5;
        8'h53: data_o = 32'h3ea6a6a7;
        8'h54: data_o = 32'h3ea8a8a9;
        8'h55: data_o = 32'h3eaaaaab;
        8'h56: data_o = 32'h3eacacad;
        8'h57: data_o = 32'h3eaeaeaf;
        8'h58: data_o = 32'h3eb0b0b1;
        8'h59: data_o = 32'h3eb2b2b3;
        8'h5a: data_o = 32'h3eb4b4b5;
        8'h5b: data_o = 32'h3eb6b6b7;
        8'h5c: data_o = 32'h3eb8b8b9;
        8'h5d: data_o = 32'h3ebababb;
        8'h5e: data_o = 32'h3ebcbcbd;
        8'h5f: data_o = 32'h3ebebebf;
        8'h60: data_o = 32'h3ec0c0c1;
        8'h61: data_o = 32'h3ec2c2c3;
        8'h62: data_o = 32'h3ec4c4c5;
        8'h63: data_o = 32'h3ec6c6c7;
        8'h64: data_o = 32'h3ec8c8c9;
        8'h65: data_o = 32'h3ecacacb;
        8'h66: data_o = 32'h3ecccccd;
        8'h67: data_o = 32'h3ecececf;
        8'h68: data_o = 32'h3ed0d0d1;
        8'h69: data_o = 32'h3ed2d2d3;
        8'h6a: data_o = 32'h3ed4d4d5;
        8'h6b: data_o = 32'h3ed6d6d7;
        8'h6c: data_o = 32'h3ed8d8d9;
        8'h6d: data_o = 32'h3edadadb;
        8'h6e: data_o = 32'h3edcdcdd;
        8'h6f: data_o = 32'h3edededf;
        8'h70: data_o = 32'h3ee0e0e1;
        8'h71: data_o = 32'h3ee2e2e3;
        8'h72: data_o = 32'h3ee4e4e5;
        8'h73: data_o = 32'h3ee6e6e7;
        8'h74: data_o = 32'h3ee8e8e9;
        8'h75: data_o = 32'h3eeaeaeb;
        8'h76: data_o = 32'h3eececed;
        8'h77: data_o = 32'h3eeeeeef;
        8'h78: data_o = 32'h3ef0f0f1;
        8'h79: data_o = 32'h3ef2f2f3;
        8'h7a: data_o = 32'h3ef4f4f5;
        8'h7b: data_o = 32'h3ef6f6f7;
        8'h7c: data_o = 32'h3ef8f8f9;
        8'h7d: data_o = 32'h3efafafb;
        8'h7e: data_o = 32'h3efcfcfd;
        8'h7f: data_o = 32'h3efefeff;
        8'h80: data_o = 32'h3f008081;
        8'h81: data_o = 32'h3f018182;
        8'h82: data_o = 32'h3f028283;
        8'h83: data_o = 32'h3f038384;
        8'h84: data_o = 32'h3f048485;
        8'h85: data_o = 32'h3f058586;
        8'h86: data_o = 32'h3f068687;
        8'h87: data_o = 32'h3f078788;
        8'h88: data_o = 32'h3f088889;
        8'h89: data_o = 32'h3f09898a;
        8'h8a: data_o = 32'h3f0a8a8b;
        8'h8b: data_o = 32'h3f0b8b8c;
        8'h8c: data_o = 32'h3f0c8c8d;
        8'h8d: data_o = 32'h3f0d8d8e;
        8'h8e: data_o = 32'h3f0e8e8f;
        8'h8f: data_o = 32'h3f0f8f90;
        8'h90: data_o = 32'h3f109091;
        8'h91: data_o = 32'h3f119192;
        8'h92: data_o = 32'h3f129293;
        8'h93: data_o = 32'h3f139394;
        8'h94: data_o = 32'h3f149495;
        8'h95: data_o = 32'h3f159596;
        8'h96: data_o = 32'h3f169697;
        8'h97: data_o = 32'h3f179798;
        8'h98: data_o = 32'h3f189899;
        8'h99: data_o = 32'h3f19999a;
        8'h9a: data_o = 32'h3f1a9a9b;
        8'h9b: data_o = 32'h3f1b9b9c;
        8'h9c: data_o = 32'h3f1c9c9d;
        8'h9d: data_o = 32'h3f1d9d9e;
        8'h9e: data_o = 32'h3f1e9e9f;
        8'h9f: data_o = 32'h3f1f9fa0;
        8'ha0: data_o = 32'h3f20a0a1;
        8'ha1: data_o = 32'h3f21a1a2;
        8'ha2: data_o = 32'h3f22a2a3;
        8'ha3: data_o = 32'h3f23a3a4;
        8'ha4: data_o = 32'h3f24a4a5;
        8'ha5: data_o = 32'h3f25a5a6;
        8'ha6: data_o = 32'h3f26a6a7;
        8'ha7: data_o = 32'h3f27a7a8;
        8'ha8: data_o = 32'h3f28a8a9;
        8'ha9: data_o = 32'h3f29a9aa;
        8'haa: data_o = 32'h3f2aaaab;
        8'hab: data_o = 32'h3f2babac;
        8'hac: data_o = 32'h3f2cacad;
        8'had: data_o = 32'h3f2dadae;
        8'hae: data_o = 32'h3f2eaeaf;
        8'haf: data_o = 32'h3f2fafb0;
        8'hb0: data_o = 32'h3f30b0b1;
        8'hb1: data_o = 32'h3f31b1b2;
        8'hb2: data_o = 32'h3f32b2b3;
        8'hb3: data_o = 32'h3f33b3b4;
        8'hb4: data_o = 32'h3f34b4b5;
        8'hb5: data_o = 32'h3f35b5b6;
        8'hb6: data_o = 32'h3f36b6b7;
        8'hb7: data_o = 32'h3f37b7b8;
        8'hb8: data_o = 32'h3f38b8b9;
        8'hb9: data_o = 32'h3f39b9ba;
        8'hba: data_o = 32'h3f3ababb;
        8'hbb: data_o = 32'h3f3bbbbc;
        8'hbc: data_o = 32'h3f3cbcbd;
        8'hbd: data_o = 32'h3f3dbdbe;
        8'hbe: data_o = 32'h3f3ebebf;
        8'hbf: data_o = 32'h3f3fbfc0;
        8'hc0: data_o = 32'h3f40c0c1;
        8'hc1: data_o = 32'h3f41c1c2;
        8'hc2: data_o = 32'h3f42c2c3;
        8'hc3: data_o = 32'h3f43c3c4;
        8'hc4: data_o = 32'h3f44c4c5;
        8'hc5: data_o = 32'h3f45c5c6;
        8'hc6: data_o = 32'h3f46c6c7;
        8'hc7: data_o = 32'h3f47c7c8;
        8'hc8: data_o = 32'h3f48c8c9;
        8'hc9: data_o = 32'h3f49c9ca;
        8'hca: data_o = 32'h3f4acacb;
        8'hcb: data_o = 32'h3f4bcbcc;
        8'hcc: data_o = 32'h3f4ccccd;
        8'hcd: data_o = 32'h3f4dcdce;
        8'hce: data_o = 32'h3f4ececf;
        8'hcf: data_o = 32'h3f4fcfd0;
        8'hd0: data_o = 32'h3f50d0d1;
        8'hd1: data_o = 32'h3f51d1d2;
        8'hd2: data_o = 32'h3f52d2d3;
        8'hd3: data_o = 32'h3f53d3d4;
        8'hd4: data_o = 32'h3f54d4d5;
        8'hd5: data_o = 32'h3f55d5d6;
        8'hd6: data_o = 32'h3f56d6d7;
        8'hd7: data_o = 32'h3f57d7d8;
        8'hd8: data_o = 32'h3f58d8d9;
        8'hd9: data_o = 32'h3f59d9da;
        8'hda: data_o = 32'h3f5adadb;
        8'hdb: data_o = 32'h3f5bdbdc;
        8'hdc: data_o = 32'h3f5cdcdd;
        8'hdd: data_o = 32'h3f5dddde;
        8'hde: data_o = 32'h3f5ededf;
        8'hdf: data_o = 32'h3f5fdfe0;
        8'he0: data_o = 32'h3f60e0e1;
        8'he1: data_o = 32'h3f61e1e2;
        8'he2: data_o = 32'h3f62e2e3;
        8'he3: data_o = 32'h3f63e3e4;
        8'he4: data_o = 32'h3f64e4e5;
        8'he5: data_o = 32'h3f65e5e6;
        8'he6: data_o = 32'h3f66e6e7;
        8'he7: data_o = 32'h3f67e7e8;
        8'he8: data_o = 32'h3f68e8e9;
        8'he9: data_o = 32'h3f69e9ea;
        8'hea: data_o = 32'h3f6aeaeb;
        8'heb: data_o = 32'h3f6bebec;
        8'hec: data_o = 32'h3f6ceced;
        8'hed: data_o = 32'h3f6dedee;
        8'hee: data_o = 32'h3f6eeeef;
        8'hef: data_o = 32'h3f6feff0;
        8'hf0: data_o = 32'h3f70f0f1;
        8'hf1: data_o = 32'h3f71f1f2;
        8'hf2: data_o = 32'h3f72f2f3;
        8'hf3: data_o = 32'h3f73f3f4;
        8'hf4: data_o = 32'h3f74f4f5;
        8'hf5: data_o = 32'h3f75f5f6;
        8'hf6: data_o = 32'h3f76f6f7;
        8'hf7: data_o = 32'h3f77f7f8;
        8'hf8: data_o = 32'h3f78f8f9;
        8'hf9: data_o = 32'h3f79f9fa;
        8'hfa: data_o = 32'h3f7afafb;
        8'hfb: data_o = 32'h3f7bfbfc;
        8'hfc: data_o = 32'h3f7cfcfd;
        8'hfd: data_o = 32'h3f7dfdfe;
        8'hfe: data_o = 32'h3f7efeff;
        8'hff: data_o = 32'h3F800000;
        default: data_o = 32'h00000000;
        endcase
    end
endmodule