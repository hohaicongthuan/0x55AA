module layer_10_featuremap_369(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba1843),
	.w1(32'h3a827d62),
	.w2(32'hbb335b03),
	.w3(32'hbbafc063),
	.w4(32'h3c86165b),
	.w5(32'hbb009541),
	.w6(32'h3c9c5c4c),
	.w7(32'hbc0e88dc),
	.w8(32'h3c0cece1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9561bf),
	.w1(32'h3b9ac94a),
	.w2(32'hbcb94c8e),
	.w3(32'h3b7939e2),
	.w4(32'hbbac5d98),
	.w5(32'h3c425637),
	.w6(32'h3b6e3454),
	.w7(32'h3acaddab),
	.w8(32'h3a35ff8e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393afdc1),
	.w1(32'hb978b7c5),
	.w2(32'hbbc46d60),
	.w3(32'h3c1b26da),
	.w4(32'h3b420d21),
	.w5(32'hbbaf4103),
	.w6(32'hbb55a22a),
	.w7(32'h3c0b4b83),
	.w8(32'hbbc1de45),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46a920),
	.w1(32'h3ba07ec3),
	.w2(32'h3c953037),
	.w3(32'hbb65b64a),
	.w4(32'h3c6f2d68),
	.w5(32'h3c29fd0f),
	.w6(32'hba66c2d9),
	.w7(32'hbb57891e),
	.w8(32'hbc09f5e2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20c0f4),
	.w1(32'hbb54efdd),
	.w2(32'h3aaf11e4),
	.w3(32'hbd3ebad2),
	.w4(32'h3b045dd8),
	.w5(32'h3bb0da8f),
	.w6(32'h3c33362f),
	.w7(32'h389d70ba),
	.w8(32'h3c0fe053),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29e43b),
	.w1(32'h3b19ec3c),
	.w2(32'h3a9e5afa),
	.w3(32'hbabfdb0f),
	.w4(32'hbb83ed11),
	.w5(32'h3c20bad0),
	.w6(32'h3b0e67d0),
	.w7(32'hbc346fab),
	.w8(32'h3c33a015),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ff23),
	.w1(32'h3be51ac2),
	.w2(32'h3a1de4f8),
	.w3(32'h3c6386df),
	.w4(32'h3d0002fc),
	.w5(32'hbdc4023a),
	.w6(32'hbb96a76e),
	.w7(32'h3b56aa61),
	.w8(32'hbb3e8afd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d03ca),
	.w1(32'h3c1ece8b),
	.w2(32'hbb2b2931),
	.w3(32'hbbd86136),
	.w4(32'h3b74d76f),
	.w5(32'h3c0428d1),
	.w6(32'h3ba4f108),
	.w7(32'hbbb65f3e),
	.w8(32'hbc22f69f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cec41be),
	.w1(32'hbdd4365f),
	.w2(32'hbc79d818),
	.w3(32'h3bbb552d),
	.w4(32'hbcae0a02),
	.w5(32'hbbda5ae4),
	.w6(32'h3c764987),
	.w7(32'hbba0e951),
	.w8(32'hba5f1944),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc970614),
	.w1(32'hbbe697fa),
	.w2(32'h3ae34f21),
	.w3(32'h39e1b44e),
	.w4(32'h3a6b9ccc),
	.w5(32'hbb29a90c),
	.w6(32'hbb37c598),
	.w7(32'h3d554671),
	.w8(32'h3bc3392a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6b695),
	.w1(32'hbb1da42c),
	.w2(32'h3a9bc56b),
	.w3(32'h3a79159e),
	.w4(32'hba712543),
	.w5(32'h3b9a923d),
	.w6(32'hbc916d76),
	.w7(32'h3b66798c),
	.w8(32'hbb8fb3cd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d18c5),
	.w1(32'hbac9a100),
	.w2(32'hbb6b243f),
	.w3(32'hbba83105),
	.w4(32'hbcc43479),
	.w5(32'h3a93eb12),
	.w6(32'hbb8f7978),
	.w7(32'h3a098110),
	.w8(32'hba059f81),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaff44),
	.w1(32'h3b8405f6),
	.w2(32'hbbcd13aa),
	.w3(32'hbc1bc633),
	.w4(32'h3aaf43e3),
	.w5(32'hb805ecb9),
	.w6(32'hbabf3f94),
	.w7(32'h3ba3e898),
	.w8(32'hbc92f2b0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdcf3b1c),
	.w1(32'h3b98f679),
	.w2(32'h3b62b3b6),
	.w3(32'h3c1555f5),
	.w4(32'h3d308df0),
	.w5(32'hbc5b0da2),
	.w6(32'hbc7f28e5),
	.w7(32'hbb4f3c65),
	.w8(32'hbc6485ec),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c008c02),
	.w1(32'hbbe914e1),
	.w2(32'h3afc5948),
	.w3(32'hbbb27a52),
	.w4(32'h3bbd01f5),
	.w5(32'h3b78820c),
	.w6(32'h3b22df40),
	.w7(32'hbb062be8),
	.w8(32'hbbfc00b3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1232a0),
	.w1(32'h3bed8abd),
	.w2(32'h3b5d7bc7),
	.w3(32'hbd498aff),
	.w4(32'h3b95832a),
	.w5(32'hba36eb5d),
	.w6(32'h3a5c1918),
	.w7(32'hbbddbc94),
	.w8(32'hbdc13308),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89d608),
	.w1(32'hbd724ed3),
	.w2(32'hbbf26a5e),
	.w3(32'hbc0947e2),
	.w4(32'h3a991a87),
	.w5(32'h3ca5fbbf),
	.w6(32'h3aa890e4),
	.w7(32'h3b16743f),
	.w8(32'h3bf5f0bb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b3f2f),
	.w1(32'h3d4da24d),
	.w2(32'h3cffd60f),
	.w3(32'hbbe9f1e7),
	.w4(32'hbcef15ca),
	.w5(32'hbbb6ca1d),
	.w6(32'h3b9a4868),
	.w7(32'hbd2332fe),
	.w8(32'hb9c4f45b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6113ed),
	.w1(32'hbcb00670),
	.w2(32'h3b671d3e),
	.w3(32'hbb44e7af),
	.w4(32'hbb4538d1),
	.w5(32'hbbf05c1b),
	.w6(32'hbb783b5b),
	.w7(32'hbc8aeb75),
	.w8(32'h3c3b2960),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe7280),
	.w1(32'h3c20f28b),
	.w2(32'h3c622b42),
	.w3(32'hbc240707),
	.w4(32'h3c12e5bf),
	.w5(32'hbb9b8606),
	.w6(32'hbac70bcb),
	.w7(32'h3c17daf7),
	.w8(32'hbbe0bd67),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8633c9),
	.w1(32'h3bc9bd46),
	.w2(32'hbbb4fa82),
	.w3(32'h3bc708b3),
	.w4(32'h3bac8e41),
	.w5(32'h3c531737),
	.w6(32'hbcc9345b),
	.w7(32'hbc18ba68),
	.w8(32'h3b9deb4c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2acfe1),
	.w1(32'hbc2028af),
	.w2(32'h3b96157b),
	.w3(32'h3b2bee78),
	.w4(32'hba5ae627),
	.w5(32'hbc374fb0),
	.w6(32'hbc7a26af),
	.w7(32'h3b7ca71a),
	.w8(32'hbab9e7b5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f60e8),
	.w1(32'h3b858b53),
	.w2(32'hbcb2a378),
	.w3(32'hb8859281),
	.w4(32'h3c6b0bf1),
	.w5(32'h3d34296e),
	.w6(32'h3b16e671),
	.w7(32'h3ab21794),
	.w8(32'h3b96df3f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20d1e3),
	.w1(32'hbbfc448b),
	.w2(32'hbc297eef),
	.w3(32'h3c168e20),
	.w4(32'hbc080bea),
	.w5(32'h3bb967f2),
	.w6(32'hbc00d929),
	.w7(32'h3bae775b),
	.w8(32'h3a15f321),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7ee35),
	.w1(32'hbb11d08e),
	.w2(32'h3bca08ae),
	.w3(32'hbb087535),
	.w4(32'hb9318dca),
	.w5(32'h3bb1dc9c),
	.w6(32'h3ae93168),
	.w7(32'hbb8397fb),
	.w8(32'h3bd0d236),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f272f),
	.w1(32'hbb3a6795),
	.w2(32'hbc2c3763),
	.w3(32'h3b5ef241),
	.w4(32'hbc193305),
	.w5(32'hb9d4f43d),
	.w6(32'hbb13de37),
	.w7(32'h3b5634f6),
	.w8(32'h3b9b6010),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a23d5),
	.w1(32'hbc1e4971),
	.w2(32'hbb5e11c1),
	.w3(32'h3b6f475c),
	.w4(32'h3bf90590),
	.w5(32'hb9cf1dcf),
	.w6(32'h3c38cbde),
	.w7(32'hbb626b96),
	.w8(32'h3c2da5ce),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38283d),
	.w1(32'hbbcdbe40),
	.w2(32'hbcf33249),
	.w3(32'h3a53d4b9),
	.w4(32'h3be8f52f),
	.w5(32'hbc814e91),
	.w6(32'h3bd595df),
	.w7(32'h3c42f0f4),
	.w8(32'h3c1c947b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a004c),
	.w1(32'h3bb272f8),
	.w2(32'hbca86e1b),
	.w3(32'hbbef998c),
	.w4(32'hbad95b5f),
	.w5(32'hbbd2d89f),
	.w6(32'h3cbec37b),
	.w7(32'hbb297e85),
	.w8(32'h3b12be1c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ff315),
	.w1(32'h3b4f39da),
	.w2(32'h3c3f13dc),
	.w3(32'h3c057cd0),
	.w4(32'h3c321a83),
	.w5(32'hbc02baab),
	.w6(32'h3c330f6e),
	.w7(32'hbbda8fe7),
	.w8(32'h3ba8b2e6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadabf1b),
	.w1(32'hbb684c4f),
	.w2(32'h3c17fb2d),
	.w3(32'hbbd121fd),
	.w4(32'h3ba01b03),
	.w5(32'hb8fdaf8b),
	.w6(32'hbbe3e059),
	.w7(32'hbc3916fa),
	.w8(32'h3c34b3f5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2af282),
	.w1(32'hbc37dab3),
	.w2(32'hbc0192ba),
	.w3(32'hbbd88e2c),
	.w4(32'h3b21d2a4),
	.w5(32'h3a850d0d),
	.w6(32'h3ab4cab2),
	.w7(32'hba98be31),
	.w8(32'hbc5468b5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cf9d8),
	.w1(32'h3c982b2c),
	.w2(32'h3c74f043),
	.w3(32'hbc1006b8),
	.w4(32'hbc55b131),
	.w5(32'hbc49fee9),
	.w6(32'hbcc2adf3),
	.w7(32'hbd25f946),
	.w8(32'hbb28d525),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affe5d7),
	.w1(32'hbcb8526c),
	.w2(32'h3aee4e65),
	.w3(32'hbc1e7265),
	.w4(32'hbc198d17),
	.w5(32'hbc4f9ba7),
	.w6(32'h387aca0d),
	.w7(32'h39f9603d),
	.w8(32'hbb307443),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c316b1a),
	.w1(32'hbbae2033),
	.w2(32'h3c646186),
	.w3(32'h39fd328e),
	.w4(32'hbbc06aea),
	.w5(32'h3b93c3fe),
	.w6(32'hbbbb3e75),
	.w7(32'h3b9cc98c),
	.w8(32'hbbe666be),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40df75),
	.w1(32'hba7b1bed),
	.w2(32'hbc20b03d),
	.w3(32'hbb027164),
	.w4(32'hb9c35a2e),
	.w5(32'h3b277473),
	.w6(32'h3af287b8),
	.w7(32'h3c545542),
	.w8(32'hbca977cb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb082adf),
	.w1(32'h3ad55f35),
	.w2(32'hbc21bc20),
	.w3(32'h3ba20c47),
	.w4(32'h3ab97565),
	.w5(32'h3c187b57),
	.w6(32'hba4e0d02),
	.w7(32'h3bbb251a),
	.w8(32'h3c110a94),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa603f7),
	.w1(32'hbace5fbd),
	.w2(32'hbcd05887),
	.w3(32'hbb2dc87d),
	.w4(32'h3c009444),
	.w5(32'h3aef6126),
	.w6(32'hbc1b9e33),
	.w7(32'h3c21ccc3),
	.w8(32'h3c456332),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a21b1f),
	.w1(32'hbab4b421),
	.w2(32'h3bbe4cf4),
	.w3(32'hbaf991c1),
	.w4(32'hbbb38122),
	.w5(32'hbc320778),
	.w6(32'hbc28abc8),
	.w7(32'h3c438f8b),
	.w8(32'hbc421774),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0503af),
	.w1(32'hbbac6305),
	.w2(32'h38e3b47b),
	.w3(32'h3915c103),
	.w4(32'h3afda398),
	.w5(32'h3c496399),
	.w6(32'h3c8e7dea),
	.w7(32'h3b665a95),
	.w8(32'hbbdf3165),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c6b6f4),
	.w1(32'hbbf30353),
	.w2(32'h3c625200),
	.w3(32'hbc1b7468),
	.w4(32'hbc058a3e),
	.w5(32'h3bd6e9c2),
	.w6(32'h3acd5dc5),
	.w7(32'hbb1d3bad),
	.w8(32'hbbde1a09),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48d799),
	.w1(32'hbbbec7b9),
	.w2(32'h3cdfae87),
	.w3(32'hbc1f1e88),
	.w4(32'h3b8c0ac2),
	.w5(32'hbc9a18ce),
	.w6(32'h3c85c1e7),
	.w7(32'h3b536caf),
	.w8(32'hbb1e1a88),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd3e3d),
	.w1(32'h39b6b468),
	.w2(32'h3c86cd82),
	.w3(32'h3b9c91cf),
	.w4(32'hbc71f280),
	.w5(32'h3c438360),
	.w6(32'hbc5a40ce),
	.w7(32'hbbcdd791),
	.w8(32'h3a0adb68),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09c573),
	.w1(32'h3b40cc77),
	.w2(32'h3c1d7da3),
	.w3(32'hbb241fb4),
	.w4(32'hbb3eb827),
	.w5(32'hbb325584),
	.w6(32'h3c2f196d),
	.w7(32'h3bf45f1e),
	.w8(32'h3a0cf734),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabfe3a),
	.w1(32'h3c8ef85d),
	.w2(32'h3c1313bb),
	.w3(32'h3c05e8cb),
	.w4(32'h3b9347b3),
	.w5(32'hbc457c42),
	.w6(32'h3cda6a68),
	.w7(32'h3c1a66f9),
	.w8(32'hba0e32de),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb697e59),
	.w1(32'hba892535),
	.w2(32'h3c968ba5),
	.w3(32'hb97b802d),
	.w4(32'h3b5af2df),
	.w5(32'h3c783c6a),
	.w6(32'hbbd74127),
	.w7(32'h3cbd6e55),
	.w8(32'hbc33d442),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb98018),
	.w1(32'hbb95e68d),
	.w2(32'hbc00fb7a),
	.w3(32'hb8174379),
	.w4(32'h3b9e7ece),
	.w5(32'h3acbf470),
	.w6(32'hbb7d1a65),
	.w7(32'hbc3b81e7),
	.w8(32'h3c7f29eb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b67dc),
	.w1(32'h3b16d0e0),
	.w2(32'h3baa6474),
	.w3(32'h3b8cc979),
	.w4(32'h3b9b37ff),
	.w5(32'h3a41f0d6),
	.w6(32'h3c5af5f7),
	.w7(32'h3c377063),
	.w8(32'h3cd534b6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5a5fc),
	.w1(32'hbb5c7f6b),
	.w2(32'h3bd8c77c),
	.w3(32'hbb462582),
	.w4(32'h3be0e3f4),
	.w5(32'h3b1531c6),
	.w6(32'h3c243ef2),
	.w7(32'hbaa733c6),
	.w8(32'h3c552a3f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad385b0),
	.w1(32'h3bc31cfd),
	.w2(32'hbd0bf925),
	.w3(32'h3c1f2c7a),
	.w4(32'hbc0ff8a7),
	.w5(32'h3b82f4f3),
	.w6(32'h3b11c880),
	.w7(32'hbb858ab9),
	.w8(32'h3a44a716),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf07d0),
	.w1(32'h3c90ad14),
	.w2(32'h3b74743f),
	.w3(32'h3b0dbae5),
	.w4(32'h3af1718f),
	.w5(32'h395f5db2),
	.w6(32'h3c0fb99d),
	.w7(32'h38a355fe),
	.w8(32'h3b18fc6e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba819a8),
	.w1(32'hbc91eeec),
	.w2(32'hbb7450cb),
	.w3(32'hbc5b76dd),
	.w4(32'hbcb6afa7),
	.w5(32'hb98afc14),
	.w6(32'hbc482133),
	.w7(32'hb99cc354),
	.w8(32'hbc724e16),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be95fac),
	.w1(32'h3c560d53),
	.w2(32'hbc5e1771),
	.w3(32'hbbdb88ce),
	.w4(32'hbaa5ecb8),
	.w5(32'hbc90f3ac),
	.w6(32'hbaab606a),
	.w7(32'h3b230f0e),
	.w8(32'hbcb4e902),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07fa3f),
	.w1(32'hbd1d41eb),
	.w2(32'hbaf9ff2a),
	.w3(32'h3bb5379d),
	.w4(32'h3c542138),
	.w5(32'h3a998756),
	.w6(32'hbb192183),
	.w7(32'h3a8d0340),
	.w8(32'h3baaf800),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab632c7),
	.w1(32'h3ac386e4),
	.w2(32'hbb39d7ed),
	.w3(32'hbc168034),
	.w4(32'h3a22d2c0),
	.w5(32'hbbb3a2d5),
	.w6(32'hbbb16497),
	.w7(32'hbc2e01f2),
	.w8(32'h393a667b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1245),
	.w1(32'hbba47721),
	.w2(32'h3c2d6d8e),
	.w3(32'h3b54fbe2),
	.w4(32'h3c37de74),
	.w5(32'h3bbe18cf),
	.w6(32'h3c1fda90),
	.w7(32'h3ae2bad2),
	.w8(32'hbb8142fd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cb482),
	.w1(32'hbbef8c49),
	.w2(32'h3c305697),
	.w3(32'h3cb10d00),
	.w4(32'h3c57a6a3),
	.w5(32'hbc0a40db),
	.w6(32'hbb9971e4),
	.w7(32'hbb9e624d),
	.w8(32'h3bb67eb0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaed3d9),
	.w1(32'h39db92fc),
	.w2(32'h39216810),
	.w3(32'hbc86f659),
	.w4(32'hbbe7bfb0),
	.w5(32'hbbeaaa69),
	.w6(32'hbbebc33f),
	.w7(32'hbbda0db3),
	.w8(32'h3b6b98da),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb51a6c),
	.w1(32'h3b2e9fa5),
	.w2(32'h3bc2f63e),
	.w3(32'h3a126d2d),
	.w4(32'hbb796157),
	.w5(32'hbc33eb17),
	.w6(32'hbb8ec985),
	.w7(32'hbc0f4454),
	.w8(32'h3b8dee75),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0214b),
	.w1(32'h3b90ebbc),
	.w2(32'hbb962230),
	.w3(32'h3ba252a2),
	.w4(32'h3c1131a6),
	.w5(32'h3b8351ce),
	.w6(32'h3be30555),
	.w7(32'h3a8a8b52),
	.w8(32'hbb0ca777),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6255d8),
	.w1(32'hbb511974),
	.w2(32'hb84c9330),
	.w3(32'h3b97f4d1),
	.w4(32'h3be93216),
	.w5(32'hbc2e5ce6),
	.w6(32'hbcad6dd2),
	.w7(32'h3c250d2a),
	.w8(32'hbb87bdd1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01ac4a),
	.w1(32'h3bd620d0),
	.w2(32'h388e7cf9),
	.w3(32'hbb59c74b),
	.w4(32'h3b543f55),
	.w5(32'h3b857ac3),
	.w6(32'hbc2fd3b5),
	.w7(32'h3b8eb373),
	.w8(32'h3ba745c7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41a4ba),
	.w1(32'hb9f10081),
	.w2(32'h3ca9c3c3),
	.w3(32'h3b5311a6),
	.w4(32'hbc39deb4),
	.w5(32'hbc3c88eb),
	.w6(32'h3c8cf847),
	.w7(32'hbc058108),
	.w8(32'h3b9ec2cd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc435142),
	.w1(32'h3cca2b67),
	.w2(32'hbc7c3152),
	.w3(32'hbb922e90),
	.w4(32'hbbc759a3),
	.w5(32'h3c1abb5d),
	.w6(32'hbc855d67),
	.w7(32'h3b2bf629),
	.w8(32'hbc380b75),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf373dd),
	.w1(32'h3ca9986d),
	.w2(32'hbb0c3900),
	.w3(32'hbb4661a7),
	.w4(32'hbc5eeeb2),
	.w5(32'h3c2a2fe4),
	.w6(32'hbc3a9e9c),
	.w7(32'h3c155479),
	.w8(32'h3b3844de),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a42f8),
	.w1(32'hb88ab8e8),
	.w2(32'hbc1c33ca),
	.w3(32'h3c996524),
	.w4(32'hbbe584d4),
	.w5(32'hbad8bc93),
	.w6(32'h3afef3f8),
	.w7(32'h3ceb1c23),
	.w8(32'hbb8ab4a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90ece9),
	.w1(32'h3aeb389f),
	.w2(32'h3bb4d9ce),
	.w3(32'h3c6429f0),
	.w4(32'hbbd57892),
	.w5(32'h3a0a14cf),
	.w6(32'hbb80584a),
	.w7(32'hbcd93319),
	.w8(32'h3aa6ddc9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28aa45),
	.w1(32'h3cb2697b),
	.w2(32'hbb553499),
	.w3(32'hbc57ba47),
	.w4(32'hbb56e554),
	.w5(32'h391967ec),
	.w6(32'hb9b3123a),
	.w7(32'h3c07097d),
	.w8(32'h3abdb83d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23b4c8),
	.w1(32'h3c42e405),
	.w2(32'h3ba87550),
	.w3(32'hbb38c6de),
	.w4(32'hb9f3395d),
	.w5(32'h3c890534),
	.w6(32'h3b9292a2),
	.w7(32'hba490047),
	.w8(32'h3ac70068),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38090f),
	.w1(32'h3c2200db),
	.w2(32'hbd0a0a94),
	.w3(32'hbb980785),
	.w4(32'hbc016f8f),
	.w5(32'hbbcafbd4),
	.w6(32'h3bd15024),
	.w7(32'hbb220dc0),
	.w8(32'h3b89f69c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0822df),
	.w1(32'h3bd7e96b),
	.w2(32'h39ed2cc8),
	.w3(32'h3aaebb6f),
	.w4(32'hbaf38cd6),
	.w5(32'h3b24cded),
	.w6(32'hbbbd1fde),
	.w7(32'h3c1b2f06),
	.w8(32'h3b0023e2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34da2f),
	.w1(32'hbc5deb4e),
	.w2(32'hbc3629be),
	.w3(32'hbc5f83ed),
	.w4(32'h3a9c2fe2),
	.w5(32'hb93d40fa),
	.w6(32'hba880ac1),
	.w7(32'h3c45038a),
	.w8(32'h3a530f8c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1ca6b),
	.w1(32'hbbb1cbd1),
	.w2(32'hbc0021cb),
	.w3(32'hbc7836ba),
	.w4(32'hbbaa7571),
	.w5(32'h3b37d285),
	.w6(32'h3b8253e0),
	.w7(32'h39e76563),
	.w8(32'hbb0be7db),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ec1e2),
	.w1(32'hba73cdfe),
	.w2(32'hba6e0537),
	.w3(32'h3ba9da37),
	.w4(32'hbb1334c0),
	.w5(32'hbac2dbf7),
	.w6(32'hbb431edd),
	.w7(32'h3b3fa31a),
	.w8(32'h3c209bd6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42adbb),
	.w1(32'h3cd2e075),
	.w2(32'h3a0ccfa7),
	.w3(32'hbc3c18e5),
	.w4(32'h3be6c9c6),
	.w5(32'h3b02b0d6),
	.w6(32'hbc7f5575),
	.w7(32'h3ca16aaa),
	.w8(32'hbbab7492),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9d8c0),
	.w1(32'hbca6ca87),
	.w2(32'hbbebe0a5),
	.w3(32'h3bd34591),
	.w4(32'h3c13583b),
	.w5(32'h3c28973e),
	.w6(32'hbc9a024d),
	.w7(32'h3cae1b10),
	.w8(32'hb9423d9b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9abc1),
	.w1(32'h3c0bfd66),
	.w2(32'hba33a9c9),
	.w3(32'hbbbcf049),
	.w4(32'hbb454691),
	.w5(32'hbc8d1a39),
	.w6(32'h3a585f22),
	.w7(32'hb99dfabb),
	.w8(32'hbbdc026b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba67c2a),
	.w1(32'h3b690bc9),
	.w2(32'h3be8a1dd),
	.w3(32'h3c8271ae),
	.w4(32'hbb905220),
	.w5(32'hba85868d),
	.w6(32'hbbc45a94),
	.w7(32'hbc2ffdb4),
	.w8(32'h3cbf5e52),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e72306),
	.w1(32'hbb07d446),
	.w2(32'hbb338cb1),
	.w3(32'hbc60024d),
	.w4(32'hbaba4bbf),
	.w5(32'h3a34a3cf),
	.w6(32'hbb2dc0ab),
	.w7(32'hbc2c7294),
	.w8(32'h3b571383),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7896b9),
	.w1(32'h3bd96e60),
	.w2(32'hbbc70df6),
	.w3(32'h399cc375),
	.w4(32'hbb340758),
	.w5(32'h3a24a823),
	.w6(32'hb9e5284e),
	.w7(32'hbc80fa5f),
	.w8(32'h3bf0e53e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb315f3b),
	.w1(32'hbb3615c8),
	.w2(32'h3c59985e),
	.w3(32'h3abeab5a),
	.w4(32'h3b1fb350),
	.w5(32'hbbfa5978),
	.w6(32'hbb7f6def),
	.w7(32'h3c0ef6ff),
	.w8(32'hbc6ceb7a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fe91c),
	.w1(32'h3c1f4fec),
	.w2(32'hbbc53d3b),
	.w3(32'h3ca17ef4),
	.w4(32'hb9c321dd),
	.w5(32'hbbaa269b),
	.w6(32'hbb9cfdad),
	.w7(32'h3b2a0c08),
	.w8(32'hbb400eb0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40cb38),
	.w1(32'hbc8bbc57),
	.w2(32'hb82eb39d),
	.w3(32'hb96ed8d4),
	.w4(32'h3b48b8f7),
	.w5(32'h3c522be4),
	.w6(32'h38d9af6f),
	.w7(32'hbc0c6244),
	.w8(32'hbb5c4fe5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27f346),
	.w1(32'h3b16de69),
	.w2(32'h3be1c92f),
	.w3(32'hbafd0e39),
	.w4(32'hbc02e25f),
	.w5(32'hbb9fd1a7),
	.w6(32'h3b32c5f8),
	.w7(32'hbbc7042a),
	.w8(32'hba871120),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fec34),
	.w1(32'hbb820f4b),
	.w2(32'hbcba83b9),
	.w3(32'h3bc2a1ae),
	.w4(32'h3a2845fb),
	.w5(32'hba06bbe8),
	.w6(32'h3b6cf3d7),
	.w7(32'hbbaf1265),
	.w8(32'h3a959130),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba154a83),
	.w1(32'hba0a0df0),
	.w2(32'hba9afaf9),
	.w3(32'h3c2f5a97),
	.w4(32'h3a5452c9),
	.w5(32'hba39835f),
	.w6(32'hbc5e4ed2),
	.w7(32'h3cdb758b),
	.w8(32'h3bb609ba),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb568cdf),
	.w1(32'h3c5fb55f),
	.w2(32'hbcd3a32f),
	.w3(32'h3b147362),
	.w4(32'hbc13c41b),
	.w5(32'hbb273bf6),
	.w6(32'h3b1eecf2),
	.w7(32'h3b927a1e),
	.w8(32'hbc2d80a4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e2e0b),
	.w1(32'h3cafd484),
	.w2(32'h3be5ba6b),
	.w3(32'hbc2a09ab),
	.w4(32'hbc075b84),
	.w5(32'h3c107f04),
	.w6(32'hbb3281d8),
	.w7(32'hbacc8c31),
	.w8(32'hbc4013c1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b052106),
	.w1(32'hbaca2440),
	.w2(32'hbc8e9a1a),
	.w3(32'hbb4a1f7e),
	.w4(32'hbbb0dfbc),
	.w5(32'hbca16573),
	.w6(32'hbc3ac75e),
	.w7(32'hbbd18fbc),
	.w8(32'hbbe478e5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27fe3f),
	.w1(32'hbc3656aa),
	.w2(32'h3be33452),
	.w3(32'hbc5359b7),
	.w4(32'hbb980411),
	.w5(32'hba2cb607),
	.w6(32'hbc59584d),
	.w7(32'h3c4872ac),
	.w8(32'h3a289953),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60a03e),
	.w1(32'hbbb631db),
	.w2(32'h3c2da65a),
	.w3(32'h37e7d6ff),
	.w4(32'h3c617419),
	.w5(32'hba4abdad),
	.w6(32'h3c3c5cad),
	.w7(32'h3a298886),
	.w8(32'hbba4ff0d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002984),
	.w1(32'hbc1dc67d),
	.w2(32'hbc2bb911),
	.w3(32'hbafa9d3c),
	.w4(32'h3b675563),
	.w5(32'hbcbf5fac),
	.w6(32'h3bace9dc),
	.w7(32'h3c6fe080),
	.w8(32'h3c1185cd),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b9652),
	.w1(32'hbb3614f1),
	.w2(32'hbb898538),
	.w3(32'hbc1b08df),
	.w4(32'h3c5e7336),
	.w5(32'hbae2c0c3),
	.w6(32'hbbf77fef),
	.w7(32'hbb94699f),
	.w8(32'hbc40fe39),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf682d6),
	.w1(32'hbcaf8987),
	.w2(32'hbc9b14c4),
	.w3(32'hbbc9763e),
	.w4(32'hbbe723d3),
	.w5(32'hbcc26e55),
	.w6(32'hbc12f5e6),
	.w7(32'hbba4d041),
	.w8(32'h3c622fc5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c72e2),
	.w1(32'hbb9496c8),
	.w2(32'hba13c212),
	.w3(32'hbb76153e),
	.w4(32'h3c87e7de),
	.w5(32'h3c2d5b21),
	.w6(32'hba94db33),
	.w7(32'hbccee102),
	.w8(32'hbbf3e041),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ced08),
	.w1(32'hbbb383a2),
	.w2(32'hbc985de7),
	.w3(32'hbb457837),
	.w4(32'h3b951e81),
	.w5(32'hbad03835),
	.w6(32'hbbaf6f4c),
	.w7(32'hbc1517e5),
	.w8(32'hbb446b04),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91baa5),
	.w1(32'h3b1630c7),
	.w2(32'h3bb0d4e7),
	.w3(32'hbb0847b4),
	.w4(32'hbb9b7226),
	.w5(32'hbc99916b),
	.w6(32'hbb7c19d7),
	.w7(32'hbbb24fb3),
	.w8(32'hb9d69aff),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820235),
	.w1(32'h3c1a2aa7),
	.w2(32'h3cc682c9),
	.w3(32'h3bdd488e),
	.w4(32'h3bfc5254),
	.w5(32'hbbb93594),
	.w6(32'hbc151631),
	.w7(32'h3c89c06b),
	.w8(32'hbc43c92e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc839cf7),
	.w1(32'hbc6ed7db),
	.w2(32'hbbbbac55),
	.w3(32'hbbd46db2),
	.w4(32'h3b29068f),
	.w5(32'h3cce3b7f),
	.w6(32'h3ad4eab9),
	.w7(32'h3b8c23ca),
	.w8(32'hbbdcf9b6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba833d6),
	.w1(32'h3baa836f),
	.w2(32'hbc07de42),
	.w3(32'hbc25fd45),
	.w4(32'h3b7f87f4),
	.w5(32'hbb835d5a),
	.w6(32'h3c078712),
	.w7(32'h3ca10614),
	.w8(32'h3b42734a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2512e3),
	.w1(32'hbb81ac10),
	.w2(32'hbb0077c2),
	.w3(32'hbaed4f40),
	.w4(32'h3c6dbf07),
	.w5(32'h3aa7d6d2),
	.w6(32'hb9153e68),
	.w7(32'h3cbd71cd),
	.w8(32'hbc3ac576),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbacd7a),
	.w1(32'h3ac34643),
	.w2(32'hbc6606c3),
	.w3(32'hba99d8aa),
	.w4(32'hbc0c4f59),
	.w5(32'h393e0edc),
	.w6(32'h3a47730a),
	.w7(32'h3bdec3d3),
	.w8(32'hbbb6e6c2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb323d),
	.w1(32'h3c6f07ed),
	.w2(32'hbcb6aa0b),
	.w3(32'hbbccf8d3),
	.w4(32'h3cc2c395),
	.w5(32'h3ace087c),
	.w6(32'h3b2d550d),
	.w7(32'h3c933e77),
	.w8(32'h3c8414e2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d1db4),
	.w1(32'h3be9753e),
	.w2(32'hba4d8a03),
	.w3(32'h3ac3ac85),
	.w4(32'hbbbea6dc),
	.w5(32'h3be6578f),
	.w6(32'hbc10818b),
	.w7(32'hba68856a),
	.w8(32'hbc86b70d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe5a26),
	.w1(32'hbb04f7d2),
	.w2(32'h3b881fc7),
	.w3(32'h3ab4dd23),
	.w4(32'h3c12b493),
	.w5(32'hbccc47b1),
	.w6(32'hba869c6a),
	.w7(32'h3bfd84aa),
	.w8(32'h3ac31ef3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40b092),
	.w1(32'h37b7c87d),
	.w2(32'h3bce60bb),
	.w3(32'h3c05eb81),
	.w4(32'h3b3b9dfd),
	.w5(32'h3b37b22f),
	.w6(32'h3b265bb3),
	.w7(32'hb7d5ea59),
	.w8(32'hbbc371af),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85538b),
	.w1(32'hbc5fc65b),
	.w2(32'hbc8ec1ca),
	.w3(32'h3c1d2fcf),
	.w4(32'hbb25fdc8),
	.w5(32'hb9bac571),
	.w6(32'h3c5bcd45),
	.w7(32'h3b8b100e),
	.w8(32'h3ad53f61),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bafd51),
	.w1(32'hb9815822),
	.w2(32'h39ea02c6),
	.w3(32'hbc2e3097),
	.w4(32'h3ac5b68e),
	.w5(32'h3ba7f927),
	.w6(32'h3bd4fac8),
	.w7(32'h3b5b082e),
	.w8(32'hbb55e002),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d69582b),
	.w1(32'hbb12d107),
	.w2(32'h3b567b79),
	.w3(32'h3b5f8d5a),
	.w4(32'hbc1872c9),
	.w5(32'hbba96549),
	.w6(32'hbb025bc6),
	.w7(32'hba187993),
	.w8(32'hbc167faf),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c00cd),
	.w1(32'h3b24c2f8),
	.w2(32'hbb13f95b),
	.w3(32'hbafa0895),
	.w4(32'h3bcdb4c3),
	.w5(32'h3bad2aed),
	.w6(32'h3ba34cda),
	.w7(32'hbac2d6a4),
	.w8(32'hbb7fb5af),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7df71),
	.w1(32'hbb614fcc),
	.w2(32'hbc07ad84),
	.w3(32'hbb3596e2),
	.w4(32'h3bbd3eb4),
	.w5(32'hbc961081),
	.w6(32'hbc9153c9),
	.w7(32'hbacd8b92),
	.w8(32'h3bf91b89),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83edc2),
	.w1(32'hbcc290b7),
	.w2(32'hbba44de1),
	.w3(32'hbb30dcd7),
	.w4(32'hbb41a005),
	.w5(32'hbaa0854f),
	.w6(32'hbbc783bc),
	.w7(32'hbc1b335b),
	.w8(32'hbc439212),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96f559),
	.w1(32'h3bb42d0a),
	.w2(32'hbc90883d),
	.w3(32'h3a91b902),
	.w4(32'h3c0e4642),
	.w5(32'h3aa99d70),
	.w6(32'h3c131ec3),
	.w7(32'h3c370c39),
	.w8(32'hbcf8fcc1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be39b1a),
	.w1(32'h3b7db1e0),
	.w2(32'h3b2d9108),
	.w3(32'h3c6cba20),
	.w4(32'h3b9a331a),
	.w5(32'hb98d3e71),
	.w6(32'h389b369d),
	.w7(32'h3c01c48c),
	.w8(32'hbbe44d0b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78cfe7),
	.w1(32'h3c07058d),
	.w2(32'h39b7e034),
	.w3(32'hbb24c0f7),
	.w4(32'h3a9a2069),
	.w5(32'h3d1b4bc6),
	.w6(32'hbaab14e9),
	.w7(32'hba156293),
	.w8(32'h3c46daef),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09c478),
	.w1(32'hbb45d888),
	.w2(32'hbb455a92),
	.w3(32'hbb742089),
	.w4(32'hbda60dcf),
	.w5(32'hba08def1),
	.w6(32'h3bd507fc),
	.w7(32'hbc15420b),
	.w8(32'hbc8951b0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca677aa),
	.w1(32'h3bdc2dce),
	.w2(32'hbc3361da),
	.w3(32'hbb628180),
	.w4(32'hbb83ce51),
	.w5(32'h3a923974),
	.w6(32'hbc074cba),
	.w7(32'h3aa92b2c),
	.w8(32'hbb1f4add),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46d757),
	.w1(32'hbbe154d6),
	.w2(32'hbbdde5e3),
	.w3(32'h3c43b0cf),
	.w4(32'hbb757cfc),
	.w5(32'hbbddf653),
	.w6(32'h3bc55b28),
	.w7(32'hbbc4e413),
	.w8(32'hbca74001),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d5e7f),
	.w1(32'h3b459255),
	.w2(32'h3c5945b1),
	.w3(32'hb9f9890d),
	.w4(32'h3b92a672),
	.w5(32'h3bf59885),
	.w6(32'h3c287a6c),
	.w7(32'h3b7b45f5),
	.w8(32'hbbae92de),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0b520),
	.w1(32'h3c87d323),
	.w2(32'h3b60e73f),
	.w3(32'hbcaff32c),
	.w4(32'h3ad11aaf),
	.w5(32'hbbee256a),
	.w6(32'h3a567d1a),
	.w7(32'hbbf21b2d),
	.w8(32'h3b943806),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b9bfc),
	.w1(32'hbc32ff14),
	.w2(32'hbc58ae6b),
	.w3(32'h3a66ba12),
	.w4(32'h39f4701d),
	.w5(32'hbc0b51cc),
	.w6(32'h3b8d1154),
	.w7(32'h3c527a9a),
	.w8(32'h3bba63cf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d346b),
	.w1(32'hb97a3468),
	.w2(32'hbc2f8ea9),
	.w3(32'hbb8360a3),
	.w4(32'h3b2aa3cd),
	.w5(32'h3bd53d9c),
	.w6(32'h3b81d08f),
	.w7(32'hbbbfe72e),
	.w8(32'h3b513860),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d0fe8),
	.w1(32'hbbde1373),
	.w2(32'h3b8de484),
	.w3(32'h3ac0c913),
	.w4(32'hbae31506),
	.w5(32'hbcac9acd),
	.w6(32'h3b38c42f),
	.w7(32'h39c7d51c),
	.w8(32'h3b8ef276),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13c107),
	.w1(32'hbb206e7e),
	.w2(32'h3bda639a),
	.w3(32'h3a9dd732),
	.w4(32'hba647bf6),
	.w5(32'h3ab1e4d5),
	.w6(32'hbc1720bd),
	.w7(32'h3bb9a82e),
	.w8(32'h3ba33a8f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab7bc7),
	.w1(32'h3b17726b),
	.w2(32'hbba5a14f),
	.w3(32'h3c0da9ba),
	.w4(32'hbaeab812),
	.w5(32'h3c08ee97),
	.w6(32'hba6df102),
	.w7(32'hbe0acab0),
	.w8(32'h3b9104c4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab535d0),
	.w1(32'h39fe1716),
	.w2(32'h3aafdc61),
	.w3(32'h3be7a7d7),
	.w4(32'hbca663ef),
	.w5(32'hbc1eb503),
	.w6(32'hbcf3619e),
	.w7(32'h39bf10df),
	.w8(32'h3b45a647),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89815),
	.w1(32'h3bf23c3b),
	.w2(32'h3c9fa363),
	.w3(32'hbadd1f39),
	.w4(32'h3b844b0f),
	.w5(32'hbcb6c85f),
	.w6(32'h3bbb54f3),
	.w7(32'hbb96178f),
	.w8(32'hbc851cb1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18767d),
	.w1(32'h3c18fd81),
	.w2(32'h3c575f46),
	.w3(32'hbc8b8f7c),
	.w4(32'h3b829554),
	.w5(32'hbd8c38e2),
	.w6(32'h3afd03cd),
	.w7(32'h3c3eb9c7),
	.w8(32'h3b88f4f2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a6cc9),
	.w1(32'hbc03b722),
	.w2(32'h3a858e04),
	.w3(32'h3b5b79e9),
	.w4(32'h3b4a18ed),
	.w5(32'h3bb8565c),
	.w6(32'hbc0bc634),
	.w7(32'h3c3c7179),
	.w8(32'hbc13fe94),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08381d),
	.w1(32'hbb264269),
	.w2(32'hbc966f70),
	.w3(32'h3557b332),
	.w4(32'h3c18bdbf),
	.w5(32'h3a5579e1),
	.w6(32'h3c169819),
	.w7(32'hbb922536),
	.w8(32'h3b2ca3b8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a517f81),
	.w1(32'h3bc793ee),
	.w2(32'h3b28f037),
	.w3(32'h3ba60a86),
	.w4(32'hbc8322d9),
	.w5(32'hbbd3b5c9),
	.w6(32'hb990b7e7),
	.w7(32'h3a74d46e),
	.w8(32'h3b8a453e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b394abf),
	.w1(32'hbcf8ab2f),
	.w2(32'hbbfca165),
	.w3(32'h39df73e0),
	.w4(32'hbb90ac2e),
	.w5(32'h3be9eaf4),
	.w6(32'hbb9fca38),
	.w7(32'hbb82c4dc),
	.w8(32'hbbd37e7a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1cb6a),
	.w1(32'h3bfd2fec),
	.w2(32'h3b340d10),
	.w3(32'h3c82df83),
	.w4(32'h3a528b3d),
	.w5(32'h3c69d698),
	.w6(32'hba386f9b),
	.w7(32'hbd0eca1c),
	.w8(32'h3b546da2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b660745),
	.w1(32'h3b7f8d8f),
	.w2(32'hbbde8bae),
	.w3(32'h3ac7e8ff),
	.w4(32'h3a62bdf1),
	.w5(32'h3b3cd294),
	.w6(32'h3bf93580),
	.w7(32'h3b7c49bf),
	.w8(32'hbbeac943),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e6568),
	.w1(32'h3a85e5de),
	.w2(32'hbc03f892),
	.w3(32'hbb465954),
	.w4(32'h3b80d00a),
	.w5(32'hbbe763c5),
	.w6(32'hbb928fcd),
	.w7(32'hbc41ca4a),
	.w8(32'hbbb1a319),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88babb),
	.w1(32'h3af4f587),
	.w2(32'h3c19d7bb),
	.w3(32'h3ba96e2f),
	.w4(32'h3b81e577),
	.w5(32'hb9d2ebdf),
	.w6(32'h3b5cdd22),
	.w7(32'h3b8f4528),
	.w8(32'h3b6b81a0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a299b98),
	.w1(32'h3beee7e0),
	.w2(32'hbca44cf2),
	.w3(32'h3999ba61),
	.w4(32'h3c0b409f),
	.w5(32'h3bcfcbb8),
	.w6(32'hbb729048),
	.w7(32'h3c509b23),
	.w8(32'hbc2288b9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26f422),
	.w1(32'hbc8ffe77),
	.w2(32'hbbb96e00),
	.w3(32'hb9e37054),
	.w4(32'hbbac74b1),
	.w5(32'h3a9dd4c4),
	.w6(32'h3bd06a2e),
	.w7(32'hba40d843),
	.w8(32'h38d175ee),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72ff1e),
	.w1(32'hba8dad7f),
	.w2(32'h3c24e90b),
	.w3(32'hbc05a77d),
	.w4(32'hb9cd5ce9),
	.w5(32'h3cac69a0),
	.w6(32'hbce09822),
	.w7(32'h3bb1f0d4),
	.w8(32'hb9b17f49),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05404e),
	.w1(32'h3b487f7d),
	.w2(32'hbbe1c1dc),
	.w3(32'hbbdac7fb),
	.w4(32'h3c96bf5c),
	.w5(32'hbad80456),
	.w6(32'h39a91e08),
	.w7(32'h3b1f9f9a),
	.w8(32'h39c93ccc),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2aca7),
	.w1(32'h3af42690),
	.w2(32'hbbe47a30),
	.w3(32'hbd2cbbec),
	.w4(32'hbc46b803),
	.w5(32'h3b508e5c),
	.w6(32'h3bac9dfa),
	.w7(32'h3bb09c82),
	.w8(32'hbc4070aa),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9a2cb),
	.w1(32'hbc93abec),
	.w2(32'hbb1c05f5),
	.w3(32'hbcca76ad),
	.w4(32'h3b7ca45f),
	.w5(32'hbbe7a179),
	.w6(32'hbb54f559),
	.w7(32'hbbf5eead),
	.w8(32'hbcb4112c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc373568),
	.w1(32'hbaae1c17),
	.w2(32'h3bf3de97),
	.w3(32'h3a9693ca),
	.w4(32'h3c2a2ecf),
	.w5(32'h3b8cd952),
	.w6(32'hbb015bd7),
	.w7(32'h3a0fee1b),
	.w8(32'h3bb6c3bc),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfeb54d),
	.w1(32'h3c0d3a17),
	.w2(32'h3b50635e),
	.w3(32'h3b625af2),
	.w4(32'hbb0051e8),
	.w5(32'hbbf11d50),
	.w6(32'hbbfaa5fd),
	.w7(32'h3b0cc68e),
	.w8(32'h3b7acb29),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909afd),
	.w1(32'hbba53f1d),
	.w2(32'h3c8665f8),
	.w3(32'h3a33bb59),
	.w4(32'hbd7a942f),
	.w5(32'h3c24ea39),
	.w6(32'hbb5b874a),
	.w7(32'h3a7e9d2d),
	.w8(32'h3a9f0339),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d467d),
	.w1(32'hbc0a51ff),
	.w2(32'h3becc6b7),
	.w3(32'hb9e3e416),
	.w4(32'hbc0a5b2e),
	.w5(32'hbbc713fc),
	.w6(32'h3be5eeb8),
	.w7(32'h3c388fed),
	.w8(32'h3aca68a3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c4aae),
	.w1(32'h3c61c5bd),
	.w2(32'hbc80324c),
	.w3(32'hbc09bc08),
	.w4(32'hbb8f99de),
	.w5(32'h3c3007bd),
	.w6(32'h3c099421),
	.w7(32'h3ba3e89d),
	.w8(32'hbbb5ae2e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b5b08),
	.w1(32'hbb0e497d),
	.w2(32'h3b624c29),
	.w3(32'hbc362c63),
	.w4(32'hbc7bf37a),
	.w5(32'hbc38fd93),
	.w6(32'hbc22e477),
	.w7(32'hbcce9efc),
	.w8(32'hbbb35f40),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07e576),
	.w1(32'hbb9cb20c),
	.w2(32'h3ba76b0b),
	.w3(32'h3aab3f8d),
	.w4(32'h3c570a04),
	.w5(32'hbc6bbab4),
	.w6(32'hbc14fbf1),
	.w7(32'hbbf4345f),
	.w8(32'h3c2f3de7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5755a),
	.w1(32'hbbfe4966),
	.w2(32'h3c2432bc),
	.w3(32'hbb9a8994),
	.w4(32'hbb4a75d3),
	.w5(32'hb99dfa1f),
	.w6(32'h3c6dd99e),
	.w7(32'hbb953a9c),
	.w8(32'h3a21aa83),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9d37f),
	.w1(32'h3af627ad),
	.w2(32'h3c75aeda),
	.w3(32'hba9b3410),
	.w4(32'h3b5d248c),
	.w5(32'hbbccb9b3),
	.w6(32'hbbb04000),
	.w7(32'h3cbe875b),
	.w8(32'hbbbd03fa),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6edb1e),
	.w1(32'h3ad06bec),
	.w2(32'h3b9f4807),
	.w3(32'h3ba3f9a3),
	.w4(32'h3b76f663),
	.w5(32'h3b7f35fc),
	.w6(32'h3d451b69),
	.w7(32'h3b8b8643),
	.w8(32'h3b563eba),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f8ac4),
	.w1(32'hbc6327e1),
	.w2(32'hbcd91f5f),
	.w3(32'h3b7b9134),
	.w4(32'h3cc47bd8),
	.w5(32'h3baed246),
	.w6(32'h3beb7384),
	.w7(32'hbc0be918),
	.w8(32'hb9ab4561),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13b6b2),
	.w1(32'hba5534bb),
	.w2(32'h3d1ccc96),
	.w3(32'hbbb927ca),
	.w4(32'hbb92925d),
	.w5(32'h3a98db09),
	.w6(32'h3b7dd7ce),
	.w7(32'hbbca1219),
	.w8(32'h3d2b9b6f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3af0c1),
	.w1(32'hbb0c6d77),
	.w2(32'h3a9ade06),
	.w3(32'h3c2451b2),
	.w4(32'hbb3c71c3),
	.w5(32'hbb7702a8),
	.w6(32'h3c101a49),
	.w7(32'hbbdcd3c7),
	.w8(32'h3bf54f2a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd2a7c),
	.w1(32'hbc4e048c),
	.w2(32'hbcefbdb8),
	.w3(32'h3c8a8f84),
	.w4(32'hbb9141de),
	.w5(32'hbaa3ab85),
	.w6(32'hbcfa613a),
	.w7(32'h3d16a775),
	.w8(32'h3bf3e9ab),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9029f96),
	.w1(32'hbb92e38d),
	.w2(32'h3b318d6f),
	.w3(32'hbc0375f2),
	.w4(32'hbae85c5d),
	.w5(32'hbc270254),
	.w6(32'hbd0e7d52),
	.w7(32'h3bdccb5b),
	.w8(32'h3a8e1189),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ac4f6),
	.w1(32'h3c78531e),
	.w2(32'h3bc75b17),
	.w3(32'h3b3248d1),
	.w4(32'h3b010dbd),
	.w5(32'h3ca0341a),
	.w6(32'hbc1231bd),
	.w7(32'h3abd307b),
	.w8(32'h3c7491f1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b314b7d),
	.w1(32'hb8549db9),
	.w2(32'h3a91d993),
	.w3(32'hbc1e956f),
	.w4(32'h3b0fb180),
	.w5(32'hba17acf6),
	.w6(32'h3b30aaa5),
	.w7(32'h3b24b732),
	.w8(32'hbba3282a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8adf71),
	.w1(32'hbc2c6a07),
	.w2(32'hbc5ec152),
	.w3(32'hb8b76743),
	.w4(32'h3c1093ab),
	.w5(32'h3ce960b2),
	.w6(32'hbb86e673),
	.w7(32'hbbb112f4),
	.w8(32'h3a3ad9fa),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9839511),
	.w1(32'h3c1257ba),
	.w2(32'h3b8e8593),
	.w3(32'h3ab26310),
	.w4(32'hbb1b47ab),
	.w5(32'hbbae856c),
	.w6(32'h3abb401e),
	.w7(32'h3bd305c1),
	.w8(32'hbbae140e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdec7e6),
	.w1(32'hbc39cd74),
	.w2(32'hbcb346c6),
	.w3(32'hba231e98),
	.w4(32'h3b28399f),
	.w5(32'h3c53d748),
	.w6(32'hbc97e802),
	.w7(32'h3be81e85),
	.w8(32'h3b3b7c13),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc317bc),
	.w1(32'h3bd34316),
	.w2(32'h3c32de47),
	.w3(32'hbc0a9f75),
	.w4(32'h3baa867b),
	.w5(32'hbc985abb),
	.w6(32'h3acf2001),
	.w7(32'h3bcc8174),
	.w8(32'hbc742a21),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9ead9),
	.w1(32'h3b5a66f2),
	.w2(32'hbb90e191),
	.w3(32'hbb2090fe),
	.w4(32'hbc254d4a),
	.w5(32'h3a5a15f1),
	.w6(32'h3c1903f8),
	.w7(32'hbbdb0764),
	.w8(32'hbac70abc),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d87a),
	.w1(32'h39dbb8f6),
	.w2(32'hbaf6a6f8),
	.w3(32'hbb19a298),
	.w4(32'hbb47c723),
	.w5(32'h3bc99e9c),
	.w6(32'hbb79a206),
	.w7(32'h399dcd2f),
	.w8(32'hbc0c6c04),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9340dc),
	.w1(32'h3ae1a6cc),
	.w2(32'h3c9f3982),
	.w3(32'hbcc822db),
	.w4(32'h3ac06a06),
	.w5(32'hbc947a38),
	.w6(32'h3bca73ee),
	.w7(32'hbb85463b),
	.w8(32'h3c87e7a0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb717583),
	.w1(32'h3b0d8f64),
	.w2(32'hbd076915),
	.w3(32'hbc13a6e9),
	.w4(32'h3b67aae8),
	.w5(32'hbc7e63d3),
	.w6(32'h3b9fbcd2),
	.w7(32'hbc2eb1bb),
	.w8(32'hbb7e6ce8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab991e0),
	.w1(32'h3bd9757c),
	.w2(32'h3c47d2a6),
	.w3(32'hbbfc7acf),
	.w4(32'hbbcf8f92),
	.w5(32'hbbea58cc),
	.w6(32'hbc9d61db),
	.w7(32'hba43a814),
	.w8(32'hbb3f2f6e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c7909),
	.w1(32'h3af30ab1),
	.w2(32'hbafc26b1),
	.w3(32'h3be90f5b),
	.w4(32'h3bad5339),
	.w5(32'h3a6353a7),
	.w6(32'h3a974f67),
	.w7(32'hbc4d0bc1),
	.w8(32'h3b0c6cb8),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3f13c),
	.w1(32'h3c75daa7),
	.w2(32'hba10a8f1),
	.w3(32'h3b2de1ed),
	.w4(32'hbb1fbe0f),
	.w5(32'h3b9f13e0),
	.w6(32'hbaf84ef4),
	.w7(32'hb8cae938),
	.w8(32'hbc819cbd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdbf03cf),
	.w1(32'hbbab3cf9),
	.w2(32'hbb6f9afb),
	.w3(32'hbb9d867c),
	.w4(32'hbaa55d2f),
	.w5(32'hbc2af911),
	.w6(32'hbbe69877),
	.w7(32'hbc747b04),
	.w8(32'h3ca6c53f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b96e09),
	.w1(32'hb79f495a),
	.w2(32'hbce53c5b),
	.w3(32'hbb656c41),
	.w4(32'h3bda1a95),
	.w5(32'hbb91cf23),
	.w6(32'hbaf061df),
	.w7(32'h3bb57df8),
	.w8(32'hbb837654),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0968af),
	.w1(32'hbcb48437),
	.w2(32'hbb0e9f83),
	.w3(32'h3b1f7242),
	.w4(32'h3c078fdb),
	.w5(32'hb8cfc31f),
	.w6(32'hbb9b01c3),
	.w7(32'h3b8ced21),
	.w8(32'h3c50ab34),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a313),
	.w1(32'hbac751ec),
	.w2(32'hbb519cc0),
	.w3(32'hbb9fd764),
	.w4(32'hbaf512aa),
	.w5(32'h3c1f2c66),
	.w6(32'h3ba6673b),
	.w7(32'hbb8f4247),
	.w8(32'hbafb2b88),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d1e66),
	.w1(32'h3c00189b),
	.w2(32'h3a46c0f2),
	.w3(32'hbc288e52),
	.w4(32'h3b4aaefc),
	.w5(32'hbc809838),
	.w6(32'h3bcd015f),
	.w7(32'h3b08ee4f),
	.w8(32'h3b538097),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaec56e),
	.w1(32'hba247c76),
	.w2(32'h3ad1c1d7),
	.w3(32'h3ad4255e),
	.w4(32'hb93c50e4),
	.w5(32'hbbf49f62),
	.w6(32'hbb031dd9),
	.w7(32'hbd0977d5),
	.w8(32'h3a8f61f5),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99254c),
	.w1(32'h3b9caa27),
	.w2(32'h3c65e99a),
	.w3(32'hbbf90c50),
	.w4(32'h3b0ab49c),
	.w5(32'hbccc8662),
	.w6(32'h3bbeda39),
	.w7(32'h3b46c3fe),
	.w8(32'h3ae2863d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6c499),
	.w1(32'h3c00c2c2),
	.w2(32'hbc093f46),
	.w3(32'hbbbd1bd5),
	.w4(32'hbba29fd5),
	.w5(32'h3a2f5309),
	.w6(32'hba9c6599),
	.w7(32'h3cb3ae91),
	.w8(32'hbba9b846),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba861ea),
	.w1(32'h3c7e937e),
	.w2(32'hbd810f43),
	.w3(32'h3ab04446),
	.w4(32'hbb831fcd),
	.w5(32'h3b7650e1),
	.w6(32'hbc19418c),
	.w7(32'hba3ecbf7),
	.w8(32'hbc4e44dd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafa756),
	.w1(32'hbcbdce58),
	.w2(32'h3c6659a3),
	.w3(32'hbbe08a87),
	.w4(32'hbbf33253),
	.w5(32'hb908ce49),
	.w6(32'h3afc014e),
	.w7(32'hbb8f971e),
	.w8(32'hbc9400e0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf966c),
	.w1(32'h3c220d85),
	.w2(32'hbb550bea),
	.w3(32'hbb26c2d8),
	.w4(32'h3b681db7),
	.w5(32'h3bf3afde),
	.w6(32'hbbfd758b),
	.w7(32'hbc7cc6dd),
	.w8(32'hbb94f723),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02b96a),
	.w1(32'h3abf906d),
	.w2(32'h3b83d9c1),
	.w3(32'hbc285f3e),
	.w4(32'h3c56a636),
	.w5(32'hbb247a89),
	.w6(32'hb950b3a5),
	.w7(32'h3c77f2df),
	.w8(32'hbb906415),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54fa42),
	.w1(32'h3c1bd201),
	.w2(32'hbae48e0c),
	.w3(32'h3c5e815f),
	.w4(32'h3ad0e671),
	.w5(32'hbbdd369b),
	.w6(32'hba5b2909),
	.w7(32'h3b2c0ffc),
	.w8(32'h3c6c67ae),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15a2d1),
	.w1(32'hbc107f3c),
	.w2(32'h3cf142d3),
	.w3(32'hbbdc283f),
	.w4(32'h3b0404f1),
	.w5(32'h39e7092e),
	.w6(32'hbb6526f0),
	.w7(32'hbbca3751),
	.w8(32'hbb933123),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba832a6b),
	.w1(32'h3ace070b),
	.w2(32'h3bcc36fe),
	.w3(32'hbc9ae6ce),
	.w4(32'hbcb09c07),
	.w5(32'h3b94b087),
	.w6(32'hbbc88315),
	.w7(32'hbb0a9d51),
	.w8(32'hbc11a852),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a9bfa),
	.w1(32'h3b5d8914),
	.w2(32'hbc1d4eb3),
	.w3(32'h3bc76892),
	.w4(32'h3c029851),
	.w5(32'h3cb0bf9a),
	.w6(32'h3b7d2c31),
	.w7(32'hbb2de823),
	.w8(32'h3b8beb61),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0557e8),
	.w1(32'h3acfae37),
	.w2(32'hbb22a6bb),
	.w3(32'h3aed60f8),
	.w4(32'h385d1a1b),
	.w5(32'h3ab95fde),
	.w6(32'hb9cd5a09),
	.w7(32'h3da15ae3),
	.w8(32'hbb8abee2),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8169e2),
	.w1(32'hbba6695b),
	.w2(32'h3c46c894),
	.w3(32'h3b541d0e),
	.w4(32'hbc95e9d6),
	.w5(32'h3b70f7c9),
	.w6(32'h3ad3eb3f),
	.w7(32'hbb5da6d2),
	.w8(32'h3b5c2800),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe00906c),
	.w1(32'h3c2405ff),
	.w2(32'h3bcfdd09),
	.w3(32'hbb811b92),
	.w4(32'hbb878caf),
	.w5(32'h3b8c0b92),
	.w6(32'hbcdcecab),
	.w7(32'hbad04d7f),
	.w8(32'hbc567a0b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc524ab5),
	.w1(32'h3b98ed77),
	.w2(32'hbc2ed566),
	.w3(32'hbb7aabee),
	.w4(32'h3c8f667d),
	.w5(32'hbb318e86),
	.w6(32'h3bf41ab8),
	.w7(32'hbb994307),
	.w8(32'h3c17bb78),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3fc34),
	.w1(32'h3bdbc012),
	.w2(32'h3b012b30),
	.w3(32'hbcc3cb89),
	.w4(32'h3b714e23),
	.w5(32'h3ba7bb11),
	.w6(32'h3aed7a21),
	.w7(32'hbc243c14),
	.w8(32'h3bf790ab),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90e260),
	.w1(32'hbbf25c5b),
	.w2(32'hbc4d3e90),
	.w3(32'hbacfb02f),
	.w4(32'hbbd829d1),
	.w5(32'hbc01776a),
	.w6(32'h3b835ca6),
	.w7(32'hbc20744e),
	.w8(32'hbd30ddf5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba651c2),
	.w1(32'hbb995dbe),
	.w2(32'hbbdd5f96),
	.w3(32'hb9cb5ef2),
	.w4(32'hbc0b14ec),
	.w5(32'hbbeb839e),
	.w6(32'h3bc178a4),
	.w7(32'h3bb68076),
	.w8(32'h3becf9fe),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a06acd),
	.w1(32'h3db62e07),
	.w2(32'hbc5f5f0d),
	.w3(32'h3b78b075),
	.w4(32'hbae32529),
	.w5(32'hbc10c953),
	.w6(32'hbc7c3c21),
	.w7(32'hbc519857),
	.w8(32'hbb179a68),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba8a72),
	.w1(32'hbc1859fd),
	.w2(32'hbc51e55f),
	.w3(32'hbc74db78),
	.w4(32'hbc04b755),
	.w5(32'h3b96bc4c),
	.w6(32'h3bc89529),
	.w7(32'hbb19d2ff),
	.w8(32'h3b36eb7b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf0ba5),
	.w1(32'hbb9b5856),
	.w2(32'hba0cdda4),
	.w3(32'hbcf16f02),
	.w4(32'hbb9bf042),
	.w5(32'h3b530718),
	.w6(32'hba3bba40),
	.w7(32'hbd59de0d),
	.w8(32'h3be5e74f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c7160),
	.w1(32'h3bd1bf84),
	.w2(32'hbc35d232),
	.w3(32'hbc401f15),
	.w4(32'hbbd0782c),
	.w5(32'hba004411),
	.w6(32'h3c1ad61f),
	.w7(32'hb95c2a74),
	.w8(32'h3bb407cd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4372b9),
	.w1(32'h3c8ce2e4),
	.w2(32'hbc8271ec),
	.w3(32'hbadff04d),
	.w4(32'h3aab5d92),
	.w5(32'hbbcb8f1d),
	.w6(32'hbac19a47),
	.w7(32'hbb780b1f),
	.w8(32'hb98a2358),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f9441),
	.w1(32'h3bd2db37),
	.w2(32'hbabf14b4),
	.w3(32'hbbc8f290),
	.w4(32'hbc1d1ab9),
	.w5(32'hbc080e40),
	.w6(32'h3a3f7deb),
	.w7(32'hbb9ced86),
	.w8(32'h39a54c63),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ba71a),
	.w1(32'hb8ffb095),
	.w2(32'h3a8fa8ef),
	.w3(32'h3afc6e12),
	.w4(32'h3bf87d85),
	.w5(32'hbbbc2957),
	.w6(32'hba76d87a),
	.w7(32'hbb3a5153),
	.w8(32'h3b984dad),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45dfba),
	.w1(32'hbb66467b),
	.w2(32'h3c94552c),
	.w3(32'hbb926f1d),
	.w4(32'hbc1f2272),
	.w5(32'hbc40b312),
	.w6(32'h3c21465f),
	.w7(32'h3c344aa1),
	.w8(32'h3bf4fd48),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f3f9c),
	.w1(32'h3a917233),
	.w2(32'hba70a3bd),
	.w3(32'h3b72d2e4),
	.w4(32'h3a8c2e31),
	.w5(32'h3cae8ff8),
	.w6(32'h3a75be7d),
	.w7(32'h3beb2bf0),
	.w8(32'h3b8e906d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98836a),
	.w1(32'hba31a9b5),
	.w2(32'hbbee9bd5),
	.w3(32'hbb0d0d7c),
	.w4(32'hbb10d664),
	.w5(32'hbc53fe99),
	.w6(32'hbb36b788),
	.w7(32'hbb6129fa),
	.w8(32'hbc2213ea),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd27551),
	.w1(32'h3a4af34f),
	.w2(32'h3c8359e1),
	.w3(32'h3b71ea7d),
	.w4(32'h3b67df50),
	.w5(32'h3ba6194c),
	.w6(32'hbc10e2ad),
	.w7(32'hbc00df26),
	.w8(32'h380457fa),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2388db),
	.w1(32'h3b470ee0),
	.w2(32'hbbe7f9f6),
	.w3(32'h3c121ba3),
	.w4(32'h3c220462),
	.w5(32'hb9e1a2ea),
	.w6(32'h3c073264),
	.w7(32'h3b84af14),
	.w8(32'h3cba0864),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac4bbf),
	.w1(32'hb8ed1f09),
	.w2(32'h3a6de6b2),
	.w3(32'hbc01ee15),
	.w4(32'hbb5e56f2),
	.w5(32'h3c9aef54),
	.w6(32'hbbdaaa7b),
	.w7(32'h3b3f5cb2),
	.w8(32'h3b8ea204),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74e518),
	.w1(32'hbc60e331),
	.w2(32'h3ab58f7c),
	.w3(32'h3b69fd59),
	.w4(32'h3c7372ff),
	.w5(32'hbbb0f559),
	.w6(32'hbc43a507),
	.w7(32'h3cc0ca49),
	.w8(32'hbb3be7c3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6c2a4),
	.w1(32'hbc683fda),
	.w2(32'h3bab761e),
	.w3(32'hbb56f515),
	.w4(32'hbc106f10),
	.w5(32'hbc2b54f5),
	.w6(32'h3be57fff),
	.w7(32'hbaf99899),
	.w8(32'h3c267071),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b958a1f),
	.w1(32'h3982a142),
	.w2(32'h3b4b1422),
	.w3(32'hbc649184),
	.w4(32'hbab63b28),
	.w5(32'hbc7c05c0),
	.w6(32'h3c139446),
	.w7(32'h3c806e9c),
	.w8(32'hbc1ab8f3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bc144),
	.w1(32'hbc9cb550),
	.w2(32'h3af978fc),
	.w3(32'hbbdcde7c),
	.w4(32'hbb0bba87),
	.w5(32'h3bc361c8),
	.w6(32'hbbcdb2ae),
	.w7(32'h3b04de63),
	.w8(32'hbb8809bd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac59845),
	.w1(32'h3bcdb5e8),
	.w2(32'h3813c3fc),
	.w3(32'hbb92bc14),
	.w4(32'hbbb8b01f),
	.w5(32'hbbe53630),
	.w6(32'h3c9fb49b),
	.w7(32'h3bd3fe78),
	.w8(32'h3b6ce0a7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80ad44),
	.w1(32'h3c3052b2),
	.w2(32'hbbd93a0d),
	.w3(32'h3ced9ba3),
	.w4(32'h3b93f777),
	.w5(32'h3c30e8ac),
	.w6(32'h3bebd8ea),
	.w7(32'hbbd4ffab),
	.w8(32'hbd0c13cf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920561),
	.w1(32'hbb87d2d4),
	.w2(32'h3c95de79),
	.w3(32'hba8a61fd),
	.w4(32'h3cdd22de),
	.w5(32'h3cb94df8),
	.w6(32'hbc24f404),
	.w7(32'h3cb9c4d9),
	.w8(32'h3a57ec56),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd913b7),
	.w1(32'h3bb3f388),
	.w2(32'h3ba7dfa4),
	.w3(32'hbb912f24),
	.w4(32'h3c791dd9),
	.w5(32'h3b899e66),
	.w6(32'hbc6a2869),
	.w7(32'h3bc90dcb),
	.w8(32'h3b55ecb2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92e0d7),
	.w1(32'h3ca73d49),
	.w2(32'h3b161bd2),
	.w3(32'hba91375f),
	.w4(32'h3a78565c),
	.w5(32'h3c15e87c),
	.w6(32'h3c8232d8),
	.w7(32'hbaf59104),
	.w8(32'hba816f4c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcde354),
	.w1(32'hbbde1b08),
	.w2(32'hbaeeedd9),
	.w3(32'h3af38e5b),
	.w4(32'hbb6dea2e),
	.w5(32'hbb996781),
	.w6(32'h3c957ee1),
	.w7(32'hb9e6f05f),
	.w8(32'h3ab78762),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7a8a2),
	.w1(32'h3b6f75f9),
	.w2(32'h39c4dd69),
	.w3(32'h3c8a2c66),
	.w4(32'hbc347207),
	.w5(32'hbbc6f12a),
	.w6(32'h3b26c422),
	.w7(32'hbc8a66dd),
	.w8(32'h3b7698d2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27163c),
	.w1(32'hbc2397c5),
	.w2(32'hbcd51a53),
	.w3(32'h3c6891a9),
	.w4(32'hbbb6bd26),
	.w5(32'hbc8f3511),
	.w6(32'h3c6f04e8),
	.w7(32'hbbb475de),
	.w8(32'hba0fb02b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb588eeb),
	.w1(32'hbc2d54a7),
	.w2(32'hbc3e488c),
	.w3(32'hbc3db991),
	.w4(32'hbc873ee9),
	.w5(32'hbc1fa64d),
	.w6(32'h3cbfca98),
	.w7(32'h3be380b5),
	.w8(32'h3b091882),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0bcb1),
	.w1(32'hbbcb52d9),
	.w2(32'hbbfecbcc),
	.w3(32'h3bcdee62),
	.w4(32'hbba09068),
	.w5(32'hbbdb0275),
	.w6(32'hbcd543ec),
	.w7(32'hbbbb0b00),
	.w8(32'h3c4a9cd9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98794a),
	.w1(32'hbb512955),
	.w2(32'hbb94c020),
	.w3(32'hbc055a42),
	.w4(32'hbc2011d8),
	.w5(32'hbb3da188),
	.w6(32'h3ac91ebd),
	.w7(32'h3b59ec89),
	.w8(32'h3ab7e6f4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dc374),
	.w1(32'h3b97b7d1),
	.w2(32'hbb6ab4b2),
	.w3(32'h3c0e2d65),
	.w4(32'h3aa2bfc0),
	.w5(32'hbba780fd),
	.w6(32'hbbb148dd),
	.w7(32'h3b01e040),
	.w8(32'h3d28d3cf),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a9f17),
	.w1(32'h3b3e9fb9),
	.w2(32'hbc8fc88f),
	.w3(32'hbb816d9e),
	.w4(32'h3b859559),
	.w5(32'h3c2ff9c7),
	.w6(32'h38d41eaf),
	.w7(32'hbc171dbe),
	.w8(32'hbb524776),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b83fe),
	.w1(32'h3c0384d8),
	.w2(32'h3aac95ee),
	.w3(32'hbc26570d),
	.w4(32'hbb3dc571),
	.w5(32'h3c2eded1),
	.w6(32'hbac96ef0),
	.w7(32'h3bba6b22),
	.w8(32'hbad76fa6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4da1e2),
	.w1(32'h395960ef),
	.w2(32'h3a83c981),
	.w3(32'hbc23d6be),
	.w4(32'h3be68f17),
	.w5(32'h3c372935),
	.w6(32'h399f4e9c),
	.w7(32'hbc4564e1),
	.w8(32'hbbb2a2d3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a22a),
	.w1(32'h3b706b2e),
	.w2(32'h3c59cd6b),
	.w3(32'h3c515420),
	.w4(32'hbbb4bea6),
	.w5(32'h3c6682d0),
	.w6(32'hbacd9a14),
	.w7(32'hbbbfc16c),
	.w8(32'hbaec64e0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab8896),
	.w1(32'hbb7b8786),
	.w2(32'h3a6a526a),
	.w3(32'hbb76d306),
	.w4(32'h3a86aee6),
	.w5(32'hbb8a45a3),
	.w6(32'h3b4b921a),
	.w7(32'h3b912319),
	.w8(32'hbbb763c7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e942),
	.w1(32'h3b226571),
	.w2(32'hbb5f6dd7),
	.w3(32'hbbf2f166),
	.w4(32'h3c581a4a),
	.w5(32'hb8f33d40),
	.w6(32'hbc59c7e9),
	.w7(32'hbc404055),
	.w8(32'h3c16c555),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbb26d),
	.w1(32'h3b2b364d),
	.w2(32'h3c0553de),
	.w3(32'hbc653f21),
	.w4(32'hbba36853),
	.w5(32'hbc8b496e),
	.w6(32'hbc334df1),
	.w7(32'h3c4bc98d),
	.w8(32'h3b205afd),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca8c6f),
	.w1(32'hbc48cc45),
	.w2(32'hbbd89d0d),
	.w3(32'h3b62290f),
	.w4(32'hbb8740c0),
	.w5(32'hbc81f32b),
	.w6(32'hbae5164b),
	.w7(32'h3c02974c),
	.w8(32'hbb9acecf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2c73),
	.w1(32'h3be18810),
	.w2(32'hbb0277fa),
	.w3(32'hbc8a0e37),
	.w4(32'h3c07046a),
	.w5(32'h3c48b41c),
	.w6(32'hbc2939f4),
	.w7(32'hbc1e4b3b),
	.w8(32'h3c68585f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc018340),
	.w1(32'hbc30cd41),
	.w2(32'h3be7b195),
	.w3(32'h3c8b11eb),
	.w4(32'hbbb53467),
	.w5(32'hbc524856),
	.w6(32'h3b1f634e),
	.w7(32'hbc33c29b),
	.w8(32'hbcaf0943),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc769a),
	.w1(32'h3b270a96),
	.w2(32'hbb88f997),
	.w3(32'hbca80f7a),
	.w4(32'h3c880465),
	.w5(32'hbb8107ce),
	.w6(32'hbb2bee2e),
	.w7(32'hbc649207),
	.w8(32'hbc468586),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb545146),
	.w1(32'h3c9b3f04),
	.w2(32'h3c8e9abc),
	.w3(32'hbcd5a70b),
	.w4(32'h3b7d3dcf),
	.w5(32'h3c6bbbfe),
	.w6(32'hb7f0234a),
	.w7(32'h3c1c9560),
	.w8(32'hba8c3c5b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500ca7),
	.w1(32'hbc5ed6bb),
	.w2(32'hbc75334d),
	.w3(32'h3c493616),
	.w4(32'hbc2e33e0),
	.w5(32'hbbb345d7),
	.w6(32'hbb109dce),
	.w7(32'hbbccfa69),
	.w8(32'h38708728),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918acd2),
	.w1(32'h3be86769),
	.w2(32'h38bca9ce),
	.w3(32'hbb2941a7),
	.w4(32'h3cedf4eb),
	.w5(32'h3a927871),
	.w6(32'hbb26629d),
	.w7(32'h3bacb57d),
	.w8(32'h3c437fbe),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14c11a),
	.w1(32'hbcd2b645),
	.w2(32'h3b198b28),
	.w3(32'hb9fca93f),
	.w4(32'hba77685f),
	.w5(32'hbc71d9aa),
	.w6(32'hbca65da9),
	.w7(32'hbc74f3a0),
	.w8(32'h3b269b54),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8511d),
	.w1(32'h3d1c2e92),
	.w2(32'h3aee258e),
	.w3(32'h3bd432db),
	.w4(32'hbbd77aeb),
	.w5(32'hbc05d7b1),
	.w6(32'h3b82953f),
	.w7(32'hbbe34826),
	.w8(32'hbb955f1d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d287e),
	.w1(32'h3c3c755f),
	.w2(32'hbb1a5fab),
	.w3(32'hbc3f8720),
	.w4(32'hbc3c60a2),
	.w5(32'hbb688ca8),
	.w6(32'hbbc3bb74),
	.w7(32'h3b889164),
	.w8(32'hbae87ae9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf41a5a),
	.w1(32'h3b222d06),
	.w2(32'h3bb5a227),
	.w3(32'h3912a827),
	.w4(32'h3bd06a55),
	.w5(32'hbaf9fb63),
	.w6(32'h3b87da8d),
	.w7(32'h3c8a0422),
	.w8(32'h3a937488),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d6f67e),
	.w1(32'h3bf85fcd),
	.w2(32'h3af4a0b5),
	.w3(32'hbc38aa08),
	.w4(32'hbb9e8409),
	.w5(32'hbc68e6a2),
	.w6(32'h393408b8),
	.w7(32'h3bb58fe3),
	.w8(32'hbc072f0b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c792b4b),
	.w1(32'h3c49b0cc),
	.w2(32'h3c87eee8),
	.w3(32'h3a821b0b),
	.w4(32'h3d1d1690),
	.w5(32'h3826c584),
	.w6(32'h3c9940a4),
	.w7(32'hbbc48d85),
	.w8(32'hbc300edc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba235b3),
	.w1(32'hbc0bcf9e),
	.w2(32'hba65a57e),
	.w3(32'h3bfa2290),
	.w4(32'h3b4742c7),
	.w5(32'hbc0a83da),
	.w6(32'hbc340a1e),
	.w7(32'h3c31153e),
	.w8(32'h3b16fb65),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21abd8),
	.w1(32'hbba9cc7b),
	.w2(32'hbab27284),
	.w3(32'hbc3697dc),
	.w4(32'h3badac4d),
	.w5(32'hbb031412),
	.w6(32'h3b1074ea),
	.w7(32'hbb44530f),
	.w8(32'h3ba9410f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb2d0e),
	.w1(32'h3bbe34da),
	.w2(32'h3aad4ff2),
	.w3(32'hbba02583),
	.w4(32'h3a04519b),
	.w5(32'hbc978666),
	.w6(32'h3b2d6691),
	.w7(32'h3bb1ac2c),
	.w8(32'h3ba20e6c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d4e64),
	.w1(32'h3bafae6a),
	.w2(32'h3b25e0c3),
	.w3(32'hba9c7337),
	.w4(32'h3a86f99f),
	.w5(32'hbb9643ba),
	.w6(32'hbc6027ec),
	.w7(32'hbba8ad70),
	.w8(32'h3ac7fb8a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d32e0),
	.w1(32'hbcb06569),
	.w2(32'hbb93153d),
	.w3(32'hbc8d7fd6),
	.w4(32'hbbf0f02d),
	.w5(32'hbc2bb30d),
	.w6(32'h3cdef5c4),
	.w7(32'hbb86b7c3),
	.w8(32'hbc3ce409),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04369f),
	.w1(32'hbb6dc7cd),
	.w2(32'h3c4a9f84),
	.w3(32'hbb2921ef),
	.w4(32'h3a8a14c0),
	.w5(32'hbb9c8423),
	.w6(32'hbba340cf),
	.w7(32'hbc273913),
	.w8(32'h3b46f512),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c939c38),
	.w1(32'hbada202d),
	.w2(32'h3aaccf36),
	.w3(32'hba4ae003),
	.w4(32'hba05be2a),
	.w5(32'hbc0978e9),
	.w6(32'hbc8db2f1),
	.w7(32'hbb434854),
	.w8(32'h3b5ef2ee),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba456300),
	.w1(32'hbbcf4078),
	.w2(32'hbbfca4b5),
	.w3(32'h3aaa6b5b),
	.w4(32'hbafa6ce0),
	.w5(32'h3935051c),
	.w6(32'hbbe5b7c0),
	.w7(32'h3b28cb99),
	.w8(32'hba87a77c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47dfe1),
	.w1(32'h3b8f6336),
	.w2(32'h3b5f47e4),
	.w3(32'hbc8116f9),
	.w4(32'h3aaa3b2d),
	.w5(32'h3be9201e),
	.w6(32'hbbfb084b),
	.w7(32'hba1ee499),
	.w8(32'hbcaf905b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8eac3a),
	.w1(32'hbb7f15d9),
	.w2(32'h3c1a4086),
	.w3(32'hbc9c13c3),
	.w4(32'h3b108a2f),
	.w5(32'hbbfe1f87),
	.w6(32'hbbbb81e2),
	.w7(32'h3a72c765),
	.w8(32'h3d18e74c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0a2e2),
	.w1(32'h3c0f5981),
	.w2(32'h3b4b89cb),
	.w3(32'hba8fe1b1),
	.w4(32'hbb6ff566),
	.w5(32'h3b478136),
	.w6(32'hbb694e08),
	.w7(32'hbbdffe26),
	.w8(32'h3bc1be57),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46a66e),
	.w1(32'h3bde68cf),
	.w2(32'hbc7e2620),
	.w3(32'hbc2c47b6),
	.w4(32'h39dce618),
	.w5(32'h3b5671ec),
	.w6(32'h3c42b6cb),
	.w7(32'hbbadd404),
	.w8(32'hbbc51d0b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1544f5),
	.w1(32'h3bdbee9a),
	.w2(32'hbbc2f5af),
	.w3(32'h3c64d7d9),
	.w4(32'hbb8dac09),
	.w5(32'h382ccc72),
	.w6(32'h3c0cfcd9),
	.w7(32'h39808f9d),
	.w8(32'hbc045bc4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b572e),
	.w1(32'hbbe27602),
	.w2(32'hbaf9f15f),
	.w3(32'hbbbf0b78),
	.w4(32'hbac4f9ca),
	.w5(32'h3ad6ae97),
	.w6(32'h3cd05272),
	.w7(32'h3aa5247b),
	.w8(32'hbb92518e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule