module layer_10_featuremap_18(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb40e5),
	.w1(32'h3c036861),
	.w2(32'h3aef5a3e),
	.w3(32'h3c7f6556),
	.w4(32'h3c5935c0),
	.w5(32'hbbbcdadf),
	.w6(32'h3c80455d),
	.w7(32'h3c6918fa),
	.w8(32'h3be88769),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c9d49),
	.w1(32'hbbae34ad),
	.w2(32'h3c3fee7c),
	.w3(32'hbb908e3f),
	.w4(32'hbb385067),
	.w5(32'h3c29d3e1),
	.w6(32'hba5922f4),
	.w7(32'hbb968f39),
	.w8(32'h3c4212dc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c542fb2),
	.w1(32'h3bf42396),
	.w2(32'h3ae1716f),
	.w3(32'h3c79bc2d),
	.w4(32'h3beac7ab),
	.w5(32'hbb34b5d9),
	.w6(32'h3c2a736c),
	.w7(32'h374ba169),
	.w8(32'hbc042a61),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba48e32),
	.w1(32'h3b8bae1d),
	.w2(32'h3bf533ae),
	.w3(32'hbb155932),
	.w4(32'hbb92720b),
	.w5(32'hbb986e34),
	.w6(32'hbbf56b00),
	.w7(32'h3b0634cd),
	.w8(32'hbbcfa5b2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89cde1),
	.w1(32'h3aeb2ff4),
	.w2(32'hbbb42ef7),
	.w3(32'hbc8e15d3),
	.w4(32'hbb99fe4f),
	.w5(32'hbb8c3633),
	.w6(32'hbbf9aecc),
	.w7(32'h3c4865b1),
	.w8(32'h398ada1b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fb497),
	.w1(32'h3b9e6998),
	.w2(32'h3b75224a),
	.w3(32'hbac8b762),
	.w4(32'h3bacf230),
	.w5(32'hb93b3593),
	.w6(32'h3a98d0a1),
	.w7(32'h3bde1768),
	.w8(32'h398eb424),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d547f),
	.w1(32'h3bf0dbd3),
	.w2(32'hbc382f90),
	.w3(32'hbc47ebb3),
	.w4(32'hba5d26fb),
	.w5(32'hbc8679cf),
	.w6(32'hbc2e15a4),
	.w7(32'h39f96435),
	.w8(32'h3b48adbd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc555b6),
	.w1(32'hbc1df26b),
	.w2(32'hbbc45a6e),
	.w3(32'hbca3a02e),
	.w4(32'hbc5b0940),
	.w5(32'hbc4efb57),
	.w6(32'hbc0eb6f1),
	.w7(32'hbb03ac18),
	.w8(32'h3aba4702),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72f42e),
	.w1(32'h3bda7a0c),
	.w2(32'h3c976170),
	.w3(32'hba3f92e3),
	.w4(32'h3c0b234c),
	.w5(32'h3cbc489e),
	.w6(32'h3c1ddc2e),
	.w7(32'h3c82b50d),
	.w8(32'h3c1186c1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b69b9),
	.w1(32'h3c5d2f6e),
	.w2(32'h3be3b31f),
	.w3(32'h3cc87fb9),
	.w4(32'h3c7f255b),
	.w5(32'h3bf47b5d),
	.w6(32'h3c135700),
	.w7(32'h3be06844),
	.w8(32'h3bbd01b8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcf71a),
	.w1(32'h3be2b99c),
	.w2(32'h3b15b4ff),
	.w3(32'h3bfcf133),
	.w4(32'h3b0d777b),
	.w5(32'hbb5a6e5a),
	.w6(32'h3b083cf2),
	.w7(32'hbb64e6f6),
	.w8(32'h3ad4a4b3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd154ae),
	.w1(32'hbb7cfd44),
	.w2(32'hbc0e81fa),
	.w3(32'h3b1271b9),
	.w4(32'h3bda7225),
	.w5(32'hbc0be10f),
	.w6(32'h3b3ec5ca),
	.w7(32'h3c1d35c5),
	.w8(32'hbbe3c650),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc229ff4),
	.w1(32'hbc0840db),
	.w2(32'h3aa33906),
	.w3(32'hbc3fd5e1),
	.w4(32'hbc252ad9),
	.w5(32'h3bdb2db0),
	.w6(32'hbc52f644),
	.w7(32'hbc24c848),
	.w8(32'h3b426419),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eaedb),
	.w1(32'hb9e8fdcc),
	.w2(32'h3b3911a9),
	.w3(32'hbba47170),
	.w4(32'hbbe01748),
	.w5(32'hbb6dfce5),
	.w6(32'hbbd27594),
	.w7(32'hbb4961cb),
	.w8(32'h3b522707),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc33439),
	.w1(32'h3cab29ef),
	.w2(32'hbbb1b3f4),
	.w3(32'h3c4c0274),
	.w4(32'h3c7c39d5),
	.w5(32'hbc0386cf),
	.w6(32'h3bd88c1e),
	.w7(32'hb8597983),
	.w8(32'h3a720994),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20d9e1),
	.w1(32'h3a9de0b0),
	.w2(32'h3bc82885),
	.w3(32'hbc23d505),
	.w4(32'hbc198f2b),
	.w5(32'h3bd97d1d),
	.w6(32'h3ac84cb6),
	.w7(32'hbace5b8e),
	.w8(32'h3b31acd2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf150be),
	.w1(32'h3b80df88),
	.w2(32'hbc21554d),
	.w3(32'h3bb594b3),
	.w4(32'hba166b53),
	.w5(32'hbc0650b5),
	.w6(32'hbb165e67),
	.w7(32'hbbc6b03f),
	.w8(32'hbc26c042),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc243053),
	.w1(32'hbc80f842),
	.w2(32'hbb45a924),
	.w3(32'hbc2ff887),
	.w4(32'h3b607c26),
	.w5(32'hbba6c569),
	.w6(32'h3c4d2d9c),
	.w7(32'h3d1fa2bf),
	.w8(32'hbb6f3c67),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca680),
	.w1(32'hba17757e),
	.w2(32'h3c58caff),
	.w3(32'hbb95dd1b),
	.w4(32'hbbdf16d0),
	.w5(32'h3c967451),
	.w6(32'h3a5254e3),
	.w7(32'hbbb298fe),
	.w8(32'h3bf02c24),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96a1c8),
	.w1(32'h3c561aed),
	.w2(32'hbbf64344),
	.w3(32'h3c9c86d6),
	.w4(32'h3c93ad7a),
	.w5(32'hbb474c21),
	.w6(32'h3c7dff65),
	.w7(32'h3c7bf46b),
	.w8(32'h3bd26cb1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadee5de),
	.w1(32'h3b8a7fb3),
	.w2(32'h3b1fe83a),
	.w3(32'h3c3ddbfd),
	.w4(32'h3c60ca7b),
	.w5(32'hbaa473d8),
	.w6(32'h3c7a9790),
	.w7(32'h3c73b400),
	.w8(32'h3a858f8e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9499c6),
	.w1(32'h3b8a25c7),
	.w2(32'h39291d95),
	.w3(32'hbb4503d1),
	.w4(32'h3a1c3be8),
	.w5(32'h3abf114f),
	.w6(32'h3b93d07b),
	.w7(32'h3c0bb177),
	.w8(32'h3c26b83d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93f7b5),
	.w1(32'h3c11a9c8),
	.w2(32'hbc46b942),
	.w3(32'h3c5366bb),
	.w4(32'h3c919753),
	.w5(32'hbc0eadfe),
	.w6(32'h3c92445e),
	.w7(32'h3cebf3cd),
	.w8(32'h3bb02560),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc655a2),
	.w1(32'h3bab57ff),
	.w2(32'h39ed38f7),
	.w3(32'h3b8a7ad6),
	.w4(32'h3c61710a),
	.w5(32'h3ab0c603),
	.w6(32'h3c3fecf4),
	.w7(32'h3c8e6b05),
	.w8(32'hb9dd81d2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dc4e2),
	.w1(32'h3ae99ec8),
	.w2(32'hbb982f34),
	.w3(32'hbbc07c31),
	.w4(32'hbb02ca9b),
	.w5(32'hbb3b6543),
	.w6(32'hbb84e9bc),
	.w7(32'hbc01eb6c),
	.w8(32'hba34470e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26224a),
	.w1(32'h3a70bb71),
	.w2(32'h3be70f5b),
	.w3(32'h3bb008da),
	.w4(32'h3b8a5dd8),
	.w5(32'h3b5d5103),
	.w6(32'h3c375c25),
	.w7(32'h3c7796d7),
	.w8(32'h3b61406f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b615753),
	.w1(32'h3b8e4dda),
	.w2(32'hbac9046f),
	.w3(32'h3a8d04ef),
	.w4(32'hbb0e569d),
	.w5(32'hbada5743),
	.w6(32'h3af71ca5),
	.w7(32'h3be1a7c2),
	.w8(32'hb88f8e0a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b8e43),
	.w1(32'hba72d6a5),
	.w2(32'h3bcade41),
	.w3(32'hb99d78cd),
	.w4(32'hbafc520d),
	.w5(32'hbbe5e026),
	.w6(32'h3aadd1d3),
	.w7(32'hbac245ed),
	.w8(32'hbb9e6bac),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ba396),
	.w1(32'h3b4eea95),
	.w2(32'hbb9d6635),
	.w3(32'hbc10fe7d),
	.w4(32'hbb887dd0),
	.w5(32'hbb1acf7d),
	.w6(32'hba43a52e),
	.w7(32'h3bd9dd22),
	.w8(32'hbb8422a1),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c3dfe),
	.w1(32'hbbf42cc3),
	.w2(32'h3cdc0f9f),
	.w3(32'hbc13a087),
	.w4(32'h3983c3b1),
	.w5(32'h3b995d79),
	.w6(32'hbc220c6e),
	.w7(32'hbbe13802),
	.w8(32'hbd089a72),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7f5cde),
	.w1(32'h3d19c1b6),
	.w2(32'hbbff10c7),
	.w3(32'h3b8bd163),
	.w4(32'h3ad04764),
	.w5(32'hbc198219),
	.w6(32'hbd81947e),
	.w7(32'hbd398fd2),
	.w8(32'hbb9e359c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57b866),
	.w1(32'hbc84ca16),
	.w2(32'hbc069a38),
	.w3(32'hbb2f1a97),
	.w4(32'hbbe238b4),
	.w5(32'hbbda02ce),
	.w6(32'h3b248946),
	.w7(32'hbb96dbb5),
	.w8(32'h3b9e9697),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306378),
	.w1(32'hbbd007d9),
	.w2(32'h3cc38ea0),
	.w3(32'hbc24bc63),
	.w4(32'hbbdd143b),
	.w5(32'h3c1057e9),
	.w6(32'h3a829e97),
	.w7(32'h3b9b04b7),
	.w8(32'hbce9a1ae),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7112a9),
	.w1(32'h3ce0a852),
	.w2(32'hbb245c1a),
	.w3(32'h3bbea7cd),
	.w4(32'hba9d87c9),
	.w5(32'h3be88f87),
	.w6(32'hbd7b18e6),
	.w7(32'hbd2e08bc),
	.w8(32'h3b96ccb6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bff95),
	.w1(32'h3b32c8f5),
	.w2(32'hbc8023eb),
	.w3(32'h3bd94dc2),
	.w4(32'hbbe9290c),
	.w5(32'hbb837cf1),
	.w6(32'hb7da493d),
	.w7(32'hbb0841f9),
	.w8(32'h3c406168),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd13686e),
	.w1(32'hbc997c52),
	.w2(32'hba234c4b),
	.w3(32'hbc30a9c1),
	.w4(32'hbbd6715c),
	.w5(32'hbbe16185),
	.w6(32'h3cd06dbb),
	.w7(32'h3c86f607),
	.w8(32'h3b2ca789),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf70caf),
	.w1(32'h3c0a910c),
	.w2(32'h3cc22a8d),
	.w3(32'hbbd4e66f),
	.w4(32'h3b408e01),
	.w5(32'h3b869e6b),
	.w6(32'h3ba0d0f6),
	.w7(32'hbb6ec06a),
	.w8(32'hbce8a1cb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d439a68),
	.w1(32'h3cf125c9),
	.w2(32'h3bf90d42),
	.w3(32'hbb83f6f4),
	.w4(32'hbbec21ce),
	.w5(32'h3bc311b1),
	.w6(32'hbd744232),
	.w7(32'hbd2ca293),
	.w8(32'hbc0634d3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c103771),
	.w1(32'h3c3a837a),
	.w2(32'h3be3cd8b),
	.w3(32'h3b12bed8),
	.w4(32'h3c2af224),
	.w5(32'hbb0a4ece),
	.w6(32'hbc57c145),
	.w7(32'hbc0653ec),
	.w8(32'h3b20c67f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c549fcc),
	.w1(32'h3bb43605),
	.w2(32'hbbdba546),
	.w3(32'h3b8fef1e),
	.w4(32'h3b83a7c8),
	.w5(32'hbbd525fd),
	.w6(32'hbb993db2),
	.w7(32'h3c0f669b),
	.w8(32'hbb603cc4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5cc23),
	.w1(32'hbb875dd4),
	.w2(32'h3b9d6803),
	.w3(32'hbc72a4a4),
	.w4(32'hbbe0a384),
	.w5(32'hbc09d644),
	.w6(32'hbbac6c85),
	.w7(32'hbbf34abd),
	.w8(32'hbbbe82e6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef745a),
	.w1(32'hbb2b47f7),
	.w2(32'h39aa13c5),
	.w3(32'hbc95a2f6),
	.w4(32'hbc127bd8),
	.w5(32'hbaff1579),
	.w6(32'hbc3302f5),
	.w7(32'hbc868a1c),
	.w8(32'hbc2e8093),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c8ff6),
	.w1(32'hba406d20),
	.w2(32'hbcdce9f1),
	.w3(32'hbb5e6245),
	.w4(32'h3b102050),
	.w5(32'hbc4b6d16),
	.w6(32'hb99e783b),
	.w7(32'hb9db2915),
	.w8(32'h3cb225b1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6719e9),
	.w1(32'hbd016ba9),
	.w2(32'h3c4f3900),
	.w3(32'hbc23b4b1),
	.w4(32'hbc1c42f0),
	.w5(32'h3afd0308),
	.w6(32'h3d49d541),
	.w7(32'h3cdbf13f),
	.w8(32'hba5933b0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b2315),
	.w1(32'h3b7c550c),
	.w2(32'h3bf34994),
	.w3(32'hbb86b9f1),
	.w4(32'hbb8c3de4),
	.w5(32'h3c272a75),
	.w6(32'hbc4ac3ed),
	.w7(32'hbadf6c2f),
	.w8(32'h3bc9b570),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b8315),
	.w1(32'h3b78a297),
	.w2(32'h39adf2f1),
	.w3(32'h3bf6f500),
	.w4(32'h3b8042b2),
	.w5(32'hbc47167f),
	.w6(32'hba8b1494),
	.w7(32'h3bdf38c9),
	.w8(32'hbafac8cf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58b6eb),
	.w1(32'hbb441959),
	.w2(32'h3c019027),
	.w3(32'hbba1b51b),
	.w4(32'hbbb9d792),
	.w5(32'h3a84af36),
	.w6(32'hbbb490ef),
	.w7(32'h3b729f84),
	.w8(32'h3b57a280),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52fbcc),
	.w1(32'h3b9fb326),
	.w2(32'hbcf1aaf3),
	.w3(32'hbb73ef2f),
	.w4(32'h39ea4e4c),
	.w5(32'hbc465a69),
	.w6(32'hbc642b8c),
	.w7(32'hbb869908),
	.w8(32'h3ccbf80e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8ac207),
	.w1(32'hbd279536),
	.w2(32'h3c8ac8de),
	.w3(32'hbc2da015),
	.w4(32'hbbf17d8f),
	.w5(32'h3caac7a5),
	.w6(32'h3d6c4583),
	.w7(32'h3d1c865a),
	.w8(32'h3b9cf75f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd9167),
	.w1(32'h3c54444f),
	.w2(32'h3a5e37f8),
	.w3(32'h3d0be299),
	.w4(32'h3c9412b6),
	.w5(32'h3be759c2),
	.w6(32'h3c40c452),
	.w7(32'h3c80a1e6),
	.w8(32'h3c020b11),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaee8d1),
	.w1(32'h3b128a70),
	.w2(32'h3b052642),
	.w3(32'hba97fc62),
	.w4(32'hbba0db5f),
	.w5(32'hbac1ca4b),
	.w6(32'h3c00a0b7),
	.w7(32'hba3384fd),
	.w8(32'h3bd777c7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb460896),
	.w1(32'h3b18a1d0),
	.w2(32'h3b9fb705),
	.w3(32'hbb81eb5d),
	.w4(32'hbb3a1593),
	.w5(32'h3c1c66d0),
	.w6(32'hbb2e4451),
	.w7(32'hbb1d9d3d),
	.w8(32'h3c044f5f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09972c),
	.w1(32'hbb7094ea),
	.w2(32'h3aa842e4),
	.w3(32'hbb90957b),
	.w4(32'hbb848b9a),
	.w5(32'hbbe35a42),
	.w6(32'hbacb4843),
	.w7(32'hbba69c75),
	.w8(32'h3b12938f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb398209),
	.w1(32'h3a661f75),
	.w2(32'hbb1160d8),
	.w3(32'hbc208ffb),
	.w4(32'hbbe55a54),
	.w5(32'hbab00a77),
	.w6(32'h3bf97acb),
	.w7(32'h3b2ab082),
	.w8(32'h3bbcf5de),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e6a7),
	.w1(32'h3af99fab),
	.w2(32'hbc0de3d6),
	.w3(32'h3c86b5be),
	.w4(32'h3ca75412),
	.w5(32'hbbb6aa89),
	.w6(32'h3c9abc64),
	.w7(32'h3ca5bbee),
	.w8(32'hbb95aa51),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72d406),
	.w1(32'hbb25e5c2),
	.w2(32'h3b111ce3),
	.w3(32'hbbf33789),
	.w4(32'hbb6dcdca),
	.w5(32'h3ba0df37),
	.w6(32'hbc30e059),
	.w7(32'hbbce0ac3),
	.w8(32'h39bbc2fa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00ee32),
	.w1(32'hbbe38519),
	.w2(32'h3c79947d),
	.w3(32'h3b8cf4f1),
	.w4(32'hbbee6056),
	.w5(32'h3bebce46),
	.w6(32'h3c070d64),
	.w7(32'hbbc216ad),
	.w8(32'hba8f0550),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62ae0f),
	.w1(32'h3c110310),
	.w2(32'hbac61386),
	.w3(32'hba1bdf2a),
	.w4(32'hbbba8eb0),
	.w5(32'hbba6fa34),
	.w6(32'hbc313021),
	.w7(32'hbc4046b4),
	.w8(32'h3c151cd1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04c6fb),
	.w1(32'hbb859fd3),
	.w2(32'h3baa7401),
	.w3(32'hbb1b54ba),
	.w4(32'hbbb4115d),
	.w5(32'hba80fba9),
	.w6(32'h3be9e207),
	.w7(32'h3b32abae),
	.w8(32'hbb675601),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade579a),
	.w1(32'hbb2e8c55),
	.w2(32'h3cc388b8),
	.w3(32'hbc4ecc11),
	.w4(32'hbb812d64),
	.w5(32'h3b879645),
	.w6(32'hbc1fedb2),
	.w7(32'hbbf65ab8),
	.w8(32'hbbe149ec),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0300f2),
	.w1(32'h3cbc7961),
	.w2(32'h3b9ecf24),
	.w3(32'h3c58569c),
	.w4(32'h3c410870),
	.w5(32'hbb9cd235),
	.w6(32'h3b305dfe),
	.w7(32'hba137e7c),
	.w8(32'hbbdd24a8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c266d52),
	.w1(32'h3c0a195b),
	.w2(32'h3b0f12a6),
	.w3(32'h3aab4096),
	.w4(32'h3c040a7e),
	.w5(32'h3b19beaf),
	.w6(32'hbc3e75de),
	.w7(32'h3a5402e3),
	.w8(32'h3b924339),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8ccf0),
	.w1(32'hbb99c2e1),
	.w2(32'hba5ad0c7),
	.w3(32'hbb776680),
	.w4(32'hbb10803f),
	.w5(32'hbc1fdfa8),
	.w6(32'h3a9e9e97),
	.w7(32'hbb8e2605),
	.w8(32'h3b1e0e47),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d0b53),
	.w1(32'h3982c9d2),
	.w2(32'h3b18277f),
	.w3(32'hbc39fb60),
	.w4(32'hbc1371e8),
	.w5(32'hbc2979a6),
	.w6(32'hba00789b),
	.w7(32'hba6d6c29),
	.w8(32'h3a485ecc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8765f),
	.w1(32'hbb3260af),
	.w2(32'h3b41af6e),
	.w3(32'hbb9f851d),
	.w4(32'hbc0f08ca),
	.w5(32'h3b1def4a),
	.w6(32'hbb109875),
	.w7(32'h3b2e05ab),
	.w8(32'h3a5b2de6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b3b3e),
	.w1(32'h3ba112f8),
	.w2(32'h3bacc0e8),
	.w3(32'h3b306a10),
	.w4(32'h3b20bf68),
	.w5(32'h3b32c2a7),
	.w6(32'h3a5e1b0a),
	.w7(32'hbae5ac8d),
	.w8(32'h3b59077f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc4031),
	.w1(32'h3c100e85),
	.w2(32'hbb4d8d99),
	.w3(32'h3b52b79d),
	.w4(32'hba105483),
	.w5(32'h3a05f853),
	.w6(32'hba8a8f7c),
	.w7(32'hbb9cc553),
	.w8(32'h3b9a6bd0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c10b5),
	.w1(32'h3ad7fa9a),
	.w2(32'h3b5fbdb1),
	.w3(32'h3b90c9bc),
	.w4(32'hbb61fda2),
	.w5(32'h3a89a643),
	.w6(32'h3baf74e3),
	.w7(32'h3b6e9a4d),
	.w8(32'hbb15282a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b757c43),
	.w1(32'hbadda01f),
	.w2(32'hbb236e35),
	.w3(32'hbbe832de),
	.w4(32'hbbedbda7),
	.w5(32'h39621a11),
	.w6(32'hbbac3abc),
	.w7(32'hbb984ff3),
	.w8(32'hb9ce3e9a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d5ac),
	.w1(32'hbb1d8ce4),
	.w2(32'h3bb6ad67),
	.w3(32'hbb211ea3),
	.w4(32'h3a591d56),
	.w5(32'hbbd6ab83),
	.w6(32'hbb84f4e5),
	.w7(32'h3b09154c),
	.w8(32'hbbef4be4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53b1e0),
	.w1(32'h3bcff638),
	.w2(32'h3b85aa36),
	.w3(32'hbb49c4da),
	.w4(32'h3c15c559),
	.w5(32'h3b8b6bfe),
	.w6(32'hbc42d207),
	.w7(32'h3b521f94),
	.w8(32'h3bbc6bd1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41c90a),
	.w1(32'h3b3a80b6),
	.w2(32'h3b1df18f),
	.w3(32'h3c05aac0),
	.w4(32'h3ab519ff),
	.w5(32'h3b3ac42e),
	.w6(32'h3c04dffd),
	.w7(32'h3af45d92),
	.w8(32'h3b9d6ace),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aec82),
	.w1(32'h3ba2e2bb),
	.w2(32'h3b4ccd2c),
	.w3(32'hba03bfd7),
	.w4(32'h3b0653ed),
	.w5(32'hbb3ec2a5),
	.w6(32'hb6759b68),
	.w7(32'h3c3a9bc4),
	.w8(32'hbc25b3ff),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beff1ca),
	.w1(32'h3c6015db),
	.w2(32'hbc943b58),
	.w3(32'hbb81ad89),
	.w4(32'h3af3c87f),
	.w5(32'hbc4c9d72),
	.w6(32'hbc4b1fa9),
	.w7(32'hbbf0d4e5),
	.w8(32'h3c38a973),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2c9a2a),
	.w1(32'hbcc454da),
	.w2(32'h3c12e715),
	.w3(32'hbc12ddcb),
	.w4(32'hbbefca89),
	.w5(32'h3badd0d5),
	.w6(32'h3d076e9f),
	.w7(32'h3c9ed566),
	.w8(32'h3b0a02e4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10d637),
	.w1(32'h3b37da3f),
	.w2(32'h3b890e5b),
	.w3(32'h3b36cc25),
	.w4(32'h3b0ef3b6),
	.w5(32'hba39057d),
	.w6(32'h3aac153b),
	.w7(32'h3a1e459f),
	.w8(32'h3b3929ed),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4550ac),
	.w1(32'h3a578736),
	.w2(32'h3b63802c),
	.w3(32'hbba5c9b7),
	.w4(32'hbc065945),
	.w5(32'hbade4eb3),
	.w6(32'hbb30799e),
	.w7(32'hbb5ca55c),
	.w8(32'h3b6a692e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64ecf8),
	.w1(32'h3b4a705a),
	.w2(32'hbb99adbe),
	.w3(32'h3b7e4835),
	.w4(32'hbb42e554),
	.w5(32'hbaf298a1),
	.w6(32'h3b1808d2),
	.w7(32'hbb5e852b),
	.w8(32'hbb6bddc6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae60f93),
	.w1(32'hbc0df1d7),
	.w2(32'hba9dfad6),
	.w3(32'h3b7e31e2),
	.w4(32'h356a4070),
	.w5(32'h39ddadff),
	.w6(32'h3ba82161),
	.w7(32'h3c319d3a),
	.w8(32'h3a010c91),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbacfbe),
	.w1(32'hba45efd0),
	.w2(32'h3ba331cd),
	.w3(32'hbb937f03),
	.w4(32'h3ae5a3f8),
	.w5(32'h3b5186fd),
	.w6(32'hbb7e1d37),
	.w7(32'hb8f0d9cc),
	.w8(32'h3bff1265),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b709dd7),
	.w1(32'h3b56e7e5),
	.w2(32'h3c3dfca4),
	.w3(32'h3a558226),
	.w4(32'h3baf4145),
	.w5(32'h3a7cec78),
	.w6(32'h39c29b0a),
	.w7(32'h3a6e0695),
	.w8(32'hbc7643ed),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07da15),
	.w1(32'h3c679a54),
	.w2(32'h3bcdcc45),
	.w3(32'h3ac2da78),
	.w4(32'hbb493fdb),
	.w5(32'h3b345bd4),
	.w6(32'hbd036135),
	.w7(32'hbcbc2457),
	.w8(32'h3bac64e7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1347b2),
	.w1(32'h3c38db5d),
	.w2(32'h3b9bdaa1),
	.w3(32'hbafe1df6),
	.w4(32'h3c3c9d89),
	.w5(32'hbc038af1),
	.w6(32'hbbb8ade0),
	.w7(32'h3c0649df),
	.w8(32'hbc1963d9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87df92),
	.w1(32'h3c2a5a3e),
	.w2(32'h3bd3f97d),
	.w3(32'hb95f81d0),
	.w4(32'h3c5b6415),
	.w5(32'h3b4551dc),
	.w6(32'hbbdbcf0e),
	.w7(32'h3c21b6a2),
	.w8(32'h3bce276c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5757ea),
	.w1(32'hbbabd79f),
	.w2(32'h3b3385f6),
	.w3(32'hbbd762dc),
	.w4(32'h3bb32a46),
	.w5(32'h3bd3ab03),
	.w6(32'h3b77a44a),
	.w7(32'h3b92f672),
	.w8(32'h3916d765),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0abc00),
	.w1(32'h3a3e2766),
	.w2(32'hb82b37a6),
	.w3(32'hbb06a5ba),
	.w4(32'h384dcd3d),
	.w5(32'h3aba4bd1),
	.w6(32'hbb02033e),
	.w7(32'hbb014b80),
	.w8(32'h3b94de2a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b162e),
	.w1(32'h3a82c636),
	.w2(32'h3b647400),
	.w3(32'hb9e0b1cc),
	.w4(32'hbb386b89),
	.w5(32'h3b3e2bb7),
	.w6(32'h3afd048f),
	.w7(32'hba9d4a59),
	.w8(32'h38fdd8e9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a320ac4),
	.w1(32'h3a85fd86),
	.w2(32'hbb7ea7c5),
	.w3(32'hba2d07ba),
	.w4(32'h3aa8aa7a),
	.w5(32'hba014c12),
	.w6(32'h3b2d050c),
	.w7(32'h3bc2304f),
	.w8(32'hbbc31e11),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29ee8c),
	.w1(32'hbbb8d95a),
	.w2(32'h3bf78bd9),
	.w3(32'hbc3d9de9),
	.w4(32'hbc0a57b2),
	.w5(32'h3bddde33),
	.w6(32'h3af553f9),
	.w7(32'hbbb3a246),
	.w8(32'hbc0557d2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c524e),
	.w1(32'h3c46ebac),
	.w2(32'h3c1a557d),
	.w3(32'h3c1d7bdb),
	.w4(32'h3c5ea2e2),
	.w5(32'h3c3f2636),
	.w6(32'hbc392725),
	.w7(32'hbbec4b7f),
	.w8(32'h3a063cea),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf80ee1),
	.w1(32'h3c39f1f5),
	.w2(32'h3c296318),
	.w3(32'h3c66e558),
	.w4(32'h3b8a7a27),
	.w5(32'h3b6fc896),
	.w6(32'h3b9afd48),
	.w7(32'hba9c2bd7),
	.w8(32'h3c82657c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd75209),
	.w1(32'h3c631c6a),
	.w2(32'hbc22a6b4),
	.w3(32'h3ba8eba3),
	.w4(32'h3bcc6c15),
	.w5(32'hbc1c12d9),
	.w6(32'h3ca2ddd8),
	.w7(32'h3c8ddb2c),
	.w8(32'hbc4516ae),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b6f77),
	.w1(32'hbc14ef56),
	.w2(32'hba1c8525),
	.w3(32'hbc5c8879),
	.w4(32'hbc1d70f5),
	.w5(32'hbbe56fa4),
	.w6(32'hbc83ca6f),
	.w7(32'hbc4cbd7a),
	.w8(32'hbb824fef),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5bc15),
	.w1(32'hbb718567),
	.w2(32'h398bd971),
	.w3(32'hbbd7cb60),
	.w4(32'hbbec52cb),
	.w5(32'hbac3905f),
	.w6(32'hbb0e0142),
	.w7(32'hbbbd14da),
	.w8(32'hbb10b880),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb396d),
	.w1(32'hbb9b5c7f),
	.w2(32'hbc2c9a5c),
	.w3(32'hbbd05632),
	.w4(32'hbc301232),
	.w5(32'hbcabda4b),
	.w6(32'hbbe328a0),
	.w7(32'h3a361466),
	.w8(32'hbc758eb4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a66c8),
	.w1(32'hbb396406),
	.w2(32'h3c1197bf),
	.w3(32'hbcc6a631),
	.w4(32'hbcad2973),
	.w5(32'h3bb2d9be),
	.w6(32'hbceb7377),
	.w7(32'hbc703865),
	.w8(32'h3b8b97e7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ecb10),
	.w1(32'h3b0e9ef4),
	.w2(32'h3b041d21),
	.w3(32'h3c388c5d),
	.w4(32'h3c2ce010),
	.w5(32'hbb69dee2),
	.w6(32'h3c275a28),
	.w7(32'h3b653a19),
	.w8(32'h3b181623),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb138e2e),
	.w1(32'hbbede3c1),
	.w2(32'hbbfd277a),
	.w3(32'hbc29a4ce),
	.w4(32'h3b18c06d),
	.w5(32'h38209930),
	.w6(32'hba224dd0),
	.w7(32'hbb2324ac),
	.w8(32'h3bc1532e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac08553),
	.w1(32'h3b7de107),
	.w2(32'h3a55cebc),
	.w3(32'h3c206d42),
	.w4(32'hbb42b12b),
	.w5(32'h3b8d9471),
	.w6(32'h3ab46fb1),
	.w7(32'hbc227605),
	.w8(32'h3c38ca13),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb284811),
	.w1(32'h3ae921f3),
	.w2(32'hbb865337),
	.w3(32'hbb1bf620),
	.w4(32'hbbd6d10d),
	.w5(32'hbbc46372),
	.w6(32'h3af9ee8a),
	.w7(32'hbc16bf29),
	.w8(32'hbb5230d7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc79f9f),
	.w1(32'hbaddc5c6),
	.w2(32'hbb1328ff),
	.w3(32'hbbab5980),
	.w4(32'hbb27771d),
	.w5(32'hbaadc59b),
	.w6(32'h3c073efa),
	.w7(32'h3bc1415b),
	.w8(32'h3b09bf1c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fc0b9),
	.w1(32'h3aee4b8c),
	.w2(32'h3a48f631),
	.w3(32'hbbbca78c),
	.w4(32'h3b35357d),
	.w5(32'hbbd7eaad),
	.w6(32'hb8393e16),
	.w7(32'h3ba841ae),
	.w8(32'hbab465bb),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89100d),
	.w1(32'hbb8b843d),
	.w2(32'h3c757a0f),
	.w3(32'hbbbbd8c9),
	.w4(32'hb8af7ff8),
	.w5(32'h3c1caca9),
	.w6(32'hbb267e4a),
	.w7(32'hba20e785),
	.w8(32'h3bd87c74),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3456a2),
	.w1(32'h3b9f2dfb),
	.w2(32'hbc29c05a),
	.w3(32'h3bd18ac7),
	.w4(32'h3bc6b922),
	.w5(32'hbb891618),
	.w6(32'h3baa5565),
	.w7(32'h3ae75c6e),
	.w8(32'h3bd41c0f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a0c76),
	.w1(32'hbb0539e9),
	.w2(32'h3b9d5c82),
	.w3(32'hbc5e5bc9),
	.w4(32'hbaba81e8),
	.w5(32'h3bb803c3),
	.w6(32'hbb48fe87),
	.w7(32'hba662891),
	.w8(32'h3bcaa2e7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6c7b4),
	.w1(32'h3b32f4d4),
	.w2(32'h3b545315),
	.w3(32'h3b60954a),
	.w4(32'h3aad9266),
	.w5(32'hba41877b),
	.w6(32'h3b85df7c),
	.w7(32'h3a43d4c5),
	.w8(32'hbae69153),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49a1c7),
	.w1(32'hb9180b60),
	.w2(32'hbbfadef9),
	.w3(32'hbb55723b),
	.w4(32'hbacb939d),
	.w5(32'hbb9753fd),
	.w6(32'hbb92d5ae),
	.w7(32'hbad04476),
	.w8(32'hbb9cc9ca),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dd508),
	.w1(32'hbbe40802),
	.w2(32'h3c38af76),
	.w3(32'hbcbffd46),
	.w4(32'hbc544f37),
	.w5(32'h3b093e6d),
	.w6(32'hbc44ce82),
	.w7(32'hbc5f2f66),
	.w8(32'h3bc76969),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27a7fc),
	.w1(32'h3b944202),
	.w2(32'h3bafa41c),
	.w3(32'h3b6b6629),
	.w4(32'h3be1caa0),
	.w5(32'h3c26db1e),
	.w6(32'h3b63552e),
	.w7(32'h3c35bd49),
	.w8(32'hba2afb50),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c024470),
	.w1(32'h3b6584e4),
	.w2(32'h3c18c73a),
	.w3(32'h3bf657b7),
	.w4(32'h3c2c955e),
	.w5(32'h3bd15d2c),
	.w6(32'h3c19bf27),
	.w7(32'h3c046a81),
	.w8(32'h3bd01fa1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee38ca),
	.w1(32'hbb9685b2),
	.w2(32'hbc06e0a0),
	.w3(32'h3b13c7d5),
	.w4(32'h3b9e2500),
	.w5(32'hbbbad78e),
	.w6(32'h3b88f03e),
	.w7(32'h3a12d4d8),
	.w8(32'hbbb5cc14),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9e6c6),
	.w1(32'h3a9fd30f),
	.w2(32'h3a06b330),
	.w3(32'hbc1bf719),
	.w4(32'hbb3304bc),
	.w5(32'hba03d6fe),
	.w6(32'hbbdda9a5),
	.w7(32'hbc1cdb57),
	.w8(32'hba311b78),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ace9d),
	.w1(32'h3ab71a90),
	.w2(32'hbb43a7df),
	.w3(32'h3b741dcf),
	.w4(32'hbab84477),
	.w5(32'hbbb38643),
	.w6(32'hbb3ac289),
	.w7(32'hbbc9a3c0),
	.w8(32'hbbd4b4c9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb6e5),
	.w1(32'hbc002f62),
	.w2(32'h3c14fb21),
	.w3(32'hbc0a25b7),
	.w4(32'hbb24a7eb),
	.w5(32'h3b2330ac),
	.w6(32'hbb590f6a),
	.w7(32'hbb38fe60),
	.w8(32'h3aee6be8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa801c3),
	.w1(32'h3bc1d189),
	.w2(32'hbc10e235),
	.w3(32'h3988eb73),
	.w4(32'hbb8fa1b0),
	.w5(32'hbbff4417),
	.w6(32'hbb836e1c),
	.w7(32'hbc3c2a73),
	.w8(32'hba27fbf5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aa870),
	.w1(32'hbbf87554),
	.w2(32'h3b543056),
	.w3(32'hbc444e27),
	.w4(32'hbc13f9ed),
	.w5(32'hbc50c844),
	.w6(32'hbbb15f63),
	.w7(32'hbbc0b277),
	.w8(32'hbb6d2cf5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ebd0e),
	.w1(32'h3aeb57aa),
	.w2(32'hbbb52e27),
	.w3(32'hbc4f7658),
	.w4(32'hbc38973c),
	.w5(32'hbc951152),
	.w6(32'hbb28eb3e),
	.w7(32'hbc0c7fbc),
	.w8(32'hbbea1c6f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32cbaa),
	.w1(32'hbc1d9aff),
	.w2(32'hbc35a099),
	.w3(32'hbcc5e639),
	.w4(32'hbc95920e),
	.w5(32'hbbf70f52),
	.w6(32'hbc240aca),
	.w7(32'hbbb0ab62),
	.w8(32'hbbbad938),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cdea3),
	.w1(32'hbc299ba6),
	.w2(32'h3b014262),
	.w3(32'hbc95a6ec),
	.w4(32'hbc6b3832),
	.w5(32'hbbbf12d0),
	.w6(32'hbbbb1acc),
	.w7(32'hbc0eadd1),
	.w8(32'h3c42573d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c8b2),
	.w1(32'h3c172e25),
	.w2(32'h3b93b20d),
	.w3(32'hbbe630ad),
	.w4(32'hbb9855ac),
	.w5(32'h3ba3c07a),
	.w6(32'h3c437088),
	.w7(32'h3c11b4e9),
	.w8(32'h3abf7560),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a4d85),
	.w1(32'hbbe28e9f),
	.w2(32'h3bc901a7),
	.w3(32'hbb01729f),
	.w4(32'hbb80d4db),
	.w5(32'hba094d1a),
	.w6(32'hbb9acdb4),
	.w7(32'hbb33d8ec),
	.w8(32'hbbf84f46),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4117db),
	.w1(32'h3bd70359),
	.w2(32'h3c6b02e4),
	.w3(32'hba6398b0),
	.w4(32'hbbc12043),
	.w5(32'h3b034080),
	.w6(32'hbc7607e6),
	.w7(32'hbc606774),
	.w8(32'hbc90d9e9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf8536e),
	.w1(32'h3c8d1f18),
	.w2(32'h3ac22e67),
	.w3(32'h3b185e32),
	.w4(32'h38d916c4),
	.w5(32'hbaaebd7b),
	.w6(32'hbcf4ea97),
	.w7(32'hbcb4ecc0),
	.w8(32'h3a10b4f3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91d189),
	.w1(32'hbc270427),
	.w2(32'hbaa6d42f),
	.w3(32'h3b484bbc),
	.w4(32'hbbb3bf95),
	.w5(32'hbc1b9e29),
	.w6(32'hba422838),
	.w7(32'hbbf74dcd),
	.w8(32'hbbc60251),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f845b),
	.w1(32'hbb2cd70f),
	.w2(32'hbb074c6b),
	.w3(32'hbbcd282f),
	.w4(32'hbb3fa0ba),
	.w5(32'h3b22650a),
	.w6(32'hbb85c0d4),
	.w7(32'hba087ae4),
	.w8(32'h3b2f07de),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4381a),
	.w1(32'hbb814402),
	.w2(32'hbbcae015),
	.w3(32'hbbfb5c26),
	.w4(32'hbbe30cd6),
	.w5(32'hbb889792),
	.w6(32'h3ab8bdca),
	.w7(32'h3aa78b84),
	.w8(32'hbbae75a7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85fabfb),
	.w1(32'hbae0a412),
	.w2(32'h3b315768),
	.w3(32'hbbcd8ad5),
	.w4(32'h3b17ea70),
	.w5(32'hbb58228b),
	.w6(32'h3b189d11),
	.w7(32'h3c3303b6),
	.w8(32'h3b08b32c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc0933),
	.w1(32'hbb1276fb),
	.w2(32'hb9a35417),
	.w3(32'h3b90275e),
	.w4(32'h3accf221),
	.w5(32'hbc757379),
	.w6(32'h3bb520ed),
	.w7(32'hbb3d4b03),
	.w8(32'hbc513db9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3b32a),
	.w1(32'h3a39b0c0),
	.w2(32'h3bc20881),
	.w3(32'hbc8fa098),
	.w4(32'hbba9c357),
	.w5(32'h3abb7203),
	.w6(32'hbc8bc4f0),
	.w7(32'hbc1dffc1),
	.w8(32'hbc58bb53),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c274b5d),
	.w1(32'h3babe01a),
	.w2(32'hbc1661e8),
	.w3(32'hbc20564a),
	.w4(32'h3aaec6ea),
	.w5(32'hbc5349ad),
	.w6(32'hbc19cd60),
	.w7(32'hb951ff1e),
	.w8(32'hbc8e91a0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5990c2),
	.w1(32'h3ba05185),
	.w2(32'hbb8fdf93),
	.w3(32'hbc9fca4f),
	.w4(32'hbc45ba0c),
	.w5(32'hbb437052),
	.w6(32'hbcb4cfab),
	.w7(32'hbc549b21),
	.w8(32'h3c36fa0d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829bb5),
	.w1(32'hbbf5bd5f),
	.w2(32'h3c6246e4),
	.w3(32'hbb8027ff),
	.w4(32'hba89314e),
	.w5(32'h3c944e0f),
	.w6(32'h3b5e9e6b),
	.w7(32'h3b0e97dd),
	.w8(32'hbc0248b8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d385e),
	.w1(32'h3c2e4794),
	.w2(32'hbb380dd5),
	.w3(32'h3c6b5433),
	.w4(32'h3c3b128d),
	.w5(32'hbbc3bab4),
	.w6(32'hbbb90e4b),
	.w7(32'hbae7add3),
	.w8(32'hbb8224e2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b414490),
	.w1(32'h3a19f347),
	.w2(32'hbc6f0ea9),
	.w3(32'h3b9082f5),
	.w4(32'h3b2a031d),
	.w5(32'hbc3cbe80),
	.w6(32'hbc069301),
	.w7(32'hbb95f681),
	.w8(32'h3c83a45c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1494cb),
	.w1(32'hbc9e559d),
	.w2(32'hbc4f8e5b),
	.w3(32'hbbf15c30),
	.w4(32'hbbf368c5),
	.w5(32'hbcbf0644),
	.w6(32'h3d0e3351),
	.w7(32'h3c94ed2f),
	.w8(32'hbba69eaf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fbca7),
	.w1(32'hbc8628f2),
	.w2(32'h39f23888),
	.w3(32'hbccdd888),
	.w4(32'hbc8a3556),
	.w5(32'h39f3e948),
	.w6(32'hbc50e938),
	.w7(32'hbbb5b0a0),
	.w8(32'hbb9543e9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d87a8),
	.w1(32'h3b0738bd),
	.w2(32'h3b90a882),
	.w3(32'hbb02b62f),
	.w4(32'hbab7d05f),
	.w5(32'hbb9440db),
	.w6(32'hba6685bf),
	.w7(32'hbbe567bd),
	.w8(32'hbb07c1b8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0f382),
	.w1(32'hbc270ebe),
	.w2(32'h3cb0fa1a),
	.w3(32'hbc534784),
	.w4(32'hbc610e06),
	.w5(32'h3c19fef7),
	.w6(32'hbc144146),
	.w7(32'hbc38663c),
	.w8(32'hbc38fcda),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2625a1),
	.w1(32'h3cdc2d73),
	.w2(32'hbb528ed4),
	.w3(32'h3be8acda),
	.w4(32'h3ba46da7),
	.w5(32'hbacd5093),
	.w6(32'hbd03ffa5),
	.w7(32'hbcaf3fe2),
	.w8(32'h3b8bdf73),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0f71),
	.w1(32'hbb8fcfb2),
	.w2(32'hbb9d12a6),
	.w3(32'hbb830ba8),
	.w4(32'hba884d14),
	.w5(32'hbc100e38),
	.w6(32'h3b563ac1),
	.w7(32'hb91ef42f),
	.w8(32'hbbc03832),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34bb86),
	.w1(32'hbc1cbc8b),
	.w2(32'hba051e52),
	.w3(32'hbbf1b2da),
	.w4(32'hbbf378e0),
	.w5(32'h3b01bc8e),
	.w6(32'hb8036cf7),
	.w7(32'hbac0f02d),
	.w8(32'hba74e738),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b952867),
	.w1(32'h3b560960),
	.w2(32'hbb350ba2),
	.w3(32'hbb6a139f),
	.w4(32'hbb2ae735),
	.w5(32'hbbbd8b9c),
	.w6(32'hbb3cbcfa),
	.w7(32'hba015437),
	.w8(32'h3ab2ef7e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a9a15),
	.w1(32'h3a64951c),
	.w2(32'hbc06953b),
	.w3(32'h3ad2d86d),
	.w4(32'hb9b274e5),
	.w5(32'hbbfc5b0c),
	.w6(32'hbb0a1c3d),
	.w7(32'h3aa39333),
	.w8(32'hbab3a330),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc222f94),
	.w1(32'hbbf89dd2),
	.w2(32'h3c81b958),
	.w3(32'hbc79dafa),
	.w4(32'hbc373f94),
	.w5(32'h3be17114),
	.w6(32'hbc4a7463),
	.w7(32'hbbc77738),
	.w8(32'hbbea87bf),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfa2a38),
	.w1(32'h3ca7ed27),
	.w2(32'h3af3f8fb),
	.w3(32'h3bee8e75),
	.w4(32'h3bc4dafd),
	.w5(32'h3a72203b),
	.w6(32'hbca3146f),
	.w7(32'hbc367166),
	.w8(32'h3b759bb5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa684d1),
	.w1(32'hbba768ed),
	.w2(32'h3ac95058),
	.w3(32'h3bb9de5b),
	.w4(32'h3aaddd7b),
	.w5(32'hbb264098),
	.w6(32'h3b6702f8),
	.w7(32'hbac4bea0),
	.w8(32'hbb6a3251),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43de5f),
	.w1(32'h3b8be84e),
	.w2(32'h3a5b8f84),
	.w3(32'h3b6fa243),
	.w4(32'h3bed17fa),
	.w5(32'hbb83c8d8),
	.w6(32'hb98e91e4),
	.w7(32'hba2f7ab4),
	.w8(32'hba251fa2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21c840),
	.w1(32'hbbaa1dca),
	.w2(32'hb865b6d7),
	.w3(32'hbc0f9dae),
	.w4(32'h3b0130f3),
	.w5(32'hb9dfef85),
	.w6(32'hbb7d1214),
	.w7(32'h3b1b4876),
	.w8(32'h3bc6249d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b140a8d),
	.w1(32'h3afa4ebb),
	.w2(32'h3bfdedd2),
	.w3(32'hba559654),
	.w4(32'h3b1947fb),
	.w5(32'h3c099f81),
	.w6(32'h3c09ee32),
	.w7(32'h3c156fa5),
	.w8(32'h3bfd666f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b683a9b),
	.w1(32'hbb1e6c1a),
	.w2(32'h3b7a8903),
	.w3(32'hba2f0f3b),
	.w4(32'hbbd36af4),
	.w5(32'hbb8aad09),
	.w6(32'h3bd7d2c6),
	.w7(32'hba83cc91),
	.w8(32'hbc4817f4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15780a),
	.w1(32'h3b432a74),
	.w2(32'h3be6bae3),
	.w3(32'hbba2e695),
	.w4(32'h3c2f2b5e),
	.w5(32'hbb8222a8),
	.w6(32'hbc457689),
	.w7(32'hbaf9e23c),
	.w8(32'hbce288da),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdab9e1),
	.w1(32'h3c286b89),
	.w2(32'h38b7b8b9),
	.w3(32'hbc12202e),
	.w4(32'hbc37d309),
	.w5(32'hbba8f773),
	.w6(32'hbd364d06),
	.w7(32'hbd0c0bac),
	.w8(32'hbb4bba9e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ff848),
	.w1(32'h3bb39893),
	.w2(32'h3b266c5d),
	.w3(32'h3a532da2),
	.w4(32'h3bc2d247),
	.w5(32'h3b60afd8),
	.w6(32'h3a4585ca),
	.w7(32'h3a79c021),
	.w8(32'hba857dbb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddf381),
	.w1(32'h3b51d31d),
	.w2(32'h3b9a59dd),
	.w3(32'hbb6c3a26),
	.w4(32'h3b82d68b),
	.w5(32'hbbc001f9),
	.w6(32'hbbe63f0e),
	.w7(32'hbb89801f),
	.w8(32'hbb03e033),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99424b),
	.w1(32'hbb6105d2),
	.w2(32'h3bc2c5f3),
	.w3(32'hbc062e5e),
	.w4(32'hbc4d233e),
	.w5(32'h3bdf65ac),
	.w6(32'h3b7a20c7),
	.w7(32'hbb73aeaa),
	.w8(32'hbb0641c8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b981bf2),
	.w1(32'h3a1fe7fa),
	.w2(32'hbae93448),
	.w3(32'hba6b5b07),
	.w4(32'h39a5d4f6),
	.w5(32'hbcaf0734),
	.w6(32'hbbf77f57),
	.w7(32'hbb6c732d),
	.w8(32'hbc9a847b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0009c),
	.w1(32'hbc632464),
	.w2(32'hbaaef677),
	.w3(32'hbc00caad),
	.w4(32'hbbc7726d),
	.w5(32'h3b65dd5f),
	.w6(32'hbafd1343),
	.w7(32'h3b566f05),
	.w8(32'h3b93d966),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974054c),
	.w1(32'h3b0b860b),
	.w2(32'hbd2b56c3),
	.w3(32'h3c0a480d),
	.w4(32'h3ba86c50),
	.w5(32'hbb9f38e7),
	.w6(32'h3bf0f845),
	.w7(32'h3aafd593),
	.w8(32'h3cae697b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda6282d),
	.w1(32'hbd889bec),
	.w2(32'hbb888963),
	.w3(32'h3cb30b36),
	.w4(32'hbc5e8eb2),
	.w5(32'hbc027e1a),
	.w6(32'h3de517dc),
	.w7(32'h3d2271f2),
	.w8(32'h3a7f1ff2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f3fd),
	.w1(32'hbb92c2e4),
	.w2(32'hbc274416),
	.w3(32'hbabddb1f),
	.w4(32'hbb061110),
	.w5(32'hba75f9aa),
	.w6(32'h3b11ab05),
	.w7(32'h37fd79a9),
	.w8(32'h3b0deddf),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd052f2),
	.w1(32'hbc058a05),
	.w2(32'hbdbcc2ff),
	.w3(32'h3bbd91d5),
	.w4(32'hbb062a9e),
	.w5(32'hbcda955e),
	.w6(32'hbbecceb9),
	.w7(32'hbaf0bc93),
	.w8(32'h3d007509),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe09260a),
	.w1(32'hbdc81356),
	.w2(32'h399d0559),
	.w3(32'h3ccaad9d),
	.w4(32'hbb2c16f4),
	.w5(32'hbad0531a),
	.w6(32'h3e2dce5d),
	.w7(32'h3da00bb7),
	.w8(32'hbb5a10e7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc249f),
	.w1(32'hbb4a8bc3),
	.w2(32'h3c9bded6),
	.w3(32'hba8b7ffb),
	.w4(32'hbbe8fd45),
	.w5(32'hbb3bcd83),
	.w6(32'hbb10d0d1),
	.w7(32'hbc10f9ec),
	.w8(32'hbc7331d8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2a3ede),
	.w1(32'h3d0f46be),
	.w2(32'hb994ce8d),
	.w3(32'hbc28a9f9),
	.w4(32'h3bf71ac2),
	.w5(32'hbb2dea31),
	.w6(32'hbd76a4f2),
	.w7(32'hbccf4199),
	.w8(32'hbc151489),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf706fd),
	.w1(32'h3bba1063),
	.w2(32'hbd814a6d),
	.w3(32'h3b9dd018),
	.w4(32'h3a044776),
	.w5(32'hbc60b24a),
	.w6(32'h3abe698c),
	.w7(32'hbbd2cbac),
	.w8(32'h3d15d35a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdc37b48),
	.w1(32'hbd7d4aaf),
	.w2(32'h3c21da82),
	.w3(32'h3d165dcf),
	.w4(32'h3c0692a8),
	.w5(32'h386529ba),
	.w6(32'h3e1b31df),
	.w7(32'h3d8d6a1a),
	.w8(32'h3bbe2d89),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13e281),
	.w1(32'h3bf2de11),
	.w2(32'hbbb3d095),
	.w3(32'hbbb8a66b),
	.w4(32'hbbbcd07c),
	.w5(32'hbc56a1f0),
	.w6(32'h3b91d7d3),
	.w7(32'h39869bc1),
	.w8(32'hbbcd4578),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d47868),
	.w1(32'h3aaeaa12),
	.w2(32'h3b370e44),
	.w3(32'hbb06dd23),
	.w4(32'hbb8a748b),
	.w5(32'hb9e234bc),
	.w6(32'hbc27f2ba),
	.w7(32'hbc512646),
	.w8(32'hbbcc6c52),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036f6c),
	.w1(32'hbb4d7c85),
	.w2(32'h3aba8729),
	.w3(32'hbb08e3cb),
	.w4(32'h39fc26c5),
	.w5(32'h3bb5362c),
	.w6(32'hbc0d4f30),
	.w7(32'hbb7bb166),
	.w8(32'hbb034e87),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ced53),
	.w1(32'h3acd6248),
	.w2(32'hbc313b60),
	.w3(32'h3b2f7fcd),
	.w4(32'h39fab6d2),
	.w5(32'hbb74bd01),
	.w6(32'hbbf9e422),
	.w7(32'hbc0874ca),
	.w8(32'hbab30904),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9fe33),
	.w1(32'hba054ef2),
	.w2(32'h3d88301d),
	.w3(32'hbbad35d0),
	.w4(32'h3b170d95),
	.w5(32'h3c945563),
	.w6(32'hbbac394d),
	.w7(32'hb916f687),
	.w8(32'hbd0aaf4d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dc87fcb),
	.w1(32'h3d8d64ab),
	.w2(32'hba8ee857),
	.w3(32'hbce2c1ff),
	.w4(32'hbbb06cb0),
	.w5(32'h399f4429),
	.w6(32'hbe1176f6),
	.w7(32'hbd8cf46b),
	.w8(32'h3a9f2f29),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd443bd),
	.w1(32'h3b94b713),
	.w2(32'h3bbe8385),
	.w3(32'h3be61720),
	.w4(32'hbb8a253d),
	.w5(32'h3bd3c9c3),
	.w6(32'h3b8102b9),
	.w7(32'h3b4a1529),
	.w8(32'h39a2d015),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978b176),
	.w1(32'h3ad25232),
	.w2(32'hbc056e88),
	.w3(32'h3c01152b),
	.w4(32'hbaa92550),
	.w5(32'hbc221fb8),
	.w6(32'h3be09acf),
	.w7(32'hba7ab46a),
	.w8(32'hbb4eea72),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936fc0),
	.w1(32'hbb2d62a2),
	.w2(32'hbb2e5e7a),
	.w3(32'h3a4ea05d),
	.w4(32'h3b8e85d6),
	.w5(32'hba8668b3),
	.w6(32'h3b009820),
	.w7(32'h3b7a4103),
	.w8(32'h3b2c25c6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10e973),
	.w1(32'h3b6eb6dc),
	.w2(32'h3d66381a),
	.w3(32'h3c0bb8f4),
	.w4(32'h3bb9376e),
	.w5(32'h3c12d0b3),
	.w6(32'hbb5470e0),
	.w7(32'hbbd0bcca),
	.w8(32'hbcfeb25f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd26957),
	.w1(32'h3daf87c1),
	.w2(32'hbb8a9ae3),
	.w3(32'hbc8e7019),
	.w4(32'h3c562542),
	.w5(32'hbb55b156),
	.w6(32'hbe09eaf3),
	.w7(32'hbd6918df),
	.w8(32'hba860663),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebf002),
	.w1(32'hbabbe004),
	.w2(32'hbb4d2ad4),
	.w3(32'h3be31591),
	.w4(32'h3a9ccb79),
	.w5(32'h3b147a80),
	.w6(32'hbaa67958),
	.w7(32'hbaf6f9b8),
	.w8(32'h3aa4bcfb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b83022),
	.w1(32'hbbc7ef16),
	.w2(32'h3b842527),
	.w3(32'h3a5e701b),
	.w4(32'h3b8e2c9b),
	.w5(32'h3b9e1f44),
	.w6(32'h3b670e63),
	.w7(32'h3bbdf8e4),
	.w8(32'h3b458c1f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0eb59c),
	.w1(32'h3be1282c),
	.w2(32'hbbd211f8),
	.w3(32'h3bfe082e),
	.w4(32'h3c3824ac),
	.w5(32'h3aa317a8),
	.w6(32'h3b579225),
	.w7(32'h3c34e58c),
	.w8(32'h3a6fcf82),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ffd70),
	.w1(32'hbc071838),
	.w2(32'hbc02d171),
	.w3(32'hbc00df14),
	.w4(32'hbc2294ee),
	.w5(32'hbc49a706),
	.w6(32'h3b1b9425),
	.w7(32'hb9826232),
	.w8(32'h38a03c71),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93aa75b),
	.w1(32'hb9a5d070),
	.w2(32'hbb5af2bd),
	.w3(32'hbc5c010c),
	.w4(32'hbbc169a8),
	.w5(32'hbb1d915e),
	.w6(32'hbb832a9f),
	.w7(32'h3bae1a95),
	.w8(32'h3b54462c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1158d),
	.w1(32'hbbca062a),
	.w2(32'hbb1f8bb3),
	.w3(32'h3aa9f7c8),
	.w4(32'h3c22cb82),
	.w5(32'hbbd1d141),
	.w6(32'hba824cba),
	.w7(32'h3a85171a),
	.w8(32'hbc46260b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62985a),
	.w1(32'hbaa65625),
	.w2(32'hbb49b82a),
	.w3(32'hbc10b2b9),
	.w4(32'hbc4fe133),
	.w5(32'hbbcf1964),
	.w6(32'hbc68b29c),
	.w7(32'hbcada08d),
	.w8(32'hbc08ec7f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd6200),
	.w1(32'hbafd1002),
	.w2(32'h3bb8e218),
	.w3(32'h3bc2509f),
	.w4(32'h3c460c2b),
	.w5(32'h3b8068ba),
	.w6(32'h3bf3db3d),
	.w7(32'h3b8b16fc),
	.w8(32'h3bc25926),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12985e),
	.w1(32'h3c3f1a94),
	.w2(32'hbb8581fe),
	.w3(32'h3b211ccf),
	.w4(32'h3a309473),
	.w5(32'hbbb29825),
	.w6(32'hba0eb886),
	.w7(32'hbc5c7f33),
	.w8(32'h3c6f7868),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb436e06),
	.w1(32'hbc952fb0),
	.w2(32'h3c8eb632),
	.w3(32'hbb0dd520),
	.w4(32'hbc37b235),
	.w5(32'h3c1f2bd3),
	.w6(32'h3cea614c),
	.w7(32'h3c767bcf),
	.w8(32'h3befc214),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96c6f8),
	.w1(32'h3c93dfaa),
	.w2(32'h3c4868aa),
	.w3(32'h3b580034),
	.w4(32'h3c67f90b),
	.w5(32'h3b59abaa),
	.w6(32'h3c037166),
	.w7(32'h3c2170f6),
	.w8(32'h3be32ddb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86bfd3),
	.w1(32'h3c0e6ec1),
	.w2(32'hba67d7c9),
	.w3(32'h3be237e0),
	.w4(32'h3b804afd),
	.w5(32'hbb1d4ce2),
	.w6(32'h3aa41eb9),
	.w7(32'h3b4f2fce),
	.w8(32'h3aa9e3b9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4c52a),
	.w1(32'h3c9d4673),
	.w2(32'h3baac810),
	.w3(32'hbb00d72b),
	.w4(32'h3c34ae06),
	.w5(32'hb9bceda8),
	.w6(32'hbb3162f1),
	.w7(32'h3a9e7e3a),
	.w8(32'h3b2246c3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba44d4d),
	.w1(32'hbb677d81),
	.w2(32'h3bf4307e),
	.w3(32'h3b519fde),
	.w4(32'h39e1d265),
	.w5(32'h3bf3f254),
	.w6(32'h3b33186b),
	.w7(32'hbb20dfdc),
	.w8(32'h3c02c45d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0735d0),
	.w1(32'h3b92b27b),
	.w2(32'hbbb6d13d),
	.w3(32'h3be14e0a),
	.w4(32'h3b014a14),
	.w5(32'hbbb09447),
	.w6(32'h3ba343c4),
	.w7(32'h3a342762),
	.w8(32'hbbcf352f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab87121),
	.w1(32'hbaee98b7),
	.w2(32'h3b19795e),
	.w3(32'h3b4070bc),
	.w4(32'hbab29afc),
	.w5(32'h3c4a1d6f),
	.w6(32'hba8557db),
	.w7(32'h3b10faf1),
	.w8(32'h3b483893),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f4a28),
	.w1(32'hbb720107),
	.w2(32'h3cb3525c),
	.w3(32'h3c34bb29),
	.w4(32'h3b7051f8),
	.w5(32'h3c8c6bd4),
	.w6(32'h3bcad0a0),
	.w7(32'h3b9d52b8),
	.w8(32'h3979a947),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1db02f),
	.w1(32'hbba16bb1),
	.w2(32'hbba83ed9),
	.w3(32'h3ad68505),
	.w4(32'hbc6d53ad),
	.w5(32'h3ab671a3),
	.w6(32'hb9cebe07),
	.w7(32'hbc073fe9),
	.w8(32'h3b9a3296),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99840d6),
	.w1(32'h3a88a8af),
	.w2(32'h3944bdd2),
	.w3(32'hba15f871),
	.w4(32'hbb7844d5),
	.w5(32'h3958a555),
	.w6(32'h3b941cc0),
	.w7(32'h3b959c17),
	.w8(32'hbbdbc672),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae762e3),
	.w1(32'hbbcd4e0d),
	.w2(32'h3c341b06),
	.w3(32'hba4874a1),
	.w4(32'hbb76cf52),
	.w5(32'h3af8017a),
	.w6(32'h3bc8920b),
	.w7(32'hbb86ee46),
	.w8(32'h3b37dd50),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbb91d),
	.w1(32'h3c4bf93c),
	.w2(32'h3c0d2608),
	.w3(32'hb9b92b6d),
	.w4(32'h3bb32e76),
	.w5(32'hbb1a5293),
	.w6(32'hbbdd30ba),
	.w7(32'h3a26b4c3),
	.w8(32'hbbdb4840),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15db4d),
	.w1(32'h3ba005fd),
	.w2(32'hbbfcc0b1),
	.w3(32'h3b42e1d9),
	.w4(32'hba8be084),
	.w5(32'h3af84b53),
	.w6(32'hbb945a2d),
	.w7(32'h3aa9f9dd),
	.w8(32'hbba8ab3f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba823c8f),
	.w1(32'hbba89fd0),
	.w2(32'hbb356a86),
	.w3(32'h3b36f64d),
	.w4(32'hbbdd4c1d),
	.w5(32'hba829b30),
	.w6(32'hba2dfda0),
	.w7(32'h3a68be97),
	.w8(32'h3b4be824),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6a9f8),
	.w1(32'hbbc8e2d3),
	.w2(32'h3be453d8),
	.w3(32'hbbb89ada),
	.w4(32'hb885e308),
	.w5(32'hba2d2a44),
	.w6(32'h39c36524),
	.w7(32'h3a96d889),
	.w8(32'hbb9caff3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67924e),
	.w1(32'h39cc5dec),
	.w2(32'h3d45d9be),
	.w3(32'h3b94bd79),
	.w4(32'h3bc9eb8c),
	.w5(32'h3c9ef3b4),
	.w6(32'hbb982932),
	.w7(32'hb8ad77b9),
	.w8(32'hbcefe9e3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9d50d2),
	.w1(32'h3d8b2528),
	.w2(32'hbab96d77),
	.w3(32'hbb9de72c),
	.w4(32'h3c891aa5),
	.w5(32'h3aa74b11),
	.w6(32'hbde896e3),
	.w7(32'hbd6d2e81),
	.w8(32'hbb93014d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85461c),
	.w1(32'h3aae74ed),
	.w2(32'hbb7d4e6a),
	.w3(32'h3b7e2343),
	.w4(32'hb9db0508),
	.w5(32'hba897f91),
	.w6(32'hbb3ce613),
	.w7(32'hbb3fa2a2),
	.w8(32'hbc2507af),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1198fe),
	.w1(32'hbc1effd2),
	.w2(32'hbb0a342c),
	.w3(32'hbbc2326e),
	.w4(32'hbb9e1150),
	.w5(32'hbad2a757),
	.w6(32'hba9a2fc4),
	.w7(32'hba65f4de),
	.w8(32'h3b8862de),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb831e20),
	.w1(32'hbb3062a5),
	.w2(32'hbba811be),
	.w3(32'h3ba6a839),
	.w4(32'hbc08a128),
	.w5(32'h39732dfe),
	.w6(32'hbacdb549),
	.w7(32'h3c1657f1),
	.w8(32'h3a57daa3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e2c2e),
	.w1(32'hba06e771),
	.w2(32'h3c1a51b9),
	.w3(32'h3b6f1f6e),
	.w4(32'hb986cecf),
	.w5(32'h3b894406),
	.w6(32'h3b5e917e),
	.w7(32'h3c0672ff),
	.w8(32'hbb1340a6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993b8ba),
	.w1(32'h3aa62c7d),
	.w2(32'hbc0793ce),
	.w3(32'hbc53843f),
	.w4(32'hbb78c2d7),
	.w5(32'hbb65f4f6),
	.w6(32'hbcae2e11),
	.w7(32'hbbccfd09),
	.w8(32'hbb71f4e6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacf6cc),
	.w1(32'hb93841e7),
	.w2(32'h3afece84),
	.w3(32'hbbabfc24),
	.w4(32'hbbb8b8dd),
	.w5(32'h3c90698c),
	.w6(32'hbb3bd4ff),
	.w7(32'h39033d0a),
	.w8(32'h3c579f93),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce28e0f),
	.w1(32'hbcebe545),
	.w2(32'hbc1d419e),
	.w3(32'h3c85c26e),
	.w4(32'hbc9b13eb),
	.w5(32'hbaf2f98e),
	.w6(32'h3d6112ad),
	.w7(32'h3b760848),
	.w8(32'h39632fbb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdec4da),
	.w1(32'h39754a3e),
	.w2(32'hbbc65439),
	.w3(32'hbba8e28d),
	.w4(32'h3c15b1ee),
	.w5(32'hbb23ee38),
	.w6(32'hba21d601),
	.w7(32'h3c3ba7a7),
	.w8(32'h3b16fde6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00c87b),
	.w1(32'hb7244213),
	.w2(32'h3aad8d72),
	.w3(32'hb8f0cbc1),
	.w4(32'hbaa762e1),
	.w5(32'hbac1a3ef),
	.w6(32'h3c0c5346),
	.w7(32'h3b874a30),
	.w8(32'h3ace380e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42a005),
	.w1(32'hb9c9b3a6),
	.w2(32'h3acd7747),
	.w3(32'h3a8472b7),
	.w4(32'hbb9b4798),
	.w5(32'h3c1e926d),
	.w6(32'h3a56f8e9),
	.w7(32'h3b446fd3),
	.w8(32'h3acdfd1b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe62a79),
	.w1(32'h3b577cc6),
	.w2(32'h3aa01fb5),
	.w3(32'hbc0b80dd),
	.w4(32'h3bb0129e),
	.w5(32'h3b22ae7f),
	.w6(32'hbc135d91),
	.w7(32'h3b7e4ae1),
	.w8(32'hbae5f9ca),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a0a88),
	.w1(32'hbaafbaae),
	.w2(32'h3c9a3a45),
	.w3(32'h3b6b51a7),
	.w4(32'h3bc11fed),
	.w5(32'h3c44fcdf),
	.w6(32'h3b078820),
	.w7(32'h3b887eb5),
	.w8(32'h3bb859b0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd47f6d),
	.w1(32'h3c9ee188),
	.w2(32'hba0e91c9),
	.w3(32'h3c1e6df3),
	.w4(32'h3b5153bb),
	.w5(32'h3b92428b),
	.w6(32'hbbdc70cf),
	.w7(32'hbc6824c9),
	.w8(32'h3a90eaea),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17908),
	.w1(32'hbbfdaed2),
	.w2(32'hbbd531ad),
	.w3(32'hbb8f1e87),
	.w4(32'hbbf4771e),
	.w5(32'hbb9fd644),
	.w6(32'hbb11c5b9),
	.w7(32'hb98e6eb6),
	.w8(32'hbc303b8e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae5a43),
	.w1(32'h3b176d3e),
	.w2(32'h3cbe1bd2),
	.w3(32'hbbb9578e),
	.w4(32'hbc413e53),
	.w5(32'h3cf95920),
	.w6(32'hbc07b9c4),
	.w7(32'hbb94e733),
	.w8(32'h3c906f9b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d098065),
	.w1(32'h3cdd2721),
	.w2(32'hbc19a06e),
	.w3(32'h3d1696e6),
	.w4(32'h3ce8f95f),
	.w5(32'hbbeea46e),
	.w6(32'h3c48b1b3),
	.w7(32'h3c06562b),
	.w8(32'hbb8edf3e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb506),
	.w1(32'hbbbf3884),
	.w2(32'h3c7e801f),
	.w3(32'hb9e263d3),
	.w4(32'hbbcb6e98),
	.w5(32'h3a8786bf),
	.w6(32'h3aafe01c),
	.w7(32'h3aa3e62f),
	.w8(32'hbc22a068),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cea7c),
	.w1(32'h3c16553d),
	.w2(32'h3d55b7c3),
	.w3(32'h3afbed68),
	.w4(32'h3a8909bb),
	.w5(32'h3cb5ab95),
	.w6(32'hbc2a1f41),
	.w7(32'hbc1091d6),
	.w8(32'hbc0517b5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6c5830),
	.w1(32'h3d1a022c),
	.w2(32'h3a12e413),
	.w3(32'hbbc50283),
	.w4(32'hbc1702ba),
	.w5(32'h3b5c2e8a),
	.w6(32'hbd6545de),
	.w7(32'hbd215534),
	.w8(32'h38871d05),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8155b49),
	.w1(32'hbba77ba3),
	.w2(32'hbbb40c29),
	.w3(32'hbb012665),
	.w4(32'hbbb0c147),
	.w5(32'hbb2c38cd),
	.w6(32'hbb6d7359),
	.w7(32'hbb837c58),
	.w8(32'hbb021c8d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11170f),
	.w1(32'hbb8b12d3),
	.w2(32'h3ab4028d),
	.w3(32'hbbbb107a),
	.w4(32'hbb9fbcca),
	.w5(32'h3adb5986),
	.w6(32'hb9dac24f),
	.w7(32'hbad9901e),
	.w8(32'hbba8d88f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbeb95),
	.w1(32'hbb05fc8c),
	.w2(32'h3a6c0d04),
	.w3(32'h3b2194d8),
	.w4(32'h3b22b965),
	.w5(32'h3a0c2bff),
	.w6(32'h39eb20d8),
	.w7(32'hbbb83dc9),
	.w8(32'hbaf2a20d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd56fe),
	.w1(32'hbbfa3251),
	.w2(32'h3b782a30),
	.w3(32'h3c35b480),
	.w4(32'h3ac56f03),
	.w5(32'h3b56e832),
	.w6(32'h3b085dce),
	.w7(32'hbb4362ec),
	.w8(32'hbb27c84c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5c73),
	.w1(32'hbb0377e8),
	.w2(32'hbbf7b392),
	.w3(32'h3ba28f69),
	.w4(32'hbbff6ffc),
	.w5(32'h3c1df5df),
	.w6(32'hba866a7c),
	.w7(32'h391d3bd2),
	.w8(32'h3c4fe626),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5e5d6),
	.w1(32'h3c638cd9),
	.w2(32'hbc2e14d5),
	.w3(32'h3abf1237),
	.w4(32'hbbea8129),
	.w5(32'hbbe993f0),
	.w6(32'h3bad44e3),
	.w7(32'hbc8b3289),
	.w8(32'hbabe0d8c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52ed31),
	.w1(32'hba8b5499),
	.w2(32'hba45a71f),
	.w3(32'h3a95cafa),
	.w4(32'hb481cb99),
	.w5(32'hbb3fb103),
	.w6(32'hbba6a5c3),
	.w7(32'hbb86996c),
	.w8(32'hbb51d523),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad62855),
	.w1(32'hbbd320a2),
	.w2(32'hbbeda8b3),
	.w3(32'hbaf44469),
	.w4(32'hbb1eb6ad),
	.w5(32'hbba862e8),
	.w6(32'hbbb8d160),
	.w7(32'h3ab68045),
	.w8(32'h37fa2d12),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc33dc7),
	.w1(32'hbba18777),
	.w2(32'hbb13eb21),
	.w3(32'hb9be56cc),
	.w4(32'h3b4af340),
	.w5(32'h3bc81243),
	.w6(32'h3b5de8c4),
	.w7(32'h3a6ace22),
	.w8(32'h3bc38918),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d407b),
	.w1(32'h3c3c204d),
	.w2(32'hbae0e3b9),
	.w3(32'h3c4484db),
	.w4(32'h3c632f43),
	.w5(32'h3b74d481),
	.w6(32'h3bf0ca11),
	.w7(32'h3b8c3474),
	.w8(32'h3c47d2ac),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12bbc6),
	.w1(32'hbb1e815c),
	.w2(32'hbc02d418),
	.w3(32'h3ac6ef97),
	.w4(32'h3bf4f5d2),
	.w5(32'hbbd502a5),
	.w6(32'h3c0cf292),
	.w7(32'h3c1fbfd2),
	.w8(32'hbbdb6368),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7003e4),
	.w1(32'h3aafacdf),
	.w2(32'hbb9db117),
	.w3(32'hbb601864),
	.w4(32'h3c408d66),
	.w5(32'hbb85bbca),
	.w6(32'h3b96d7ec),
	.w7(32'h3bd457d0),
	.w8(32'hbc43b5ba),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb37172),
	.w1(32'hba273b5a),
	.w2(32'hbba51c0c),
	.w3(32'h39622176),
	.w4(32'h3a4af42c),
	.w5(32'hbb7695f2),
	.w6(32'hbb5f0e60),
	.w7(32'hbbc93d85),
	.w8(32'h3bfce3d5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb583c1a),
	.w1(32'h39144554),
	.w2(32'hbbdd3bc4),
	.w3(32'hbc5936ef),
	.w4(32'hbc427bf0),
	.w5(32'h3a33f052),
	.w6(32'hbbc9c87c),
	.w7(32'hbbcd1024),
	.w8(32'h3b8f3449),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dcc6be),
	.w1(32'hbb596022),
	.w2(32'h3ace4cc6),
	.w3(32'hbbb5e497),
	.w4(32'h3ba9bd93),
	.w5(32'h3aa1e92b),
	.w6(32'h3b80b834),
	.w7(32'h3b3a1923),
	.w8(32'h3b0974af),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc092ea),
	.w1(32'h3bac9110),
	.w2(32'hbbf41e50),
	.w3(32'h3b233b7c),
	.w4(32'h3bb8b997),
	.w5(32'hbb5a25bd),
	.w6(32'hbac4079e),
	.w7(32'h3aecb823),
	.w8(32'h3a8ba8bb),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc348212),
	.w1(32'hbc2f7010),
	.w2(32'hbb967260),
	.w3(32'hbbc9f180),
	.w4(32'hbb915487),
	.w5(32'hb82d3aae),
	.w6(32'hbb79f914),
	.w7(32'hba77e87e),
	.w8(32'h3b62ca8a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68cc70),
	.w1(32'h3b6cb3b9),
	.w2(32'hbbeb7206),
	.w3(32'h38165e5f),
	.w4(32'h3ba170e0),
	.w5(32'h3b0fc717),
	.w6(32'h3b8a467c),
	.w7(32'h3afc7b23),
	.w8(32'hbbd2758e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52029e),
	.w1(32'hbbf3be2e),
	.w2(32'hbba1726b),
	.w3(32'h3b1a1f59),
	.w4(32'hbb57f74f),
	.w5(32'hbb89ff74),
	.w6(32'hbc362c7f),
	.w7(32'hbb7071eb),
	.w8(32'hbbc3ad4d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8cd76),
	.w1(32'hbb877b5f),
	.w2(32'hbb8ff9ae),
	.w3(32'hbaa09557),
	.w4(32'hb94b30fa),
	.w5(32'hbc42128b),
	.w6(32'hbaab806b),
	.w7(32'h3b1b8c0f),
	.w8(32'hbc4bbb6e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4c8f),
	.w1(32'hbb0a987e),
	.w2(32'hbbc0e904),
	.w3(32'hbc1e2b47),
	.w4(32'hbc4cc38b),
	.w5(32'hbc1f09e7),
	.w6(32'hbc61bfde),
	.w7(32'hbc54719d),
	.w8(32'h3afd3d48),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc645316),
	.w1(32'hbc61769a),
	.w2(32'hba660797),
	.w3(32'hbc8fdbd9),
	.w4(32'hbc8d49df),
	.w5(32'hbb17609e),
	.w6(32'h3b416fb6),
	.w7(32'h3b4a1c22),
	.w8(32'hbbc532c9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6985a6),
	.w1(32'hbb911f22),
	.w2(32'hbc01b0d7),
	.w3(32'hbbedb2e4),
	.w4(32'hbc081ad6),
	.w5(32'hbc5e4ea9),
	.w6(32'hbbaa36cf),
	.w7(32'hbbd6c283),
	.w8(32'hbaff39cd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ec30b),
	.w1(32'hbc339eb4),
	.w2(32'h3b938d42),
	.w3(32'hbcacf79c),
	.w4(32'hbca1efc4),
	.w5(32'hbafc9571),
	.w6(32'hbba81873),
	.w7(32'hbb602883),
	.w8(32'h3b44498d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb935eab),
	.w1(32'hbb43d782),
	.w2(32'hbb7b848e),
	.w3(32'hbc1abdd0),
	.w4(32'hbbdbea2f),
	.w5(32'hbbf49a88),
	.w6(32'hba5b5f54),
	.w7(32'h3c520a42),
	.w8(32'h3a8fd23c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc227a56),
	.w1(32'hbaba1b2a),
	.w2(32'hbab92737),
	.w3(32'hbbbf1049),
	.w4(32'hbb0b8ee0),
	.w5(32'h39088647),
	.w6(32'hba53902a),
	.w7(32'hbbd768e3),
	.w8(32'hbafcf0d8),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70b0a1),
	.w1(32'hbb06934d),
	.w2(32'hbbc18422),
	.w3(32'hba8b229a),
	.w4(32'hba869e58),
	.w5(32'hbb30b3d1),
	.w6(32'h3bd3865c),
	.w7(32'h394be4cc),
	.w8(32'h3c2b98e2),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5551af),
	.w1(32'hbc2f0c86),
	.w2(32'hbc9eaed4),
	.w3(32'h3b9d8f98),
	.w4(32'h3bdd1e2f),
	.w5(32'hbc0c4281),
	.w6(32'h3cf38f55),
	.w7(32'h3cae2bb9),
	.w8(32'h3bf588c8),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0361a0),
	.w1(32'hbcc6cd88),
	.w2(32'hbb3e8500),
	.w3(32'h3bfb15bb),
	.w4(32'hbb82dba6),
	.w5(32'h399b2f46),
	.w6(32'h3d47c1fe),
	.w7(32'h3c9a5444),
	.w8(32'hbc0465fb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b476674),
	.w1(32'hbb7f1e97),
	.w2(32'hbc04af73),
	.w3(32'h3b53ece9),
	.w4(32'hbb4e729e),
	.w5(32'hbc4a6a1d),
	.w6(32'h3b97fd7b),
	.w7(32'h38f3a319),
	.w8(32'hbb3503af),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43cd62),
	.w1(32'hbb776c08),
	.w2(32'h3ba1ee07),
	.w3(32'hbc43813a),
	.w4(32'hbba2a6a1),
	.w5(32'h3c12de84),
	.w6(32'hbb40f217),
	.w7(32'h3bda56d0),
	.w8(32'h39becca1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad56a2a),
	.w1(32'hb93631bd),
	.w2(32'hba7eeefb),
	.w3(32'hbb87ed09),
	.w4(32'h3a6aa5b1),
	.w5(32'h3b08394c),
	.w6(32'h3b71f14b),
	.w7(32'h3c1817a7),
	.w8(32'h3b863c9e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35be92),
	.w1(32'h3826f141),
	.w2(32'hba944c8a),
	.w3(32'hbbe6af38),
	.w4(32'h394fe204),
	.w5(32'hbaa13a8b),
	.w6(32'h3be98862),
	.w7(32'h3bad3de2),
	.w8(32'h3bdf6e3c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b9c8),
	.w1(32'h38cf23b7),
	.w2(32'hbb4ba8c2),
	.w3(32'hbb004275),
	.w4(32'h3aad498a),
	.w5(32'hb9b5e085),
	.w6(32'h3ac36fa7),
	.w7(32'h3a7b5d5c),
	.w8(32'h3b0a1e35),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule