module layer_8_featuremap_81(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ee1b6),
	.w1(32'h3b861354),
	.w2(32'hba295464),
	.w3(32'hb919f372),
	.w4(32'h3ae8cda1),
	.w5(32'hba5d5bac),
	.w6(32'hba36f514),
	.w7(32'h3aaa5cf3),
	.w8(32'hba44c1d5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a1f34),
	.w1(32'hb9747d11),
	.w2(32'h3b0c5aab),
	.w3(32'h3a5bddcf),
	.w4(32'h3af38641),
	.w5(32'h3b3e1d34),
	.w6(32'h3b289be8),
	.w7(32'h3accfef2),
	.w8(32'h3b1e3663),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0028be),
	.w1(32'hbafe8360),
	.w2(32'hba915f7a),
	.w3(32'hb9db0755),
	.w4(32'h3a85781a),
	.w5(32'h3a08e9e6),
	.w6(32'h3aac055f),
	.w7(32'h3b1bd19c),
	.w8(32'h3937c71c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0703),
	.w1(32'hb7a63a70),
	.w2(32'hba1ee187),
	.w3(32'h3b7af2ca),
	.w4(32'h3b34c322),
	.w5(32'h3a53e6a4),
	.w6(32'h3b1b1d8b),
	.w7(32'h3a4bbcca),
	.w8(32'h39abd77d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd5443),
	.w1(32'h3a5d34b4),
	.w2(32'h3adf9f95),
	.w3(32'h3a2cc751),
	.w4(32'h3aa2767b),
	.w5(32'h3b2370db),
	.w6(32'h3a56a628),
	.w7(32'h3aaf52f3),
	.w8(32'h3b1e002d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11fc4e),
	.w1(32'hbb8c265d),
	.w2(32'h3a2e6004),
	.w3(32'hba1405e4),
	.w4(32'hb97fa233),
	.w5(32'h3b6f5649),
	.w6(32'h3a7f3027),
	.w7(32'h3a41d7c6),
	.w8(32'h3bbfd0f2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7682873),
	.w1(32'h37312c32),
	.w2(32'hb76516c8),
	.w3(32'hb6b948de),
	.w4(32'h37d54945),
	.w5(32'h36a8896e),
	.w6(32'hb7bd8b4c),
	.w7(32'h36fd61fd),
	.w8(32'hb72860c7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4975b5),
	.w1(32'h3b4aaae6),
	.w2(32'h3a7ee197),
	.w3(32'h3bc7d18e),
	.w4(32'h3bbbede4),
	.w5(32'h3b417295),
	.w6(32'h3ba0b01a),
	.w7(32'h3b3693bb),
	.w8(32'h3a1d3354),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71ada7),
	.w1(32'h3b2e310b),
	.w2(32'h3b2f0f34),
	.w3(32'h3b39af49),
	.w4(32'h3b915f63),
	.w5(32'h3a4ebe8a),
	.w6(32'h3b00cdc9),
	.w7(32'h3b84b699),
	.w8(32'h3b107ddc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00f057),
	.w1(32'h3b3ae17e),
	.w2(32'h37350e6e),
	.w3(32'h3ad1ed96),
	.w4(32'h3ad0fee6),
	.w5(32'hbaefa341),
	.w6(32'hba2f2e5e),
	.w7(32'hba81adac),
	.w8(32'hbb6d8db6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a737844),
	.w1(32'h3adc1ec9),
	.w2(32'hbb7e464c),
	.w3(32'h3b0569c6),
	.w4(32'h3b860b08),
	.w5(32'hbaab019f),
	.w6(32'h39c2ccea),
	.w7(32'h3b1c8c31),
	.w8(32'hbae14cb6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06ca24),
	.w1(32'h3b4909f8),
	.w2(32'h3ad7c0d7),
	.w3(32'h39bc53fb),
	.w4(32'h3ad98f54),
	.w5(32'h3a9abfbb),
	.w6(32'hbade3110),
	.w7(32'hbb25eeca),
	.w8(32'hbb1a51b6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9121e6d),
	.w1(32'h3a016586),
	.w2(32'h3acc439b),
	.w3(32'h3ad0c2b2),
	.w4(32'h3aba482d),
	.w5(32'h3a3b6d75),
	.w6(32'h3b0f081c),
	.w7(32'h3b05fd82),
	.w8(32'h3ab6af41),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39815393),
	.w1(32'h39f154d4),
	.w2(32'h3984199b),
	.w3(32'h393b95a0),
	.w4(32'h39c589f7),
	.w5(32'h3968616b),
	.w6(32'h37c7b8e7),
	.w7(32'h3949623c),
	.w8(32'h38e016ef),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377c077e),
	.w1(32'h3807c649),
	.w2(32'h37992a4b),
	.w3(32'h380bfcc6),
	.w4(32'h386fcace),
	.w5(32'h37ddb61f),
	.w6(32'h37842baf),
	.w7(32'h383a9a95),
	.w8(32'h3799df4c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397faf6e),
	.w1(32'h399dd41f),
	.w2(32'h39728d90),
	.w3(32'h395725a7),
	.w4(32'h39827dea),
	.w5(32'h3948cc92),
	.w6(32'h3932d003),
	.w7(32'h397f3de9),
	.w8(32'h396e7030),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ab4c4),
	.w1(32'h3aa218ed),
	.w2(32'h36858f48),
	.w3(32'h39e00499),
	.w4(32'h3af76b66),
	.w5(32'h39198fee),
	.w6(32'h3acd3e71),
	.w7(32'h3b3f6c13),
	.w8(32'h3b13ba41),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a859406),
	.w1(32'hb9a09ccc),
	.w2(32'hbab49719),
	.w3(32'h3ab81899),
	.w4(32'hb9cae28b),
	.w5(32'hba9bf54c),
	.w6(32'h3a392bed),
	.w7(32'hbafeae34),
	.w8(32'hbb657e53),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f9f64),
	.w1(32'h3bf472b4),
	.w2(32'hbc859dc0),
	.w3(32'h3c1eefd4),
	.w4(32'h3c343352),
	.w5(32'hbba4a172),
	.w6(32'hbbcbc2a9),
	.w7(32'hbb941dea),
	.w8(32'hbc94bc7e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c63d4),
	.w1(32'h3ba1b80f),
	.w2(32'h3bb2a110),
	.w3(32'hba90870b),
	.w4(32'hba337e88),
	.w5(32'h3b8be21d),
	.w6(32'hbb16621d),
	.w7(32'hba82356b),
	.w8(32'h3810b7ce),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad039dc),
	.w1(32'h3b6a508f),
	.w2(32'h3b6b8c2d),
	.w3(32'hbb3a0a48),
	.w4(32'h3af65df9),
	.w5(32'h3ba91a2f),
	.w6(32'hbb960f1c),
	.w7(32'hb9e54184),
	.w8(32'h3b9a53f0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90233dc),
	.w1(32'hba9dfb8f),
	.w2(32'h3b4a6f67),
	.w3(32'h3aa9199e),
	.w4(32'h3a3f2c15),
	.w5(32'h3b7650fd),
	.w6(32'h3b264843),
	.w7(32'h3a81e432),
	.w8(32'h3b30abb0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dc84c),
	.w1(32'h3be82b5a),
	.w2(32'hbbbb1760),
	.w3(32'hbadd1003),
	.w4(32'h3befacb2),
	.w5(32'hbabedf5a),
	.w6(32'hbb32b240),
	.w7(32'h3b7fad44),
	.w8(32'hbb9997de),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06ffb6),
	.w1(32'h3a012ee5),
	.w2(32'h3aa0afd9),
	.w3(32'hbaf7b699),
	.w4(32'hba86f2e8),
	.w5(32'hba8c4b72),
	.w6(32'hba0e5a56),
	.w7(32'h3aa48f15),
	.w8(32'h3abf718a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e1a76),
	.w1(32'h3ab67417),
	.w2(32'h3abae763),
	.w3(32'h39fcebc5),
	.w4(32'h3aa29017),
	.w5(32'h3a8e7b20),
	.w6(32'h3a9b610a),
	.w7(32'h3aa6e39b),
	.w8(32'h3ad39d0d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb472ff9),
	.w1(32'h3b6b9948),
	.w2(32'h3a748a3f),
	.w3(32'h3a577ec1),
	.w4(32'h3ba6e479),
	.w5(32'h3ba7e7cc),
	.w6(32'hba9b258f),
	.w7(32'h3b6d881a),
	.w8(32'h3b406137),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994df72),
	.w1(32'hb9a4cb95),
	.w2(32'hb9ee9656),
	.w3(32'hb9734caf),
	.w4(32'hb9508b97),
	.w5(32'hb9ae1f21),
	.w6(32'hb9673658),
	.w7(32'hb9391962),
	.w8(32'hb9ae5e17),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d28de5d),
	.w1(32'h3d4c2cc2),
	.w2(32'h3d1beb58),
	.w3(32'h3cee7cb0),
	.w4(32'h3d0ff347),
	.w5(32'h3d56da0c),
	.w6(32'h3cf43be4),
	.w7(32'h3c15d98a),
	.w8(32'h3ce39217),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a209b0),
	.w1(32'h3b04d556),
	.w2(32'hb96753bf),
	.w3(32'h3b210206),
	.w4(32'h3b554dee),
	.w5(32'h3a72cb29),
	.w6(32'hba53120b),
	.w7(32'h37c55662),
	.w8(32'hba56e6a3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9549851),
	.w1(32'h39cd3f52),
	.w2(32'h3ad70d37),
	.w3(32'h3a4aba9b),
	.w4(32'h3abdbca4),
	.w5(32'h3af96837),
	.w6(32'h3a3a4117),
	.w7(32'h3a8ee55b),
	.w8(32'h3b029772),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0437d0),
	.w1(32'hbae4fc82),
	.w2(32'hbabe5784),
	.w3(32'hbad8a24f),
	.w4(32'hba741db8),
	.w5(32'hba4d6d38),
	.w6(32'hbb09f3bf),
	.w7(32'hbadc6bc5),
	.w8(32'hba5d0859),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aaf0c),
	.w1(32'hb9cfe373),
	.w2(32'h3b27664d),
	.w3(32'hbb2a9b82),
	.w4(32'hba7a4e98),
	.w5(32'h3b436f76),
	.w6(32'hba57640a),
	.w7(32'h3986ea50),
	.w8(32'h3b4e91db),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3864806a),
	.w1(32'h382c8f15),
	.w2(32'hb81a504a),
	.w3(32'h37cff87b),
	.w4(32'h379cb23e),
	.w5(32'hb85216f3),
	.w6(32'h3641e15b),
	.w7(32'hb6ac4a15),
	.w8(32'hb85e62b5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d51341),
	.w1(32'h380fad03),
	.w2(32'hb790a384),
	.w3(32'h378c9ea4),
	.w4(32'h378f1140),
	.w5(32'hb6182740),
	.w6(32'h35bb715d),
	.w7(32'h36cf0d7a),
	.w8(32'hb7ade962),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20dcb1),
	.w1(32'hbae58070),
	.w2(32'h3a360fbb),
	.w3(32'hbb5a4231),
	.w4(32'hbbbb906f),
	.w5(32'hbb43cfa1),
	.w6(32'hbb0760f0),
	.w7(32'hbb77eaf2),
	.w8(32'hbb22e338),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b443dc3),
	.w1(32'h3b891d10),
	.w2(32'hbac6b2b9),
	.w3(32'h3b51f50e),
	.w4(32'h3b248579),
	.w5(32'h39a402a4),
	.w6(32'h38beaad2),
	.w7(32'hb9838fc4),
	.w8(32'hbb17435b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39697e5b),
	.w1(32'h3950e1c9),
	.w2(32'h38e2ac62),
	.w3(32'h394f1378),
	.w4(32'h3943ceff),
	.w5(32'h38f72eda),
	.w6(32'h3932cca3),
	.w7(32'h3916e18c),
	.w8(32'h3906184c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d8c82),
	.w1(32'hb84c1ba6),
	.w2(32'h3b0f2718),
	.w3(32'h3a526f70),
	.w4(32'h3a96bcdf),
	.w5(32'h3b0eca56),
	.w6(32'h39aff902),
	.w7(32'h3a6a37e4),
	.w8(32'h3afc13bf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c694a),
	.w1(32'h38bb13bd),
	.w2(32'h39685748),
	.w3(32'hb72e1998),
	.w4(32'h3946fbc6),
	.w5(32'h39659df7),
	.w6(32'h382eb1a8),
	.w7(32'h3947e5bb),
	.w8(32'h38e978b1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f14dc3),
	.w1(32'hb9b30068),
	.w2(32'hb9f9679b),
	.w3(32'hb9c8b1e7),
	.w4(32'h390405ce),
	.w5(32'hb9c00b28),
	.w6(32'h379f2be4),
	.w7(32'h39e5294a),
	.w8(32'hb961240a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d673b6),
	.w1(32'h3a84c34c),
	.w2(32'h3afafc54),
	.w3(32'h3bc30e48),
	.w4(32'h3b67067e),
	.w5(32'h3b93f984),
	.w6(32'h3ad6126e),
	.w7(32'hba5dad0a),
	.w8(32'h3b2cd678),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5f4a4),
	.w1(32'h3b1eb8bb),
	.w2(32'h39672a21),
	.w3(32'h3abb6cdb),
	.w4(32'h3aebd95c),
	.w5(32'hb9ae0681),
	.w6(32'h3a8ddf57),
	.w7(32'h3a09ed4e),
	.w8(32'hbb1caa7e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f23d9),
	.w1(32'hba93095e),
	.w2(32'h3a0f1359),
	.w3(32'hba8dfdc8),
	.w4(32'hb9ec1c89),
	.w5(32'hba0cbe6d),
	.w6(32'hbaa339ee),
	.w7(32'hb92ef028),
	.w8(32'h38ffcdeb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5866ee),
	.w1(32'h3a7a685f),
	.w2(32'hb746e2dd),
	.w3(32'hb8f37020),
	.w4(32'h3b208afc),
	.w5(32'h3acffcfb),
	.w6(32'h387b08b6),
	.w7(32'h3a25ef0c),
	.w8(32'h39972151),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f04c1),
	.w1(32'h3bacb584),
	.w2(32'hbb0c845b),
	.w3(32'h3b71fc94),
	.w4(32'h3c01c91b),
	.w5(32'h3add7aae),
	.w6(32'h3991f812),
	.w7(32'h3b0e5c45),
	.w8(32'hbb27aef4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7063c3),
	.w1(32'h3b81c73e),
	.w2(32'h39bc0f9e),
	.w3(32'h3b1ecaa2),
	.w4(32'h3b44b990),
	.w5(32'h3a035ea0),
	.w6(32'h3aa151f5),
	.w7(32'hb91c6e28),
	.w8(32'hbb270445),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb757278b),
	.w1(32'hb7a5039a),
	.w2(32'hba75e4af),
	.w3(32'h39ba1ddb),
	.w4(32'h398edf4f),
	.w5(32'hba68a6e3),
	.w6(32'h3aa5e666),
	.w7(32'h3a3afd88),
	.w8(32'hb9e193b8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390365f3),
	.w1(32'h3c06c494),
	.w2(32'h3b16bb90),
	.w3(32'h3b2b0030),
	.w4(32'h3bf3c36f),
	.w5(32'h3b931854),
	.w6(32'h3a6472b7),
	.w7(32'h3b419473),
	.w8(32'h3a6cc126),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c96c4),
	.w1(32'hb914689c),
	.w2(32'hba85abb0),
	.w3(32'h3a943880),
	.w4(32'h39944311),
	.w5(32'h39311cb6),
	.w6(32'h39d72148),
	.w7(32'hb9a20e2b),
	.w8(32'hba591957),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e90a6),
	.w1(32'h392ec98b),
	.w2(32'hbb402544),
	.w3(32'h3ab5a9e4),
	.w4(32'h3b2aa77b),
	.w5(32'hba80446a),
	.w6(32'h398fe589),
	.w7(32'hb92b8679),
	.w8(32'hbb0a79b2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe47be0),
	.w1(32'hbb07caf7),
	.w2(32'h3bf67754),
	.w3(32'hbb51d87f),
	.w4(32'hb978c58a),
	.w5(32'h3c0e5ce7),
	.w6(32'hbb773e32),
	.w7(32'hbadf8d76),
	.w8(32'h3bc2eebb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba05437),
	.w1(32'hba9ea882),
	.w2(32'hbbfbf543),
	.w3(32'h3c0f785d),
	.w4(32'h3c1cf094),
	.w5(32'h388a5977),
	.w6(32'hbb31696d),
	.w7(32'h3a8273c0),
	.w8(32'hbbbeb7df),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e3d4a),
	.w1(32'h3a8b0c5c),
	.w2(32'hbb48851d),
	.w3(32'h3b9b6d7e),
	.w4(32'h3b3b6e5d),
	.w5(32'hbaa2b6d7),
	.w6(32'hba5cb209),
	.w7(32'h3b08cc34),
	.w8(32'h3aa81dbe),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5e9a2),
	.w1(32'h3ba66bd9),
	.w2(32'h3a5e50c9),
	.w3(32'h3abbdfea),
	.w4(32'h3a6dfc99),
	.w5(32'hbb3c0517),
	.w6(32'hbad0ba2b),
	.w7(32'hbaa00d8c),
	.w8(32'hbbc435c9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abc941),
	.w1(32'hb99fe3b9),
	.w2(32'hbb02df46),
	.w3(32'h39e5d665),
	.w4(32'hb9db02f2),
	.w5(32'hbad5d3e2),
	.w6(32'h3a6b75f9),
	.w7(32'hb99dbba9),
	.w8(32'h3a75d86a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f794),
	.w1(32'h3c2b4925),
	.w2(32'h3b838ddc),
	.w3(32'h3b21e8fd),
	.w4(32'h3bb82851),
	.w5(32'h3b88f9c0),
	.w6(32'h3b9478f6),
	.w7(32'h3b6c7765),
	.w8(32'hbb8f4487),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8fa8c),
	.w1(32'hb9beca67),
	.w2(32'hbaa5aa61),
	.w3(32'hba565211),
	.w4(32'hbaa33bf3),
	.w5(32'hbb8d918f),
	.w6(32'hb9e21ae4),
	.w7(32'h3a181036),
	.w8(32'hbaf899e9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa814f0),
	.w1(32'h395b04ab),
	.w2(32'hbbd8b095),
	.w3(32'h3baa6d41),
	.w4(32'h3b505e38),
	.w5(32'hbb3de8ff),
	.w6(32'h3b3dbb8a),
	.w7(32'hba4c0072),
	.w8(32'hbb16716a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a110a9c),
	.w1(32'h3b5eddd7),
	.w2(32'h3a9d52fe),
	.w3(32'h3ac69cfa),
	.w4(32'h3babac73),
	.w5(32'h3b4ce759),
	.w6(32'h3b2a4081),
	.w7(32'h3bae001d),
	.w8(32'h3b4330fe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02558d),
	.w1(32'h3b188392),
	.w2(32'h3a8f9a43),
	.w3(32'h3b245c6c),
	.w4(32'h3a997d7a),
	.w5(32'h3a786635),
	.w6(32'h3b473afe),
	.w7(32'h3b1bfe3b),
	.w8(32'h3abaea09),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc9d63),
	.w1(32'hba971111),
	.w2(32'h3a804df2),
	.w3(32'hb9044a1e),
	.w4(32'h3ab89508),
	.w5(32'h399d31f1),
	.w6(32'hb907e8eb),
	.w7(32'h39da0f49),
	.w8(32'h398340bf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e12e2),
	.w1(32'hb9a75f6e),
	.w2(32'hba1d74ff),
	.w3(32'hb8f02884),
	.w4(32'h39c8be4f),
	.w5(32'hb98aa2f5),
	.w6(32'h37ffe7d6),
	.w7(32'hb95d2690),
	.w8(32'h3abbc8c3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47d451),
	.w1(32'h3bbd39cc),
	.w2(32'h3b225608),
	.w3(32'h3bac4fac),
	.w4(32'h3bbeb560),
	.w5(32'h3b630ed4),
	.w6(32'h3b05c844),
	.w7(32'h3b1f89f5),
	.w8(32'hba4ae0e7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1177e6),
	.w1(32'h3b1ab85a),
	.w2(32'h3a1feac5),
	.w3(32'h3aec0e30),
	.w4(32'h3baa8b73),
	.w5(32'h3b726813),
	.w6(32'h3aab9427),
	.w7(32'h3aca06e2),
	.w8(32'h3811299d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba901a9f),
	.w1(32'h38b7d502),
	.w2(32'h3a305225),
	.w3(32'hba9f24d2),
	.w4(32'h3a960aa0),
	.w5(32'h3acf479c),
	.w6(32'hb9ab4e73),
	.w7(32'h3ab0b159),
	.w8(32'h3aadbb85),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac907cd),
	.w1(32'h3a7db8ca),
	.w2(32'hba47f62c),
	.w3(32'h3b0701d1),
	.w4(32'h3b12d708),
	.w5(32'h3aa3c68c),
	.w6(32'h3a7d9a24),
	.w7(32'h3aa32135),
	.w8(32'h396eb32a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d205e),
	.w1(32'hba64e079),
	.w2(32'h3ad02b0c),
	.w3(32'h3a0f8cfa),
	.w4(32'h3b59eece),
	.w5(32'h3b6f857d),
	.w6(32'h3a893d39),
	.w7(32'h3b5aa84f),
	.w8(32'h3a90820b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7725e6),
	.w1(32'h3ad6c5c1),
	.w2(32'h39defec4),
	.w3(32'h3a828b6d),
	.w4(32'h3a1e47e0),
	.w5(32'h3a66f083),
	.w6(32'hbaa5b0ec),
	.w7(32'hbb060917),
	.w8(32'hba85e121),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d0e504),
	.w1(32'hb951c228),
	.w2(32'h3905fe98),
	.w3(32'hb9314910),
	.w4(32'hb8c142fa),
	.w5(32'h397b7f83),
	.w6(32'hb7a6fa62),
	.w7(32'h3871572d),
	.w8(32'h3a72680a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2121e6),
	.w1(32'h3c3444f9),
	.w2(32'h3a49e7c4),
	.w3(32'h3b981c14),
	.w4(32'h3c506b33),
	.w5(32'h3bc57a89),
	.w6(32'h3b9a56e5),
	.w7(32'h3c497d0d),
	.w8(32'h3b690fad),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9673669),
	.w1(32'hb878b876),
	.w2(32'h388a00d2),
	.w3(32'hba230728),
	.w4(32'hb98e0ee2),
	.w5(32'h38c40000),
	.w6(32'hb9c55bd0),
	.w7(32'hb9ad597a),
	.w8(32'hb97a11e4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d4151),
	.w1(32'h3a3d06df),
	.w2(32'h3b01900a),
	.w3(32'hbad99c96),
	.w4(32'hb7901740),
	.w5(32'h3ac9bb39),
	.w6(32'h3afdcd59),
	.w7(32'h3b6ef48f),
	.w8(32'h3b861fe0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3fe38),
	.w1(32'h39a71d55),
	.w2(32'h399459a0),
	.w3(32'h39b2ee7b),
	.w4(32'h39a29a74),
	.w5(32'h3a1cbba2),
	.w6(32'h39f947fd),
	.w7(32'h39a91560),
	.w8(32'hba9311e7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e576a4),
	.w1(32'h3b3f7a2e),
	.w2(32'h36846910),
	.w3(32'h3abda6f5),
	.w4(32'h3a99cd37),
	.w5(32'hb96d6c5d),
	.w6(32'hbaa96e1b),
	.w7(32'hbb903edb),
	.w8(32'hba3278f6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c03ccd),
	.w1(32'hba17ba7b),
	.w2(32'hb9d0c9c0),
	.w3(32'hb9d30ce6),
	.w4(32'hb9f4ca2d),
	.w5(32'hb9eb3f3a),
	.w6(32'hba38cd3d),
	.w7(32'hba2602b1),
	.w8(32'h391b5154),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae258fb),
	.w1(32'h3a370455),
	.w2(32'hb9df821c),
	.w3(32'h3b06696b),
	.w4(32'h3b07dbf3),
	.w5(32'h397b8f47),
	.w6(32'h3a4a5555),
	.w7(32'h3b5350f5),
	.w8(32'h3b3af445),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a231b),
	.w1(32'hb911b95d),
	.w2(32'hb7b3eb33),
	.w3(32'hb954a02b),
	.w4(32'hb8d9678e),
	.w5(32'hb5cc74d7),
	.w6(32'hb97867aa),
	.w7(32'hb99f1cb5),
	.w8(32'h3a5dfe3d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42ba4a),
	.w1(32'h3bcece98),
	.w2(32'hb9542685),
	.w3(32'h3b9d0844),
	.w4(32'h3be26f84),
	.w5(32'h3b289642),
	.w6(32'h3b5fd042),
	.w7(32'h3bb1f98c),
	.w8(32'hb9cf5c26),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801d48),
	.w1(32'h3ba56f9d),
	.w2(32'h3aa11f9e),
	.w3(32'h3b73fa0d),
	.w4(32'h3b10a868),
	.w5(32'h3a471f45),
	.w6(32'h3ac40fb2),
	.w7(32'h3997154a),
	.w8(32'hbb4c9a1b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b9659),
	.w1(32'h38bf2c69),
	.w2(32'h38178728),
	.w3(32'hb9b542c2),
	.w4(32'hb80f4574),
	.w5(32'hb8ac1f43),
	.w6(32'hb8279b47),
	.w7(32'hb90cb605),
	.w8(32'hba13bb7b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ad903),
	.w1(32'hbaa8ab3d),
	.w2(32'hba8f27c0),
	.w3(32'hba02964a),
	.w4(32'hba1e43d2),
	.w5(32'hbafea038),
	.w6(32'h3820b8f6),
	.w7(32'h3a2a0cf9),
	.w8(32'hb8bd7ecb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ecddd2),
	.w1(32'hba817eb1),
	.w2(32'hba7b2fc6),
	.w3(32'hb9d807cb),
	.w4(32'h3a1201e1),
	.w5(32'hb9863898),
	.w6(32'h3b260565),
	.w7(32'h3b717d61),
	.w8(32'h3b497fd5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387431a0),
	.w1(32'h3b6a7f47),
	.w2(32'h3a7d1119),
	.w3(32'h3b685437),
	.w4(32'h3bd40a4f),
	.w5(32'h3b91ad2e),
	.w6(32'h3a93f26f),
	.w7(32'h3b37c9bb),
	.w8(32'h3a8181a8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c59b3),
	.w1(32'h3ba3f143),
	.w2(32'h3b80c96c),
	.w3(32'h3c50f6ed),
	.w4(32'h3a74c242),
	.w5(32'h3b8a3411),
	.w6(32'h3b092e55),
	.w7(32'hbb89f19c),
	.w8(32'h3ac8dd03),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b306faa),
	.w1(32'h3c28077e),
	.w2(32'h3ab8ffe7),
	.w3(32'h3c0ef1ec),
	.w4(32'h3c6bfdf5),
	.w5(32'h3c03b99f),
	.w6(32'h3adee517),
	.w7(32'h3b9312cf),
	.w8(32'hba2c1b51),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a378c53),
	.w1(32'h3a99476b),
	.w2(32'hbb092e65),
	.w3(32'h3af571bc),
	.w4(32'h3b7f6667),
	.w5(32'hbaae9a5e),
	.w6(32'h3a2ba470),
	.w7(32'h3b748f72),
	.w8(32'hb9ec726b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db55a2),
	.w1(32'hb9c1b98b),
	.w2(32'hb9840d29),
	.w3(32'h39cb173c),
	.w4(32'hb91c481c),
	.w5(32'h39df93ac),
	.w6(32'hb90f9395),
	.w7(32'hb9522620),
	.w8(32'hb9ea845b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec9d26),
	.w1(32'hb99a41a3),
	.w2(32'h3984c2fc),
	.w3(32'hb9986aac),
	.w4(32'hb94f1933),
	.w5(32'h3705ca18),
	.w6(32'hb9a605f2),
	.w7(32'hb8eb08e8),
	.w8(32'hb957101e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b93a6),
	.w1(32'h3ad80b4a),
	.w2(32'h39b895d1),
	.w3(32'h3a812bf3),
	.w4(32'h3a9fd6ed),
	.w5(32'h3a15c300),
	.w6(32'h39814d39),
	.w7(32'hba1521b1),
	.w8(32'h3a075709),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac60005),
	.w1(32'h3b4afca5),
	.w2(32'h3b10db41),
	.w3(32'h3b4577b1),
	.w4(32'h3b60eb00),
	.w5(32'h3b1354e0),
	.w6(32'h3ab3c152),
	.w7(32'h3b531e8d),
	.w8(32'h3b139ecb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea225c),
	.w1(32'h3b130941),
	.w2(32'h3a9e41ef),
	.w3(32'h3b3b8903),
	.w4(32'h3b4b04c5),
	.w5(32'h3b19015c),
	.w6(32'h3b0741c6),
	.w7(32'h3b470d64),
	.w8(32'h3b3439ae),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba626627),
	.w1(32'hb974adef),
	.w2(32'hb9998066),
	.w3(32'hba906798),
	.w4(32'hb8508a18),
	.w5(32'h3883c97f),
	.w6(32'hbac02223),
	.w7(32'hb9f7b985),
	.w8(32'hbaa97bcb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c704),
	.w1(32'hbab9beb8),
	.w2(32'hbada44d1),
	.w3(32'hba96bf05),
	.w4(32'hba8901dd),
	.w5(32'hbb9a6b7f),
	.w6(32'h3a9cbb43),
	.w7(32'h3a055e04),
	.w8(32'h3a81bfe6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba634cb9),
	.w1(32'h3a85663a),
	.w2(32'h383ff489),
	.w3(32'h3928629f),
	.w4(32'h3acea89c),
	.w5(32'h39c3b165),
	.w6(32'hba749bb0),
	.w7(32'h3784eddc),
	.w8(32'hba0d2828),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdf0a9),
	.w1(32'h3aa72c8b),
	.w2(32'h3afb64e8),
	.w3(32'h3b00ab9b),
	.w4(32'h3acd0d42),
	.w5(32'h3abdb680),
	.w6(32'h3a780b73),
	.w7(32'h3a836254),
	.w8(32'h3adb37a6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25fae0),
	.w1(32'h3addc373),
	.w2(32'hba711a28),
	.w3(32'hbb1b7ede),
	.w4(32'h3a9c921f),
	.w5(32'h39d236aa),
	.w6(32'hbb8a90d1),
	.w7(32'hbabfa433),
	.w8(32'hbb04eee4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c9b77),
	.w1(32'h3bfcab79),
	.w2(32'h3bb08705),
	.w3(32'h3ba99c6b),
	.w4(32'h3be81ff4),
	.w5(32'h3b43c34e),
	.w6(32'h3a853efe),
	.w7(32'h3b90f713),
	.w8(32'h3b0d6119),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bf793),
	.w1(32'h39702862),
	.w2(32'hbaa5a0a7),
	.w3(32'hb86e6277),
	.w4(32'hba6b6066),
	.w5(32'h38280cb7),
	.w6(32'h3ac07865),
	.w7(32'h3a962f63),
	.w8(32'h3a3b376a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39811416),
	.w1(32'h3a11f79e),
	.w2(32'h3a9303e1),
	.w3(32'hb92442cc),
	.w4(32'h39876e91),
	.w5(32'h393f222c),
	.w6(32'h3a801f87),
	.w7(32'h3ae6fbe9),
	.w8(32'hb7d8b332),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95eb03d),
	.w1(32'hb92263eb),
	.w2(32'h3994eab3),
	.w3(32'hb9ada3e6),
	.w4(32'h38356145),
	.w5(32'h3957e908),
	.w6(32'hb62d6230),
	.w7(32'h38882e83),
	.w8(32'h396dc008),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af321e),
	.w1(32'h39aab230),
	.w2(32'hb9ccfede),
	.w3(32'h3a0d595d),
	.w4(32'h396f3f35),
	.w5(32'hb98d48f9),
	.w6(32'hb78d97b8),
	.w7(32'hba144b2a),
	.w8(32'h39b0d05d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ece4d7),
	.w1(32'h38f580a9),
	.w2(32'h3a2da51a),
	.w3(32'h378f1f48),
	.w4(32'h3a9b4f2f),
	.w5(32'h3ac494c9),
	.w6(32'h3a19fae5),
	.w7(32'h3ac19141),
	.w8(32'h3ab77c69),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dbe54),
	.w1(32'h3ae80fce),
	.w2(32'h3aae3a89),
	.w3(32'h39c62d99),
	.w4(32'h3a8cb914),
	.w5(32'h396cae16),
	.w6(32'h3b12f2d2),
	.w7(32'h3b1d638e),
	.w8(32'h39b7ba2d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c456c),
	.w1(32'hbb0a437c),
	.w2(32'hba7d2a53),
	.w3(32'hba8f7580),
	.w4(32'hbb51065e),
	.w5(32'hbb5304c9),
	.w6(32'h3a6662ab),
	.w7(32'hba22bdcf),
	.w8(32'hba451674),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba178193),
	.w1(32'hbab66e09),
	.w2(32'hba0b63dd),
	.w3(32'hba8db176),
	.w4(32'hbaff4a09),
	.w5(32'hba555556),
	.w6(32'h388f7517),
	.w7(32'hba6dbb5e),
	.w8(32'hba82ce1f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb347cb7),
	.w1(32'h3af8f47e),
	.w2(32'h3a4632be),
	.w3(32'h3b2fe467),
	.w4(32'h3bc2332c),
	.w5(32'hbba5c0df),
	.w6(32'h3b99b11e),
	.w7(32'h3c30442d),
	.w8(32'h3a3941fe),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2925e5),
	.w1(32'h3c2ea1ee),
	.w2(32'h3c8e2ecf),
	.w3(32'hbb9116b9),
	.w4(32'hbc4d33cb),
	.w5(32'h3bbd18da),
	.w6(32'hb8c17536),
	.w7(32'hbc542658),
	.w8(32'hbaf657de),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd757f8),
	.w1(32'hbab6dc6b),
	.w2(32'h3b79220c),
	.w3(32'h3a385051),
	.w4(32'h3b11b048),
	.w5(32'hbb47c2a4),
	.w6(32'hbb65b300),
	.w7(32'h3b685abf),
	.w8(32'hbabf3d36),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813023),
	.w1(32'hb9acdb61),
	.w2(32'h3a85ee74),
	.w3(32'hbb2383e0),
	.w4(32'hbb414a40),
	.w5(32'hbbb9e9ae),
	.w6(32'hbb545c69),
	.w7(32'hb9ea1dd0),
	.w8(32'h3b4bcb0e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57e4ef),
	.w1(32'hba9adaa0),
	.w2(32'hbb4f7855),
	.w3(32'hba2ab0d6),
	.w4(32'h3ab9959d),
	.w5(32'hbb2c9bd4),
	.w6(32'h3b36b51c),
	.w7(32'h3b0ef744),
	.w8(32'hbcb55bad),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2317b8),
	.w1(32'hbb2f85a6),
	.w2(32'hbc3f7ac6),
	.w3(32'hbc55bf67),
	.w4(32'hbbba7d84),
	.w5(32'h3be1d430),
	.w6(32'hbc5b581f),
	.w7(32'hbc8078df),
	.w8(32'hbc32b206),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6f0ed),
	.w1(32'h3a75b13b),
	.w2(32'h3c06159d),
	.w3(32'hba0686c8),
	.w4(32'h3b9cc686),
	.w5(32'h3b1ae716),
	.w6(32'hbc22932d),
	.w7(32'hbb1918e4),
	.w8(32'h3c99b7ae),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc57d3c),
	.w1(32'hbc0aca95),
	.w2(32'hbcc78848),
	.w3(32'h3b311837),
	.w4(32'hbca848b1),
	.w5(32'hbcb7688a),
	.w6(32'h3c21c009),
	.w7(32'hbbb9fb2d),
	.w8(32'hbb79d913),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1be2b),
	.w1(32'hbb934420),
	.w2(32'hba0a5cbf),
	.w3(32'hbb3bfc5f),
	.w4(32'hbad3c1d7),
	.w5(32'hbbb76ba4),
	.w6(32'hbb7f5551),
	.w7(32'h39553903),
	.w8(32'hbb109bd1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ae432),
	.w1(32'h3b028732),
	.w2(32'h3b692bf7),
	.w3(32'h3afbc83d),
	.w4(32'h3babb981),
	.w5(32'h3b241a3e),
	.w6(32'h3a8aaab6),
	.w7(32'h3b30f732),
	.w8(32'hbbb19596),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd732c9),
	.w1(32'h3bdc5f4e),
	.w2(32'h3c03c7ed),
	.w3(32'h3a664efd),
	.w4(32'h3c0e11e3),
	.w5(32'h3a1b94fe),
	.w6(32'h3a814764),
	.w7(32'h3b9bcca0),
	.w8(32'hbc1974c4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f5959),
	.w1(32'h3c8b4ef6),
	.w2(32'hbc8ee052),
	.w3(32'h3a892631),
	.w4(32'h3bc0df38),
	.w5(32'hbc94799b),
	.w6(32'h3c93787a),
	.w7(32'hbb75794e),
	.w8(32'h3c40d2f3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c536669),
	.w1(32'hbb8556df),
	.w2(32'hbc2efea8),
	.w3(32'h3c088692),
	.w4(32'hbb49b666),
	.w5(32'hbbcfaecf),
	.w6(32'h3c1ec6da),
	.w7(32'h3b8a460a),
	.w8(32'hbba4a31a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e682),
	.w1(32'hbbed3c47),
	.w2(32'h3b85fb48),
	.w3(32'hbc953d96),
	.w4(32'hbc02933a),
	.w5(32'h3c05fc7c),
	.w6(32'hbc32cfef),
	.w7(32'hbc7f0fb9),
	.w8(32'h3c4bbc70),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cb39d),
	.w1(32'hbbfc53db),
	.w2(32'h389dbe62),
	.w3(32'h3b1fcc10),
	.w4(32'hbc063d3b),
	.w5(32'h3ace0c96),
	.w6(32'h3abcafb5),
	.w7(32'hbb61039c),
	.w8(32'hbabe9076),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47857c),
	.w1(32'hbc005337),
	.w2(32'hbc4e56c7),
	.w3(32'hbc3061b0),
	.w4(32'hbc93eaf6),
	.w5(32'hbc23544b),
	.w6(32'hbcac2d5f),
	.w7(32'hbc5d7054),
	.w8(32'h3b1c31e5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06ebf3),
	.w1(32'hba177306),
	.w2(32'h3cfb76bc),
	.w3(32'hba9d5731),
	.w4(32'h3accc6d8),
	.w5(32'h3c815b51),
	.w6(32'hbc7e80a3),
	.w7(32'hbbd25300),
	.w8(32'hbaeadd36),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ab46b),
	.w1(32'h3a7e925e),
	.w2(32'h3b209971),
	.w3(32'h39d2af02),
	.w4(32'hbb57a778),
	.w5(32'hbbf13f82),
	.w6(32'hbbc81470),
	.w7(32'hbb94d113),
	.w8(32'hbbe63388),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb15dd),
	.w1(32'h3ac10206),
	.w2(32'hb8dd53ab),
	.w3(32'hbc1a2412),
	.w4(32'hbbd3834f),
	.w5(32'h3ba67cd5),
	.w6(32'hbbf6c90b),
	.w7(32'hbb6fa241),
	.w8(32'hbc830937),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb9ad9),
	.w1(32'h3b53ad10),
	.w2(32'hbc0900be),
	.w3(32'hbc4febf7),
	.w4(32'hbc1a7f2e),
	.w5(32'hbbc5a2a8),
	.w6(32'hbcafa0aa),
	.w7(32'hbb89bf07),
	.w8(32'hbaee2cf1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc982e2a),
	.w1(32'h3abf1545),
	.w2(32'h3b92f9a0),
	.w3(32'hbc149d63),
	.w4(32'hbbc2303b),
	.w5(32'hbbeaaf69),
	.w6(32'hbbaeee24),
	.w7(32'h3ab0aa30),
	.w8(32'hbb31e197),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2097b8),
	.w1(32'hbb53c730),
	.w2(32'h3be3250e),
	.w3(32'h3b208738),
	.w4(32'h3afcec41),
	.w5(32'h3acb9fca),
	.w6(32'h3a177e52),
	.w7(32'h3bf0d27d),
	.w8(32'h3c2c91e3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd28e5f),
	.w1(32'h3bed7451),
	.w2(32'h3c83b5f6),
	.w3(32'h3bd8bbb3),
	.w4(32'hbc1aa1c0),
	.w5(32'hbc5018ac),
	.w6(32'h3c014703),
	.w7(32'h3bc67d9d),
	.w8(32'h3aba11ea),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule