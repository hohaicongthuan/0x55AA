module layer_10_featuremap_23(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f5b06),
	.w1(32'h3b5aed29),
	.w2(32'h3d17da32),
	.w3(32'h3b6d7d51),
	.w4(32'h3c17cfed),
	.w5(32'h3cb1ab48),
	.w6(32'h3ad5ee2f),
	.w7(32'h3c38780d),
	.w8(32'hbc64e2e0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cce2385),
	.w1(32'h3c2e2222),
	.w2(32'hbc7a5799),
	.w3(32'h3cddc482),
	.w4(32'h3d1261cc),
	.w5(32'h3c579103),
	.w6(32'hbc34016c),
	.w7(32'h3bdde658),
	.w8(32'h3b95d722),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2e362f),
	.w1(32'hbd021aa3),
	.w2(32'h3b4fd143),
	.w3(32'h3bf64178),
	.w4(32'h3c254445),
	.w5(32'h38e343d5),
	.w6(32'h3c6d6c5d),
	.w7(32'h3cbe5a6c),
	.w8(32'hb8a23720),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99c26a),
	.w1(32'hbad609ce),
	.w2(32'hbc7ff7b3),
	.w3(32'h3c1f42af),
	.w4(32'h3adcec26),
	.w5(32'hbc3156e0),
	.w6(32'hba5ce547),
	.w7(32'h3b12d961),
	.w8(32'hbc1e0db6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a98b8),
	.w1(32'hbaa69bea),
	.w2(32'h3b267a5c),
	.w3(32'hbc17b2ad),
	.w4(32'hbb9a89f8),
	.w5(32'hbc6ae9dc),
	.w6(32'hbc29fbd2),
	.w7(32'hbc26a719),
	.w8(32'hbc1f85b9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecdca5),
	.w1(32'hbc346c24),
	.w2(32'hbb680c58),
	.w3(32'hbc30729f),
	.w4(32'h3b235d74),
	.w5(32'hbbb6268b),
	.w6(32'hbb926ba7),
	.w7(32'h3b0fb9c5),
	.w8(32'hbb3726a0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932ba0a),
	.w1(32'hba72138c),
	.w2(32'hbc54cf28),
	.w3(32'hbc0e68a7),
	.w4(32'hbc0af3bf),
	.w5(32'hbc3f3075),
	.w6(32'hbc0b8657),
	.w7(32'hbbb76f46),
	.w8(32'h3b076468),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a43f2),
	.w1(32'hbccc9282),
	.w2(32'hbcbf6b9f),
	.w3(32'hbcc7470b),
	.w4(32'hbc9fd432),
	.w5(32'hbc1f6844),
	.w6(32'hbc563f4e),
	.w7(32'hbcbc9222),
	.w8(32'hbb03327f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53f791),
	.w1(32'hbad4037b),
	.w2(32'h3afbd66b),
	.w3(32'hbc8b4a53),
	.w4(32'hbbbf7d26),
	.w5(32'hbba3403c),
	.w6(32'h3be68979),
	.w7(32'h3af0417b),
	.w8(32'hb9266a67),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe1ffc),
	.w1(32'h3ba34a05),
	.w2(32'hbc2ef797),
	.w3(32'h3a7f1b8f),
	.w4(32'hbbbd5200),
	.w5(32'hbbf2dc4d),
	.w6(32'hbc9075da),
	.w7(32'hbc722858),
	.w8(32'hbc8c0506),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b883ac5),
	.w1(32'h3ba3b73b),
	.w2(32'hbae1c440),
	.w3(32'h3b2e37c5),
	.w4(32'h3b9ddde5),
	.w5(32'h3bd92db5),
	.w6(32'hb9ebee50),
	.w7(32'h3aa36cb5),
	.w8(32'hbb847591),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b833e),
	.w1(32'h3b864a31),
	.w2(32'hbc09fc68),
	.w3(32'h3c6e1f6b),
	.w4(32'hbbd05e73),
	.w5(32'hbbfc9f22),
	.w6(32'hbbe1c1e0),
	.w7(32'h3bc89931),
	.w8(32'hbb5d4f0c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba361415),
	.w1(32'hbb961672),
	.w2(32'hbc11c753),
	.w3(32'h3a62b6b1),
	.w4(32'hb92ccaca),
	.w5(32'hbb3caf80),
	.w6(32'hbb9fc194),
	.w7(32'hbb288a34),
	.w8(32'hbc5627f2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be397a9),
	.w1(32'h3bb15972),
	.w2(32'hbcdaf30f),
	.w3(32'h3b2a860f),
	.w4(32'h3ba15220),
	.w5(32'hbc700735),
	.w6(32'h3bd76b7d),
	.w7(32'h3b55b0d7),
	.w8(32'hbc18c295),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc851bc4),
	.w1(32'hbab4e3b7),
	.w2(32'h38c50465),
	.w3(32'hbbfa285c),
	.w4(32'hba977108),
	.w5(32'h3c182229),
	.w6(32'h3b275dcd),
	.w7(32'hbbd9fb64),
	.w8(32'h351de030),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03464),
	.w1(32'h3a836813),
	.w2(32'hbc36265c),
	.w3(32'hb9008669),
	.w4(32'h3c3457b2),
	.w5(32'hba82bce5),
	.w6(32'hbc37b1da),
	.w7(32'hbb2ca81e),
	.w8(32'hbbebe1b7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46267c),
	.w1(32'h3b1d881b),
	.w2(32'hbb9bc6b1),
	.w3(32'h3b873fec),
	.w4(32'h3bc916fc),
	.w5(32'hb84100fb),
	.w6(32'h3b7b778b),
	.w7(32'h3ba5851f),
	.w8(32'h3b695394),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc883c88),
	.w1(32'hbc8ae6e9),
	.w2(32'hbca6e969),
	.w3(32'hbc67ee22),
	.w4(32'hbc05fe21),
	.w5(32'hbb8b991a),
	.w6(32'hbc4cbd39),
	.w7(32'hba65914b),
	.w8(32'hbc6c81de),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0cd90),
	.w1(32'h3b0f89e1),
	.w2(32'hbc83d889),
	.w3(32'h3b915bc6),
	.w4(32'h3ada595f),
	.w5(32'hbc1c1660),
	.w6(32'hbba51fa8),
	.w7(32'hbafde1b8),
	.w8(32'hbbbca956),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84c5d6),
	.w1(32'hbc40ddb1),
	.w2(32'h3940f4a6),
	.w3(32'hbc3c8bfc),
	.w4(32'hbc30659e),
	.w5(32'hbbab6234),
	.w6(32'h3bc1158a),
	.w7(32'hba95c45b),
	.w8(32'h3b2b4652),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db6709),
	.w1(32'hbb7718c4),
	.w2(32'h3ae24546),
	.w3(32'hbc18f582),
	.w4(32'hbc481a29),
	.w5(32'h3c0a203d),
	.w6(32'h3aa5181e),
	.w7(32'hb7e1379c),
	.w8(32'h3a0b4339),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51677c),
	.w1(32'h3c43475b),
	.w2(32'h3a6ba495),
	.w3(32'h3b494302),
	.w4(32'hbb1b59ec),
	.w5(32'h3a217fae),
	.w6(32'h3a31f83c),
	.w7(32'hbad4a0e9),
	.w8(32'h3b333452),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4545f0),
	.w1(32'hbc45e321),
	.w2(32'hbced1fd0),
	.w3(32'hbbf221ab),
	.w4(32'hbc0ea4f5),
	.w5(32'hbc56da29),
	.w6(32'hbced37dd),
	.w7(32'hbc1886ee),
	.w8(32'hbd011b62),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9195b5),
	.w1(32'h39820811),
	.w2(32'hbc11a100),
	.w3(32'h3bb62137),
	.w4(32'h3b7dd54b),
	.w5(32'hbbc3369a),
	.w6(32'hbbc8fc42),
	.w7(32'hbba287d6),
	.w8(32'hbc311fd4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c785b01),
	.w1(32'h3cba2344),
	.w2(32'h3bf7054b),
	.w3(32'h3c7914a8),
	.w4(32'h3c6d06e3),
	.w5(32'h3b8af0ca),
	.w6(32'h3bb4f770),
	.w7(32'h3bd863c0),
	.w8(32'hbb8be331),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bf10c),
	.w1(32'hbb2a3380),
	.w2(32'hbbb1f7a9),
	.w3(32'hbbbcb354),
	.w4(32'h3bb320d5),
	.w5(32'hbbb7d589),
	.w6(32'hbac77600),
	.w7(32'hbbb0f6c2),
	.w8(32'hbc0d3db3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf66114),
	.w1(32'h3c22d3cf),
	.w2(32'hb91d7638),
	.w3(32'hbb928a5c),
	.w4(32'h3b0ee591),
	.w5(32'h394e5550),
	.w6(32'hbbe2ee3a),
	.w7(32'h3a79399d),
	.w8(32'hb9e1d879),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d866cdf),
	.w1(32'hbc1b212d),
	.w2(32'hbcc4783c),
	.w3(32'h3d2e1c23),
	.w4(32'hbc9d18e4),
	.w5(32'hbcb05f27),
	.w6(32'h3d5f3810),
	.w7(32'hbbad5418),
	.w8(32'hbb886835),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ed22a),
	.w1(32'h3c079cc7),
	.w2(32'hbb38eee2),
	.w3(32'h3c08bd64),
	.w4(32'h3b0642f1),
	.w5(32'h3baa1161),
	.w6(32'h3a5a72f0),
	.w7(32'hbbfc5604),
	.w8(32'h3b64123b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d575b27),
	.w1(32'h3c1e204b),
	.w2(32'h3b12e375),
	.w3(32'h3d17899e),
	.w4(32'hbb5eaf33),
	.w5(32'hbc41f53a),
	.w6(32'h3cd25955),
	.w7(32'hbbe20736),
	.w8(32'hbc86881d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba658a84),
	.w1(32'hbb2b95fc),
	.w2(32'h37935f4c),
	.w3(32'hb8e96c6d),
	.w4(32'hba3e32cc),
	.w5(32'hbc59b2ce),
	.w6(32'hbadffea9),
	.w7(32'hbb13622a),
	.w8(32'hbbe88295),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9202b5),
	.w1(32'h3b014f9a),
	.w2(32'h3c1c4876),
	.w3(32'hbc4db34b),
	.w4(32'hbb1a14f4),
	.w5(32'h3bb8c936),
	.w6(32'hba514d92),
	.w7(32'hbb81ce31),
	.w8(32'hbc1d57e7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb97c),
	.w1(32'hba3afd7e),
	.w2(32'hbc0c0544),
	.w3(32'h3b76c496),
	.w4(32'hbbe3bc98),
	.w5(32'hbbdeab1c),
	.w6(32'hbca6cea0),
	.w7(32'hbcd6b216),
	.w8(32'hbc467496),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab4fc4),
	.w1(32'hba837046),
	.w2(32'h3a829bef),
	.w3(32'hb64391a2),
	.w4(32'h3ac35aa3),
	.w5(32'h3c116c17),
	.w6(32'hbb6ccbbf),
	.w7(32'hbbe6cd37),
	.w8(32'h3c9182af),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c132b07),
	.w1(32'h3c5d6b5d),
	.w2(32'h39f5c614),
	.w3(32'h3ced933a),
	.w4(32'h3d2a4777),
	.w5(32'h3b1f4434),
	.w6(32'h3d25a22d),
	.w7(32'h3ca71892),
	.w8(32'h3a795ea9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0836b0),
	.w1(32'hba87efb9),
	.w2(32'hbbb5c071),
	.w3(32'h3a8b3fb1),
	.w4(32'hbb99c190),
	.w5(32'h3c4a4b16),
	.w6(32'hbb8964a0),
	.w7(32'hbb8905eb),
	.w8(32'h3b141b3e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa05480),
	.w1(32'h3c966f43),
	.w2(32'h3a2c3b88),
	.w3(32'hba1b03e6),
	.w4(32'h3b278d1e),
	.w5(32'h3bcb30f4),
	.w6(32'hbcdd2b74),
	.w7(32'h3b393cc8),
	.w8(32'h3b9649c4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce54e9e),
	.w1(32'h3bae692c),
	.w2(32'h3c288f68),
	.w3(32'h3ce14737),
	.w4(32'h3c411489),
	.w5(32'h3c9864ce),
	.w6(32'h3ccb0cb4),
	.w7(32'h3a8692f7),
	.w8(32'hbc3c4ae3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8a951b),
	.w1(32'h3c61fe6a),
	.w2(32'hbbbfd47f),
	.w3(32'h3d74b981),
	.w4(32'hbc860673),
	.w5(32'hbcb9687a),
	.w6(32'h3d120e37),
	.w7(32'hbd188660),
	.w8(32'hbca7ea0b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad6026),
	.w1(32'h3a4aa064),
	.w2(32'h3bbf13ca),
	.w3(32'h3a76f0eb),
	.w4(32'h3be9b7ba),
	.w5(32'h3b404c2d),
	.w6(32'h3b83e0dd),
	.w7(32'h3c472198),
	.w8(32'hba8c91a7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bb3d4),
	.w1(32'h3b262310),
	.w2(32'hbbd5ca87),
	.w3(32'h3b584a6b),
	.w4(32'hbac5babf),
	.w5(32'hbc0aee30),
	.w6(32'hbad6382c),
	.w7(32'hbc3e9f8a),
	.w8(32'h3818b4b3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b1eb6),
	.w1(32'hbb9dfc43),
	.w2(32'hbbda939e),
	.w3(32'hbb1c86b8),
	.w4(32'hb9ef6bf9),
	.w5(32'h3b87d2f8),
	.w6(32'hbb9e64b3),
	.w7(32'hbb14c0fe),
	.w8(32'h3c1b453a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e0936),
	.w1(32'h3bf6572b),
	.w2(32'hbb5bc3be),
	.w3(32'h3c180021),
	.w4(32'h3c31b665),
	.w5(32'hbb43763b),
	.w6(32'hba68b4e6),
	.w7(32'hbb0c6dcf),
	.w8(32'h3891e6f6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86972a),
	.w1(32'hbbc87841),
	.w2(32'hbb9c6198),
	.w3(32'hbba36b3e),
	.w4(32'hbb642ece),
	.w5(32'hbc4eef96),
	.w6(32'hbbf20541),
	.w7(32'hbb921f0c),
	.w8(32'hbca68ec9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59d6b1),
	.w1(32'h3c2cb5c2),
	.w2(32'hbc8dc91d),
	.w3(32'h3c25ed3b),
	.w4(32'h3bcfc5bd),
	.w5(32'hbcaaf1db),
	.w6(32'h3b00a317),
	.w7(32'hbaa13d3a),
	.w8(32'hbb4cdbb6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03e9f7),
	.w1(32'h3bb5c34e),
	.w2(32'hbbac107b),
	.w3(32'h3c851c1b),
	.w4(32'h3c64f4f2),
	.w5(32'hba94e917),
	.w6(32'hba47bb74),
	.w7(32'h3aa98322),
	.w8(32'hbbe6437a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3eb67),
	.w1(32'hb78f64d9),
	.w2(32'hbbaaea46),
	.w3(32'h3c09d998),
	.w4(32'h3c2c7937),
	.w5(32'h38a97150),
	.w6(32'hbb952081),
	.w7(32'hbbb13736),
	.w8(32'hbc4e81b8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae34efc),
	.w1(32'hbb1f7fb0),
	.w2(32'hbca1793e),
	.w3(32'hbaacdb1d),
	.w4(32'hbc17bf2e),
	.w5(32'hbc2eb612),
	.w6(32'hbceaed85),
	.w7(32'hbced6c50),
	.w8(32'hbc763dc6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1080be),
	.w1(32'h3ad48b8f),
	.w2(32'hbc22bd25),
	.w3(32'hba0140b5),
	.w4(32'h3ab867a4),
	.w5(32'hbc889d34),
	.w6(32'h3aa1700f),
	.w7(32'h3b03ad71),
	.w8(32'h3c5982e6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1ca8e),
	.w1(32'h3a4791ed),
	.w2(32'hbb4d0370),
	.w3(32'hbb99c937),
	.w4(32'h3c8a2c56),
	.w5(32'hbba1287c),
	.w6(32'h3cb0b443),
	.w7(32'h3c9c07e5),
	.w8(32'hbbc2d046),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9c7e9),
	.w1(32'h3a8e6790),
	.w2(32'hbb1bd65e),
	.w3(32'h3af18d0d),
	.w4(32'h3b951183),
	.w5(32'hbc99ca13),
	.w6(32'h3b94aba7),
	.w7(32'hbb3dabd8),
	.w8(32'hbcc03b9e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc496184),
	.w1(32'hbc821b18),
	.w2(32'hbc16cc3b),
	.w3(32'hbc9ba8fb),
	.w4(32'hbc73d332),
	.w5(32'hbb0c8fa6),
	.w6(32'hbca0077b),
	.w7(32'hbb0d613c),
	.w8(32'hbb8f8bc2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5aa183),
	.w1(32'h3bccd3bf),
	.w2(32'hbb59bee2),
	.w3(32'h3bf825e9),
	.w4(32'hb9f8e022),
	.w5(32'hbbd9e562),
	.w6(32'hba371de3),
	.w7(32'hbc1463d0),
	.w8(32'hbbb7cf97),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51aa50),
	.w1(32'hbc7e3fa6),
	.w2(32'hbcee4605),
	.w3(32'hbcb028b4),
	.w4(32'hbc38ba65),
	.w5(32'hbc7d53a8),
	.w6(32'hbc7e8676),
	.w7(32'hbc452bfb),
	.w8(32'hbc6d91c7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37c766),
	.w1(32'hbbb3d84a),
	.w2(32'h3aa2c8f9),
	.w3(32'hbbb062cb),
	.w4(32'hbaf2845e),
	.w5(32'hbb07d201),
	.w6(32'h3bb6d9d2),
	.w7(32'h3cb735cf),
	.w8(32'hbb25ea67),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37be43),
	.w1(32'hbb508ae6),
	.w2(32'hbc190752),
	.w3(32'hbb602de9),
	.w4(32'h3a7d5dac),
	.w5(32'hbc2a12ed),
	.w6(32'h3b8d29be),
	.w7(32'h3b38d6d8),
	.w8(32'h3a34b3cb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69be62),
	.w1(32'h3bb8eec4),
	.w2(32'h3b09bade),
	.w3(32'h3bdfaf19),
	.w4(32'h3bdf27cf),
	.w5(32'hbbaf01c1),
	.w6(32'h3bda8f35),
	.w7(32'h3b2b6c17),
	.w8(32'hbb85c3ad),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67f8ee),
	.w1(32'h3b553cc1),
	.w2(32'h3a638267),
	.w3(32'h3a3d56cc),
	.w4(32'h3c1415b3),
	.w5(32'hbb53e3e1),
	.w6(32'h3b922e7b),
	.w7(32'h3bb6448c),
	.w8(32'hbc0e4feb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06d695),
	.w1(32'hbb919821),
	.w2(32'h39adda32),
	.w3(32'h3a768ccb),
	.w4(32'hbbbe67b3),
	.w5(32'hbbda57cd),
	.w6(32'hbb560538),
	.w7(32'hbc1d1739),
	.w8(32'h39fbc5be),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2bbb4),
	.w1(32'h3b319d5d),
	.w2(32'hbb074b26),
	.w3(32'hbada7567),
	.w4(32'h3c22182b),
	.w5(32'h3b39b21c),
	.w6(32'h3c615dfb),
	.w7(32'h3b990752),
	.w8(32'h3c371680),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a6670),
	.w1(32'h3b6e0611),
	.w2(32'hbbca2928),
	.w3(32'h3c0de34d),
	.w4(32'h3bf6c309),
	.w5(32'hbad3f5fc),
	.w6(32'h3b063815),
	.w7(32'h3b10abd6),
	.w8(32'hbb8cedcc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f5949),
	.w1(32'hbc24c752),
	.w2(32'hbc44e912),
	.w3(32'hbc014440),
	.w4(32'hbbf92ebd),
	.w5(32'hbbd7a5e1),
	.w6(32'hbbbf8ddb),
	.w7(32'hbbe289ae),
	.w8(32'hbbc361c2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06befb),
	.w1(32'hba1cb25f),
	.w2(32'hba358264),
	.w3(32'hbb8cb1d3),
	.w4(32'h3aad9014),
	.w5(32'h3b571dc3),
	.w6(32'h3b180c1b),
	.w7(32'hbbca8319),
	.w8(32'h3aca8566),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b485c32),
	.w1(32'h3be67071),
	.w2(32'hb9a8bd2a),
	.w3(32'h3c6ce10e),
	.w4(32'h3c6abbdf),
	.w5(32'hbb9f6349),
	.w6(32'h3bb2be1c),
	.w7(32'hbb93a8b7),
	.w8(32'h3b97ff7c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beec5f7),
	.w1(32'h3c0391dd),
	.w2(32'h3b24ff9c),
	.w3(32'h3bf4ab09),
	.w4(32'h3bbc9d2c),
	.w5(32'hb73f564c),
	.w6(32'h3adf96e3),
	.w7(32'h3a24e0ab),
	.w8(32'hbb5eabef),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ce25c),
	.w1(32'hbb1d67a1),
	.w2(32'h3b397ced),
	.w3(32'hbaf3fe1d),
	.w4(32'hba3c8e41),
	.w5(32'h3b13e909),
	.w6(32'hbbb0ec1e),
	.w7(32'hbb21106c),
	.w8(32'h3b8c9f0d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a72bf),
	.w1(32'h3c26a2f4),
	.w2(32'hbc0e5fb0),
	.w3(32'h3b3530f2),
	.w4(32'h3bb69ddf),
	.w5(32'hbb0b2aa2),
	.w6(32'hbbb6b5ba),
	.w7(32'hbb50cfbe),
	.w8(32'hbc01cfae),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3c659),
	.w1(32'hbc299012),
	.w2(32'hbc13a5e8),
	.w3(32'h3b9d9e24),
	.w4(32'h3c31ccc3),
	.w5(32'hbbb6d42a),
	.w6(32'hbcbf0ea2),
	.w7(32'hbc6bd968),
	.w8(32'hbce3e502),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2656d7),
	.w1(32'hbbafa98e),
	.w2(32'hbc8bdc9c),
	.w3(32'hbc35532c),
	.w4(32'hbb90aa38),
	.w5(32'hbb6dc45e),
	.w6(32'hbcc40d3f),
	.w7(32'hbbde32d3),
	.w8(32'hbc9bb99f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf2fc50),
	.w1(32'h3c433d80),
	.w2(32'h3bc05b96),
	.w3(32'h3c9a18fb),
	.w4(32'h3c73bf54),
	.w5(32'h3c5cb01f),
	.w6(32'h3bff7b0b),
	.w7(32'hbb6d1c7e),
	.w8(32'hbc2b796a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa94da7),
	.w1(32'h3b398652),
	.w2(32'h3a389c4a),
	.w3(32'hbbc5f7dd),
	.w4(32'h3b3e23e7),
	.w5(32'hba388498),
	.w6(32'hbbfd7963),
	.w7(32'h3c01ff59),
	.w8(32'hbbfb1338),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3cc9a),
	.w1(32'hba0302c4),
	.w2(32'hbac9bb8d),
	.w3(32'h3b5f7475),
	.w4(32'h3bc72463),
	.w5(32'h3af4861b),
	.w6(32'hbba61f55),
	.w7(32'hbb89b2bf),
	.w8(32'h3c18a78d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad773d6),
	.w1(32'hbbdaefd7),
	.w2(32'h3b98e97a),
	.w3(32'h3ae71dc9),
	.w4(32'hbba3dab7),
	.w5(32'hbbf97d86),
	.w6(32'hbbd83d32),
	.w7(32'hbc8a1107),
	.w8(32'hbc609337),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d76186),
	.w1(32'h3ba3a3ab),
	.w2(32'hbbc0ed97),
	.w3(32'hbbb6395a),
	.w4(32'hbba3bb0a),
	.w5(32'hbaa84896),
	.w6(32'h39da1ea9),
	.w7(32'h3b879d90),
	.w8(32'hbb4ae5a7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05706),
	.w1(32'h3afafdf7),
	.w2(32'hbb3fb027),
	.w3(32'hbabb362d),
	.w4(32'h3b1a1a7a),
	.w5(32'hbc36cdd6),
	.w6(32'hba1b5028),
	.w7(32'h3b85d8d8),
	.w8(32'hbc304a2e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39799c),
	.w1(32'hbc06380f),
	.w2(32'hbbb96148),
	.w3(32'hbc4b3e87),
	.w4(32'hbc798ace),
	.w5(32'hbbe583f7),
	.w6(32'hbc8b61ec),
	.w7(32'hbc7df273),
	.w8(32'hbb1c60eb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81076e),
	.w1(32'hbbc6148a),
	.w2(32'hbb3c7838),
	.w3(32'hbaeb411c),
	.w4(32'hbc103342),
	.w5(32'hbbb64855),
	.w6(32'hbc851f84),
	.w7(32'hbc229d0e),
	.w8(32'h3b862dc9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddebb0),
	.w1(32'h3c386cfe),
	.w2(32'hbb29b122),
	.w3(32'h3c329885),
	.w4(32'h3cb6fbf9),
	.w5(32'hbc0e7350),
	.w6(32'h3c113307),
	.w7(32'hbb8dce33),
	.w8(32'hbba473da),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08fc38),
	.w1(32'h3c0a2cc7),
	.w2(32'hbbead214),
	.w3(32'hbc06ae40),
	.w4(32'h3c715540),
	.w5(32'hbb761b54),
	.w6(32'h3bb0c92c),
	.w7(32'h3c008f5a),
	.w8(32'hbbd17479),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d0dc5),
	.w1(32'h3b1c153f),
	.w2(32'hbbca0782),
	.w3(32'h3b0e86f4),
	.w4(32'h3b4c328d),
	.w5(32'hbbe4b066),
	.w6(32'hbbbbe9ef),
	.w7(32'hbbaf4f2f),
	.w8(32'hbc250be0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbe28f),
	.w1(32'hbbb94ae6),
	.w2(32'hbb286def),
	.w3(32'hbc43d59e),
	.w4(32'hbb94b836),
	.w5(32'hb9f4f0ba),
	.w6(32'hbc39c34a),
	.w7(32'h3b807a63),
	.w8(32'hbbc7c97d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ec577),
	.w1(32'hb9123e00),
	.w2(32'hbb9db7c7),
	.w3(32'h3b178118),
	.w4(32'hbae70dc4),
	.w5(32'h3bc06ffc),
	.w6(32'hbbca3803),
	.w7(32'hbbf1d1ef),
	.w8(32'hbb36b244),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6cc838),
	.w1(32'h3ca1a98b),
	.w2(32'hbb1619ab),
	.w3(32'h3c335534),
	.w4(32'h3c3a32aa),
	.w5(32'h3b397328),
	.w6(32'h3c11e78f),
	.w7(32'h3b96c044),
	.w8(32'hbb1cc911),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc207015),
	.w1(32'hbc0358c0),
	.w2(32'hbb3f9224),
	.w3(32'hbaa3507d),
	.w4(32'hba217632),
	.w5(32'h3b08e82f),
	.w6(32'hbbb1d82f),
	.w7(32'hbb94cb8b),
	.w8(32'hba88ef3c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b486a2c),
	.w1(32'h3afcba37),
	.w2(32'hb9e5fc5b),
	.w3(32'h3b9421e5),
	.w4(32'h3b41e131),
	.w5(32'h3cb3f32a),
	.w6(32'h3ace6006),
	.w7(32'hb85fd910),
	.w8(32'h3cbf87eb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca704e8),
	.w1(32'h3cddafc2),
	.w2(32'h3b395712),
	.w3(32'h3d3fc1cf),
	.w4(32'h3c248414),
	.w5(32'h3891f0ce),
	.w6(32'h3c8e5f03),
	.w7(32'hbc8e7fd5),
	.w8(32'hbb611cb8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae544c2),
	.w1(32'h3b8f3221),
	.w2(32'h3b0e33ae),
	.w3(32'h3a828499),
	.w4(32'h3c4bacd3),
	.w5(32'h3b8246ee),
	.w6(32'hbb9e10f4),
	.w7(32'hbb059591),
	.w8(32'hbb443755),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996f64b),
	.w1(32'h3a768eda),
	.w2(32'h3b44534b),
	.w3(32'hb8c703a4),
	.w4(32'h3ae39d3d),
	.w5(32'hbb1c5be1),
	.w6(32'hbab47215),
	.w7(32'h391cdc1e),
	.w8(32'hba92e66f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90435c9),
	.w1(32'hbbc06d1d),
	.w2(32'h38fae083),
	.w3(32'hbb3b8380),
	.w4(32'hbadd3aae),
	.w5(32'h3c8a8fa9),
	.w6(32'hbba26e39),
	.w7(32'hbc114bdd),
	.w8(32'h3c7fb438),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99c75a),
	.w1(32'h3ba763b7),
	.w2(32'hb984b16b),
	.w3(32'h3bdfb787),
	.w4(32'h3c8fa14e),
	.w5(32'hbbce844d),
	.w6(32'h3a9a9405),
	.w7(32'hbbbe14e8),
	.w8(32'hbc7ace1a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95edf2),
	.w1(32'hb96cfebf),
	.w2(32'hba24cd0a),
	.w3(32'hba7ac8aa),
	.w4(32'hbc425431),
	.w5(32'hbc0bd19f),
	.w6(32'h3c51bafd),
	.w7(32'h3bba51f4),
	.w8(32'hbb7f1cf5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc383dd5),
	.w1(32'h3b2afd74),
	.w2(32'hbb7330df),
	.w3(32'hbb59e726),
	.w4(32'hbb857e37),
	.w5(32'hbb233cb0),
	.w6(32'hbc555ce9),
	.w7(32'h39cc933b),
	.w8(32'hbc1f95f8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6591b),
	.w1(32'hbafa7a11),
	.w2(32'h3b657cad),
	.w3(32'h390d990c),
	.w4(32'hbc08a5aa),
	.w5(32'hbbe91a41),
	.w6(32'hbb5fc232),
	.w7(32'hbc4f6fc6),
	.w8(32'hbbe118c2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07bd7d),
	.w1(32'h3c06b9ec),
	.w2(32'hbc1f6069),
	.w3(32'h3afe643d),
	.w4(32'h3c647469),
	.w5(32'h3b9a4392),
	.w6(32'hbbf5b508),
	.w7(32'h3b21e252),
	.w8(32'hbc90593b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962a897),
	.w1(32'hba833f6c),
	.w2(32'h3c4673c2),
	.w3(32'hbc393ddc),
	.w4(32'hbc05924c),
	.w5(32'h3b8a5024),
	.w6(32'hbc39224c),
	.w7(32'hbbace53c),
	.w8(32'h3ade802a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb07a0),
	.w1(32'h3999091f),
	.w2(32'hbbbf6019),
	.w3(32'h3c3e127b),
	.w4(32'h3bb339dc),
	.w5(32'hbc4a1f3d),
	.w6(32'h3cb782d8),
	.w7(32'hbc629413),
	.w8(32'hbc4e2a2e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c2192),
	.w1(32'hbb9b31ca),
	.w2(32'h3bd944e7),
	.w3(32'hbba85b9b),
	.w4(32'h3c51bd26),
	.w5(32'hbb3136a9),
	.w6(32'h3b8d5ab1),
	.w7(32'h3c65c98a),
	.w8(32'h3b0c52e6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be19680),
	.w1(32'hbb651906),
	.w2(32'hbcc4639e),
	.w3(32'h3c1443e3),
	.w4(32'h3c7bf2f3),
	.w5(32'hbc8f1e25),
	.w6(32'hbabab674),
	.w7(32'hba996d63),
	.w8(32'hbc506e0f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b9a67),
	.w1(32'hba4c238f),
	.w2(32'hbbd12b8d),
	.w3(32'hbada1449),
	.w4(32'h3c8ce495),
	.w5(32'hbbbd8ba3),
	.w6(32'h3c7f0a5f),
	.w7(32'h3ade30e7),
	.w8(32'hbc3eeedd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b9daa),
	.w1(32'hbb00edfe),
	.w2(32'hbc652263),
	.w3(32'hbc4b041e),
	.w4(32'hbbdf9528),
	.w5(32'hbac67daf),
	.w6(32'hbd038f30),
	.w7(32'h3aa0cbdd),
	.w8(32'h3ba7aee3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c1878),
	.w1(32'h3bb6aae5),
	.w2(32'h3abca76b),
	.w3(32'h3bc22755),
	.w4(32'h3c37204e),
	.w5(32'h3a77e17a),
	.w6(32'h3bbb38f5),
	.w7(32'hbb8fcc44),
	.w8(32'h39d4d4dd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c659558),
	.w1(32'h3c7da828),
	.w2(32'hbc185b94),
	.w3(32'h3ca150a0),
	.w4(32'h3ca0eaf9),
	.w5(32'hbb2e3205),
	.w6(32'h3bbf042c),
	.w7(32'hbbae3ea0),
	.w8(32'hbc0438d2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e00f6),
	.w1(32'h3bc2a914),
	.w2(32'hbb1b255e),
	.w3(32'h3c5c1e52),
	.w4(32'h3c8af167),
	.w5(32'h3c0e8bcf),
	.w6(32'h3c30ff1b),
	.w7(32'h3c0a909a),
	.w8(32'hbb643356),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ab33b),
	.w1(32'hba9189d5),
	.w2(32'hba068553),
	.w3(32'hbc0f9ef4),
	.w4(32'hb91a434c),
	.w5(32'h3b94aad1),
	.w6(32'hbab0e9b6),
	.w7(32'h3bcb4b06),
	.w8(32'h3ba1b22d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d7baa),
	.w1(32'h3c5e60b3),
	.w2(32'hbc53eefb),
	.w3(32'h3b94edaa),
	.w4(32'h3bce66f7),
	.w5(32'hbc364eb7),
	.w6(32'hbc39b7e5),
	.w7(32'hbc34dee9),
	.w8(32'hbb8a243b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b113797),
	.w1(32'h3b8fbe7f),
	.w2(32'hbbadae19),
	.w3(32'h3b6aab29),
	.w4(32'h3c195b01),
	.w5(32'hbbe555a6),
	.w6(32'h3baea5ac),
	.w7(32'hbb2743cf),
	.w8(32'hbbdb5507),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1029e1),
	.w1(32'h3b720495),
	.w2(32'h3aa3e72c),
	.w3(32'h3b48160f),
	.w4(32'h3baabbe3),
	.w5(32'h3b6612b3),
	.w6(32'h3b3ddd4d),
	.w7(32'h383236d7),
	.w8(32'hbbbdfce0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd71e9),
	.w1(32'hbb575b34),
	.w2(32'hb9a16450),
	.w3(32'hbbb143bf),
	.w4(32'hbb8e4d66),
	.w5(32'h3be90fe0),
	.w6(32'hbc02939b),
	.w7(32'hbc38779e),
	.w8(32'h3a525a65),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61ffcd),
	.w1(32'hba1190bf),
	.w2(32'hbc39f8ab),
	.w3(32'hbb0c83e6),
	.w4(32'h397a99a0),
	.w5(32'hbc89a32c),
	.w6(32'hbc84870b),
	.w7(32'hbc1b88b9),
	.w8(32'hbbfe426c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9973b75),
	.w1(32'h3a992946),
	.w2(32'hba8abd15),
	.w3(32'hba63bf58),
	.w4(32'h3c6c727f),
	.w5(32'h3c1d29b4),
	.w6(32'h3c8234d0),
	.w7(32'hbaac5bc6),
	.w8(32'hbbbe00df),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61c1ea),
	.w1(32'h36515430),
	.w2(32'hbbcae881),
	.w3(32'h3cb7a79d),
	.w4(32'h3bc3e008),
	.w5(32'hbbaedfa3),
	.w6(32'h3caeafd8),
	.w7(32'h3bb343b9),
	.w8(32'h3c077e2d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bb273),
	.w1(32'h3c6f7203),
	.w2(32'hbab05901),
	.w3(32'h3ca6679b),
	.w4(32'h3cacb395),
	.w5(32'h3a924e1d),
	.w6(32'h3c500b42),
	.w7(32'hb8d1391b),
	.w8(32'hbc8421b6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ada6f),
	.w1(32'hbc177da3),
	.w2(32'h3be423f5),
	.w3(32'hbc2d0bc1),
	.w4(32'hbc6dabf2),
	.w5(32'h3b9df474),
	.w6(32'hbcceedad),
	.w7(32'hbc82fbd4),
	.w8(32'h3c050cab),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc735ce2),
	.w1(32'hbb07bd0d),
	.w2(32'hbc433d28),
	.w3(32'hbc088c50),
	.w4(32'h3c75b570),
	.w5(32'hbb96d675),
	.w6(32'hbbb1d9b2),
	.w7(32'hbbf5cb19),
	.w8(32'h3c6d9883),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b04b6),
	.w1(32'h3c3f83b4),
	.w2(32'h3a2f6a61),
	.w3(32'h3c8057a3),
	.w4(32'h3d36afb9),
	.w5(32'h3af8585f),
	.w6(32'h3cfdc4cc),
	.w7(32'h3d0b52d2),
	.w8(32'hbb7670b3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be16910),
	.w1(32'h3bbfff6c),
	.w2(32'h3b5f62b9),
	.w3(32'h3b303963),
	.w4(32'hbae9b8b3),
	.w5(32'h3bc939c9),
	.w6(32'h3b38f92d),
	.w7(32'hbb1c1e1e),
	.w8(32'h3b44714a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef13f1),
	.w1(32'hbb5b6206),
	.w2(32'hbb474422),
	.w3(32'hbb513195),
	.w4(32'hb7c1b227),
	.w5(32'h3b25bea5),
	.w6(32'hbba71228),
	.w7(32'h3bc320ab),
	.w8(32'h3a94f3c6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb857a814),
	.w1(32'h3b38cc66),
	.w2(32'h3a7dc90a),
	.w3(32'h3b236bd6),
	.w4(32'h3aeba24a),
	.w5(32'hbc26a187),
	.w6(32'h3b37f25d),
	.w7(32'hbbb2f179),
	.w8(32'hbabc0c39),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a566f7a),
	.w1(32'h3c1469b2),
	.w2(32'h3b168f63),
	.w3(32'h3bafe2af),
	.w4(32'hbb764d5b),
	.w5(32'h3a8ec8c2),
	.w6(32'hbc1e4738),
	.w7(32'hbc84db89),
	.w8(32'h387ef73f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f38f5),
	.w1(32'h3c52f3fd),
	.w2(32'hbc413cb6),
	.w3(32'h3c65600c),
	.w4(32'h3c924dc6),
	.w5(32'hba589307),
	.w6(32'h3bd4ca9d),
	.w7(32'hbbcb91e0),
	.w8(32'hbc0d42a6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb398888),
	.w1(32'hbb5710ba),
	.w2(32'hb99ad005),
	.w3(32'h3b3da92a),
	.w4(32'h3b471994),
	.w5(32'h3981e60a),
	.w6(32'hb94a3a4f),
	.w7(32'hbbb8f706),
	.w8(32'hbb13e21f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af06df),
	.w1(32'h39b13545),
	.w2(32'h37b1cb61),
	.w3(32'h3b22f895),
	.w4(32'hbab18028),
	.w5(32'hbaeaaec6),
	.w6(32'hbb6e6a82),
	.w7(32'hbbadae42),
	.w8(32'hbb8dff58),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62c886),
	.w1(32'h3b4edc80),
	.w2(32'hbb025f47),
	.w3(32'h3c5bf130),
	.w4(32'h3bb6764f),
	.w5(32'hbc0ee9f9),
	.w6(32'h3c28f744),
	.w7(32'hbb8b7b29),
	.w8(32'hbc8e1dfb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ac0d7),
	.w1(32'h3ae00074),
	.w2(32'hbaec1f30),
	.w3(32'hbb26df43),
	.w4(32'h3cc2c2c6),
	.w5(32'h3b49038c),
	.w6(32'h3c669f7d),
	.w7(32'h3c6db71e),
	.w8(32'h3b2971d1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9134d1a),
	.w1(32'h3b6cb76f),
	.w2(32'hbbe88922),
	.w3(32'h3b5343ef),
	.w4(32'h3b35c78d),
	.w5(32'hbc6f0901),
	.w6(32'h3b267621),
	.w7(32'hbb76af2c),
	.w8(32'hbcb426da),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98b8ed),
	.w1(32'hbc9b1c9c),
	.w2(32'hbbc7d085),
	.w3(32'hbcba4419),
	.w4(32'hbc8d0f37),
	.w5(32'h3b9b204e),
	.w6(32'hbc8662d5),
	.w7(32'h3a2578bf),
	.w8(32'h3b9fe97b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f1b6c),
	.w1(32'hbba37126),
	.w2(32'hbb930a3e),
	.w3(32'hbb1d13a2),
	.w4(32'hbc0f52ea),
	.w5(32'hbb586efe),
	.w6(32'hbb98d8f2),
	.w7(32'hbc4da83e),
	.w8(32'h3992e684),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d1436),
	.w1(32'hbc9ae630),
	.w2(32'hbbc8a930),
	.w3(32'h3bfb35f5),
	.w4(32'hbc01817a),
	.w5(32'h3b768c58),
	.w6(32'hbc3c5929),
	.w7(32'hbc241a69),
	.w8(32'hbc21ecc0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b095),
	.w1(32'h3a26e67d),
	.w2(32'hbbee0611),
	.w3(32'h3bdba8e2),
	.w4(32'h3b6453c1),
	.w5(32'hbc3250b0),
	.w6(32'hbc8b186b),
	.w7(32'hbc786132),
	.w8(32'hbc855401),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae6ff4),
	.w1(32'hbba09cb5),
	.w2(32'h3bfc93d3),
	.w3(32'hbc8181d5),
	.w4(32'hbbbaba6c),
	.w5(32'h3c00916f),
	.w6(32'hbc204a0b),
	.w7(32'hbbbdf8ff),
	.w8(32'hbb3786b2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae2615),
	.w1(32'hbb80add0),
	.w2(32'h3969617f),
	.w3(32'hbb3c628f),
	.w4(32'hbc4b2a3a),
	.w5(32'hbb824024),
	.w6(32'hbca88e02),
	.w7(32'hbb6e6390),
	.w8(32'hbbb89cb1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b32d8),
	.w1(32'hbb2c6de9),
	.w2(32'h3ae44fad),
	.w3(32'hbac0deb9),
	.w4(32'h3c1469ba),
	.w5(32'h3cb9c786),
	.w6(32'h3bb2ebef),
	.w7(32'h3bc28743),
	.w8(32'h3c893ed3),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8eaec4),
	.w1(32'h3cbeee40),
	.w2(32'h3a7b0580),
	.w3(32'h3d1e8489),
	.w4(32'h3c48c393),
	.w5(32'hba3896b9),
	.w6(32'h3b5ac30c),
	.w7(32'hbc05ac9c),
	.w8(32'hbbd38b88),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05b7ce),
	.w1(32'h3b5898a4),
	.w2(32'hbc1a3086),
	.w3(32'hba95e457),
	.w4(32'h3bc16fc6),
	.w5(32'hbb540102),
	.w6(32'h3bbda663),
	.w7(32'h3ba71840),
	.w8(32'hbbbc5d18),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005f03),
	.w1(32'hbb5ac314),
	.w2(32'hbcc86a9d),
	.w3(32'hbb9dc033),
	.w4(32'hbb154828),
	.w5(32'hbc2361ba),
	.w6(32'hbbffe417),
	.w7(32'hbb1ce8ef),
	.w8(32'hbc1feefd),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf37c8a),
	.w1(32'h3c2d29ab),
	.w2(32'h3b3e1887),
	.w3(32'h3c007cf3),
	.w4(32'h3c987a19),
	.w5(32'hbb903df4),
	.w6(32'h3c71f0cf),
	.w7(32'hbb421c55),
	.w8(32'hbc8dae96),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc187b89),
	.w1(32'hbbb5a638),
	.w2(32'hb8f992f4),
	.w3(32'hbbb5292f),
	.w4(32'hbbc53fe0),
	.w5(32'h3c5453fe),
	.w6(32'hbca53726),
	.w7(32'hbc95044c),
	.w8(32'h3bc5e3ff),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf55d85),
	.w1(32'h3845a8f5),
	.w2(32'hbbd44a66),
	.w3(32'h3c049efd),
	.w4(32'hbbaddb63),
	.w5(32'hbb859ec2),
	.w6(32'hbb7000f8),
	.w7(32'h3b0b2c72),
	.w8(32'hbbc16f11),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5e60e),
	.w1(32'h3b6a97d4),
	.w2(32'h3c06e2f4),
	.w3(32'hb8d6abbc),
	.w4(32'h3bcdc7a7),
	.w5(32'h3c57409c),
	.w6(32'hbc1fd7a4),
	.w7(32'hbb0c2152),
	.w8(32'hbba7a708),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9d2e8),
	.w1(32'h3ae091fc),
	.w2(32'h3b0a0d85),
	.w3(32'h3b8960bd),
	.w4(32'h3bf1cf5a),
	.w5(32'hbaac52ee),
	.w6(32'hbbc3c80c),
	.w7(32'hbb85cf06),
	.w8(32'hbb22c0b1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66d136),
	.w1(32'h3afbafc6),
	.w2(32'hbaa328ab),
	.w3(32'h3a3a74a7),
	.w4(32'h3b48fb8b),
	.w5(32'h3ad93da9),
	.w6(32'h3ad9a380),
	.w7(32'h3b6104aa),
	.w8(32'hbc030c0f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d37b93a),
	.w1(32'h3b062a14),
	.w2(32'hba98c973),
	.w3(32'h3cff1727),
	.w4(32'hb91031ea),
	.w5(32'hbcb45cd5),
	.w6(32'h3d363aa0),
	.w7(32'hbc0390ee),
	.w8(32'hbc986dc7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe59a3b),
	.w1(32'hbc2b374b),
	.w2(32'h3a6e5c78),
	.w3(32'hbc70a67d),
	.w4(32'hbc3b16fe),
	.w5(32'h395fcd7a),
	.w6(32'hbc109d1f),
	.w7(32'hbb326262),
	.w8(32'h3b0c8dcf),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ad17f),
	.w1(32'hbb470246),
	.w2(32'h3b73ece3),
	.w3(32'hba145cdb),
	.w4(32'hba82b87c),
	.w5(32'h3a4ef1e9),
	.w6(32'h3bbcb8e6),
	.w7(32'h3b2dd504),
	.w8(32'hb9d06e1a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b129e59),
	.w1(32'h3893abe2),
	.w2(32'h3ba166d2),
	.w3(32'hba127367),
	.w4(32'hba1e9e21),
	.w5(32'h3b57ae29),
	.w6(32'h388677f0),
	.w7(32'h3a3bf173),
	.w8(32'hbb3753f8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb709bb4),
	.w1(32'hb85e1bda),
	.w2(32'hbb834fad),
	.w3(32'hbbadd6b6),
	.w4(32'hba98a350),
	.w5(32'hbbfb7ce0),
	.w6(32'hbc12f322),
	.w7(32'hbba33c81),
	.w8(32'hbb489449),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa14b2),
	.w1(32'h3b8389e2),
	.w2(32'h3c23b556),
	.w3(32'h3768a079),
	.w4(32'h3c2e8f4b),
	.w5(32'h3c546ea5),
	.w6(32'h39cde411),
	.w7(32'h3ad99faa),
	.w8(32'hbc7acf4f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c423d80),
	.w1(32'h3b8143bb),
	.w2(32'h3b812322),
	.w3(32'hbadedd87),
	.w4(32'hbb30d8ab),
	.w5(32'h3af11246),
	.w6(32'hbc4dc643),
	.w7(32'hbc40ef67),
	.w8(32'hbc6c073d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d72dd),
	.w1(32'hbb887aa1),
	.w2(32'hbb7c1f3f),
	.w3(32'hbbeced4d),
	.w4(32'hbc14006e),
	.w5(32'hba05fe25),
	.w6(32'hbc5757dc),
	.w7(32'hbb5915a4),
	.w8(32'h3a406090),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d4e46),
	.w1(32'h3c12c1a5),
	.w2(32'hbbaa9d24),
	.w3(32'h3c188166),
	.w4(32'h3ba7372a),
	.w5(32'h3b0b80ee),
	.w6(32'hbb19b7e4),
	.w7(32'hb9d610fa),
	.w8(32'hbc730838),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2ce30),
	.w1(32'h3b66566e),
	.w2(32'h3a853913),
	.w3(32'h3c2cb216),
	.w4(32'hbaa99f56),
	.w5(32'h3b3d385d),
	.w6(32'hbc4d2b1b),
	.w7(32'hbc7be2a1),
	.w8(32'hbb6003b5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c45c9),
	.w1(32'h3bce43c8),
	.w2(32'hbae7177d),
	.w3(32'h3a1154e5),
	.w4(32'hbafba0e8),
	.w5(32'h3a8ae0c0),
	.w6(32'hbbf9c650),
	.w7(32'hbb70c6a7),
	.w8(32'h3aa52e6a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2417da),
	.w1(32'h3b8b43e9),
	.w2(32'hbc5ebfa6),
	.w3(32'h3cf608a2),
	.w4(32'h3c097bbc),
	.w5(32'hbc463c67),
	.w6(32'h3d328a0b),
	.w7(32'h3c4b800f),
	.w8(32'hbc9e3e04),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd57400),
	.w1(32'h3b26e1eb),
	.w2(32'hbb9751fd),
	.w3(32'hbc2d66fe),
	.w4(32'hbc5c859c),
	.w5(32'hbb3052fa),
	.w6(32'hbc831732),
	.w7(32'hbcafdbcf),
	.w8(32'hbb98ed2b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cf0f7),
	.w1(32'hbb125878),
	.w2(32'h3afb44fa),
	.w3(32'hbbb6d4ad),
	.w4(32'hba1830c0),
	.w5(32'h3b2d7ce1),
	.w6(32'hba41e957),
	.w7(32'hbc35c906),
	.w8(32'h3abb4637),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c584cb8),
	.w1(32'h3b67c564),
	.w2(32'hbb20fea9),
	.w3(32'h3c861cdb),
	.w4(32'h3bc203c7),
	.w5(32'hbb8eebcb),
	.w6(32'h3c2d7e03),
	.w7(32'h3ad29496),
	.w8(32'hbbd03b0d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda65e8),
	.w1(32'hbbcb1079),
	.w2(32'hba8b8fe3),
	.w3(32'hbbf5c4d0),
	.w4(32'h3b5b2832),
	.w5(32'hbb7cf157),
	.w6(32'hbbb2bb19),
	.w7(32'h3a935020),
	.w8(32'hbc1d8313),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982eda),
	.w1(32'h3bb5bb74),
	.w2(32'h3b97f54d),
	.w3(32'h3c6cf78c),
	.w4(32'h3b725470),
	.w5(32'h3b432a6e),
	.w6(32'h3c78786c),
	.w7(32'h3bbb8cf5),
	.w8(32'h3a7e3578),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3997e),
	.w1(32'h3be069c0),
	.w2(32'hbbbf8965),
	.w3(32'h3b03b822),
	.w4(32'h3b5e2b8d),
	.w5(32'hbb33e637),
	.w6(32'h3b0a07e2),
	.w7(32'h3b733e49),
	.w8(32'hbb167080),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfcb78),
	.w1(32'h3a4d184c),
	.w2(32'hbc02fa86),
	.w3(32'hbb438a1d),
	.w4(32'hbb958d0b),
	.w5(32'hbb54f284),
	.w6(32'hbbd055b8),
	.w7(32'hb984db6d),
	.w8(32'hb9f42d92),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2cdf),
	.w1(32'hb91effcf),
	.w2(32'hbc21cd89),
	.w3(32'hbc161a50),
	.w4(32'hbb2a3068),
	.w5(32'hbaa1abd4),
	.w6(32'hbc195bea),
	.w7(32'hbc01d80c),
	.w8(32'hbbadfde0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7515c8),
	.w1(32'h3b6a61da),
	.w2(32'hbb76be43),
	.w3(32'h3acc3c7a),
	.w4(32'h3b9e3a82),
	.w5(32'h3b172232),
	.w6(32'h3b41ccef),
	.w7(32'h3bb653cc),
	.w8(32'h3c7d6ec2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47d02c),
	.w1(32'h3bbdbf63),
	.w2(32'hbb46ab87),
	.w3(32'h3c9a5660),
	.w4(32'hbbbe6e9d),
	.w5(32'hbb8e20f0),
	.w6(32'h3c293002),
	.w7(32'hbbb1070e),
	.w8(32'hbc0abdbc),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb066007),
	.w1(32'h3988d28e),
	.w2(32'hbbccecae),
	.w3(32'hbb9c5ec4),
	.w4(32'hbbbbb6a0),
	.w5(32'h3a8d76f7),
	.w6(32'hbbbcaa30),
	.w7(32'hbb736522),
	.w8(32'hbc25bd01),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3dcc2),
	.w1(32'hbaad8718),
	.w2(32'hbc8b3b27),
	.w3(32'hbc09f1da),
	.w4(32'hbc1a9ab9),
	.w5(32'hbc91c5d1),
	.w6(32'h3b5ec0df),
	.w7(32'h3c1d3716),
	.w8(32'hbc974311),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab24ac),
	.w1(32'h3bddf7d2),
	.w2(32'hbbefa203),
	.w3(32'h3b93369d),
	.w4(32'h3c3e3869),
	.w5(32'hbb3052d1),
	.w6(32'h3b9444c0),
	.w7(32'h3c04ae16),
	.w8(32'hbbe34c67),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43e61f),
	.w1(32'h3b8fe1f0),
	.w2(32'hbc3233e2),
	.w3(32'hbbfa233e),
	.w4(32'hba3ad058),
	.w5(32'hba8b2592),
	.w6(32'hbbd491f5),
	.w7(32'hba96cc44),
	.w8(32'hbc01c52c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e8709),
	.w1(32'h39bee5d1),
	.w2(32'h3acec59f),
	.w3(32'h3baacc33),
	.w4(32'h3c2d85c7),
	.w5(32'h3b0dee61),
	.w6(32'h3c0d5231),
	.w7(32'hb8d9e73a),
	.w8(32'h3bb4b5e4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf4711),
	.w1(32'hba5dd402),
	.w2(32'hbca304a3),
	.w3(32'h3a214153),
	.w4(32'hbacd88cf),
	.w5(32'hbc8af6f3),
	.w6(32'hbbf0bfff),
	.w7(32'hbc2fba25),
	.w8(32'hbcc27332),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973a4d),
	.w1(32'h39a1c4f5),
	.w2(32'hb7ad30cd),
	.w3(32'hbc8f13e7),
	.w4(32'hbc58a64a),
	.w5(32'h3c5980ff),
	.w6(32'hbc4e02a7),
	.w7(32'hbc988158),
	.w8(32'h3bfbbac0),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9acfc2),
	.w1(32'h3c75a42c),
	.w2(32'h3ac78714),
	.w3(32'h3cf81b1d),
	.w4(32'h3c8d529c),
	.w5(32'hbab3d4b8),
	.w6(32'h3c50a028),
	.w7(32'h3b302d82),
	.w8(32'hbc10b6cd),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c826b43),
	.w1(32'h3a37bf0c),
	.w2(32'hbb319a45),
	.w3(32'h3c37f7f1),
	.w4(32'hba88fa0e),
	.w5(32'hbc4bb617),
	.w6(32'h3c09cb3a),
	.w7(32'hba891a87),
	.w8(32'hbc1b17e6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4094ee),
	.w1(32'hbc39039e),
	.w2(32'hbc0b992a),
	.w3(32'h3a9eb210),
	.w4(32'h39e24b44),
	.w5(32'h3b39d63a),
	.w6(32'hbb36129b),
	.w7(32'hbbea45d2),
	.w8(32'hbb79b27c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70ec2b),
	.w1(32'h3bb203b2),
	.w2(32'hbc20c559),
	.w3(32'h3c8d3f48),
	.w4(32'h3c6d96d2),
	.w5(32'hbc350cfb),
	.w6(32'h3c164ac3),
	.w7(32'hbba4c15f),
	.w8(32'hbc6078ee),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc993628),
	.w1(32'hba94b4cf),
	.w2(32'hbc0f8872),
	.w3(32'hbcb77a14),
	.w4(32'hbcb343bc),
	.w5(32'h3b83ebb8),
	.w6(32'hbc6241a2),
	.w7(32'hbca0c2fb),
	.w8(32'hbbe01253),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92e107),
	.w1(32'h3be2ad44),
	.w2(32'hbaa97f1d),
	.w3(32'h3c4c049b),
	.w4(32'hbae67cac),
	.w5(32'hbb38b401),
	.w6(32'hbab8f502),
	.w7(32'hbb828390),
	.w8(32'hbb33f889),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a24ec),
	.w1(32'h3b2fb749),
	.w2(32'h3921683e),
	.w3(32'h3be2af91),
	.w4(32'h3c021737),
	.w5(32'h3bccd1d1),
	.w6(32'h3a2cdafd),
	.w7(32'h3b31bc92),
	.w8(32'hbae10082),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c146e40),
	.w1(32'h3b80703e),
	.w2(32'h3b274dcf),
	.w3(32'h3c7137a0),
	.w4(32'h3b3b609e),
	.w5(32'h3c79c58a),
	.w6(32'h3acf3887),
	.w7(32'h3a807bad),
	.w8(32'h3beb9321),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c71a6),
	.w1(32'h3be017aa),
	.w2(32'h3c0a0b48),
	.w3(32'h3b335543),
	.w4(32'hbb0924e7),
	.w5(32'hbb3133b9),
	.w6(32'hbbfa4436),
	.w7(32'h3a807fe7),
	.w8(32'hbc2d6d72),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d4752),
	.w1(32'h3b7e3487),
	.w2(32'h3ba4d0ee),
	.w3(32'h3ab88025),
	.w4(32'h3c4979e6),
	.w5(32'h3bfd9725),
	.w6(32'h3b8e62e5),
	.w7(32'h3c6514ee),
	.w8(32'h3c399b4d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f4fc4),
	.w1(32'h3c68d953),
	.w2(32'hbb664aed),
	.w3(32'h3ad50489),
	.w4(32'h3c181111),
	.w5(32'hbb30d080),
	.w6(32'hbc1d2cd0),
	.w7(32'h3be7b2b7),
	.w8(32'hbbaebfd7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a4169),
	.w1(32'h3af92aeb),
	.w2(32'h3bd76613),
	.w3(32'h3bd79100),
	.w4(32'h3a9dcc3d),
	.w5(32'hbb6965f1),
	.w6(32'hbacb5a9c),
	.w7(32'hbadb7230),
	.w8(32'hbc6231b9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e4db2),
	.w1(32'hba09f9de),
	.w2(32'hbc225328),
	.w3(32'h3acea129),
	.w4(32'hbb0c0075),
	.w5(32'hbc62b461),
	.w6(32'h3b6c0328),
	.w7(32'hbaa01898),
	.w8(32'hbc0a072d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0985d5),
	.w1(32'hbc44f4c4),
	.w2(32'hbae07bf8),
	.w3(32'hbca474ff),
	.w4(32'hbc6db9a7),
	.w5(32'h3c495809),
	.w6(32'hbbb8f9b1),
	.w7(32'hbc586edf),
	.w8(32'hbbce08e1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95ebdd),
	.w1(32'h3b5c275b),
	.w2(32'hbc2a71c2),
	.w3(32'hbb928ef0),
	.w4(32'h3b44f120),
	.w5(32'hbbe0a88a),
	.w6(32'hbb95541f),
	.w7(32'h3b66b518),
	.w8(32'hbc4b72cb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a4bc),
	.w1(32'h3a859e6a),
	.w2(32'hbc181cbd),
	.w3(32'hbb79499c),
	.w4(32'h3aab9bfe),
	.w5(32'hbb8e5a43),
	.w6(32'hbbce8fa1),
	.w7(32'hba2589b8),
	.w8(32'h3c9bf9f2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d6868),
	.w1(32'h3b344192),
	.w2(32'h3c0708ab),
	.w3(32'h3a788ba6),
	.w4(32'h387a4d81),
	.w5(32'h3bb0461c),
	.w6(32'h3c92a86a),
	.w7(32'h3c940599),
	.w8(32'hb9edfa14),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d76f1),
	.w1(32'h3b4ed097),
	.w2(32'hbc9fc8b4),
	.w3(32'h3c36b4f0),
	.w4(32'h3c544215),
	.w5(32'hbc2b3e27),
	.w6(32'hbc011a1d),
	.w7(32'h3b966e51),
	.w8(32'hbc83ff6f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0096c),
	.w1(32'h3b15438d),
	.w2(32'hbbdff725),
	.w3(32'h3c85f71f),
	.w4(32'hb9152636),
	.w5(32'h3b3f58d7),
	.w6(32'h3cc68f62),
	.w7(32'h3c0eb1ab),
	.w8(32'hbb3124a1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52d1dc),
	.w1(32'h3c3953f6),
	.w2(32'h3c33a3f6),
	.w3(32'h3c4b2ce7),
	.w4(32'h3c1b050b),
	.w5(32'h3c88aa42),
	.w6(32'h3c2ffbdf),
	.w7(32'hbb3779d7),
	.w8(32'h3bde6e9f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d1c11),
	.w1(32'h3c2a0e05),
	.w2(32'h3b3a8548),
	.w3(32'h3d0fc475),
	.w4(32'h3cee1508),
	.w5(32'h3c161a54),
	.w6(32'h3cb480c3),
	.w7(32'h3cc50286),
	.w8(32'h3b5366df),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a9cd),
	.w1(32'h3a26ee53),
	.w2(32'hbbee7f3e),
	.w3(32'h3bee132e),
	.w4(32'h3b2753d4),
	.w5(32'hbb604134),
	.w6(32'h3be24f1f),
	.w7(32'h3b5ab13d),
	.w8(32'hbbf53ff2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba47aab),
	.w1(32'h3aa74e63),
	.w2(32'hb98c9d24),
	.w3(32'hbbe1b355),
	.w4(32'hbb2f29ba),
	.w5(32'hba94682a),
	.w6(32'hbb605184),
	.w7(32'hbb6c7330),
	.w8(32'h3a013722),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae05625),
	.w1(32'h3ab8c19e),
	.w2(32'hbb315c10),
	.w3(32'hba2ca4c2),
	.w4(32'hbb912aec),
	.w5(32'hbbc3f941),
	.w6(32'hba924a5b),
	.w7(32'h3b00d500),
	.w8(32'hbba5c4bb),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be79c8),
	.w1(32'h39f8ad9f),
	.w2(32'hbc575687),
	.w3(32'h3a711ef3),
	.w4(32'h3bcc82f2),
	.w5(32'hbd176e01),
	.w6(32'hbb9d47be),
	.w7(32'hb8a4910d),
	.w8(32'hbd15fd58),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1118ec),
	.w1(32'hbcfbadef),
	.w2(32'h3a9c7ec5),
	.w3(32'hbd88e0ab),
	.w4(32'hbd446665),
	.w5(32'h3ca82558),
	.w6(32'hbd568790),
	.w7(32'hbd05ea30),
	.w8(32'h3c4d9a6e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c390977),
	.w1(32'h3c26e0a8),
	.w2(32'h3ba15624),
	.w3(32'h3cf8f238),
	.w4(32'h3cb7ec1e),
	.w5(32'h3a83cc67),
	.w6(32'h3c650195),
	.w7(32'h3c7c995c),
	.w8(32'h3b085a92),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c585456),
	.w1(32'h3b829a2d),
	.w2(32'hbc640776),
	.w3(32'h3c133aaf),
	.w4(32'h3af2a5dd),
	.w5(32'hbc72160e),
	.w6(32'h3a62d483),
	.w7(32'hbb18b764),
	.w8(32'hbca7b6bb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c0b7e),
	.w1(32'hbbeefda3),
	.w2(32'hbc128423),
	.w3(32'h3a84706e),
	.w4(32'hba91bbb0),
	.w5(32'hbbec0b96),
	.w6(32'hbabbc069),
	.w7(32'hbc18ff3a),
	.w8(32'h39f4db2b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e6f6a),
	.w1(32'hbbc958b8),
	.w2(32'hbd07552f),
	.w3(32'hbb3d84c6),
	.w4(32'hbc121412),
	.w5(32'hbd1da70b),
	.w6(32'h3abc28ea),
	.w7(32'h3ae1eed6),
	.w8(32'hbc804911),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3f345a),
	.w1(32'hbcbbb54d),
	.w2(32'hbc4d2e17),
	.w3(32'hbda5f780),
	.w4(32'hbd8694ae),
	.w5(32'h3b8a4da7),
	.w6(32'hbd65f225),
	.w7(32'hbd6fb738),
	.w8(32'hb99e3ff5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83db23),
	.w1(32'h3c2353bf),
	.w2(32'h3aecc010),
	.w3(32'h3d90b46c),
	.w4(32'h3d73c1ab),
	.w5(32'hbaa00634),
	.w6(32'h3d3388aa),
	.w7(32'h3d017e78),
	.w8(32'h37f97ea2),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ecd3e),
	.w1(32'h3ba3c5f7),
	.w2(32'h3b4159f2),
	.w3(32'h3b1b25e8),
	.w4(32'h3b2c3b2b),
	.w5(32'h3ae6a66a),
	.w6(32'hbbb6ad27),
	.w7(32'hbb7359b3),
	.w8(32'hbb3913e3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfd27c),
	.w1(32'h3b983e43),
	.w2(32'h3bb0b2f2),
	.w3(32'h3c0fb570),
	.w4(32'h3c0c247d),
	.w5(32'h3cc733a4),
	.w6(32'h3ace1955),
	.w7(32'hba8d183d),
	.w8(32'h3c47159d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c569c4f),
	.w1(32'h3c3e4512),
	.w2(32'h3bda5403),
	.w3(32'h3d4929bb),
	.w4(32'h3d1012db),
	.w5(32'h3c6be6d7),
	.w6(32'h3d287a23),
	.w7(32'h3cbe19a9),
	.w8(32'hb9692557),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c42cb),
	.w1(32'h3c0ecdcd),
	.w2(32'h3b340111),
	.w3(32'h3d076d4e),
	.w4(32'h3cc32ab0),
	.w5(32'h3c08f238),
	.w6(32'h3ce1dd36),
	.w7(32'h3c949d2a),
	.w8(32'h3becc5d8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d845e),
	.w1(32'h3aa25f83),
	.w2(32'hbb2e0b35),
	.w3(32'h3c995573),
	.w4(32'h38ca766c),
	.w5(32'hbb567b30),
	.w6(32'h3c42aa91),
	.w7(32'hbb7a5875),
	.w8(32'hbc1899b9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bace31f),
	.w1(32'hba54f78a),
	.w2(32'hbc2af25a),
	.w3(32'h3bdc5b9b),
	.w4(32'hbb02b08d),
	.w5(32'hbb58577d),
	.w6(32'hb8e5e502),
	.w7(32'hbb99584b),
	.w8(32'hbab3c117),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c5614),
	.w1(32'h3bf11c9d),
	.w2(32'hbbf5b5e2),
	.w3(32'h3b40a90c),
	.w4(32'h39cd6f1b),
	.w5(32'hbb660e50),
	.w6(32'hbbaf784b),
	.w7(32'hbba8160c),
	.w8(32'hbc4ffddd),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85b172),
	.w1(32'hbac607b8),
	.w2(32'hbb834fd3),
	.w3(32'hba949de9),
	.w4(32'hbb4a356e),
	.w5(32'h3b46d78c),
	.w6(32'h3a888a1d),
	.w7(32'hbb487689),
	.w8(32'h39fcc3ee),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15c706),
	.w1(32'h3b12dcca),
	.w2(32'h3c1f50bb),
	.w3(32'hbcc48b05),
	.w4(32'hbcc399ff),
	.w5(32'h3a581e9a),
	.w6(32'hbc9e1f09),
	.w7(32'hbc19c34a),
	.w8(32'h3c5da4c0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b8efb),
	.w1(32'hbb84d38c),
	.w2(32'hbc944067),
	.w3(32'h3c6ef92e),
	.w4(32'h3bf1f781),
	.w5(32'hbcafb77c),
	.w6(32'hbc4d9121),
	.w7(32'h3a5e331b),
	.w8(32'hbc869571),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc216e8a),
	.w1(32'hbc2a1798),
	.w2(32'hbc5b2fce),
	.w3(32'hbd2368f4),
	.w4(32'hbcda3d17),
	.w5(32'hbc3cfa3d),
	.w6(32'hbd11e11c),
	.w7(32'hbd00b8d8),
	.w8(32'hbcc3a8c0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a1092),
	.w1(32'hbbff668f),
	.w2(32'hb99c24d0),
	.w3(32'hbc641416),
	.w4(32'hbb2c991d),
	.w5(32'h3ba666f6),
	.w6(32'hbc82fa71),
	.w7(32'hbb079e69),
	.w8(32'hbaa75c06),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed4a3),
	.w1(32'hbb37ac74),
	.w2(32'h3c27fd00),
	.w3(32'h3a536a10),
	.w4(32'hbc4a54c1),
	.w5(32'h3ac9a256),
	.w6(32'hb9ab0173),
	.w7(32'hbb8c9cf8),
	.w8(32'h3b28772b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39838015),
	.w1(32'hba1148ab),
	.w2(32'h3c0be808),
	.w3(32'h3a406912),
	.w4(32'hbacf4c91),
	.w5(32'h3c793545),
	.w6(32'hbb899016),
	.w7(32'hba737b85),
	.w8(32'h3bb4944e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c463999),
	.w1(32'h3b87771a),
	.w2(32'hbbba705f),
	.w3(32'h3bc911c5),
	.w4(32'h3b9a90b3),
	.w5(32'hbc67d756),
	.w6(32'h3b38ad5b),
	.w7(32'h3c4a4e37),
	.w8(32'hbbcc804a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe29719),
	.w1(32'hbb97cde8),
	.w2(32'hbc33bd7e),
	.w3(32'hbcc91f8e),
	.w4(32'hbc7c58a4),
	.w5(32'hbcadd408),
	.w6(32'hbd07f86f),
	.w7(32'hbc1f27c6),
	.w8(32'hbbf1e598),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb643aae),
	.w1(32'h3b8bb9c8),
	.w2(32'hbcbda246),
	.w3(32'h3b36a4a5),
	.w4(32'h3bc18920),
	.w5(32'hbc28045c),
	.w6(32'hbb6055fd),
	.w7(32'hbb81676c),
	.w8(32'hbc815525),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc217d5d),
	.w1(32'hbbe394cc),
	.w2(32'h3b18d5d9),
	.w3(32'hba3ef93a),
	.w4(32'hbb14adf4),
	.w5(32'hbaf005e9),
	.w6(32'hbc3e71ae),
	.w7(32'hbabb64ad),
	.w8(32'hbbf52e0c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2d194),
	.w1(32'h3bcfa41c),
	.w2(32'h3b86a842),
	.w3(32'h3c4020b5),
	.w4(32'hbab6c54a),
	.w5(32'hbb900c96),
	.w6(32'h3c1dc26c),
	.w7(32'hbba7c04d),
	.w8(32'hbc285cb6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ffeca),
	.w1(32'h3b87d6cd),
	.w2(32'h3ae9c0dd),
	.w3(32'h3c485a91),
	.w4(32'h3c0558e8),
	.w5(32'h3c867288),
	.w6(32'h3c10e2ca),
	.w7(32'hb9235365),
	.w8(32'h3b89a7f9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51e14e),
	.w1(32'h3c68cd51),
	.w2(32'hbafad1b4),
	.w3(32'h3cb24eba),
	.w4(32'h3ca74cbf),
	.w5(32'h3bc093df),
	.w6(32'h3c7ef000),
	.w7(32'h3c163e5a),
	.w8(32'h3b28d741),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cbe33),
	.w1(32'h3c087b98),
	.w2(32'h3b60483d),
	.w3(32'h3c3b5db8),
	.w4(32'h3c5b322f),
	.w5(32'h3c1f679d),
	.w6(32'h3c2004bd),
	.w7(32'hbb8fb177),
	.w8(32'hb9f4a15f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18b376),
	.w1(32'h3c0b50b3),
	.w2(32'h3c676a03),
	.w3(32'h3c2e407b),
	.w4(32'h3b85a235),
	.w5(32'h3cdba4a8),
	.w6(32'h3bbe59a7),
	.w7(32'h3b4a3733),
	.w8(32'h3c2e0f6b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c732d5b),
	.w1(32'h3c8ca468),
	.w2(32'h3c1608bc),
	.w3(32'h3d20144e),
	.w4(32'h3cc45730),
	.w5(32'h3c9f1afb),
	.w6(32'h3ca54343),
	.w7(32'h3cb949c1),
	.w8(32'h3c170623),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e38b5),
	.w1(32'h3baac43b),
	.w2(32'hbc3127ba),
	.w3(32'h3cb7b613),
	.w4(32'h3c524019),
	.w5(32'hbc4cf487),
	.w6(32'h3c89ac4c),
	.w7(32'h3be6dd6e),
	.w8(32'hbc19b386),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6d452),
	.w1(32'h3b7a6221),
	.w2(32'hbc7e29b6),
	.w3(32'hbc09a395),
	.w4(32'h3c92f882),
	.w5(32'hbc309451),
	.w6(32'hbc3f6fee),
	.w7(32'h3a52384a),
	.w8(32'hbc1e6cd4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d12b0),
	.w1(32'hbbe07f5d),
	.w2(32'hbc44537a),
	.w3(32'hbcb00d70),
	.w4(32'hbc8039d4),
	.w5(32'hbcb4510a),
	.w6(32'hbbb7e7e1),
	.w7(32'hbc4034bb),
	.w8(32'hbc9171b6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889f46),
	.w1(32'hbb03075d),
	.w2(32'hbb8310d8),
	.w3(32'hbce84855),
	.w4(32'hbc9f74a8),
	.w5(32'hbae44ca5),
	.w6(32'hbc2cb964),
	.w7(32'hbc0122f7),
	.w8(32'hbbe048cf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71ecf6),
	.w1(32'hba72cc54),
	.w2(32'hbc00c26e),
	.w3(32'hbb90ea0a),
	.w4(32'hbbe55ebc),
	.w5(32'hbbae55ff),
	.w6(32'hbcb06cd3),
	.w7(32'hbbfd11ac),
	.w8(32'hbc2965df),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392be3),
	.w1(32'h3b9e380c),
	.w2(32'hba99ab3e),
	.w3(32'h3b045867),
	.w4(32'h3b8f9468),
	.w5(32'hbc2de512),
	.w6(32'hbc0dc9d9),
	.w7(32'hbb197ef6),
	.w8(32'hbb99c0d7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ed9df),
	.w1(32'hba18e427),
	.w2(32'h3a8be156),
	.w3(32'hbca112b3),
	.w4(32'hbc979e43),
	.w5(32'h3b2f5cfc),
	.w6(32'hbc4319a5),
	.w7(32'hbc30e109),
	.w8(32'h3b8d4741),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85c14c),
	.w1(32'h3bd43551),
	.w2(32'h39de3ee1),
	.w3(32'h3b5f0fa5),
	.w4(32'h3a2594ba),
	.w5(32'h3affd7f8),
	.w6(32'hbb7437ab),
	.w7(32'hba235768),
	.w8(32'h3a6eea73),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a431e14),
	.w1(32'h3ad75c34),
	.w2(32'hba865aa5),
	.w3(32'hbb087898),
	.w4(32'hbbbe11e9),
	.w5(32'h3bb82c5e),
	.w6(32'hba92d66c),
	.w7(32'h3ac1abb7),
	.w8(32'h3b582c88),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82b8a9),
	.w1(32'h3b0179f2),
	.w2(32'hbba81401),
	.w3(32'h3bb67ca3),
	.w4(32'h3c0f047f),
	.w5(32'hbc82e43a),
	.w6(32'h3b9454f0),
	.w7(32'h3b7fdcf8),
	.w8(32'hbc68a9e7),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71e591),
	.w1(32'hbbb2c516),
	.w2(32'hbbb0f85f),
	.w3(32'hbcf5c789),
	.w4(32'hbc799f4c),
	.w5(32'hbba55a3f),
	.w6(32'hbc8e5e36),
	.w7(32'hbca8e463),
	.w8(32'h3b78d7db),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc80b33),
	.w1(32'h3a595a5a),
	.w2(32'h3ca91523),
	.w3(32'hbc512f59),
	.w4(32'hbc2a0597),
	.w5(32'h3cdf2fff),
	.w6(32'hbb017a6c),
	.w7(32'hbb7ec58b),
	.w8(32'h3ca27e5f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb7bbf),
	.w1(32'h3ca58986),
	.w2(32'h3b85395d),
	.w3(32'h3d443f85),
	.w4(32'h3d0657b7),
	.w5(32'h3b89b947),
	.w6(32'h3d011b4e),
	.w7(32'h3c92ac14),
	.w8(32'hb9d7505b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d5110),
	.w1(32'h3ba14473),
	.w2(32'hbc473912),
	.w3(32'h3a005fe9),
	.w4(32'hbbbd62e9),
	.w5(32'hbb98ee36),
	.w6(32'h3bb1791b),
	.w7(32'h3b13632c),
	.w8(32'hbbeae100),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc6d1c),
	.w1(32'hbad00133),
	.w2(32'h39c78e6e),
	.w3(32'h3b114779),
	.w4(32'h3a69b8a9),
	.w5(32'h3c1a4e97),
	.w6(32'hbbdb1bc8),
	.w7(32'hbc1eb8d5),
	.w8(32'hb8013ceb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c826c8c),
	.w1(32'h3be00f0c),
	.w2(32'hbc3ab738),
	.w3(32'h3cb030ec),
	.w4(32'h3c53ed17),
	.w5(32'hbbe0aced),
	.w6(32'h3b98905d),
	.w7(32'hb9efb6b6),
	.w8(32'hbc15505a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf33bd),
	.w1(32'hbba416aa),
	.w2(32'h3ba4a94e),
	.w3(32'hba8b0f24),
	.w4(32'hbc088b1f),
	.w5(32'hbae89239),
	.w6(32'h3b788a6a),
	.w7(32'hbbc6e959),
	.w8(32'h3b341c3d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d125a),
	.w1(32'h3aedfa30),
	.w2(32'hbc313faf),
	.w3(32'h3b7b4ac7),
	.w4(32'h3bbf4e51),
	.w5(32'hbc1d637c),
	.w6(32'h3b9787b6),
	.w7(32'h3bbb224b),
	.w8(32'hbc45c6c9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b385646),
	.w1(32'h3bf673a4),
	.w2(32'hb95709e3),
	.w3(32'h3af2f073),
	.w4(32'hbad8e2ea),
	.w5(32'hbba1bbb0),
	.w6(32'h3b8815b3),
	.w7(32'h3aacb62b),
	.w8(32'h3bc6f4b9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace81ab),
	.w1(32'hb88c930a),
	.w2(32'h3bf42e20),
	.w3(32'hbacd40a0),
	.w4(32'h3a851132),
	.w5(32'h3be7aba1),
	.w6(32'h3b548f43),
	.w7(32'h3bcd8213),
	.w8(32'h3c51036f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2534c),
	.w1(32'h3a2e44c3),
	.w2(32'hbc80bdce),
	.w3(32'h3c13cc87),
	.w4(32'h3accc1a9),
	.w5(32'hbcb988ad),
	.w6(32'h3bdb515c),
	.w7(32'h3c0b5b01),
	.w8(32'hbc995524),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12c3cc),
	.w1(32'hbbf99363),
	.w2(32'h3c8053e9),
	.w3(32'hbcd6a472),
	.w4(32'hbcdc3b4e),
	.w5(32'h3cbd4e00),
	.w6(32'hbca44a27),
	.w7(32'hbc547e23),
	.w8(32'h3c8778e2),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac27ba),
	.w1(32'h3bfb8d1d),
	.w2(32'hbb764a51),
	.w3(32'h3d51be12),
	.w4(32'h3d049c11),
	.w5(32'hbb47f789),
	.w6(32'h3cef3bb0),
	.w7(32'h3ccd6f4f),
	.w8(32'hba9bafbc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbacd6b),
	.w1(32'hbb7f5b2c),
	.w2(32'hbbf9969d),
	.w3(32'hbbc6c888),
	.w4(32'hba82c528),
	.w5(32'hbbf862f9),
	.w6(32'hbaf4f886),
	.w7(32'h3b443ba3),
	.w8(32'hbb297482),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25576b),
	.w1(32'hbb1bf270),
	.w2(32'h3ae98bc3),
	.w3(32'hbbac2409),
	.w4(32'hbb110ea8),
	.w5(32'h3c69ec0d),
	.w6(32'hb94fc5bc),
	.w7(32'hbadfd091),
	.w8(32'h3c0dbffa),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18adc7),
	.w1(32'hb832942c),
	.w2(32'hbb9a0abc),
	.w3(32'h3ca7ae2f),
	.w4(32'hbb90ecc4),
	.w5(32'hbbceb1a9),
	.w6(32'h3c9c549c),
	.w7(32'h3a85bb32),
	.w8(32'hbb33a73a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd6d40),
	.w1(32'hba947260),
	.w2(32'h3c0d97c0),
	.w3(32'hba5ec821),
	.w4(32'h3b1d21f7),
	.w5(32'h3bd5d9f1),
	.w6(32'hba2bed4e),
	.w7(32'h3aa70701),
	.w8(32'hb79c9303),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b916608),
	.w1(32'h3bf30573),
	.w2(32'hbcf4ed7e),
	.w3(32'h3bb10c8f),
	.w4(32'h3c5760e4),
	.w5(32'hbcda4847),
	.w6(32'h3bd89cdd),
	.w7(32'h3bc8a34d),
	.w8(32'hbcbeb42d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ff5d6),
	.w1(32'hbcdf76c2),
	.w2(32'hbca7f7d2),
	.w3(32'hbd933062),
	.w4(32'hbd62b6cd),
	.w5(32'hbd39a04b),
	.w6(32'hbd4d9f80),
	.w7(32'hbd0bbda1),
	.w8(32'hbd1eb49e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd251897),
	.w1(32'hbcff6470),
	.w2(32'h3af49889),
	.w3(32'hbdc76cd7),
	.w4(32'hbd859528),
	.w5(32'h3be198b2),
	.w6(32'hbda2a386),
	.w7(32'hbd4e4e4b),
	.w8(32'hbbac7a96),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule