module layer_10_featuremap_440(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e783d7),
	.w1(32'hb6460aa2),
	.w2(32'h39da1abf),
	.w3(32'hb9ebf9dd),
	.w4(32'h3a1eaedb),
	.w5(32'h3aba55cd),
	.w6(32'hb92ef0a6),
	.w7(32'h39f86f9a),
	.w8(32'h3a71b539),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8251f7),
	.w1(32'hbb1d6c58),
	.w2(32'hbb40d9d1),
	.w3(32'hb9b831fe),
	.w4(32'hb9e420f7),
	.w5(32'hbaba1977),
	.w6(32'hb964d9b6),
	.w7(32'h3a844d59),
	.w8(32'hba808dd2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39218ab9),
	.w1(32'hbb2027ce),
	.w2(32'hba921c8a),
	.w3(32'h38a4a814),
	.w4(32'hbb2ccf88),
	.w5(32'hbb1b5791),
	.w6(32'h38b168db),
	.w7(32'hba320674),
	.w8(32'hb970e72d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffde40),
	.w1(32'h3acab69a),
	.w2(32'h3ac79455),
	.w3(32'hbaf7c8d6),
	.w4(32'h3b043fc2),
	.w5(32'h3a80f097),
	.w6(32'hbaff6cf0),
	.w7(32'h3a03d814),
	.w8(32'hba818d46),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9864863),
	.w1(32'h3a562d91),
	.w2(32'h3a0fe9fe),
	.w3(32'hb92dc083),
	.w4(32'h3a1c99a6),
	.w5(32'h398252e0),
	.w6(32'h36c8b2ca),
	.w7(32'hba156995),
	.w8(32'h380385d9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43c762),
	.w1(32'hb909d6aa),
	.w2(32'hba92354f),
	.w3(32'h3724fe7b),
	.w4(32'hb9c9ad47),
	.w5(32'hbaef86fe),
	.w6(32'h39309791),
	.w7(32'hba1b68b6),
	.w8(32'hbab24b59),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae5c2a),
	.w1(32'h3b316b6b),
	.w2(32'h3b6f0174),
	.w3(32'hbb078967),
	.w4(32'h3a6a3f09),
	.w5(32'h3bcb0f0e),
	.w6(32'h3a6046fc),
	.w7(32'h37d93acc),
	.w8(32'h3af28f6e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88caaa),
	.w1(32'h3c0863c0),
	.w2(32'hba41e77e),
	.w3(32'h3c59ac5d),
	.w4(32'h3b606b9a),
	.w5(32'hb8c1dcea),
	.w6(32'h3c8887e9),
	.w7(32'h3bbbdcc2),
	.w8(32'hbb67c946),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c663f6),
	.w1(32'h39a703ea),
	.w2(32'h3b096944),
	.w3(32'hb8cbd53c),
	.w4(32'h3a2ed1f9),
	.w5(32'h3b341a52),
	.w6(32'h3a632eee),
	.w7(32'h3a22d20d),
	.w8(32'h3b0de70e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4de8b2),
	.w1(32'hbae27f8a),
	.w2(32'hbb4c7e40),
	.w3(32'h3b3751f9),
	.w4(32'h3a7b5a3a),
	.w5(32'h3b11c3df),
	.w6(32'h3bc85c07),
	.w7(32'h39e0950e),
	.w8(32'h3a61bf5c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fd898),
	.w1(32'hba3bff1a),
	.w2(32'h3743c74f),
	.w3(32'hb8970330),
	.w4(32'hb8eab3cb),
	.w5(32'h3a7dd26c),
	.w6(32'hb9fb3732),
	.w7(32'hbaf1f2c8),
	.w8(32'hbaaa5040),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bfc74),
	.w1(32'h3af2780b),
	.w2(32'h3a909649),
	.w3(32'hbb87156e),
	.w4(32'h3b260a1c),
	.w5(32'h3b33b240),
	.w6(32'hbb10f40f),
	.w7(32'hba99cbfd),
	.w8(32'hb92b5ad4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d1fc5),
	.w1(32'hb9a3216b),
	.w2(32'hbb0b95b0),
	.w3(32'h3ab123f9),
	.w4(32'hb9475c98),
	.w5(32'h3aa568b4),
	.w6(32'h3b69e889),
	.w7(32'h3a0dd085),
	.w8(32'h3a2112d9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95d7b3),
	.w1(32'h3ad15877),
	.w2(32'h3afe30e8),
	.w3(32'h3aaae4d4),
	.w4(32'h3a93b06f),
	.w5(32'hb9cd8049),
	.w6(32'h3a35cf72),
	.w7(32'hb9c85742),
	.w8(32'h3761f8da),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9bbfa),
	.w1(32'hbb6db46a),
	.w2(32'hbb73b85d),
	.w3(32'h3ae74a52),
	.w4(32'h37af8f9c),
	.w5(32'hbb196e8f),
	.w6(32'h3b0f06b1),
	.w7(32'h3a0472b6),
	.w8(32'hbacc158a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a71c1),
	.w1(32'hbb10b069),
	.w2(32'hba9b224c),
	.w3(32'h3b5bdd09),
	.w4(32'h3b682b04),
	.w5(32'hbb083c09),
	.w6(32'h3bb0a5dc),
	.w7(32'h3b2b6be2),
	.w8(32'h39cb719e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b29e3),
	.w1(32'hb95d9fce),
	.w2(32'hb95c7ec5),
	.w3(32'hb9de7d63),
	.w4(32'h3a2431bd),
	.w5(32'h38d6d905),
	.w6(32'hb7891eb3),
	.w7(32'hb9c1adae),
	.w8(32'hb9cc648f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58beeb),
	.w1(32'h3c22cdec),
	.w2(32'h3c0ee1e9),
	.w3(32'h3c68019f),
	.w4(32'h3c01b4c6),
	.w5(32'h3b3f0539),
	.w6(32'h3c86feaa),
	.w7(32'h3b8a194d),
	.w8(32'hbb15a67b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d2c45),
	.w1(32'h3b4d6c47),
	.w2(32'h3a428882),
	.w3(32'h3b827da6),
	.w4(32'h3afa2c1d),
	.w5(32'h3a9908e4),
	.w6(32'h3bebdae5),
	.w7(32'h3b3af35a),
	.w8(32'h3a68a2c3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b7632),
	.w1(32'hb9f69c67),
	.w2(32'h3996d3a3),
	.w3(32'h399a33a3),
	.w4(32'hba929254),
	.w5(32'hb9f26128),
	.w6(32'h3974f81c),
	.w7(32'hba57bd74),
	.w8(32'hba9bfdb8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994cf77),
	.w1(32'hb88881da),
	.w2(32'hb9cc8f32),
	.w3(32'h3a14353d),
	.w4(32'hb84dead6),
	.w5(32'hbadef67c),
	.w6(32'h3aa61bb3),
	.w7(32'hb93d009d),
	.w8(32'hbab18457),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91969ac),
	.w1(32'hb985a020),
	.w2(32'hb9c69636),
	.w3(32'hbae2509c),
	.w4(32'hba08a1fa),
	.w5(32'hb9249d61),
	.w6(32'hbb09a9d7),
	.w7(32'h3a0653a8),
	.w8(32'h39b6797a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabfcde),
	.w1(32'h3c50a2a4),
	.w2(32'hb603a9ca),
	.w3(32'h3cbc66f8),
	.w4(32'h3c26348e),
	.w5(32'hba5f7c44),
	.w6(32'h3cd9f154),
	.w7(32'h3c3f9f84),
	.w8(32'h3a0282d4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77a461),
	.w1(32'hbb32152a),
	.w2(32'hbbbe3bdb),
	.w3(32'hba7ef5a5),
	.w4(32'hbae21d1a),
	.w5(32'hbb8138bb),
	.w6(32'h3b02ea5e),
	.w7(32'h39a69ed7),
	.w8(32'hb9fba07c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ed7c),
	.w1(32'hbb695fef),
	.w2(32'hbba23e90),
	.w3(32'hbbc9a2ff),
	.w4(32'hbb098611),
	.w5(32'hbb3bc3dd),
	.w6(32'hbb11f565),
	.w7(32'h3bd36b92),
	.w8(32'h3b92838b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74e0be),
	.w1(32'h3ab5e86b),
	.w2(32'h3a0bdfe5),
	.w3(32'hba9e891e),
	.w4(32'h3a9236de),
	.w5(32'hbae01bd8),
	.w6(32'hb9ee4b9d),
	.w7(32'h3a94b0fb),
	.w8(32'h39c139d6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a998643),
	.w1(32'h3ab25231),
	.w2(32'h3a74b70f),
	.w3(32'h3aa4751c),
	.w4(32'h3afa6044),
	.w5(32'h3a4f3e40),
	.w6(32'h3ae68e67),
	.w7(32'h3a8fd07b),
	.w8(32'h3a09fa3f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394963b4),
	.w1(32'hbb27f0b4),
	.w2(32'h3b022483),
	.w3(32'hbba575e1),
	.w4(32'hbaa8dff9),
	.w5(32'h3c021a74),
	.w6(32'hbbcb2efc),
	.w7(32'hbbac3e15),
	.w8(32'h3a53b197),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9e2da),
	.w1(32'h3a202037),
	.w2(32'h3a8aa12d),
	.w3(32'hbaeedee0),
	.w4(32'hb7c7e317),
	.w5(32'h3ac3dad7),
	.w6(32'hbb581403),
	.w7(32'hbb0ced77),
	.w8(32'hbaaf23ce),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f5f72),
	.w1(32'hbb2d5c8c),
	.w2(32'hbb284179),
	.w3(32'hbb8dedc4),
	.w4(32'h3a5c8b44),
	.w5(32'h3a3581ab),
	.w6(32'hbbbe3e9a),
	.w7(32'hba3ba777),
	.w8(32'h3a5010e5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28c514),
	.w1(32'hbacbb1f1),
	.w2(32'hbad4e4a7),
	.w3(32'h39ee8aa6),
	.w4(32'hbac78bc0),
	.w5(32'hba69f0f7),
	.w6(32'hb97af6d5),
	.w7(32'hba4de199),
	.w8(32'hba604fbc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfa78a),
	.w1(32'hb8f65d40),
	.w2(32'h38aed845),
	.w3(32'hb9f94e2d),
	.w4(32'h398fac9b),
	.w5(32'h38d09992),
	.w6(32'hb9e35c1a),
	.w7(32'h3a2b7cb6),
	.w8(32'hb592d7c5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af77566),
	.w1(32'hbab2e8c2),
	.w2(32'hbb3737a3),
	.w3(32'h3ac6d347),
	.w4(32'hbaab9ccf),
	.w5(32'hbb2a759c),
	.w6(32'h3b62f6a1),
	.w7(32'h39ffbef4),
	.w8(32'hbad77068),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c3f38),
	.w1(32'hba938e87),
	.w2(32'hbb1f3c77),
	.w3(32'hbb251359),
	.w4(32'hba292f3c),
	.w5(32'hba8d242e),
	.w6(32'h38db5e7a),
	.w7(32'h3ab42609),
	.w8(32'hb8e05e1e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba109817),
	.w1(32'hbac1fd7c),
	.w2(32'hbac89011),
	.w3(32'hb9dd8f86),
	.w4(32'hbae212fd),
	.w5(32'hbb5b82d4),
	.w6(32'hb9d576d6),
	.w7(32'hb9d9220f),
	.w8(32'hba4c9de3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16f285),
	.w1(32'h3b3d3f64),
	.w2(32'h3911e7b0),
	.w3(32'h3b15fe87),
	.w4(32'h3b01a150),
	.w5(32'h3a83913b),
	.w6(32'h3b863d59),
	.w7(32'h3b148594),
	.w8(32'h39eb46fc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57d0ad),
	.w1(32'h3abd78c3),
	.w2(32'hbb969810),
	.w3(32'h3b29e6c5),
	.w4(32'h3b663814),
	.w5(32'hbbda2e47),
	.w6(32'h3c5eb6b0),
	.w7(32'h3bf42fac),
	.w8(32'hbbb72a99),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5edd2d),
	.w1(32'hbb418071),
	.w2(32'hbb8802c2),
	.w3(32'hbbf6a810),
	.w4(32'hbaca6dbb),
	.w5(32'hbac3ec4a),
	.w6(32'hbc11332d),
	.w7(32'h3af295b0),
	.w8(32'hba869b86),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba10244),
	.w1(32'hbb602cbe),
	.w2(32'h39c059f8),
	.w3(32'hbc41aecf),
	.w4(32'hba318090),
	.w5(32'h3c0217a0),
	.w6(32'hbc740b09),
	.w7(32'hbb1e3ee5),
	.w8(32'h3b8ff1c4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa73d29),
	.w1(32'hba724c1e),
	.w2(32'hbac6e1ce),
	.w3(32'hbb065ced),
	.w4(32'hb97f469e),
	.w5(32'hba520847),
	.w6(32'hbac5863e),
	.w7(32'h3a8d37b4),
	.w8(32'hb98732f5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6c5a6),
	.w1(32'h39696745),
	.w2(32'h3a08550d),
	.w3(32'h3a3194d1),
	.w4(32'hb89ab492),
	.w5(32'h3a13fe4b),
	.w6(32'h39809490),
	.w7(32'h3906b24c),
	.w8(32'h3a59964e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9595dd),
	.w1(32'hb9ba15ae),
	.w2(32'hb98b44e1),
	.w3(32'h3a100ef5),
	.w4(32'hba173919),
	.w5(32'h38f39ec1),
	.w6(32'h391638c2),
	.w7(32'hba56765c),
	.w8(32'h38e6d64e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1311c1),
	.w1(32'h3a1d1daa),
	.w2(32'hba396e1b),
	.w3(32'hba066518),
	.w4(32'h39ceb88e),
	.w5(32'hb96711cb),
	.w6(32'hb98eae75),
	.w7(32'h3a16a6a5),
	.w8(32'hbaddf3d8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4aa910),
	.w1(32'hba5d3083),
	.w2(32'h3b5d2eaf),
	.w3(32'h3b0f524f),
	.w4(32'h3ab2ec1c),
	.w5(32'h3992242e),
	.w6(32'h3b392782),
	.w7(32'hbb422d48),
	.w8(32'h3ab36298),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c86b69),
	.w1(32'hba38473c),
	.w2(32'hbac6d697),
	.w3(32'hb9951552),
	.w4(32'h39744bd1),
	.w5(32'h3b0c4599),
	.w6(32'h3b126b7d),
	.w7(32'h3b58e47f),
	.w8(32'h3b4b97a2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b115f30),
	.w1(32'hbb828ea9),
	.w2(32'hbc03e095),
	.w3(32'hb9ae5701),
	.w4(32'hbb125508),
	.w5(32'hbb580121),
	.w6(32'h3bbc1669),
	.w7(32'h3b3afe8a),
	.w8(32'h38f9fe2f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbe1b6),
	.w1(32'h3b584608),
	.w2(32'h38e9b8ce),
	.w3(32'h3b81d27d),
	.w4(32'h3b6f0a03),
	.w5(32'hbace0dd6),
	.w6(32'h3c25f9fc),
	.w7(32'h3b94e2f5),
	.w8(32'h3b15cf72),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d9a85),
	.w1(32'h3c39ca08),
	.w2(32'h3bdda55a),
	.w3(32'h3c33ec4c),
	.w4(32'h3b4ec4d2),
	.w5(32'h3a5966c4),
	.w6(32'h3c957936),
	.w7(32'h3b8a979a),
	.w8(32'hbb8257c0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a8fcc),
	.w1(32'h38b7f920),
	.w2(32'h3ae0bc09),
	.w3(32'hbb2885e4),
	.w4(32'hb9938685),
	.w5(32'hba313fcd),
	.w6(32'hbb01fe8d),
	.w7(32'hb8c0d0d1),
	.w8(32'h3ac7944d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c8cdc),
	.w1(32'h3af502b7),
	.w2(32'h3b5cbe24),
	.w3(32'h3b094a12),
	.w4(32'h3af8a05c),
	.w5(32'h3ada6726),
	.w6(32'h3b135ddc),
	.w7(32'h3b53237b),
	.w8(32'h3b72238f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56bb7b),
	.w1(32'hba60c2f4),
	.w2(32'hba7817a2),
	.w3(32'hb91b3cb7),
	.w4(32'hbafe1b4e),
	.w5(32'h3862ce99),
	.w6(32'hba582444),
	.w7(32'hba80e089),
	.w8(32'h3a60bda6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1faa36),
	.w1(32'h3b140d59),
	.w2(32'h3ab7dbcd),
	.w3(32'h3b3088da),
	.w4(32'h3abaea53),
	.w5(32'h3ad4a4f1),
	.w6(32'h3b29a229),
	.w7(32'h3b2ca827),
	.w8(32'h3b22ebdc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0be625),
	.w1(32'h3af22524),
	.w2(32'h3acd1231),
	.w3(32'h3b0edb3b),
	.w4(32'h3a58a317),
	.w5(32'hba221118),
	.w6(32'h3b70ffe8),
	.w7(32'h3ac44330),
	.w8(32'h3a2281d4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b9047),
	.w1(32'h3c02da04),
	.w2(32'h3b1fba12),
	.w3(32'h3c04a113),
	.w4(32'h3b6f98b3),
	.w5(32'hba308ed5),
	.w6(32'h3c73b6f4),
	.w7(32'h3bcb7c77),
	.w8(32'hbac839e6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b599b),
	.w1(32'h3b50ee7d),
	.w2(32'h3b75b39e),
	.w3(32'h3a5ba286),
	.w4(32'h3a59dd65),
	.w5(32'h3b14681d),
	.w6(32'h3a807dbc),
	.w7(32'h3ab56f48),
	.w8(32'h3af31a7e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946f832),
	.w1(32'h3a43339b),
	.w2(32'h3a3580cb),
	.w3(32'h3a5943c2),
	.w4(32'h3a5bb4dd),
	.w5(32'hb9ecd6b8),
	.w6(32'h39c891e1),
	.w7(32'h3a0be35c),
	.w8(32'hba965011),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08fefd),
	.w1(32'hba006216),
	.w2(32'hbaa3bfa1),
	.w3(32'h3a197dc6),
	.w4(32'h39340bdf),
	.w5(32'hba2e6bc8),
	.w6(32'hb906d9e3),
	.w7(32'hb969a7ce),
	.w8(32'hba83ed1e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba985346),
	.w1(32'h3a13b6f8),
	.w2(32'h39c81321),
	.w3(32'hba4767f0),
	.w4(32'h39363937),
	.w5(32'h3a85f74e),
	.w6(32'hbab48622),
	.w7(32'hb9430f57),
	.w8(32'h399b6ffc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2086d),
	.w1(32'hba237234),
	.w2(32'hba8f31d8),
	.w3(32'h38e0c016),
	.w4(32'hb9fd8e81),
	.w5(32'hba7406dd),
	.w6(32'hb7eb0be8),
	.w7(32'hb972002a),
	.w8(32'hba24ce32),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab94f1c),
	.w1(32'h3a27189c),
	.w2(32'h3a71c57f),
	.w3(32'hbadd6a19),
	.w4(32'h395d7308),
	.w5(32'h3a81a44c),
	.w6(32'hbabbb223),
	.w7(32'h3a89c203),
	.w8(32'h3ac471e5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407f02),
	.w1(32'h3b7f593a),
	.w2(32'h3b0c32e1),
	.w3(32'h3b830426),
	.w4(32'h3b5cac10),
	.w5(32'h3aa906c7),
	.w6(32'h3bbc7559),
	.w7(32'h3b51a9d6),
	.w8(32'h3b45fd0c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08da89),
	.w1(32'h3a874a0e),
	.w2(32'h3b4119e3),
	.w3(32'h3bbb3ad0),
	.w4(32'h3ad9784b),
	.w5(32'h3b45d235),
	.w6(32'h3b6b5a8e),
	.w7(32'hb9d2d127),
	.w8(32'h3b1a757a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9987064),
	.w1(32'h3a20a9ab),
	.w2(32'hb86d829c),
	.w3(32'hba655870),
	.w4(32'h3a3dbd84),
	.w5(32'h39316ce4),
	.w6(32'hba566e92),
	.w7(32'h39d79b69),
	.w8(32'hba545cbe),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fc008),
	.w1(32'hb8befc52),
	.w2(32'hb909c6b2),
	.w3(32'hba457b0d),
	.w4(32'h3a1871bb),
	.w5(32'h3a4e05cc),
	.w6(32'hba758f24),
	.w7(32'h3a2efd62),
	.w8(32'h3a8121f6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921a3a8),
	.w1(32'h3a93cd7d),
	.w2(32'h3a172261),
	.w3(32'h39c8bb70),
	.w4(32'h3acaee1c),
	.w5(32'h39d9a59f),
	.w6(32'h39cf6ed1),
	.w7(32'h3ad1c566),
	.w8(32'h3a6bdabf),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9263f6),
	.w1(32'hb9d53b00),
	.w2(32'hb9c72636),
	.w3(32'h3ab95a72),
	.w4(32'hb6cce826),
	.w5(32'hb895944b),
	.w6(32'h3ad44eb0),
	.w7(32'hba255932),
	.w8(32'hb819121a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a288938),
	.w1(32'hbc143ab1),
	.w2(32'hbc014b67),
	.w3(32'hba4e1563),
	.w4(32'hbbbf6f03),
	.w5(32'hbba1ca0c),
	.w6(32'h3b9519e9),
	.w7(32'hbbd7d988),
	.w8(32'hbc0a43d6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6c098),
	.w1(32'hbb7a3258),
	.w2(32'hbb9f5605),
	.w3(32'hb9371582),
	.w4(32'hbb678091),
	.w5(32'hbb993100),
	.w6(32'h3b88c707),
	.w7(32'h3b22e547),
	.w8(32'h3b532965),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10b901),
	.w1(32'h3b8bb2d8),
	.w2(32'h3b5623b2),
	.w3(32'h3b97452e),
	.w4(32'hb9708abd),
	.w5(32'h3ab5a27f),
	.w6(32'h3b608ef4),
	.w7(32'h3aa8333d),
	.w8(32'h3b42df41),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba723901),
	.w1(32'h3b8eaeba),
	.w2(32'h3bab9776),
	.w3(32'hbbae945b),
	.w4(32'h3bbe4510),
	.w5(32'h3d00fef8),
	.w6(32'h39a8e7d6),
	.w7(32'h3c2e795d),
	.w8(32'h3cb8929b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b02c5),
	.w1(32'hbb203e0f),
	.w2(32'hbb8d7efd),
	.w3(32'h3cbb6cd4),
	.w4(32'h3b76913e),
	.w5(32'hbc6ed021),
	.w6(32'h3bb33322),
	.w7(32'hbaf04897),
	.w8(32'h3abd18b2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bec24),
	.w1(32'h3b51b47d),
	.w2(32'hbbd68c0f),
	.w3(32'hbb36aa20),
	.w4(32'h39a441ef),
	.w5(32'hbc359f9d),
	.w6(32'h39d7b77d),
	.w7(32'hba461e83),
	.w8(32'hba369762),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb381af2),
	.w1(32'hb958df10),
	.w2(32'h3c4ae709),
	.w3(32'hbbbbb593),
	.w4(32'h3b8d0f16),
	.w5(32'h3c504ee0),
	.w6(32'hbc284158),
	.w7(32'h3a96e439),
	.w8(32'h3c071d1f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15543b),
	.w1(32'hb99b48c4),
	.w2(32'h3a8fe84f),
	.w3(32'h3b50e27f),
	.w4(32'hbbb25b30),
	.w5(32'h39e38604),
	.w6(32'h3b9ece5d),
	.w7(32'h3a6321bd),
	.w8(32'h3afa2086),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada3139),
	.w1(32'h3bbf7350),
	.w2(32'hbacbbc81),
	.w3(32'h3b595c9e),
	.w4(32'h398c2a67),
	.w5(32'hba14a27f),
	.w6(32'h3ad91b68),
	.w7(32'h3bcebfca),
	.w8(32'h39fa86d3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3c66d),
	.w1(32'h3c39d1f4),
	.w2(32'h3ba36ea5),
	.w3(32'hba857bbc),
	.w4(32'h3c0e6274),
	.w5(32'h3be2ec3a),
	.w6(32'h3af50130),
	.w7(32'h3c0eb411),
	.w8(32'h3c291464),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69d156),
	.w1(32'h3c441cc5),
	.w2(32'h3c2b4b51),
	.w3(32'h3cae2d38),
	.w4(32'h3c52feb5),
	.w5(32'h3c39843a),
	.w6(32'h3c92adfc),
	.w7(32'h3bd4c542),
	.w8(32'hbb917975),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a8109),
	.w1(32'hbb8a342b),
	.w2(32'hbbc97ec6),
	.w3(32'hbbf500f7),
	.w4(32'h3b522e39),
	.w5(32'hbba25f11),
	.w6(32'hbb74baa1),
	.w7(32'hbba7bbc8),
	.w8(32'h3b85d3dc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf26dcd),
	.w1(32'h3c00ab8d),
	.w2(32'hbb78212d),
	.w3(32'h3b917eed),
	.w4(32'h3b38b4f2),
	.w5(32'hbbbb5f0b),
	.w6(32'h3b2c565b),
	.w7(32'hbabdbef2),
	.w8(32'h3b2378af),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3143c2),
	.w1(32'hba0af7f1),
	.w2(32'h3b2442a7),
	.w3(32'hbb57bd33),
	.w4(32'hbb3594ee),
	.w5(32'h3c299ceb),
	.w6(32'h3b305f55),
	.w7(32'hba81f331),
	.w8(32'hbc190f3e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745c1e),
	.w1(32'h3a143c6a),
	.w2(32'hbaf16384),
	.w3(32'hbc3adcc4),
	.w4(32'hbb5489c8),
	.w5(32'hbae7d2b3),
	.w6(32'hbc2cacee),
	.w7(32'hbb07a469),
	.w8(32'h3b181428),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41f2fb),
	.w1(32'h3bce8103),
	.w2(32'h38f382d9),
	.w3(32'h3c55ab19),
	.w4(32'h3b921e37),
	.w5(32'hbc3d7a50),
	.w6(32'h3c909824),
	.w7(32'h3b9a9a13),
	.w8(32'hbbb0980a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8cbd7),
	.w1(32'h3956f983),
	.w2(32'h3b9e292d),
	.w3(32'hbaac38bb),
	.w4(32'hba067642),
	.w5(32'h3b315226),
	.w6(32'hb976bea7),
	.w7(32'hbbc61544),
	.w8(32'hbb036d04),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7b8cb),
	.w1(32'hbb5191eb),
	.w2(32'hbb3e5d37),
	.w3(32'h3b0216df),
	.w4(32'hb982cf58),
	.w5(32'hbb645935),
	.w6(32'hbb2709a2),
	.w7(32'hbc284adc),
	.w8(32'hb9925ea7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52da76),
	.w1(32'hbbadb11c),
	.w2(32'hbae0a59e),
	.w3(32'hba82527a),
	.w4(32'hbad9029d),
	.w5(32'hbc055842),
	.w6(32'hbbc9c415),
	.w7(32'h3a7b724c),
	.w8(32'hbb02e147),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7735c),
	.w1(32'h3c5df6e9),
	.w2(32'h3beba448),
	.w3(32'hbb8718db),
	.w4(32'h3c74567d),
	.w5(32'h3ba44fff),
	.w6(32'hbad8b9ac),
	.w7(32'h3bf29906),
	.w8(32'hb8867d3a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c009a19),
	.w1(32'hbb822848),
	.w2(32'hbac7f940),
	.w3(32'h3b51b0f9),
	.w4(32'h3a72da02),
	.w5(32'h3a9eba42),
	.w6(32'h39dd344a),
	.w7(32'h3b9f860e),
	.w8(32'hbab0f87b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd37b1),
	.w1(32'hbbc6ec25),
	.w2(32'h3b9a6ebc),
	.w3(32'hbc17923c),
	.w4(32'hbabfeb2b),
	.w5(32'hba7871fb),
	.w6(32'hbbe6d561),
	.w7(32'h399d6c62),
	.w8(32'hbbfa6782),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8733e9),
	.w1(32'h3b27af61),
	.w2(32'hbbe60337),
	.w3(32'hbb441c3c),
	.w4(32'h3b97e4b1),
	.w5(32'h3b34495f),
	.w6(32'hbbd37cad),
	.w7(32'hbbc1f555),
	.w8(32'hbc104e9b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5d248),
	.w1(32'hba0bffc9),
	.w2(32'hbbbd3755),
	.w3(32'h3bc72e93),
	.w4(32'h3bf87c12),
	.w5(32'hbc7a64b4),
	.w6(32'h3cbcc44f),
	.w7(32'h3c0c5ab4),
	.w8(32'hbb92bb19),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910912),
	.w1(32'h3be6e376),
	.w2(32'h3ba296ca),
	.w3(32'hbbe09ce0),
	.w4(32'h3bc8b238),
	.w5(32'hbbea8053),
	.w6(32'h39bd426c),
	.w7(32'h3b996909),
	.w8(32'hba858d91),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29eb55),
	.w1(32'h3ba060ae),
	.w2(32'h3b99aea8),
	.w3(32'h3c2c7738),
	.w4(32'hbb642c85),
	.w5(32'h3ae914b8),
	.w6(32'h3c0e8810),
	.w7(32'hbb7d42f5),
	.w8(32'hba949637),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb815927),
	.w1(32'hbba46f66),
	.w2(32'hbb76799d),
	.w3(32'hbb12b8c8),
	.w4(32'hbae04353),
	.w5(32'h3ad19ad7),
	.w6(32'h3b6d7789),
	.w7(32'hbba697b8),
	.w8(32'hbb62daf1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb509d0),
	.w1(32'hbb930edd),
	.w2(32'hba9df30b),
	.w3(32'h3c1dba7f),
	.w4(32'hbb5c9881),
	.w5(32'h3b077a7f),
	.w6(32'h3c39b6b3),
	.w7(32'hba1b437c),
	.w8(32'h3ba9acc0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd28d1b),
	.w1(32'h3bb35711),
	.w2(32'hbbb8799d),
	.w3(32'h3c04c40f),
	.w4(32'h398c6d57),
	.w5(32'hbc38fbf5),
	.w6(32'h3bb29ca5),
	.w7(32'h3bb67bf7),
	.w8(32'hbb83744e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4124f),
	.w1(32'h39a59849),
	.w2(32'hbae6f6bd),
	.w3(32'hbc6cba9d),
	.w4(32'hb9040354),
	.w5(32'h3b9b7938),
	.w6(32'h39f1d8db),
	.w7(32'hbba773c9),
	.w8(32'h38f820c2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6123e),
	.w1(32'h39b9a01a),
	.w2(32'hbb39839e),
	.w3(32'hbba3d7f3),
	.w4(32'h399bf69c),
	.w5(32'hbc7c8956),
	.w6(32'hbc2c34d4),
	.w7(32'h3ae0ec5f),
	.w8(32'h3aca77b8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269a94),
	.w1(32'h3a5e97ae),
	.w2(32'hbb49dc3f),
	.w3(32'h3bc7105f),
	.w4(32'h3c034c2f),
	.w5(32'hbb992a4c),
	.w6(32'h3b7af87b),
	.w7(32'h3c356207),
	.w8(32'h3b9fd219),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a3ebb),
	.w1(32'h38e81998),
	.w2(32'h3bd180a8),
	.w3(32'hbbc4e3dc),
	.w4(32'h397f9fd9),
	.w5(32'hbb8c93cf),
	.w6(32'h3bbd38cd),
	.w7(32'h3aa073e4),
	.w8(32'h3c953423),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cb5b1),
	.w1(32'h3c36a518),
	.w2(32'h3a74c42c),
	.w3(32'h3d0a3cb3),
	.w4(32'h3c3a61bf),
	.w5(32'hba6e6239),
	.w6(32'h3cb588fa),
	.w7(32'h3c4cac92),
	.w8(32'hbc02e4b6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd343d),
	.w1(32'hbbe00be9),
	.w2(32'hbbf7fb67),
	.w3(32'hbc205828),
	.w4(32'hbbbba3e1),
	.w5(32'hbc53e1a4),
	.w6(32'hbbf19b4b),
	.w7(32'h39a1c49d),
	.w8(32'hbbb97d02),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7312f),
	.w1(32'hbb1bd3d1),
	.w2(32'hbc015abc),
	.w3(32'hbc598909),
	.w4(32'h3c0ecf0a),
	.w5(32'hbaa913f8),
	.w6(32'hbbeb56f1),
	.w7(32'h3bc61588),
	.w8(32'h3b0f0b01),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad16730),
	.w1(32'h3ba53ce9),
	.w2(32'h3ad8622c),
	.w3(32'hba4ce4b6),
	.w4(32'hb8a982a9),
	.w5(32'h368a0bc0),
	.w6(32'h3ae2c588),
	.w7(32'h3bb3f566),
	.w8(32'h3baa5620),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1edcf),
	.w1(32'hbaa8de5c),
	.w2(32'hbbbd683f),
	.w3(32'h3b4c40aa),
	.w4(32'h3b8554c7),
	.w5(32'hbbaac60c),
	.w6(32'hbb46f0d1),
	.w7(32'hba0abfe1),
	.w8(32'h3bd0bd6f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c761b2e),
	.w1(32'h3ca5bf28),
	.w2(32'h3c9757e6),
	.w3(32'h3b92c37b),
	.w4(32'h3c4a304c),
	.w5(32'h3b87d15f),
	.w6(32'h3cbe2c8c),
	.w7(32'h3c091d88),
	.w8(32'hb978ce4c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae65713),
	.w1(32'h3c309191),
	.w2(32'h3bd7b783),
	.w3(32'hbbcc666c),
	.w4(32'h3bb46210),
	.w5(32'h39ecd2b1),
	.w6(32'hba2d08b6),
	.w7(32'h3b779e6c),
	.w8(32'h3970c593),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a069a2b),
	.w1(32'hbb219f66),
	.w2(32'h3bbeed17),
	.w3(32'h3a2f657d),
	.w4(32'h3b9fa0dd),
	.w5(32'hba348465),
	.w6(32'hbaa2baf3),
	.w7(32'hba84c5ed),
	.w8(32'h3baf6d62),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a3738),
	.w1(32'h3aa00a8e),
	.w2(32'hba677178),
	.w3(32'hbab03e89),
	.w4(32'hbb13a2b5),
	.w5(32'hbc68a00f),
	.w6(32'hbb153f05),
	.w7(32'hba92d77d),
	.w8(32'hbba2bf57),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa5f14),
	.w1(32'hbb472397),
	.w2(32'hbb293371),
	.w3(32'h3cca5355),
	.w4(32'h39e0183a),
	.w5(32'hbba05b3a),
	.w6(32'h3c55d3a8),
	.w7(32'h3badd5b2),
	.w8(32'h3c9b25bc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfd953),
	.w1(32'hbbc47838),
	.w2(32'hbb977bee),
	.w3(32'h3bbdfa51),
	.w4(32'h3b3fc2a7),
	.w5(32'h3b8e6670),
	.w6(32'h3a91af00),
	.w7(32'h3ad3c6fa),
	.w8(32'hbc215885),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25e248),
	.w1(32'hbb8d14fa),
	.w2(32'hbb87f617),
	.w3(32'hbc11455f),
	.w4(32'hbc7ad469),
	.w5(32'hbc1bb53b),
	.w6(32'hbc08c7ea),
	.w7(32'hbb9edd68),
	.w8(32'hbad87da0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed6d78),
	.w1(32'h3ba2120c),
	.w2(32'h3b9183fa),
	.w3(32'h3b325951),
	.w4(32'h3bc11e29),
	.w5(32'hbc4d86af),
	.w6(32'hbc175a8d),
	.w7(32'h3b7e65b3),
	.w8(32'hbc13697e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f245a),
	.w1(32'h3b8c164b),
	.w2(32'h3ac6a76e),
	.w3(32'h3b92a9d3),
	.w4(32'h3c3c3648),
	.w5(32'h3bd69c5a),
	.w6(32'hbb44fe25),
	.w7(32'h3c243054),
	.w8(32'h3bba87a1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6276d3),
	.w1(32'h3b4005e2),
	.w2(32'h3bdb7a70),
	.w3(32'h3c2ce6c0),
	.w4(32'h3ba2ed58),
	.w5(32'h3ae1b7a7),
	.w6(32'h3c318a00),
	.w7(32'h3b04119e),
	.w8(32'hbc4cf7d8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1c6b3),
	.w1(32'hbb4bc65c),
	.w2(32'h3c49a5eb),
	.w3(32'h3b309eb5),
	.w4(32'hbbcf9610),
	.w5(32'h3ceb5bf0),
	.w6(32'h3ba7e596),
	.w7(32'h3ad35a95),
	.w8(32'h3c3deeef),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb8f5c),
	.w1(32'h3aba5e33),
	.w2(32'hbafd33b9),
	.w3(32'h3ab7a5b3),
	.w4(32'h3a9d97e4),
	.w5(32'hbb86557d),
	.w6(32'h3b76dc21),
	.w7(32'hb9bbc8f0),
	.w8(32'h3b29dd33),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83580e),
	.w1(32'hbc237aa1),
	.w2(32'hb9619826),
	.w3(32'h3acecdb2),
	.w4(32'hbbbe8d4b),
	.w5(32'h3c9f167a),
	.w6(32'h38c9a20e),
	.w7(32'hbb20ec4c),
	.w8(32'h3c06fb89),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7a683),
	.w1(32'hbbffbd9c),
	.w2(32'hbabccfb4),
	.w3(32'hbbecbb4c),
	.w4(32'hbb8f1010),
	.w5(32'hbbc10daf),
	.w6(32'hbb9b1156),
	.w7(32'h3aa4509d),
	.w8(32'h3c0de7ce),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be727b8),
	.w1(32'hbc000ce9),
	.w2(32'hbaaf5c44),
	.w3(32'h3aa5ecfb),
	.w4(32'hbbf01b6f),
	.w5(32'hbbc9ae89),
	.w6(32'h3b83ffcd),
	.w7(32'hbb71f047),
	.w8(32'hbb161b74),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc289798),
	.w1(32'hbb11b7af),
	.w2(32'hbb47d340),
	.w3(32'hbbd11d42),
	.w4(32'hbadecceb),
	.w5(32'hbc0f9a4e),
	.w6(32'hbbf7c0bb),
	.w7(32'h3b37d776),
	.w8(32'hbaa53bd7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32af46),
	.w1(32'hbb93f9cf),
	.w2(32'hbb65497b),
	.w3(32'h3ba93d6d),
	.w4(32'hbb437c05),
	.w5(32'h3bc2930c),
	.w6(32'hbc068b98),
	.w7(32'hbc3edbc9),
	.w8(32'hbc0a40b2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb648431),
	.w1(32'h3ba1a253),
	.w2(32'hbb3f9ed2),
	.w3(32'hbb9721f8),
	.w4(32'h3ac7cebf),
	.w5(32'hbab10471),
	.w6(32'h3b73ddfe),
	.w7(32'h3bc944f7),
	.w8(32'h3cb49cc8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf1724),
	.w1(32'h39950fd7),
	.w2(32'h3afdfdbb),
	.w3(32'h3c877e16),
	.w4(32'h3bada34c),
	.w5(32'h39bc889c),
	.w6(32'h3b825906),
	.w7(32'h3a89d779),
	.w8(32'h3b80c675),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c58323),
	.w1(32'h3acd4d0a),
	.w2(32'hbaaa53ff),
	.w3(32'h3b10aa65),
	.w4(32'h3b916bf3),
	.w5(32'h3b145525),
	.w6(32'hbb28731b),
	.w7(32'hba6ba35f),
	.w8(32'hba791699),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ec896),
	.w1(32'hbae284fd),
	.w2(32'hbb1a45a4),
	.w3(32'h3b4c773d),
	.w4(32'h3b29e609),
	.w5(32'hbbd49577),
	.w6(32'hba440896),
	.w7(32'hba7e1188),
	.w8(32'hbb5259c1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe70f30),
	.w1(32'hbbab7fbf),
	.w2(32'h3b2db82d),
	.w3(32'hbc087190),
	.w4(32'h3b0927de),
	.w5(32'h3b44179e),
	.w6(32'hbc2dd69b),
	.w7(32'h3a35d954),
	.w8(32'hba55ee04),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21ac27),
	.w1(32'hbb303c16),
	.w2(32'h3a2c1cdb),
	.w3(32'hbc3a597a),
	.w4(32'hbb3592b8),
	.w5(32'hbc99e06c),
	.w6(32'hbb6f216d),
	.w7(32'h3b14965a),
	.w8(32'h3a8158a3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b4a54),
	.w1(32'hb91ca321),
	.w2(32'hbbb3f49d),
	.w3(32'h3b878184),
	.w4(32'hbb8810eb),
	.w5(32'h3bcff49c),
	.w6(32'h3c1eaa91),
	.w7(32'hbbca47fc),
	.w8(32'h39cdb468),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c892),
	.w1(32'hbb4cd4ca),
	.w2(32'hbb94d980),
	.w3(32'h390feb69),
	.w4(32'hbb68298a),
	.w5(32'hbb58bdde),
	.w6(32'h3b37786e),
	.w7(32'hba915e61),
	.w8(32'hbb9ec81a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a2ec0),
	.w1(32'h3b2b8d40),
	.w2(32'h3bf4cb14),
	.w3(32'hba3e9100),
	.w4(32'h3b097582),
	.w5(32'h3968b91e),
	.w6(32'h3ad84f39),
	.w7(32'h3a0bb2b0),
	.w8(32'h3b83700d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9d8fe),
	.w1(32'h3a7fcb79),
	.w2(32'h3aa60bef),
	.w3(32'h3b4adc4a),
	.w4(32'hbb80ba8d),
	.w5(32'hbc031daf),
	.w6(32'h3bc405a2),
	.w7(32'hbba3c736),
	.w8(32'hbbc2d1e1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb780433),
	.w1(32'h3bb9631a),
	.w2(32'hbba56869),
	.w3(32'hbbaee919),
	.w4(32'h3b80cd53),
	.w5(32'h3ba0deb0),
	.w6(32'hbc13181a),
	.w7(32'hbb523978),
	.w8(32'h3ba820df),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa526b5),
	.w1(32'hbba32df6),
	.w2(32'hbbb3f312),
	.w3(32'h3bff480f),
	.w4(32'hbbfd1d8a),
	.w5(32'hbc375cc9),
	.w6(32'h3ba4a8df),
	.w7(32'hba8eace5),
	.w8(32'hb96f9f88),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba38295),
	.w1(32'hbc8d62e9),
	.w2(32'hbc27c099),
	.w3(32'hbae93f41),
	.w4(32'h3a484e80),
	.w5(32'h3cd4e63e),
	.w6(32'h3b68f69c),
	.w7(32'hbb5bfe1f),
	.w8(32'h3b5d021b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c205173),
	.w1(32'h3c231208),
	.w2(32'hbae4baad),
	.w3(32'h3a02b4dc),
	.w4(32'h3ba7d7ba),
	.w5(32'hbc061d2a),
	.w6(32'h3c81a04f),
	.w7(32'h3b9ff1d4),
	.w8(32'hbb057588),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b035d),
	.w1(32'hbc16d0f0),
	.w2(32'hbb0d441b),
	.w3(32'hbb41df2a),
	.w4(32'hbb7cd47c),
	.w5(32'hbbac97d5),
	.w6(32'hbb54e9cb),
	.w7(32'hbb98064e),
	.w8(32'hb9c7999d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07faf0),
	.w1(32'h3c29b61b),
	.w2(32'h3b53f2de),
	.w3(32'h3c4b1ab3),
	.w4(32'h3bfd4828),
	.w5(32'hbb94b312),
	.w6(32'h3baafcfd),
	.w7(32'h3c4644f9),
	.w8(32'h3c0e263f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47cd66),
	.w1(32'h3c31f28f),
	.w2(32'h3c04f9da),
	.w3(32'h3c35f7b4),
	.w4(32'h3baff66a),
	.w5(32'hbb3dd6e1),
	.w6(32'h3c808894),
	.w7(32'hba251284),
	.w8(32'hbc133a25),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55e980),
	.w1(32'hbbc3aafe),
	.w2(32'hbb2bb97b),
	.w3(32'h3aa4fdd1),
	.w4(32'hbbc5b06a),
	.w5(32'h3b0d68dd),
	.w6(32'h3a93f8da),
	.w7(32'hbb08fc24),
	.w8(32'h3b1d52ce),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54925b),
	.w1(32'hbb153bbf),
	.w2(32'hbc1edf9f),
	.w3(32'h395b8ee3),
	.w4(32'hbb52528c),
	.w5(32'hbbf76fa2),
	.w6(32'h3baf973b),
	.w7(32'hbb375724),
	.w8(32'hbc0313ff),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb0928),
	.w1(32'hbbd7ac03),
	.w2(32'h3b18cd0c),
	.w3(32'hbb904a98),
	.w4(32'h3b258bef),
	.w5(32'hbc369246),
	.w6(32'hbb8a3fe4),
	.w7(32'hbb9f904c),
	.w8(32'h3bc33beb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf6339),
	.w1(32'h3a1b8632),
	.w2(32'h3b64cd16),
	.w3(32'h3b7b07c9),
	.w4(32'hbbd28bc1),
	.w5(32'h3c0d6123),
	.w6(32'hbaa07174),
	.w7(32'hbad67b2f),
	.w8(32'h3c11d8c8),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b8bd),
	.w1(32'hbb80313e),
	.w2(32'h3b265376),
	.w3(32'h3b89dfe6),
	.w4(32'h3be93cb5),
	.w5(32'hbb235588),
	.w6(32'h3b2e581b),
	.w7(32'h3ade40e9),
	.w8(32'h3b33016e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c40fe),
	.w1(32'hbb735c26),
	.w2(32'hbaa55b12),
	.w3(32'h3a317de3),
	.w4(32'h3b0eb8bf),
	.w5(32'hbc05835e),
	.w6(32'hb95e7176),
	.w7(32'hbbac071e),
	.w8(32'hbac79ca3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3875c08a),
	.w1(32'h3afc931f),
	.w2(32'hba7cea18),
	.w3(32'h3a6f736e),
	.w4(32'h3b3f5e42),
	.w5(32'hbc182bfc),
	.w6(32'hbba1564f),
	.w7(32'hbaa3125e),
	.w8(32'hbc1682cb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ab8a),
	.w1(32'hba727539),
	.w2(32'hbb52a636),
	.w3(32'hbc0cd106),
	.w4(32'hbb85cc02),
	.w5(32'hbb79e5b5),
	.w6(32'hbc2073df),
	.w7(32'hbba5b820),
	.w8(32'h3b1257dc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af56c),
	.w1(32'hbba0fc84),
	.w2(32'hbbceb570),
	.w3(32'h3b8cdaf8),
	.w4(32'h3b1f3de1),
	.w5(32'hbc36fab1),
	.w6(32'h3bc1cdac),
	.w7(32'hba29463b),
	.w8(32'hbb382b97),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa69c84),
	.w1(32'hbb49b235),
	.w2(32'hbb06b5ef),
	.w3(32'hba9f3069),
	.w4(32'h3b79ed24),
	.w5(32'hbbf5e8a8),
	.w6(32'h3a3fa88f),
	.w7(32'h3b5cd20c),
	.w8(32'hbc5bdc65),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7b288),
	.w1(32'hbabaec0f),
	.w2(32'h3c0a36a6),
	.w3(32'h393368df),
	.w4(32'h3b4c603f),
	.w5(32'h3c800252),
	.w6(32'hbc0648a1),
	.w7(32'hbb864aff),
	.w8(32'h3b40a26c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923d469),
	.w1(32'hbb816edf),
	.w2(32'h3beb2a5c),
	.w3(32'hbb1e5e3e),
	.w4(32'h3bca2af9),
	.w5(32'h3ca43dbb),
	.w6(32'h3be4da38),
	.w7(32'h3b34b9c1),
	.w8(32'h3c9b8719),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb77b2),
	.w1(32'hbba3eaf3),
	.w2(32'hbbac6823),
	.w3(32'hbb755005),
	.w4(32'h3ab88fd6),
	.w5(32'h3d1d44af),
	.w6(32'h3bcd7728),
	.w7(32'h3a5b38b8),
	.w8(32'h3cbcd2a1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b673785),
	.w1(32'h3bef21ec),
	.w2(32'hb9db28fd),
	.w3(32'h3c84256d),
	.w4(32'h3c9ed11e),
	.w5(32'hbbbde181),
	.w6(32'h3b3146f7),
	.w7(32'h3bf6e9ba),
	.w8(32'hbbabc6d8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c4a32),
	.w1(32'h3b0c0cf1),
	.w2(32'h3cc0aa81),
	.w3(32'hbb73068a),
	.w4(32'hbb454cad),
	.w5(32'h3cdaa5fc),
	.w6(32'hbc3ea5a4),
	.w7(32'h3aca9ab4),
	.w8(32'h3cb0894c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7e902),
	.w1(32'h3a7fed01),
	.w2(32'h3ca160ae),
	.w3(32'hbb2e4320),
	.w4(32'h3b9807d7),
	.w5(32'h3d48bd46),
	.w6(32'hbb0e37f9),
	.w7(32'h3a46a4ad),
	.w8(32'h3cd82053),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8275ad),
	.w1(32'h3bce75a2),
	.w2(32'hbaf55e22),
	.w3(32'h3cb4b14d),
	.w4(32'hbc008eb1),
	.w5(32'hbbb08a53),
	.w6(32'h3bb116bf),
	.w7(32'hbb4afff6),
	.w8(32'h3bbcf7aa),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d01fd),
	.w1(32'h3c0d8a72),
	.w2(32'h3b50c5cb),
	.w3(32'h3bb70b95),
	.w4(32'h3bf50388),
	.w5(32'h3a1cb447),
	.w6(32'h3c22b466),
	.w7(32'h3bed6cca),
	.w8(32'h3bcd4545),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c252933),
	.w1(32'h3c44c4da),
	.w2(32'h3c7a690b),
	.w3(32'h3c5d1412),
	.w4(32'h3b4f4db2),
	.w5(32'h3c68354a),
	.w6(32'h3aa1a84e),
	.w7(32'hbb59c370),
	.w8(32'h3aa27273),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b555e),
	.w1(32'h3b3859f2),
	.w2(32'hbbed9bf7),
	.w3(32'hbbeedcf1),
	.w4(32'h3b7ca975),
	.w5(32'hbc07de3c),
	.w6(32'h3a91e257),
	.w7(32'h3b0419d5),
	.w8(32'hbaabd9a6),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa09a65),
	.w1(32'h3bc18ef7),
	.w2(32'hba25ce46),
	.w3(32'hbc0158f7),
	.w4(32'hbbcb5208),
	.w5(32'h3992a9ab),
	.w6(32'hbb357843),
	.w7(32'h3a86ee50),
	.w8(32'hbb89abf5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc02c6),
	.w1(32'h3a1532ff),
	.w2(32'h3b874a5f),
	.w3(32'hbc17ec78),
	.w4(32'h38c31c6f),
	.w5(32'hba64d0f7),
	.w6(32'hbc567288),
	.w7(32'hbaa0cb7f),
	.w8(32'h3b50f05e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a85e),
	.w1(32'hbbac5655),
	.w2(32'hbb54536e),
	.w3(32'h3b252d05),
	.w4(32'hbb788549),
	.w5(32'hbc2e96c8),
	.w6(32'h3ab04875),
	.w7(32'hba222294),
	.w8(32'hbb45163c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06abb5),
	.w1(32'h3a5a8934),
	.w2(32'h392425af),
	.w3(32'hbac5fee1),
	.w4(32'h3a91851e),
	.w5(32'h39d3cd03),
	.w6(32'h3babd70e),
	.w7(32'hbbb80f48),
	.w8(32'h3c01cb50),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01dbcc),
	.w1(32'hbbef715d),
	.w2(32'hbb28af51),
	.w3(32'h3b928ea1),
	.w4(32'hbc07beb0),
	.w5(32'hbaba6c44),
	.w6(32'hbbf00124),
	.w7(32'hbbc2690d),
	.w8(32'h3c0b62b4),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4573eb),
	.w1(32'hba278866),
	.w2(32'hbc0abec9),
	.w3(32'h3b8b3170),
	.w4(32'h3a9e1ecc),
	.w5(32'hbc104b21),
	.w6(32'h3a359f0a),
	.w7(32'hba68509a),
	.w8(32'h3aa55022),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37a714),
	.w1(32'h37d5585c),
	.w2(32'h3a4a0fc5),
	.w3(32'hbbdf3457),
	.w4(32'hbb8e8c6e),
	.w5(32'h3b62ccd8),
	.w6(32'h37c9cd3f),
	.w7(32'hba2ca50b),
	.w8(32'h3beb36da),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bed67),
	.w1(32'h3aeed2f9),
	.w2(32'h3b321339),
	.w3(32'hbb4969c9),
	.w4(32'h3b087a7e),
	.w5(32'h3b7c830e),
	.w6(32'hbb3bf823),
	.w7(32'hbbcfd13a),
	.w8(32'h3bcaf6d6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1ba7f),
	.w1(32'hb989f499),
	.w2(32'hbb07e6e6),
	.w3(32'hb89e01a4),
	.w4(32'h3ae27b3b),
	.w5(32'hb9896dcd),
	.w6(32'h3ad35dec),
	.w7(32'hba5c162c),
	.w8(32'hbac4d660),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb7970),
	.w1(32'h3b8223d2),
	.w2(32'h3b1d5142),
	.w3(32'hbbc0f882),
	.w4(32'hbb1b14d0),
	.w5(32'h3bda9ab9),
	.w6(32'hbb8d9d43),
	.w7(32'hbac5a3a9),
	.w8(32'h3bbdcf56),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef0a66),
	.w1(32'hba03910d),
	.w2(32'hbb68fdaf),
	.w3(32'h3cbd09af),
	.w4(32'hbacb1041),
	.w5(32'h3ae6d648),
	.w6(32'h3c88a41c),
	.w7(32'hbc0791d0),
	.w8(32'hbb444895),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb414a53),
	.w1(32'hbb2cd794),
	.w2(32'h3b528d85),
	.w3(32'h3af97020),
	.w4(32'h3b1f40b0),
	.w5(32'hba5a75d5),
	.w6(32'hbb975ba1),
	.w7(32'hbb1162f9),
	.w8(32'h3b6b5b88),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2c52d),
	.w1(32'hbaa28bb8),
	.w2(32'hbbae4360),
	.w3(32'h3b149f71),
	.w4(32'h3a080e23),
	.w5(32'hbbcffbd6),
	.w6(32'hbb839158),
	.w7(32'hbb68aff9),
	.w8(32'h3b9f8e30),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1440f),
	.w1(32'hbb978666),
	.w2(32'hbbc3bbe0),
	.w3(32'h3bb61277),
	.w4(32'hbb4c6cb8),
	.w5(32'h3b22ad3b),
	.w6(32'h3bab385b),
	.w7(32'hbb980e1f),
	.w8(32'hbc38984e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75049d),
	.w1(32'hbb42c31b),
	.w2(32'hba835738),
	.w3(32'hba4aa480),
	.w4(32'hba572b54),
	.w5(32'hbb136041),
	.w6(32'h3a2f53dc),
	.w7(32'hbb9d8492),
	.w8(32'h3c26cb3b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4c8cb),
	.w1(32'hba38c5f8),
	.w2(32'hbbb8374a),
	.w3(32'h3b139d43),
	.w4(32'h3b95e34b),
	.w5(32'hbcaa5e58),
	.w6(32'h3ba8ae5c),
	.w7(32'hbb5626bd),
	.w8(32'hbb964454),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5e8de),
	.w1(32'hbab22c09),
	.w2(32'h3c23b0ba),
	.w3(32'hba28b05b),
	.w4(32'h3ba522ea),
	.w5(32'h3b9bb3a9),
	.w6(32'h3b40eead),
	.w7(32'h39ee4b90),
	.w8(32'h3a864499),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb7792),
	.w1(32'h3b9bbf45),
	.w2(32'h3a035ff2),
	.w3(32'h3aab84be),
	.w4(32'h3bb4e094),
	.w5(32'hbc26f6ba),
	.w6(32'hbb1202a5),
	.w7(32'h3b26fafb),
	.w8(32'h3b85cdc6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8b9f),
	.w1(32'h3a1e65ce),
	.w2(32'h3b24b9e2),
	.w3(32'h38c578d5),
	.w4(32'hbbdf6bdd),
	.w5(32'h3be94b74),
	.w6(32'h3b51649f),
	.w7(32'hbbd065a9),
	.w8(32'h3b8caefe),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996b8d8),
	.w1(32'h3b16c956),
	.w2(32'h3b8ecaf6),
	.w3(32'h3a18c154),
	.w4(32'h3a3d546e),
	.w5(32'hba845991),
	.w6(32'hba4a4bd5),
	.w7(32'hb9a4050a),
	.w8(32'hbaa20a32),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a1349),
	.w1(32'h3c0aa8b8),
	.w2(32'h3c251d7d),
	.w3(32'h3bcc0a48),
	.w4(32'h3c072be6),
	.w5(32'h3b63188c),
	.w6(32'h39db1bfa),
	.w7(32'h3b039454),
	.w8(32'h3b89cd77),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11adfc),
	.w1(32'h3c208be4),
	.w2(32'h3a8d18ee),
	.w3(32'hbb93be0b),
	.w4(32'h3c04ca63),
	.w5(32'hbb31869e),
	.w6(32'h3aeb5352),
	.w7(32'h3bcaddd9),
	.w8(32'h3ab12b34),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16d0c1),
	.w1(32'hbbba5869),
	.w2(32'hbaa0cb9a),
	.w3(32'hbba36995),
	.w4(32'hbc228999),
	.w5(32'hb9b9820c),
	.w6(32'hbb42e32d),
	.w7(32'h3a4fefe3),
	.w8(32'h3af8ef6c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93d855),
	.w1(32'hbbc24429),
	.w2(32'h3be39113),
	.w3(32'h3acd3d61),
	.w4(32'hbc25ff5e),
	.w5(32'hbb0a7800),
	.w6(32'h3b134390),
	.w7(32'hbc0bc685),
	.w8(32'h3b8a7c3b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa971c),
	.w1(32'hbac33615),
	.w2(32'h3b7173cd),
	.w3(32'h3b270b28),
	.w4(32'h3a7695d1),
	.w5(32'hbaf83ad1),
	.w6(32'h3b0304ba),
	.w7(32'h3ba7350f),
	.w8(32'h3c023938),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca76e),
	.w1(32'h3b93b79c),
	.w2(32'h3b8401c6),
	.w3(32'hbbab8cbc),
	.w4(32'h3c2a54a0),
	.w5(32'h3bfa6471),
	.w6(32'h3861656c),
	.w7(32'hb9a7514c),
	.w8(32'h3c8699b1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6df4),
	.w1(32'h3bad02c0),
	.w2(32'h3b173ccf),
	.w3(32'hbae98af8),
	.w4(32'hbb3aca1c),
	.w5(32'hbb0bdb8c),
	.w6(32'h3bfc824f),
	.w7(32'hbb9dc8e8),
	.w8(32'h3a90bdd8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dac22),
	.w1(32'hbae6eda9),
	.w2(32'hbb0ba096),
	.w3(32'hbb0f9f2e),
	.w4(32'h3ad913d2),
	.w5(32'hba810759),
	.w6(32'h3c17d9cf),
	.w7(32'h3b5e8473),
	.w8(32'hbb866af4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b637e09),
	.w1(32'hba864b01),
	.w2(32'hba979742),
	.w3(32'h3c016e81),
	.w4(32'h399b45d6),
	.w5(32'h3c315aad),
	.w6(32'hb919aae6),
	.w7(32'h39826e7a),
	.w8(32'hbb2b1669),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe0580),
	.w1(32'h39916f1f),
	.w2(32'h3cad7e6e),
	.w3(32'h3c102a6d),
	.w4(32'h3b075a15),
	.w5(32'h3c8b09b8),
	.w6(32'h3c5e03c2),
	.w7(32'h3c1871cc),
	.w8(32'hba3daa77),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb3bbc),
	.w1(32'hbc07c3c7),
	.w2(32'h3c58899c),
	.w3(32'h3b8ce746),
	.w4(32'hbc0c02c4),
	.w5(32'hbb8b05ae),
	.w6(32'hbb8c1d61),
	.w7(32'hbc1b099b),
	.w8(32'h3c0f6037),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8859b8),
	.w1(32'h3b30ab0e),
	.w2(32'h38a98596),
	.w3(32'h3c13b508),
	.w4(32'h3bb24865),
	.w5(32'hbc03dbfa),
	.w6(32'h3abc6392),
	.w7(32'h3b9acbd3),
	.w8(32'hbb4ca02e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4ce39),
	.w1(32'h3aee6427),
	.w2(32'hbaa05c3a),
	.w3(32'h3c048705),
	.w4(32'h3bcf471a),
	.w5(32'h3ac2570a),
	.w6(32'h3bfc0bcc),
	.w7(32'h3b1f3830),
	.w8(32'hbb5c7a57),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2efed),
	.w1(32'h38f47a31),
	.w2(32'hbb0fc7d4),
	.w3(32'hbc45a80a),
	.w4(32'hb9bcc776),
	.w5(32'hbaeb49a6),
	.w6(32'hbbecf21a),
	.w7(32'h3a48251c),
	.w8(32'hbb07956c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca5fe5),
	.w1(32'hbb5bf4c5),
	.w2(32'h3b16add5),
	.w3(32'hbb808344),
	.w4(32'hbb2ae20d),
	.w5(32'h3adc07a8),
	.w6(32'h3a141bc2),
	.w7(32'hbc114964),
	.w8(32'hba3d5b2f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5448c),
	.w1(32'hbbabe286),
	.w2(32'hbb213418),
	.w3(32'h3bc1e3e4),
	.w4(32'hbb8fff54),
	.w5(32'h3c3d6288),
	.w6(32'h3beb1264),
	.w7(32'hbb9571b6),
	.w8(32'h3a821db2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb066aaf),
	.w1(32'h3b9a676e),
	.w2(32'h3c389ffc),
	.w3(32'h3a5ff9e3),
	.w4(32'h3b3284b4),
	.w5(32'hb9faaf93),
	.w6(32'h3b7b0440),
	.w7(32'h3b1d01ba),
	.w8(32'h3c1800bb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fd756),
	.w1(32'h3b29eb14),
	.w2(32'h3c5103c0),
	.w3(32'hbbd8ca89),
	.w4(32'h3ca823f4),
	.w5(32'hbbe4e617),
	.w6(32'hbb6f7dbe),
	.w7(32'h3be5b7f6),
	.w8(32'h3c4f9a3d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbccae),
	.w1(32'h3b19b407),
	.w2(32'h3b048090),
	.w3(32'h3c093cdd),
	.w4(32'hbb49e52c),
	.w5(32'hbaaa6857),
	.w6(32'h39352d26),
	.w7(32'h39df396c),
	.w8(32'h3af1d61b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e11be),
	.w1(32'hbc19dd10),
	.w2(32'hbc8badfb),
	.w3(32'hbab8e5aa),
	.w4(32'hbb3de427),
	.w5(32'hbc0e3993),
	.w6(32'h3aba1f9b),
	.w7(32'hbbb726a4),
	.w8(32'h3a29b234),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4576d7),
	.w1(32'hbbc3efd7),
	.w2(32'h3b233a39),
	.w3(32'h3bb589ce),
	.w4(32'hb969e2f6),
	.w5(32'h3c0b5b6f),
	.w6(32'h3b1e40f6),
	.w7(32'h3b78eacf),
	.w8(32'h3af3481b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c427779),
	.w1(32'h3b3756f4),
	.w2(32'h3b9296f8),
	.w3(32'h3b74bc20),
	.w4(32'hba8938fc),
	.w5(32'h3c683643),
	.w6(32'h3bc22f46),
	.w7(32'h3b5c6839),
	.w8(32'hbb3ea5f4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0730f2),
	.w1(32'h3c58bd2c),
	.w2(32'hbb9e1c13),
	.w3(32'h3bdb4cb5),
	.w4(32'h3be27811),
	.w5(32'hbba1facf),
	.w6(32'h3b090706),
	.w7(32'h3a3bac18),
	.w8(32'hbc039d78),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bb921),
	.w1(32'hba9fb1a3),
	.w2(32'hbb63ba6a),
	.w3(32'h3c1fe022),
	.w4(32'h3a38a851),
	.w5(32'hbab8c2e9),
	.w6(32'hbbcb1c54),
	.w7(32'h3b4fad13),
	.w8(32'hbb8576dc),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8c89a),
	.w1(32'hbb06fdd4),
	.w2(32'hbc4d1dc7),
	.w3(32'hbae71905),
	.w4(32'hbb22fa83),
	.w5(32'h3af1664d),
	.w6(32'h3b8971e9),
	.w7(32'hbb545ff3),
	.w8(32'hbb4a0129),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc229777),
	.w1(32'hba236079),
	.w2(32'hbb253e91),
	.w3(32'hbb36c9c5),
	.w4(32'h3a96629d),
	.w5(32'h3b996419),
	.w6(32'hbb74bc6d),
	.w7(32'h3c0cff10),
	.w8(32'h3bdd1d66),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7764),
	.w1(32'h3bfaa556),
	.w2(32'h3c34105f),
	.w3(32'h3ab375f3),
	.w4(32'h3c1c58af),
	.w5(32'h3be2896a),
	.w6(32'h3b70254c),
	.w7(32'h3bedca18),
	.w8(32'h3a98b832),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c8fc1),
	.w1(32'hbc5f43cc),
	.w2(32'hbc0583c1),
	.w3(32'hba9995ca),
	.w4(32'hbc7d5364),
	.w5(32'hbbbb6713),
	.w6(32'hbb7b4ca2),
	.w7(32'hbc6831e9),
	.w8(32'h3a49cf6c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb279c16),
	.w1(32'hbba112fb),
	.w2(32'hbbc68e34),
	.w3(32'hbbda0fca),
	.w4(32'h388f3559),
	.w5(32'hbbcdd2c6),
	.w6(32'h39221853),
	.w7(32'h3b3a787a),
	.w8(32'h3b157470),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7783852),
	.w1(32'hbb8c69a7),
	.w2(32'hbc23e7ff),
	.w3(32'h3b8ebb7b),
	.w4(32'hbc06e3f9),
	.w5(32'hbb340589),
	.w6(32'h3b8feb01),
	.w7(32'hbbb1b8ca),
	.w8(32'hbb83227d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4ce2c),
	.w1(32'h3b343cdf),
	.w2(32'hbb895f72),
	.w3(32'hbb92db66),
	.w4(32'h3bd8ac83),
	.w5(32'hbc589cf7),
	.w6(32'hbb1ac65e),
	.w7(32'h3c364549),
	.w8(32'h3ba983c3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c093269),
	.w1(32'hbb8643e9),
	.w2(32'hbb12f23a),
	.w3(32'h3bf7490b),
	.w4(32'hbb107929),
	.w5(32'h3a94e7c7),
	.w6(32'h3b66cb91),
	.w7(32'hbb17f4b1),
	.w8(32'hbb357676),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59f98e),
	.w1(32'hba89cf31),
	.w2(32'h3a5c196e),
	.w3(32'hbb083e43),
	.w4(32'h3bc180d5),
	.w5(32'h3baef82f),
	.w6(32'hbbcd70d1),
	.w7(32'h3b437755),
	.w8(32'hba97518c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab60c04),
	.w1(32'hb9c0e721),
	.w2(32'hbc09df0a),
	.w3(32'hbb8e8b3e),
	.w4(32'hbafb0f68),
	.w5(32'h399d9c72),
	.w6(32'hbb0225c2),
	.w7(32'hbbe885cd),
	.w8(32'hbc4e130e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15cf88),
	.w1(32'h3b402b99),
	.w2(32'hbb16dd72),
	.w3(32'h3a9a3776),
	.w4(32'h3b2b47f9),
	.w5(32'hbbd637eb),
	.w6(32'h3bdae9e6),
	.w7(32'h3aa3adf0),
	.w8(32'hba5bc0ca),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9bde3),
	.w1(32'hbc10996c),
	.w2(32'h3c10c80d),
	.w3(32'hbba7ece7),
	.w4(32'h3b96d8c8),
	.w5(32'h3b91dcc5),
	.w6(32'hbb2d10f7),
	.w7(32'h3c1a0a09),
	.w8(32'h3aa83c3d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1899a1),
	.w1(32'hbbfcb12d),
	.w2(32'hbbd06a2b),
	.w3(32'h3af07e22),
	.w4(32'hbc52c2de),
	.w5(32'hbc303074),
	.w6(32'h3a7c41fa),
	.w7(32'hbc27e241),
	.w8(32'hba943c57),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb629ede),
	.w1(32'hba1fcb8b),
	.w2(32'hbb8cb50c),
	.w3(32'h3af99ec5),
	.w4(32'h3b2cdf9c),
	.w5(32'hba823a03),
	.w6(32'h3abbaf60),
	.w7(32'h3ab7cbdb),
	.w8(32'h3aae5321),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f2a69),
	.w1(32'hbbab41ff),
	.w2(32'h3b6e5195),
	.w3(32'hbb0c4bc4),
	.w4(32'h3b3ec208),
	.w5(32'hbc2e5efe),
	.w6(32'hbb883714),
	.w7(32'hbc075f5e),
	.w8(32'hbc0cbef2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba861),
	.w1(32'h3bb42ce3),
	.w2(32'h3c0f7ca1),
	.w3(32'hbc0d5724),
	.w4(32'h3b9ccf17),
	.w5(32'h39e7f621),
	.w6(32'hba07f59c),
	.w7(32'hb9361632),
	.w8(32'h3ad0ee3e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeea72a),
	.w1(32'hbbb29cb6),
	.w2(32'h3abe1938),
	.w3(32'hbacec0fd),
	.w4(32'h3ab01c0a),
	.w5(32'hbb3e47dc),
	.w6(32'h3c1c3f43),
	.w7(32'h3a83db31),
	.w8(32'hbbcd1580),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd04693),
	.w1(32'hbb048b69),
	.w2(32'hbba2b311),
	.w3(32'h3ba4cfc0),
	.w4(32'hba39d1e9),
	.w5(32'h3c0ac15f),
	.w6(32'h3c631701),
	.w7(32'hbba8896c),
	.w8(32'hbbed4ba2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8e5db),
	.w1(32'h3bc19682),
	.w2(32'hba01024f),
	.w3(32'hbbe70637),
	.w4(32'h3bab0275),
	.w5(32'hbbcb0dc9),
	.w6(32'hbbd6e567),
	.w7(32'h3ae6e7a1),
	.w8(32'hbaef0c70),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bd279),
	.w1(32'h3bb5a5ee),
	.w2(32'hbb19707c),
	.w3(32'hbc1e80df),
	.w4(32'h3bfa9ecd),
	.w5(32'hbbd81bdf),
	.w6(32'hbab16d84),
	.w7(32'h3c11c6d0),
	.w8(32'h3b5c1743),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d12442),
	.w1(32'hbb5a8ca1),
	.w2(32'hbaae9722),
	.w3(32'hbb13bfb6),
	.w4(32'hbbda2e3b),
	.w5(32'hb9070e0c),
	.w6(32'h3b8764c5),
	.w7(32'hbbc3cc5d),
	.w8(32'h3998d95b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39faf277),
	.w1(32'hbb9a4fbb),
	.w2(32'hbb1e3f79),
	.w3(32'hbb1931c7),
	.w4(32'hb96b54ce),
	.w5(32'h3c2d5d68),
	.w6(32'hb9d11ef3),
	.w7(32'hba9e1cce),
	.w8(32'h3768e286),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb320fdc),
	.w1(32'hbb0cd756),
	.w2(32'hb8c1e4f7),
	.w3(32'h3a0fdab2),
	.w4(32'h3b526375),
	.w5(32'h3c5ecb7a),
	.w6(32'hbb31ab09),
	.w7(32'h3ba6afaa),
	.w8(32'hba653837),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c1355),
	.w1(32'h3caafed8),
	.w2(32'h3cfccb31),
	.w3(32'h3b44a9e6),
	.w4(32'h3c6d7285),
	.w5(32'h3cc5e4e2),
	.w6(32'h3a9ce480),
	.w7(32'h3bd0b645),
	.w8(32'h3c092572),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97130b),
	.w1(32'h3c730033),
	.w2(32'h3cf68970),
	.w3(32'hbb04a961),
	.w4(32'h3d148de0),
	.w5(32'h3c111d29),
	.w6(32'h3c006bab),
	.w7(32'hbaad18a6),
	.w8(32'h3af5752b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b41ab),
	.w1(32'h3bf22de2),
	.w2(32'h3a963fe1),
	.w3(32'h3bab76fb),
	.w4(32'hbc163cdf),
	.w5(32'hbc35f449),
	.w6(32'h3b119325),
	.w7(32'hbb544c16),
	.w8(32'hbab6e36d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb619e9),
	.w1(32'hbb85d46a),
	.w2(32'h397c06ff),
	.w3(32'hbc1fde8f),
	.w4(32'hbad090a8),
	.w5(32'h3a4e4f8f),
	.w6(32'h3ab5f7ec),
	.w7(32'hba7a1df7),
	.w8(32'h3b41744b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d3e38d),
	.w1(32'hbac085a9),
	.w2(32'h3b111071),
	.w3(32'hbb107e6e),
	.w4(32'hbb2f0aae),
	.w5(32'h3be2925d),
	.w6(32'h3b53ee7a),
	.w7(32'hb978a869),
	.w8(32'hbb458eef),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbd130),
	.w1(32'h3bec82b4),
	.w2(32'hba895375),
	.w3(32'h3bb810cd),
	.w4(32'h3b97ee4f),
	.w5(32'h3b798b30),
	.w6(32'h3c87a9e5),
	.w7(32'h3bef0f68),
	.w8(32'h3b913bad),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a94ab),
	.w1(32'h3979a662),
	.w2(32'h3b454648),
	.w3(32'h3c0d4b80),
	.w4(32'h3ad5122e),
	.w5(32'h3bc7625b),
	.w6(32'h3b1e10ef),
	.w7(32'hb9500aba),
	.w8(32'h3bb784fc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad24158),
	.w1(32'hbbc795ef),
	.w2(32'hbb0b3ef1),
	.w3(32'hba9d6871),
	.w4(32'h3ad682ce),
	.w5(32'h3b716822),
	.w6(32'hb95f3d98),
	.w7(32'h3bcaac46),
	.w8(32'h3b8bdb17),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90bc41),
	.w1(32'h3bfaae18),
	.w2(32'h3a88fbbb),
	.w3(32'h3ac71d1f),
	.w4(32'h3b7ff80b),
	.w5(32'hbc1121c5),
	.w6(32'h3c34f8a9),
	.w7(32'hbb5396f3),
	.w8(32'hbb9297b7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9346c5),
	.w1(32'hbc198ddc),
	.w2(32'hbb36ee35),
	.w3(32'hb77c1dc3),
	.w4(32'h38aed93e),
	.w5(32'h3bb86e5b),
	.w6(32'hbb389d64),
	.w7(32'h39e463d6),
	.w8(32'hbb2e3d9c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a169f),
	.w1(32'hba479a5b),
	.w2(32'hbaacbc80),
	.w3(32'h3b164ebd),
	.w4(32'hba78be2f),
	.w5(32'h3b2e72bf),
	.w6(32'h3a0b4f35),
	.w7(32'hbc80ef12),
	.w8(32'h3a6ebdb9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a61ac),
	.w1(32'h3ba2a21e),
	.w2(32'h3b430fb9),
	.w3(32'h3b81b0e1),
	.w4(32'h387f78b7),
	.w5(32'h3ad888b4),
	.w6(32'h39946b3a),
	.w7(32'hba53f088),
	.w8(32'hba4c5823),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65980e),
	.w1(32'hbb907785),
	.w2(32'hbb9ac319),
	.w3(32'hbbd49aac),
	.w4(32'hbb8372a7),
	.w5(32'hbaf09be8),
	.w6(32'h3af1c465),
	.w7(32'hbb624ea0),
	.w8(32'h3a9ed780),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee6ea8),
	.w1(32'h3b7332de),
	.w2(32'h3cb81e5d),
	.w3(32'hbb1cf6be),
	.w4(32'h3cbe4f28),
	.w5(32'h3c239ba8),
	.w6(32'h3c1712ac),
	.w7(32'hbbdedfa6),
	.w8(32'hbc117efe),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfca47e),
	.w1(32'hbb45ea18),
	.w2(32'hba8e2120),
	.w3(32'h3ab92a51),
	.w4(32'h3b3561fb),
	.w5(32'hbbd868e4),
	.w6(32'h3b7d7c1a),
	.w7(32'hbc0134b5),
	.w8(32'hbbd35570),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd4468),
	.w1(32'hba214234),
	.w2(32'h3becd2dd),
	.w3(32'h3b7c6a0c),
	.w4(32'hbb1deb47),
	.w5(32'hbb5ded14),
	.w6(32'h3c056a34),
	.w7(32'h3b88e0bc),
	.w8(32'hbbda6a63),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d3078),
	.w1(32'hbbf86a3c),
	.w2(32'hbc11a80a),
	.w3(32'hbb03f924),
	.w4(32'hbaaea5d3),
	.w5(32'h39b59193),
	.w6(32'h3b8fb2bd),
	.w7(32'hbb022ff3),
	.w8(32'h3baef398),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b6a61),
	.w1(32'h3bd6a9f5),
	.w2(32'hbb21b957),
	.w3(32'h3c4dbffa),
	.w4(32'hbbdcd27c),
	.w5(32'hbc28880b),
	.w6(32'h3bcf19c6),
	.w7(32'hba7ef55e),
	.w8(32'hbbf2ce4a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb15b87),
	.w1(32'h3bc45e97),
	.w2(32'hbbc9b133),
	.w3(32'hbba157d6),
	.w4(32'hbb7acc16),
	.w5(32'hbba082c9),
	.w6(32'hba8d5f30),
	.w7(32'hbbff4d33),
	.w8(32'hbb4f9258),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb724f4a),
	.w1(32'hbb008bae),
	.w2(32'h3bc091a4),
	.w3(32'hbaab328f),
	.w4(32'hbb29a3ca),
	.w5(32'h3be92c6b),
	.w6(32'hbb48e7ce),
	.w7(32'h3ab5961f),
	.w8(32'hbbd8100c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a998f),
	.w1(32'h3c0db72c),
	.w2(32'h3c0992b2),
	.w3(32'hbbac9fc9),
	.w4(32'h3b945cd5),
	.w5(32'hbba49d0f),
	.w6(32'hbbb2b94a),
	.w7(32'h3b27fd7f),
	.w8(32'h3a227e43),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba063e0),
	.w1(32'hbb7bcd27),
	.w2(32'hbbebbbb4),
	.w3(32'hba99f2f4),
	.w4(32'hbc0199d3),
	.w5(32'hb9aa88dd),
	.w6(32'h3bf31bea),
	.w7(32'hbb00e613),
	.w8(32'hbb198554),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939151a),
	.w1(32'hb84c2a85),
	.w2(32'h39dcdae1),
	.w3(32'hbba73dc0),
	.w4(32'hbb82caa1),
	.w5(32'h3bbb1fb5),
	.w6(32'hbaf42cb9),
	.w7(32'h3b168d40),
	.w8(32'h3bdfbfbb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dd2b6),
	.w1(32'hbb699c17),
	.w2(32'h3ad247c7),
	.w3(32'h3ad7cb74),
	.w4(32'hb9a18652),
	.w5(32'hbb84a068),
	.w6(32'h3ba92a2d),
	.w7(32'hbb0dfa53),
	.w8(32'hbb113277),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5ee8),
	.w1(32'hbc0736ad),
	.w2(32'hb80368c8),
	.w3(32'h3ad64ddb),
	.w4(32'h3af085db),
	.w5(32'hbc1a5d7d),
	.w6(32'hbb5d91df),
	.w7(32'hbb053994),
	.w8(32'h3ac94519),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8a4e2),
	.w1(32'hbbccb3be),
	.w2(32'hbb3f6ea2),
	.w3(32'hbb2f0a1b),
	.w4(32'hbbcd1a6b),
	.w5(32'h3bc5a690),
	.w6(32'hbb2a5058),
	.w7(32'h395424cd),
	.w8(32'h3b86512d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49bceb),
	.w1(32'h39d00762),
	.w2(32'hbb344764),
	.w3(32'h3bb86181),
	.w4(32'hba831ce0),
	.w5(32'hbc03decc),
	.w6(32'h3ac813d5),
	.w7(32'h3b76672d),
	.w8(32'hbbaafeed),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32cff2),
	.w1(32'hbb25a84b),
	.w2(32'hba781e9a),
	.w3(32'hbb418f13),
	.w4(32'hbbff781c),
	.w5(32'hba87167b),
	.w6(32'hbbcb561b),
	.w7(32'hbb4bfb13),
	.w8(32'hbb1b3a34),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74d8a2),
	.w1(32'hbb11896f),
	.w2(32'hbb241baf),
	.w3(32'h3afb7377),
	.w4(32'hba4777da),
	.w5(32'h3c0abea3),
	.w6(32'h3bf9723e),
	.w7(32'hbbe91eb0),
	.w8(32'h3a84afee),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f6de5),
	.w1(32'hbba5b0f2),
	.w2(32'hbc250d55),
	.w3(32'h3ba44406),
	.w4(32'hbc400762),
	.w5(32'hbc92409a),
	.w6(32'h3b107c38),
	.w7(32'hbc2e99cb),
	.w8(32'hbc111dbb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ceaef),
	.w1(32'hbb70aca8),
	.w2(32'h3a82cede),
	.w3(32'hbc1544cd),
	.w4(32'h3a769d1f),
	.w5(32'h3cb53499),
	.w6(32'h3bd9a48c),
	.w7(32'h3c8798a0),
	.w8(32'h3cb32078),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule