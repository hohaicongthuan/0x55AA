module layer_8_featuremap_86(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8777f),
	.w1(32'h3d30c2a1),
	.w2(32'hbbaff923),
	.w3(32'h3d4f16b3),
	.w4(32'h3d913c6e),
	.w5(32'hbc986353),
	.w6(32'hbc352dee),
	.w7(32'h3b3b4945),
	.w8(32'hbc9abfe6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc6993),
	.w1(32'h3b46f8cc),
	.w2(32'h3c6d35d7),
	.w3(32'hbc63ce9d),
	.w4(32'h39c9d8a3),
	.w5(32'hbc867b65),
	.w6(32'h3d2dc907),
	.w7(32'hbce6ce7c),
	.w8(32'h3d2b0c76),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce565da),
	.w1(32'hbc2aa5cd),
	.w2(32'h3b0ca601),
	.w3(32'hbb3fdcff),
	.w4(32'h3b081a6b),
	.w5(32'hbcc8ba60),
	.w6(32'h3ae89859),
	.w7(32'h3baff7db),
	.w8(32'h3bc99a0a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c302091),
	.w1(32'hbc414e79),
	.w2(32'hbbe297f9),
	.w3(32'hbce1248c),
	.w4(32'h3bf7e760),
	.w5(32'hbbddf392),
	.w6(32'hbbbf41c4),
	.w7(32'hbb706110),
	.w8(32'h3cedeb25),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d030eea),
	.w1(32'hbc4022a8),
	.w2(32'hbb98d59b),
	.w3(32'h3cc7cab1),
	.w4(32'hbc7bbd96),
	.w5(32'hbb04b181),
	.w6(32'hbc1dbfac),
	.w7(32'h3c7c453a),
	.w8(32'hba9fefbe),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf43b6f),
	.w1(32'h3c95b15d),
	.w2(32'hbce9609d),
	.w3(32'h3c754f89),
	.w4(32'h3c2823aa),
	.w5(32'hb9aca0b0),
	.w6(32'hbc2546ed),
	.w7(32'h3b81dda8),
	.w8(32'h3c037316),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fca38),
	.w1(32'hbb9b5f51),
	.w2(32'h3acac5dd),
	.w3(32'hbc4381f2),
	.w4(32'hbbcd14b8),
	.w5(32'h3b7ab3d0),
	.w6(32'h3cb200c5),
	.w7(32'hbd398e2d),
	.w8(32'hbcce01ee),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddefb9),
	.w1(32'h3c910e5b),
	.w2(32'hbcd3c262),
	.w3(32'h3d051241),
	.w4(32'h3b3d32a6),
	.w5(32'h3b9649de),
	.w6(32'h3ced1fd1),
	.w7(32'h3d21b350),
	.w8(32'h3bd03c59),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e4e6a),
	.w1(32'hbd07081a),
	.w2(32'h3a8185ee),
	.w3(32'h3bd09362),
	.w4(32'hbbccb4eb),
	.w5(32'h3c00be06),
	.w6(32'h3b1ae602),
	.w7(32'hbc42f2b9),
	.w8(32'hbd037fc0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b8bd8),
	.w1(32'h3d23d6ed),
	.w2(32'hbcc7c6c2),
	.w3(32'hbcd39ff1),
	.w4(32'hbd1e3e63),
	.w5(32'hbbc09835),
	.w6(32'hbc6c1eb2),
	.w7(32'h3738adec),
	.w8(32'hbb27d913),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc84308),
	.w1(32'hbc9aa606),
	.w2(32'hbb8fa33b),
	.w3(32'h3b0c1c16),
	.w4(32'h3cc5a386),
	.w5(32'h3c8e9507),
	.w6(32'hbc859026),
	.w7(32'h3bc353ae),
	.w8(32'h3b014767),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86914e),
	.w1(32'h3ccb0fd5),
	.w2(32'hbb99e0eb),
	.w3(32'h3c78dc0c),
	.w4(32'h3b64f29e),
	.w5(32'hbc3e5152),
	.w6(32'hba43a348),
	.w7(32'hbc8ee4c8),
	.w8(32'hbcb7ad07),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1faff5),
	.w1(32'hbc2f0891),
	.w2(32'h3d3fd334),
	.w3(32'h3b19826e),
	.w4(32'h3b167972),
	.w5(32'hb9b4da02),
	.w6(32'hbc1f3502),
	.w7(32'h3c15a618),
	.w8(32'hbbbd565e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c97ce),
	.w1(32'hba1ed3cc),
	.w2(32'hbd67c348),
	.w3(32'hbc75f87c),
	.w4(32'hbc3cbecb),
	.w5(32'h3a19ffaf),
	.w6(32'hbd1c0c7d),
	.w7(32'h39a570b9),
	.w8(32'h3d03eb54),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7508c),
	.w1(32'h3dd20b09),
	.w2(32'hbc2ed30a),
	.w3(32'h3beba066),
	.w4(32'h3d5c0d65),
	.w5(32'hbc800e0f),
	.w6(32'hbbd89e10),
	.w7(32'h3ca72dec),
	.w8(32'hbd198dfe),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d138eb5),
	.w1(32'hbbc011d7),
	.w2(32'hbd16e9ec),
	.w3(32'h3d205a63),
	.w4(32'hbd1bf6e9),
	.w5(32'h3c19ecc7),
	.w6(32'h3cbacfa6),
	.w7(32'hb8323790),
	.w8(32'hbbe54179),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c3ca4),
	.w1(32'hbab3aac3),
	.w2(32'h3c3637a8),
	.w3(32'h3ae2aea8),
	.w4(32'h3c345fd7),
	.w5(32'hbc2c7b3f),
	.w6(32'hbbb28f34),
	.w7(32'hbb699a85),
	.w8(32'h3cd7f2a2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1c0d4),
	.w1(32'hbb412c71),
	.w2(32'h3afcecd2),
	.w3(32'hbc049e2d),
	.w4(32'h3c92f56b),
	.w5(32'hbc4221d6),
	.w6(32'hbcb64ae9),
	.w7(32'hbc0de8c4),
	.w8(32'h3c8d8e43),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1dba7),
	.w1(32'h3ce1e463),
	.w2(32'hbbddf05a),
	.w3(32'hbc9bde42),
	.w4(32'hb883f175),
	.w5(32'h3c2e92b8),
	.w6(32'h3c1871b1),
	.w7(32'hbd191c88),
	.w8(32'hbd690671),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a808021),
	.w1(32'hbcc38f75),
	.w2(32'hbbd84d7c),
	.w3(32'h3c58eef1),
	.w4(32'h3d0c34da),
	.w5(32'h3b210714),
	.w6(32'hbbaf6e9f),
	.w7(32'hbb0d1f69),
	.w8(32'h3c84e8b3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d29d753),
	.w1(32'h3cea59a0),
	.w2(32'h3c50979b),
	.w3(32'hbbd797b8),
	.w4(32'h3cd9f13e),
	.w5(32'h3c9d09fe),
	.w6(32'hbcbc71d7),
	.w7(32'h3c40b1bc),
	.w8(32'hbbfb5f84),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd96bf7),
	.w1(32'hbc993730),
	.w2(32'h3b31af3b),
	.w3(32'h3be8a279),
	.w4(32'h3c3b4354),
	.w5(32'h3bdf1cae),
	.w6(32'h3c33062e),
	.w7(32'hbcb9d4ba),
	.w8(32'h3cd452cc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00f182),
	.w1(32'hbb224aad),
	.w2(32'hb9dc6700),
	.w3(32'hbcb42e31),
	.w4(32'h3d0f3806),
	.w5(32'h3cff607d),
	.w6(32'h3c3ec73f),
	.w7(32'h3ca7e39a),
	.w8(32'hbc9d2cd3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd39cb2),
	.w1(32'hbc9ea751),
	.w2(32'hbc4e4207),
	.w3(32'hbc9be905),
	.w4(32'h3d30b3ba),
	.w5(32'hbd037d95),
	.w6(32'hbb8b64b7),
	.w7(32'h3a0c71df),
	.w8(32'hbd47f290),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f8a85),
	.w1(32'hbc66177e),
	.w2(32'h3d07ebb7),
	.w3(32'hbc61b548),
	.w4(32'h3c0051c8),
	.w5(32'hbb8c5f68),
	.w6(32'h3d47aaf6),
	.w7(32'hbbc4e472),
	.w8(32'h3b3ae2f0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6dac6d),
	.w1(32'h3caf2b5b),
	.w2(32'h3b96f4f9),
	.w3(32'h3bb4a1ff),
	.w4(32'h3c013180),
	.w5(32'h3caf30a9),
	.w6(32'h3ba9ad33),
	.w7(32'h3bdea3ed),
	.w8(32'h3d01dd56),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0ed77),
	.w1(32'h3aca690a),
	.w2(32'hbbb30498),
	.w3(32'hbc01455a),
	.w4(32'hbb0c7c85),
	.w5(32'h3b973062),
	.w6(32'hbb932e06),
	.w7(32'h3c8d86dc),
	.w8(32'h3d011c03),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2be9fb),
	.w1(32'h3c8630cd),
	.w2(32'h3c875f28),
	.w3(32'hbc0a8cab),
	.w4(32'h3dd7ea23),
	.w5(32'h3d3a28ef),
	.w6(32'hbd01a870),
	.w7(32'h3c82fb03),
	.w8(32'h3c9cafcb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce52b8e),
	.w1(32'hbb9e872c),
	.w2(32'h3caa7c59),
	.w3(32'h3d6dca6f),
	.w4(32'h3bdc8d3a),
	.w5(32'h3cae6046),
	.w6(32'h3ac28263),
	.w7(32'h3c535301),
	.w8(32'h3cccdf80),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46c5e0),
	.w1(32'hbc0eeda0),
	.w2(32'h3bbe3357),
	.w3(32'hbcf8833b),
	.w4(32'h3be60ac5),
	.w5(32'h3be7bcb9),
	.w6(32'hbbe2de6f),
	.w7(32'h3c64fc75),
	.w8(32'hbc4120f5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22e7c0),
	.w1(32'h3d6a979c),
	.w2(32'hbbb1ff66),
	.w3(32'h3ab49a9b),
	.w4(32'h3b5c6a0c),
	.w5(32'hbbe4ecd8),
	.w6(32'hba79dc02),
	.w7(32'h3c06959d),
	.w8(32'hbbdde170),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf1998),
	.w1(32'hbca7ba2b),
	.w2(32'h3cb397fd),
	.w3(32'h3c99a209),
	.w4(32'hbc98a17f),
	.w5(32'hbcf98880),
	.w6(32'h38039bb7),
	.w7(32'h3cb233a5),
	.w8(32'hbad2e8a9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc594aa1),
	.w1(32'h3cc94858),
	.w2(32'hbba88f35),
	.w3(32'hbbf85144),
	.w4(32'hbb9fe8f6),
	.w5(32'hbc8da2c9),
	.w6(32'hbc18b7a1),
	.w7(32'hbbe0dab3),
	.w8(32'h3c8b4967),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc956d73),
	.w1(32'h3bb63290),
	.w2(32'hba9f7e32),
	.w3(32'hbcac235a),
	.w4(32'hbc1b7f54),
	.w5(32'h3d38c15b),
	.w6(32'hbc785fb3),
	.w7(32'hbc09d212),
	.w8(32'hbadcf1d1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4b55d),
	.w1(32'hbccec475),
	.w2(32'h3c31916e),
	.w3(32'h3be187b7),
	.w4(32'h3c460bf9),
	.w5(32'hbbe4c85c),
	.w6(32'hbc93b8ef),
	.w7(32'hba907b5d),
	.w8(32'hbbc9eb52),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefa715),
	.w1(32'h3ca39ab2),
	.w2(32'h3c1ce6b4),
	.w3(32'h3bf68f51),
	.w4(32'hbc303278),
	.w5(32'h3af2fb6d),
	.w6(32'hbbc17aaf),
	.w7(32'hbb40316f),
	.w8(32'h3b79a187),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbded97),
	.w1(32'hbc97b509),
	.w2(32'h3c243d1f),
	.w3(32'h3b8d923d),
	.w4(32'h3c1c0f47),
	.w5(32'hbb749d97),
	.w6(32'hbb9ff0ed),
	.w7(32'h3b551074),
	.w8(32'hbbed293f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad4002),
	.w1(32'hbb17a336),
	.w2(32'hbc95d93f),
	.w3(32'hba5d1a6a),
	.w4(32'h3a549f57),
	.w5(32'h3d0e4ea5),
	.w6(32'h3bcc6fc7),
	.w7(32'hbc6491ef),
	.w8(32'hbcb91a63),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd169c9a),
	.w1(32'h3bbb0407),
	.w2(32'h3c76f187),
	.w3(32'hbd2394e4),
	.w4(32'hbcf06f7b),
	.w5(32'h3b7d7bc7),
	.w6(32'h3c5a9d55),
	.w7(32'hbb950dc7),
	.w8(32'h3c733ca3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf79a4c),
	.w1(32'h3b9b007f),
	.w2(32'hbae2ad9c),
	.w3(32'h3bb61e61),
	.w4(32'h3ca39433),
	.w5(32'h3a009267),
	.w6(32'hbb8decb0),
	.w7(32'h3b8aad0b),
	.w8(32'hba3e8fb4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dc78c),
	.w1(32'h3cbb34be),
	.w2(32'h383307f4),
	.w3(32'h3be7781e),
	.w4(32'h3c3bd00f),
	.w5(32'h3c96f635),
	.w6(32'h3bd2b81a),
	.w7(32'h3c84ab0c),
	.w8(32'h3c1041f1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0c293),
	.w1(32'hbc8ee74f),
	.w2(32'hbcb36814),
	.w3(32'h3d79464f),
	.w4(32'hbcaa6a9a),
	.w5(32'h3c0395b3),
	.w6(32'hbc03baac),
	.w7(32'h3b1c0027),
	.w8(32'hbcf85dae),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fd746),
	.w1(32'hbc23749b),
	.w2(32'h3c1d1cc9),
	.w3(32'h3d83ba74),
	.w4(32'hbd414385),
	.w5(32'hbc6a5517),
	.w6(32'h3c4f619f),
	.w7(32'hbc6019c0),
	.w8(32'hbb4b46e1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74850c),
	.w1(32'hbb73cf4a),
	.w2(32'h3c514571),
	.w3(32'h3c8bb99b),
	.w4(32'h3c1a5b88),
	.w5(32'h3c40757c),
	.w6(32'hbbd7cf0b),
	.w7(32'hba2a0a63),
	.w8(32'h3da6e98f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc8647),
	.w1(32'hbb0a84bc),
	.w2(32'hbc329696),
	.w3(32'hbc862b75),
	.w4(32'h3bb5ca75),
	.w5(32'h3c23e53a),
	.w6(32'hbc147443),
	.w7(32'h3c2b426e),
	.w8(32'hbc83f1aa),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0779b6),
	.w1(32'h3beb1994),
	.w2(32'hbc06cd84),
	.w3(32'hbbac234e),
	.w4(32'hbc36fec1),
	.w5(32'hbcc3acb1),
	.w6(32'hbbc6ac82),
	.w7(32'hbc3be76c),
	.w8(32'h39cd930a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02ef3f),
	.w1(32'hbcd9790d),
	.w2(32'hbb8de4dd),
	.w3(32'hbc160267),
	.w4(32'hbc4055be),
	.w5(32'hbcc379cd),
	.w6(32'hba569206),
	.w7(32'hbc1504c6),
	.w8(32'h3bb9ece4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7c9d8),
	.w1(32'h3b6d5798),
	.w2(32'h3a07c5b1),
	.w3(32'hbc283c54),
	.w4(32'h3c91b327),
	.w5(32'hbccbc3e2),
	.w6(32'h3bf77b19),
	.w7(32'h3c3151ee),
	.w8(32'hbd0ee8f4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d1809),
	.w1(32'hbbade942),
	.w2(32'h3bf84a93),
	.w3(32'h3bb6b2b4),
	.w4(32'hba1ed7f8),
	.w5(32'hbc9e0fb6),
	.w6(32'h3c2aac69),
	.w7(32'hbd390652),
	.w8(32'h3c14c15c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2f1a7),
	.w1(32'hbbe9b30c),
	.w2(32'hbb9ae4e9),
	.w3(32'h3ca80fae),
	.w4(32'hbc8ea7b3),
	.w5(32'h3c8f0638),
	.w6(32'h3b5f20db),
	.w7(32'h3c22cf50),
	.w8(32'hbac1a194),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc977b4f),
	.w1(32'hbc6be4ba),
	.w2(32'hbbc02e79),
	.w3(32'h3ba4ed5c),
	.w4(32'hbb7a76b3),
	.w5(32'h3cbbb143),
	.w6(32'hbd0edb92),
	.w7(32'hbca15426),
	.w8(32'hbc63c035),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd32f13),
	.w1(32'hbc26ed5f),
	.w2(32'hbca149b5),
	.w3(32'hbbea3a99),
	.w4(32'hbb89c320),
	.w5(32'h3c615d1d),
	.w6(32'hbb50cd16),
	.w7(32'h3c35afbd),
	.w8(32'hbc43e064),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f4901),
	.w1(32'hbb97aceb),
	.w2(32'h3a0c6532),
	.w3(32'hbd133bb5),
	.w4(32'h3c58e8cf),
	.w5(32'h3b9cd4b5),
	.w6(32'hbc9be9c2),
	.w7(32'h3da3def4),
	.w8(32'h3c906966),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4ef5e),
	.w1(32'hbc847fa2),
	.w2(32'h3ceebec6),
	.w3(32'h3c42968c),
	.w4(32'h3b8232d8),
	.w5(32'h3b8a48a3),
	.w6(32'h3befe60c),
	.w7(32'h3c011671),
	.w8(32'h3b589ea3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd17a4eb),
	.w1(32'hbb01a59f),
	.w2(32'h3bdf655b),
	.w3(32'h3bbcbc08),
	.w4(32'h3b6b5a46),
	.w5(32'h3c052b51),
	.w6(32'hbc1363f8),
	.w7(32'hbca66824),
	.w8(32'h3d0ed637),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc007c76),
	.w1(32'hbc781a75),
	.w2(32'h3c47b3c8),
	.w3(32'hbbfd052a),
	.w4(32'h3b8770ac),
	.w5(32'h3cc18829),
	.w6(32'h3d0dea67),
	.w7(32'h3af0065c),
	.w8(32'hbc1afc3e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd22a87),
	.w1(32'h3d10020f),
	.w2(32'h3bfd1913),
	.w3(32'hbc35752b),
	.w4(32'h3b06b09f),
	.w5(32'hbc63c66d),
	.w6(32'h3b0b8cd1),
	.w7(32'hbc5d2d92),
	.w8(32'hba8aa4ce),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9e1f1),
	.w1(32'h3ca009ac),
	.w2(32'hbcace4e4),
	.w3(32'h3c9d0ce5),
	.w4(32'hbb3230b6),
	.w5(32'h3c7d9f65),
	.w6(32'hbd8efa09),
	.w7(32'h3cd0ccdc),
	.w8(32'h3b559f7c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07f248),
	.w1(32'h3c9ceb75),
	.w2(32'h3c832d73),
	.w3(32'hbc82d77e),
	.w4(32'h3c4d22cd),
	.w5(32'hbcdbbe5e),
	.w6(32'h3c4af6b7),
	.w7(32'h3ca78e2a),
	.w8(32'hbbd63fa2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8c6d),
	.w1(32'h3c388537),
	.w2(32'h3c10aa4e),
	.w3(32'h3b3809f4),
	.w4(32'hbafd2fc1),
	.w5(32'h38afba06),
	.w6(32'h3cbddda9),
	.w7(32'hbcfd7560),
	.w8(32'hbc34032e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc644300),
	.w1(32'h3c095f54),
	.w2(32'h3c960f68),
	.w3(32'hbd2141e3),
	.w4(32'hbc0b8346),
	.w5(32'hbd8d8b9a),
	.w6(32'hbb14ca40),
	.w7(32'h3cec8971),
	.w8(32'hbb68c597),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea934),
	.w1(32'hbd833bf0),
	.w2(32'h3c2b31f3),
	.w3(32'h3c527551),
	.w4(32'hbca3bd4f),
	.w5(32'hbbdba446),
	.w6(32'hbcc1703d),
	.w7(32'hbd29c14d),
	.w8(32'h39683e25),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac6e0e),
	.w1(32'hbbbe86d5),
	.w2(32'h3ab878e4),
	.w3(32'h3cb0f32c),
	.w4(32'h3c1dd59b),
	.w5(32'hbc32e9c7),
	.w6(32'h3ce7a6d4),
	.w7(32'h3cabd88f),
	.w8(32'hbca6f67a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd00f377),
	.w1(32'h3ccd79a3),
	.w2(32'hbb3aba60),
	.w3(32'h3c046c4b),
	.w4(32'hbd20d206),
	.w5(32'hbd0ab8c0),
	.w6(32'h3cb38d0d),
	.w7(32'h3ca44b3c),
	.w8(32'hbcfcd6ef),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d420d),
	.w1(32'hbbc8c687),
	.w2(32'h3d32b07d),
	.w3(32'hbc68bec4),
	.w4(32'h3dd5b0bf),
	.w5(32'h3d2c7fdd),
	.w6(32'h3bf0b8ec),
	.w7(32'hbd9311ca),
	.w8(32'h3ce6c71d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef129a),
	.w1(32'h3cdfeca7),
	.w2(32'hbc514c7c),
	.w3(32'h3ce582b8),
	.w4(32'h3a13c7a6),
	.w5(32'hbd8d0211),
	.w6(32'h3c2b552a),
	.w7(32'h3c38f2c4),
	.w8(32'h3c034f66),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a006f),
	.w1(32'hbd4fee73),
	.w2(32'h3bb1fdd4),
	.w3(32'hbd72f708),
	.w4(32'h3b4070e0),
	.w5(32'h3c141088),
	.w6(32'hbd8b43f4),
	.w7(32'h3d1e68a3),
	.w8(32'hbc459345),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21ce4d),
	.w1(32'h3c9cfeb7),
	.w2(32'hbbb7a925),
	.w3(32'h3c85edbb),
	.w4(32'h3c8e1b32),
	.w5(32'h3b273add),
	.w6(32'hbc77bbbf),
	.w7(32'h3bff5127),
	.w8(32'hbc86ac97),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93b7d5),
	.w1(32'hbbff18ba),
	.w2(32'hbbb11b63),
	.w3(32'h3c39b114),
	.w4(32'hbb6dc09b),
	.w5(32'hbd886d57),
	.w6(32'h3c9f511b),
	.w7(32'h3c333cac),
	.w8(32'h3b3c9340),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d804d),
	.w1(32'h392289a3),
	.w2(32'hbb79f668),
	.w3(32'h3c1d9270),
	.w4(32'h3d0f9f4b),
	.w5(32'h3d04cec1),
	.w6(32'h3cf86a7a),
	.w7(32'hbb091487),
	.w8(32'h3dab119f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b629),
	.w1(32'hbaa61356),
	.w2(32'h3caf2c68),
	.w3(32'h398a0bbb),
	.w4(32'hbb29d6dc),
	.w5(32'hbc242ff0),
	.w6(32'h3ba3417d),
	.w7(32'hbda1fa6c),
	.w8(32'hbd2c8e9e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9482a3),
	.w1(32'hbb6ef572),
	.w2(32'hbc459f4f),
	.w3(32'h3c2e2388),
	.w4(32'h3b14daef),
	.w5(32'h3a4f0a01),
	.w6(32'hbce2d7a2),
	.w7(32'hbd5d8188),
	.w8(32'hbc3022bd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80abf9),
	.w1(32'hbd0ccc26),
	.w2(32'hbc7e3193),
	.w3(32'hba6abcc6),
	.w4(32'h3c79aa6f),
	.w5(32'hbba434bb),
	.w6(32'h3ce78c21),
	.w7(32'h3bef8f28),
	.w8(32'h3ca5830b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2184d4),
	.w1(32'hbbb16345),
	.w2(32'hbbb3cee4),
	.w3(32'h3d27e925),
	.w4(32'h3c4cf893),
	.w5(32'hbc119a22),
	.w6(32'h3c045f6c),
	.w7(32'hbc8b302e),
	.w8(32'hbc01509c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc258a2d),
	.w1(32'h3b6ae0ed),
	.w2(32'h3c6c3842),
	.w3(32'h3c4f01a5),
	.w4(32'h3c260311),
	.w5(32'hbcf78247),
	.w6(32'h3d14adcc),
	.w7(32'hbb83b713),
	.w8(32'hbce57916),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7669c),
	.w1(32'h3c162548),
	.w2(32'hbb3d6dc5),
	.w3(32'hbb856a39),
	.w4(32'h3d0ddfb9),
	.w5(32'h3d1533c4),
	.w6(32'hbbd3906b),
	.w7(32'hbd0fed45),
	.w8(32'hbb24f89e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5744a5),
	.w1(32'h3c08fb20),
	.w2(32'hbb3d0290),
	.w3(32'h3ba4aedc),
	.w4(32'h3c983954),
	.w5(32'hbb3c8fbc),
	.w6(32'hbb8c4bfd),
	.w7(32'h3c363431),
	.w8(32'h3cb91a61),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6fdb4),
	.w1(32'hbbf23555),
	.w2(32'hbd092f78),
	.w3(32'hbc750fb0),
	.w4(32'h3b8aaa9c),
	.w5(32'h3c5f8fb7),
	.w6(32'hbd1f74b2),
	.w7(32'h3b31151e),
	.w8(32'h3cbf1b64),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ef869),
	.w1(32'h3ca05a19),
	.w2(32'hbcc2c2ed),
	.w3(32'h3bb6cba0),
	.w4(32'hbb945509),
	.w5(32'hbc8fe932),
	.w6(32'h3b802445),
	.w7(32'hbc852b90),
	.w8(32'h3cecc3c3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe195bd),
	.w1(32'h3b6eb7d7),
	.w2(32'h3a9b27e6),
	.w3(32'hbc4e4a15),
	.w4(32'hbab16298),
	.w5(32'hbc0b067c),
	.w6(32'hbc818b8e),
	.w7(32'h3b3e8633),
	.w8(32'hbc05ed9e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91c788),
	.w1(32'hbc3ae2bf),
	.w2(32'h3d82aabb),
	.w3(32'h3b73fef7),
	.w4(32'h3a951158),
	.w5(32'hbca1874c),
	.w6(32'hbc13f51d),
	.w7(32'h3c590890),
	.w8(32'h3b164752),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f2dcf),
	.w1(32'hbc8b3175),
	.w2(32'hbb4de0ba),
	.w3(32'hbb28dda9),
	.w4(32'h3d36d1f4),
	.w5(32'h3ce1b538),
	.w6(32'hbbae8c18),
	.w7(32'hbba34b8d),
	.w8(32'hbb12a773),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20692e),
	.w1(32'h3b19cdc3),
	.w2(32'h3d0f187e),
	.w3(32'hbc442153),
	.w4(32'h3c3bed6e),
	.w5(32'hbc3c2fda),
	.w6(32'h3b3a5744),
	.w7(32'h3c37181e),
	.w8(32'h3ca528d8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa7b5b),
	.w1(32'h3b802851),
	.w2(32'hbbc2f1b7),
	.w3(32'h3b4abd46),
	.w4(32'hbc6a4515),
	.w5(32'h3cbac115),
	.w6(32'h3c26cea4),
	.w7(32'hbaa01183),
	.w8(32'h3c415864),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d010420),
	.w1(32'h3bcd0062),
	.w2(32'h3c5c4995),
	.w3(32'h3c9ea0c3),
	.w4(32'h3d185171),
	.w5(32'h3c2f91c3),
	.w6(32'h3c349739),
	.w7(32'h3c08b836),
	.w8(32'h3d5eaacd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adae709),
	.w1(32'h3ba28263),
	.w2(32'h3c27c6c2),
	.w3(32'h3c17c260),
	.w4(32'hbc054a13),
	.w5(32'hbc0c47ba),
	.w6(32'hbc60472f),
	.w7(32'h3cc6fbef),
	.w8(32'h3bd48769),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd799f),
	.w1(32'hbba4ed30),
	.w2(32'h3c6da4ac),
	.w3(32'hbb31fb7c),
	.w4(32'hbc2690f0),
	.w5(32'hbc9f7a3e),
	.w6(32'hbb804f6f),
	.w7(32'h3c81b395),
	.w8(32'h3bd55ac8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb834750),
	.w1(32'h3b1d5178),
	.w2(32'h3c2a3b95),
	.w3(32'hbc828479),
	.w4(32'hbd89027a),
	.w5(32'hba758175),
	.w6(32'h3bd6b10b),
	.w7(32'hbc49aa5a),
	.w8(32'hbb95384b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d035fa3),
	.w1(32'hbcf90d9b),
	.w2(32'h3d752cc6),
	.w3(32'hbd1cf078),
	.w4(32'hba61cd71),
	.w5(32'hbbbeadeb),
	.w6(32'h3c17717f),
	.w7(32'h3d132bfa),
	.w8(32'hbbce5b39),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b865622),
	.w1(32'h3b7930df),
	.w2(32'h3c6b4cf0),
	.w3(32'h3ca37f35),
	.w4(32'hbd45e474),
	.w5(32'hbbd4771e),
	.w6(32'hbcd1e399),
	.w7(32'h3c142f32),
	.w8(32'h3ca7900a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46339f),
	.w1(32'h3b9702dd),
	.w2(32'h3ce2c37a),
	.w3(32'hbc31d034),
	.w4(32'hb9913ee6),
	.w5(32'hbce7d525),
	.w6(32'hbc7c46c4),
	.w7(32'hbc4d1ad0),
	.w8(32'h3c80196b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce61ce6),
	.w1(32'hbc4efd33),
	.w2(32'h3c19b85b),
	.w3(32'h3b553c69),
	.w4(32'hbc630318),
	.w5(32'h3cd5613b),
	.w6(32'h3aa2f0f7),
	.w7(32'hbc9b6a72),
	.w8(32'hbca8d53e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36a634),
	.w1(32'hbbf0f6a1),
	.w2(32'h3c96c638),
	.w3(32'hbc6d149e),
	.w4(32'hbd2c7862),
	.w5(32'hbc8cb101),
	.w6(32'hbae0046e),
	.w7(32'h3c91561e),
	.w8(32'h3ccbcb2b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0817b1),
	.w1(32'hbc0fd3dd),
	.w2(32'h3c7475de),
	.w3(32'h3ca206a6),
	.w4(32'h3abb586f),
	.w5(32'h3c9df14a),
	.w6(32'h3b51f581),
	.w7(32'hbc6a4f98),
	.w8(32'hbd7813f7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c848f7e),
	.w1(32'hbbf268e6),
	.w2(32'h3cf0debf),
	.w3(32'hbb1302f3),
	.w4(32'h3cc6ba16),
	.w5(32'hbc3f7fa1),
	.w6(32'hbcdf6e69),
	.w7(32'h3cadb314),
	.w8(32'hbc0f51f3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8aab3b),
	.w1(32'hbc5fe6e9),
	.w2(32'h3c2b3fea),
	.w3(32'hbd0c610e),
	.w4(32'h3ba6c0b6),
	.w5(32'hbcfa3882),
	.w6(32'h3ca69a99),
	.w7(32'hbbffbb22),
	.w8(32'hbb1a7f98),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59ca7f),
	.w1(32'h3ce4cbda),
	.w2(32'h3b403b87),
	.w3(32'h3d11cfd9),
	.w4(32'hbaf0af21),
	.w5(32'hba078563),
	.w6(32'hbca77e80),
	.w7(32'h3c6126e2),
	.w8(32'hbc37369b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd162cc4),
	.w1(32'h3b45625a),
	.w2(32'hbc065867),
	.w3(32'hbba124f8),
	.w4(32'hbc6fa78b),
	.w5(32'h3c3d6d57),
	.w6(32'hbc93e13a),
	.w7(32'hb935e632),
	.w8(32'hbc986262),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad75c),
	.w1(32'h3c56491b),
	.w2(32'hbc1e40c0),
	.w3(32'hbaaa87ec),
	.w4(32'hbc1ef9c9),
	.w5(32'h3b84b0fc),
	.w6(32'h3c4c5977),
	.w7(32'hbc4643e8),
	.w8(32'h3c00c02f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5c591),
	.w1(32'hb8384909),
	.w2(32'hbc38fcbb),
	.w3(32'h3cd2412d),
	.w4(32'h3c00bba8),
	.w5(32'hb9625931),
	.w6(32'hbca27de4),
	.w7(32'hbc020031),
	.w8(32'h3b07d9ab),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd18e316),
	.w1(32'hbbba5dd5),
	.w2(32'hba97d82c),
	.w3(32'hbb12d43f),
	.w4(32'hbb3c7322),
	.w5(32'h3b75bde2),
	.w6(32'h3b2fbaec),
	.w7(32'h3b8da821),
	.w8(32'h3ab2fd1c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0edd17),
	.w1(32'h3a3192a9),
	.w2(32'h39a027c0),
	.w3(32'hbb313d93),
	.w4(32'hbc7d7b00),
	.w5(32'h3abef87c),
	.w6(32'h3d313c36),
	.w7(32'h3b795bdc),
	.w8(32'hbb237661),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16e30f),
	.w1(32'hbbd3d4be),
	.w2(32'hbba81399),
	.w3(32'hbc17afec),
	.w4(32'h3ac725ff),
	.w5(32'h3cbcec45),
	.w6(32'h3c57c300),
	.w7(32'h3c91fc0d),
	.w8(32'hbc489a1e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc029ec8),
	.w1(32'hbb12693f),
	.w2(32'h3cc38c79),
	.w3(32'hbc890470),
	.w4(32'h3ca7f2cd),
	.w5(32'h3b864da3),
	.w6(32'hba037c29),
	.w7(32'h3a0a3ec6),
	.w8(32'h3ca1af17),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa135e),
	.w1(32'h3b8e1368),
	.w2(32'h3b2ca821),
	.w3(32'h3c70cbf6),
	.w4(32'hbc101226),
	.w5(32'h3bbae1f1),
	.w6(32'hbb96f876),
	.w7(32'h3b3ac242),
	.w8(32'h3b989022),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad284e),
	.w1(32'hba0ea33a),
	.w2(32'hbc17fefe),
	.w3(32'h3a8d15d8),
	.w4(32'h3ce5138b),
	.w5(32'h3d35cac3),
	.w6(32'h3b2564f3),
	.w7(32'h3c3b2a02),
	.w8(32'hbc1aa385),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ca807),
	.w1(32'h3c147a13),
	.w2(32'h3c8ad558),
	.w3(32'h3d938d96),
	.w4(32'hbc16c779),
	.w5(32'h3a698c28),
	.w6(32'h3c798253),
	.w7(32'h3c40ade6),
	.w8(32'hbbd35b89),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a943b02),
	.w1(32'hbc633963),
	.w2(32'h3c05148d),
	.w3(32'hbca26492),
	.w4(32'h3b836bee),
	.w5(32'hbbfffe17),
	.w6(32'h3d1ca8a8),
	.w7(32'h3b993552),
	.w8(32'h3c522ff9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e3ac7),
	.w1(32'hbc00135b),
	.w2(32'hbbaf6f80),
	.w3(32'hbc1daa1b),
	.w4(32'h3ca19946),
	.w5(32'h3c3b667f),
	.w6(32'hbc2a10e8),
	.w7(32'hbae6ca49),
	.w8(32'hbabe361e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40017b),
	.w1(32'hbb4652bf),
	.w2(32'h3bbefe88),
	.w3(32'h3cdddba2),
	.w4(32'h3cc18bf7),
	.w5(32'h3b810a9c),
	.w6(32'hbb1b5418),
	.w7(32'h3c896e12),
	.w8(32'h3c7e20aa),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad06bda),
	.w1(32'hb92c8c50),
	.w2(32'hbb8c4ccd),
	.w3(32'h38a0f618),
	.w4(32'h3be9b1ce),
	.w5(32'h3b314edc),
	.w6(32'hbc144001),
	.w7(32'hbb5fbf47),
	.w8(32'hbc35cdd3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc2892),
	.w1(32'h3bafffc5),
	.w2(32'h3b8220dc),
	.w3(32'h3b6288b5),
	.w4(32'hbb6cb934),
	.w5(32'hbc28c6ab),
	.w6(32'h3c9b1dcf),
	.w7(32'hbc6716c9),
	.w8(32'hbb8a6fbc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bbbcd),
	.w1(32'hbb6f6fd9),
	.w2(32'hbbaa68f7),
	.w3(32'h3c9038b6),
	.w4(32'hbc197e4b),
	.w5(32'h3ca9de58),
	.w6(32'hba5a773b),
	.w7(32'hbba3c982),
	.w8(32'hbb73c4de),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a6823),
	.w1(32'hbd061c38),
	.w2(32'hbc67f78a),
	.w3(32'h3b7ab8a7),
	.w4(32'h3bc5fc4f),
	.w5(32'h3c252561),
	.w6(32'hbb1d31f8),
	.w7(32'hbb4a4606),
	.w8(32'h3c3f391a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbeb45),
	.w1(32'h3c187bab),
	.w2(32'h3bf26cd7),
	.w3(32'hbc21eaee),
	.w4(32'h3c283aee),
	.w5(32'h3c62c5d4),
	.w6(32'h3cbdd528),
	.w7(32'h3c10513d),
	.w8(32'h3b74b943),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c183117),
	.w1(32'h3d7da5c1),
	.w2(32'h3b9b4cf7),
	.w3(32'h3c2df167),
	.w4(32'hbb7c00d0),
	.w5(32'h3ab36033),
	.w6(32'h3cbf72fd),
	.w7(32'h3cb939a8),
	.w8(32'hbc2828a1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a2c03),
	.w1(32'h3bdf496e),
	.w2(32'hbc35fa7b),
	.w3(32'h3c3c1085),
	.w4(32'h3b75ea6f),
	.w5(32'hbcb4ec9d),
	.w6(32'h3c0e7ea7),
	.w7(32'h3b1dcd81),
	.w8(32'h3c29a46c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1536d6),
	.w1(32'h3bfb8b0b),
	.w2(32'h3c7fd61f),
	.w3(32'hbad76d08),
	.w4(32'h3c39c58c),
	.w5(32'hbb57033c),
	.w6(32'hbc9c9669),
	.w7(32'h3c48a775),
	.w8(32'hbc4b7ae9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3541bb),
	.w1(32'hb99f8c83),
	.w2(32'h3bbd6d56),
	.w3(32'hbbc225c8),
	.w4(32'hbb8ab08f),
	.w5(32'hbad7418b),
	.w6(32'hbb30c4ad),
	.w7(32'h3d1ab734),
	.w8(32'h3c64324b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff130c),
	.w1(32'h3bc34c14),
	.w2(32'h3c9fccbf),
	.w3(32'hbbd1ed06),
	.w4(32'h3bbb8d44),
	.w5(32'hbc21b8d7),
	.w6(32'h3b54b220),
	.w7(32'hbbfea16c),
	.w8(32'hbc86d8c3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c3367),
	.w1(32'hb9f15875),
	.w2(32'h3c70921f),
	.w3(32'hbb7ac725),
	.w4(32'h3ca413f3),
	.w5(32'h3cebec4d),
	.w6(32'hbab925e2),
	.w7(32'h3aa226c3),
	.w8(32'h3cf52287),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcab15b),
	.w1(32'h3c8898c6),
	.w2(32'h3c4b666a),
	.w3(32'hbc17e45a),
	.w4(32'h3b4e7551),
	.w5(32'h3c14b307),
	.w6(32'hbc0f7121),
	.w7(32'hbc2205da),
	.w8(32'hbb432bb4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caca734),
	.w1(32'hbc9c90c7),
	.w2(32'hbc6b2be3),
	.w3(32'hbc515834),
	.w4(32'h3bbe4a8c),
	.w5(32'h3d02de63),
	.w6(32'hbbbc0539),
	.w7(32'hbb0d20b2),
	.w8(32'hbc13ce1b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c3d9f),
	.w1(32'h3ad96ef0),
	.w2(32'h3c838246),
	.w3(32'h3c9d3833),
	.w4(32'h3ca7cdb3),
	.w5(32'h3bfd0b10),
	.w6(32'h3ad4d52e),
	.w7(32'hbbd12df4),
	.w8(32'hbb08c44b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cce7852),
	.w1(32'hbbccb2b4),
	.w2(32'hbc4c523c),
	.w3(32'h3c839167),
	.w4(32'hbc25d6b2),
	.w5(32'h3c519459),
	.w6(32'hbc20dc0e),
	.w7(32'h399d3852),
	.w8(32'h3c87834e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e2abe),
	.w1(32'h3c40763d),
	.w2(32'hba922b35),
	.w3(32'h3c5a33f0),
	.w4(32'h3b85d7d8),
	.w5(32'h3b8ea297),
	.w6(32'hbbf7c436),
	.w7(32'hbab7f014),
	.w8(32'h39f1adbf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1909fc),
	.w1(32'h3ccb7c8b),
	.w2(32'h3c9aa7cc),
	.w3(32'h3bbfb798),
	.w4(32'hbc32900d),
	.w5(32'hbb8262fe),
	.w6(32'h3b6e89d3),
	.w7(32'hbba826d2),
	.w8(32'h3b218a01),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc613cb5),
	.w1(32'h3c49603f),
	.w2(32'hb9b84a05),
	.w3(32'hbb8f1d31),
	.w4(32'hbd2e016a),
	.w5(32'h3ad89cdd),
	.w6(32'hbd382822),
	.w7(32'h3ce0f5a7),
	.w8(32'h3c1f1c66),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule