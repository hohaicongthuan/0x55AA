module layer_6_featuremap_124(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb485555),
	.w1(32'hbca072fc),
	.w2(32'hbca30c70),
	.w3(32'hbc8f389a),
	.w4(32'hbc90b238),
	.w5(32'hbc946716),
	.w6(32'hbc9a0db3),
	.w7(32'hbc9b4fd4),
	.w8(32'hbc8c7a31),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9eef7e),
	.w1(32'hbb9239f1),
	.w2(32'hbb8f1567),
	.w3(32'h3a535754),
	.w4(32'h3af2a7d3),
	.w5(32'h3a06a156),
	.w6(32'h39ec81c0),
	.w7(32'hb8899af0),
	.w8(32'hba6ba67e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54ef61),
	.w1(32'hb9372491),
	.w2(32'h3baccf10),
	.w3(32'hb9ffc212),
	.w4(32'h39e7c41f),
	.w5(32'h3bf84345),
	.w6(32'hbbf6f64a),
	.w7(32'hbaf83a0c),
	.w8(32'h3c602480),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c977c8b),
	.w1(32'hba352049),
	.w2(32'hbab93785),
	.w3(32'hb92e1f9e),
	.w4(32'hb8a62719),
	.w5(32'hbb807c13),
	.w6(32'h3a6114d0),
	.w7(32'h3aecbc54),
	.w8(32'hbba1b680),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097a3a),
	.w1(32'hbb9a10d9),
	.w2(32'hb9effbd3),
	.w3(32'hbac11363),
	.w4(32'h3b9271ea),
	.w5(32'hbb889735),
	.w6(32'h3b0d942c),
	.w7(32'h3c1fd73f),
	.w8(32'h3bc18c5d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86054a),
	.w1(32'h3c84ec3e),
	.w2(32'h3c83f225),
	.w3(32'h3c37f525),
	.w4(32'h3c5f0266),
	.w5(32'h3c20a13d),
	.w6(32'h3c9a0a87),
	.w7(32'h3caca9d8),
	.w8(32'h3c8f44d1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f0a42),
	.w1(32'hbbca7260),
	.w2(32'hbbf447ac),
	.w3(32'hbbaf7f11),
	.w4(32'hbc12c46d),
	.w5(32'hbba4a9bb),
	.w6(32'hbc151945),
	.w7(32'hbc49e10c),
	.w8(32'hbc36182b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb84eb8),
	.w1(32'hbcb10606),
	.w2(32'hbc9a5beb),
	.w3(32'h3b59f722),
	.w4(32'h3c514d9d),
	.w5(32'h3bf9225f),
	.w6(32'hbc1497ba),
	.w7(32'hbb8e4cf4),
	.w8(32'hbb412705),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64f9e),
	.w1(32'hbbb29bde),
	.w2(32'hbb0fd5cf),
	.w3(32'h3a890438),
	.w4(32'h3b952097),
	.w5(32'h3ac4d671),
	.w6(32'h3b6e170d),
	.w7(32'h3b576e5c),
	.w8(32'hbb93e717),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f6ba3),
	.w1(32'h3c8e7c4d),
	.w2(32'h3cc70acf),
	.w3(32'h3c9a2319),
	.w4(32'h3ccb8b85),
	.w5(32'h3c8e9920),
	.w6(32'h3cde981e),
	.w7(32'h3d10c72d),
	.w8(32'h3cca9967),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29d79f),
	.w1(32'hba53488a),
	.w2(32'hbb7d4b8a),
	.w3(32'hbbe2de14),
	.w4(32'hbbd761b0),
	.w5(32'hbb35fd01),
	.w6(32'h3aeddf20),
	.w7(32'hbaf9ef3a),
	.w8(32'hbaa4896a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4862d0),
	.w1(32'hbc229b19),
	.w2(32'hbc1ab74e),
	.w3(32'h3b139311),
	.w4(32'h3b76f169),
	.w5(32'h3ba56ea1),
	.w6(32'h3a5d9817),
	.w7(32'h39fcb3eb),
	.w8(32'h3b11b46c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1936f7),
	.w1(32'h3c215ccb),
	.w2(32'h3c3f10fa),
	.w3(32'h3c2b1b41),
	.w4(32'h3c434030),
	.w5(32'h3c1616f5),
	.w6(32'h3c09f8c3),
	.w7(32'h3c01e657),
	.w8(32'h3bdb0229),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82eb69),
	.w1(32'hbc89c71d),
	.w2(32'hbc2abaae),
	.w3(32'hbc303628),
	.w4(32'hbc80ed44),
	.w5(32'hbc066b05),
	.w6(32'hbca64823),
	.w7(32'hbc407068),
	.w8(32'hbc565a3e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ff060),
	.w1(32'hbb2d559c),
	.w2(32'h3a99ca4f),
	.w3(32'hbb92cf0f),
	.w4(32'hbaa0bd4d),
	.w5(32'hbb8ca5c6),
	.w6(32'hbb1e9102),
	.w7(32'hbb298928),
	.w8(32'hbb27e001),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44ebe),
	.w1(32'hba743306),
	.w2(32'h3b8a24b5),
	.w3(32'hbb4f7218),
	.w4(32'h3a104ca4),
	.w5(32'hb8ba5a7f),
	.w6(32'h3a85eefa),
	.w7(32'h3b992dcb),
	.w8(32'h3b9267c4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a140a0b),
	.w1(32'hbbf537db),
	.w2(32'hbc71f530),
	.w3(32'hbb659ef3),
	.w4(32'hbc3078c5),
	.w5(32'hbc8a861e),
	.w6(32'h38d288e0),
	.w7(32'hbc1cd7a7),
	.w8(32'hbc862268),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc471578),
	.w1(32'h3b868a66),
	.w2(32'h3c0aedeb),
	.w3(32'h3bfdf8ad),
	.w4(32'h3c51fc52),
	.w5(32'h3c12411e),
	.w6(32'h3c2769f5),
	.w7(32'h3c71cb21),
	.w8(32'h3c176664),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64120d),
	.w1(32'hba2c1e2e),
	.w2(32'h3aa1c5c7),
	.w3(32'hbaf7108b),
	.w4(32'h3add9ccf),
	.w5(32'hbbecf610),
	.w6(32'h3c02130d),
	.w7(32'h3c518327),
	.w8(32'h39e02c28),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b2f04),
	.w1(32'h3bdf3e67),
	.w2(32'h3b5a4f60),
	.w3(32'h3bb5066d),
	.w4(32'h3bddcb93),
	.w5(32'h3b9feff1),
	.w6(32'h3c0707a2),
	.w7(32'h3c451965),
	.w8(32'h3bce147f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5368ce),
	.w1(32'hba6ec6db),
	.w2(32'hbb056ca3),
	.w3(32'hbacd7544),
	.w4(32'hbb390636),
	.w5(32'h3a4bc2c0),
	.w6(32'hbb17f1c6),
	.w7(32'hbb5414e1),
	.w8(32'hbafe8fab),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07ed03),
	.w1(32'h3b0c6072),
	.w2(32'h3b9f1e26),
	.w3(32'hba2d1b1a),
	.w4(32'hb9b50020),
	.w5(32'hb911c1dd),
	.w6(32'h3b253f84),
	.w7(32'h3ac8531a),
	.w8(32'h3a8fc013),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9a17),
	.w1(32'h3c162a9c),
	.w2(32'hbba7b2ae),
	.w3(32'h3c13b305),
	.w4(32'hba392b44),
	.w5(32'hbbdbe417),
	.w6(32'h3c630f6c),
	.w7(32'h3b0bc44c),
	.w8(32'hbc36a3ee),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ea139),
	.w1(32'h3c0ea2ad),
	.w2(32'h3c2149aa),
	.w3(32'hbaaa7a5c),
	.w4(32'hbbdcc7a5),
	.w5(32'hbc0bed67),
	.w6(32'h3bee8c6a),
	.w7(32'h3ae3e371),
	.w8(32'hbb7517b5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be41004),
	.w1(32'h3b553eb8),
	.w2(32'h3bb2a5b7),
	.w3(32'h3ba9d521),
	.w4(32'h3bf01c24),
	.w5(32'hba954036),
	.w6(32'h3b260392),
	.w7(32'h3c7d933a),
	.w8(32'h3b43ef46),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44be56),
	.w1(32'h3c410b7e),
	.w2(32'h3c40933c),
	.w3(32'h3c07d743),
	.w4(32'h3bd862a7),
	.w5(32'h3bb8e127),
	.w6(32'h3c50f7e6),
	.w7(32'h3c4a303a),
	.w8(32'h3c40fe38),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11032d),
	.w1(32'h3a7980ca),
	.w2(32'h3b9883c4),
	.w3(32'h3a5453fe),
	.w4(32'h3b11bbef),
	.w5(32'hbb61421c),
	.w6(32'h3c2325e0),
	.w7(32'h3c8f64c8),
	.w8(32'h3ba3af0e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d8709),
	.w1(32'h3bd16d8d),
	.w2(32'h3bcdb5df),
	.w3(32'h3bd64bc3),
	.w4(32'h3bb5ae29),
	.w5(32'h3bd0a855),
	.w6(32'h3befaa74),
	.w7(32'h3bcebf74),
	.w8(32'h3bc99784),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb86f0b),
	.w1(32'hbc11b454),
	.w2(32'hbc37067d),
	.w3(32'hbc07fb71),
	.w4(32'hbc226868),
	.w5(32'hbc0d2c4e),
	.w6(32'hbc2d8128),
	.w7(32'hbc563afc),
	.w8(32'hbc3a2071),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00ce81),
	.w1(32'h3b04f8e9),
	.w2(32'h3c1a2b4d),
	.w3(32'h3be11bb7),
	.w4(32'h3bae9b45),
	.w5(32'h3bee5542),
	.w6(32'h3bf2ca89),
	.w7(32'h3c06c4b8),
	.w8(32'h3bd75da8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03ccac),
	.w1(32'h3bd0bfdb),
	.w2(32'h3ca0ad2b),
	.w3(32'hbc04a499),
	.w4(32'hbb01215d),
	.w5(32'hbc2923ea),
	.w6(32'hbb021d0d),
	.w7(32'h3c11ed04),
	.w8(32'h3be5c962),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8759db),
	.w1(32'hbbcddf29),
	.w2(32'h3a79eefe),
	.w3(32'hb91fa706),
	.w4(32'h3ab1c8c0),
	.w5(32'hbba32bcd),
	.w6(32'h3b88f32d),
	.w7(32'h3bcf3e6f),
	.w8(32'h3b237051),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb26b),
	.w1(32'h3c117852),
	.w2(32'h3c8ca748),
	.w3(32'h3c177d39),
	.w4(32'h3bffa1d8),
	.w5(32'h3bf91499),
	.w6(32'h3c454dbe),
	.w7(32'h3c5eaafa),
	.w8(32'h3c11e2a0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ba9d9),
	.w1(32'h3af7c6bc),
	.w2(32'hbbaa2884),
	.w3(32'hb8e7a70d),
	.w4(32'hbc12641e),
	.w5(32'hbb9df196),
	.w6(32'h3b29eb8e),
	.w7(32'hbc0b1594),
	.w8(32'hbb4d97ca),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7579),
	.w1(32'h3c193edc),
	.w2(32'h3c3ddb20),
	.w3(32'h3b95a831),
	.w4(32'h3be189c5),
	.w5(32'h3b6edd30),
	.w6(32'h3c20af54),
	.w7(32'h3c4692db),
	.w8(32'h3c19c2ca),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b206b),
	.w1(32'hbbc2a68e),
	.w2(32'hbabc78e0),
	.w3(32'h3b97253d),
	.w4(32'h3ac4dc7a),
	.w5(32'hbb59adf0),
	.w6(32'hbc674989),
	.w7(32'hbaee64dc),
	.w8(32'h3bd9d206),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983229e),
	.w1(32'h3c1ca65e),
	.w2(32'h3c7fd00a),
	.w3(32'h3b53aab3),
	.w4(32'h3bd49906),
	.w5(32'h3b18ee25),
	.w6(32'h3c26458b),
	.w7(32'h3c88be76),
	.w8(32'h3c8350a9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41469b),
	.w1(32'hbb57f999),
	.w2(32'hbb1147b3),
	.w3(32'hbbb386dc),
	.w4(32'hbba767f1),
	.w5(32'hbba92439),
	.w6(32'hbb8dd1ee),
	.w7(32'hbb84142b),
	.w8(32'hbb3998e2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306b2b),
	.w1(32'hbabbb53e),
	.w2(32'hbbc71fd7),
	.w3(32'hbb8b2d8b),
	.w4(32'hbc23feab),
	.w5(32'hbc22ff9f),
	.w6(32'hbc317f7a),
	.w7(32'hbc95527a),
	.w8(32'hbc493230),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99d02c),
	.w1(32'hbb949838),
	.w2(32'h3b3e1d54),
	.w3(32'hbc7fcdb1),
	.w4(32'hbc3c4240),
	.w5(32'hbc49f19d),
	.w6(32'hbba16f47),
	.w7(32'hbbdbf73c),
	.w8(32'h3bb8d663),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5f910),
	.w1(32'hbacc7d88),
	.w2(32'hbc4766b9),
	.w3(32'h3ae456de),
	.w4(32'hbb0213b8),
	.w5(32'hbc6c3ce0),
	.w6(32'h3b886ad2),
	.w7(32'hbc311b93),
	.w8(32'hbc8da432),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a5795),
	.w1(32'h3b687672),
	.w2(32'h3b85a7e2),
	.w3(32'h3acb83fe),
	.w4(32'h3a704706),
	.w5(32'h3a31cb6e),
	.w6(32'h3b79f48c),
	.w7(32'h3b7e3868),
	.w8(32'h3ab6360d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a616f0d),
	.w1(32'hbab2a435),
	.w2(32'h3b2c189b),
	.w3(32'hbac1e25c),
	.w4(32'h3a49ba14),
	.w5(32'hbb4ef619),
	.w6(32'h3aed350c),
	.w7(32'h3baae36d),
	.w8(32'hb90ddbd8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06f246),
	.w1(32'h3b2e6355),
	.w2(32'h3b868a0a),
	.w3(32'h3a2ff50d),
	.w4(32'h3af4c802),
	.w5(32'h3b1507e3),
	.w6(32'h3bf31b3b),
	.w7(32'h3c1d5f20),
	.w8(32'h3bf3ce97),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdf097),
	.w1(32'h395e0256),
	.w2(32'hb9f2e754),
	.w3(32'h395d5598),
	.w4(32'h391733f4),
	.w5(32'h382973ee),
	.w6(32'hba757805),
	.w7(32'hbad79cfb),
	.w8(32'hba8f030d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabceb70),
	.w1(32'h3c71892f),
	.w2(32'h3c31e116),
	.w3(32'h3c380487),
	.w4(32'h3c1d1ec4),
	.w5(32'h3c07bf4c),
	.w6(32'h3cab060c),
	.w7(32'h3c9739b9),
	.w8(32'h3c4f4313),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae88275),
	.w1(32'hbc0df290),
	.w2(32'hbbfe684f),
	.w3(32'h3a980175),
	.w4(32'h3b2288a5),
	.w5(32'hbc2410c7),
	.w6(32'hbacb89d1),
	.w7(32'hb991f81f),
	.w8(32'hbc37b1c5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc885a4a),
	.w1(32'h3c5479b6),
	.w2(32'h3c0d72a6),
	.w3(32'h3b881c1e),
	.w4(32'h3c004615),
	.w5(32'h3b33c832),
	.w6(32'h3c305c24),
	.w7(32'h3c89db33),
	.w8(32'h3c105f11),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae1e73),
	.w1(32'h3c418f59),
	.w2(32'h3c3b8042),
	.w3(32'h3bf16a8c),
	.w4(32'h3c0019b3),
	.w5(32'h3c42fd24),
	.w6(32'h3bfff68c),
	.w7(32'h3be29e85),
	.w8(32'h3c3d15d6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52a577),
	.w1(32'h3b358ce8),
	.w2(32'hbb947b12),
	.w3(32'h3b843a1b),
	.w4(32'h3aa895aa),
	.w5(32'hbbbe79fa),
	.w6(32'h3b6bf32c),
	.w7(32'h3baa2801),
	.w8(32'h3bae8e1b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8258f0),
	.w1(32'h3b780fba),
	.w2(32'h3ac86e0b),
	.w3(32'h3b840a0a),
	.w4(32'h3ab5d2ab),
	.w5(32'h3b7a28ca),
	.w6(32'h3ae1e42d),
	.w7(32'hbaaf5965),
	.w8(32'hbabf6770),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17af51),
	.w1(32'h3b15e78f),
	.w2(32'h3abaf06f),
	.w3(32'h3a084707),
	.w4(32'hbb561099),
	.w5(32'hbaba1159),
	.w6(32'h3a38ecf4),
	.w7(32'hbbac53fa),
	.w8(32'hb8fa8ca0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b779bb7),
	.w1(32'h3c06af7e),
	.w2(32'hba725db2),
	.w3(32'h3c27f2f0),
	.w4(32'h3b9745f4),
	.w5(32'h3babff55),
	.w6(32'h3c10bc53),
	.w7(32'h3a757538),
	.w8(32'hba554008),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9695),
	.w1(32'hbd13ce75),
	.w2(32'hbd54f1e2),
	.w3(32'hbd10e3ff),
	.w4(32'hbd43d111),
	.w5(32'hbd000163),
	.w6(32'hbd541ba6),
	.w7(32'hbd8fd454),
	.w8(32'hbd51b17f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1e5d1b),
	.w1(32'h3b155841),
	.w2(32'hba6e0cbe),
	.w3(32'h3bc5310a),
	.w4(32'h3b9133ef),
	.w5(32'h3b936f26),
	.w6(32'h3b64b88f),
	.w7(32'h3acd767e),
	.w8(32'hba1a4bc3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84658d),
	.w1(32'h3bd474f4),
	.w2(32'hba699de9),
	.w3(32'hbbb442e2),
	.w4(32'hbaded8b2),
	.w5(32'hbbd5e409),
	.w6(32'h3b6c97d3),
	.w7(32'hbbe558b7),
	.w8(32'hbc7f7657),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e3768),
	.w1(32'hbc417674),
	.w2(32'h3b000217),
	.w3(32'hbc08a870),
	.w4(32'hbb56fe27),
	.w5(32'h3bef3385),
	.w6(32'hbc898093),
	.w7(32'hbaf4b8e4),
	.w8(32'h3c73c26e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c147005),
	.w1(32'h3be39bd1),
	.w2(32'h3bf89b8b),
	.w3(32'h3bb0e6f8),
	.w4(32'h3c3dc754),
	.w5(32'hbc715b1b),
	.w6(32'h3c6eec36),
	.w7(32'h3bb2bc17),
	.w8(32'hbc83a06f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67841a),
	.w1(32'h3ab3701d),
	.w2(32'hbba42f91),
	.w3(32'h3b36d8b8),
	.w4(32'hbb0d9da8),
	.w5(32'hbbacaa17),
	.w6(32'h3b6678f8),
	.w7(32'hbb4cf684),
	.w8(32'hbc080e61),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0f5c4),
	.w1(32'hbc0ecce2),
	.w2(32'hbcaaf42a),
	.w3(32'hbc92b8d1),
	.w4(32'hbd0f582f),
	.w5(32'hbd09dca5),
	.w6(32'hbc80eb98),
	.w7(32'hbd22158e),
	.w8(32'hbc4567de),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f9046),
	.w1(32'h3c7bc7b9),
	.w2(32'h3c210d53),
	.w3(32'h3c3e5d87),
	.w4(32'h3c10d31d),
	.w5(32'hbb8c0e26),
	.w6(32'h3c9652d9),
	.w7(32'h3c30ab0f),
	.w8(32'hbc640976),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080225),
	.w1(32'h3c9c313b),
	.w2(32'h3c414519),
	.w3(32'h3c3240a0),
	.w4(32'h3b5d09e8),
	.w5(32'hbcafad7a),
	.w6(32'h3cd39047),
	.w7(32'h3ba00028),
	.w8(32'hbcb9e4ff),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca642ce),
	.w1(32'h3c149187),
	.w2(32'hbc826ada),
	.w3(32'hbc259de0),
	.w4(32'hbc12ed1d),
	.w5(32'h3c13902b),
	.w6(32'h3c22e06a),
	.w7(32'hbc354577),
	.w8(32'h3be75837),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b567311),
	.w1(32'h3ca7a7e4),
	.w2(32'h3bc5d035),
	.w3(32'h3c8ed788),
	.w4(32'h3c4b015c),
	.w5(32'hbc664b81),
	.w6(32'h3d06eeea),
	.w7(32'h3c647e78),
	.w8(32'hbcbeb193),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule