module layer_8_featuremap_211(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcebf3),
	.w1(32'h3a308292),
	.w2(32'h39b52606),
	.w3(32'hbb3e10ac),
	.w4(32'h3b5cb833),
	.w5(32'hbba1c734),
	.w6(32'hbc36472c),
	.w7(32'hbc1a1597),
	.w8(32'h39c0dcfb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbe5b9),
	.w1(32'h3cc52022),
	.w2(32'h3b655976),
	.w3(32'hbc291293),
	.w4(32'h3c7610f9),
	.w5(32'hb78f55ba),
	.w6(32'h3c7ba924),
	.w7(32'h3bc3ad46),
	.w8(32'hbc09c36d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd52f1a),
	.w1(32'h3b3afdc4),
	.w2(32'h3c0fca68),
	.w3(32'hbc931664),
	.w4(32'h3b7a02d5),
	.w5(32'h3b3a5736),
	.w6(32'h3aa1ff23),
	.w7(32'h3bc3bdb8),
	.w8(32'h3ba16685),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e642),
	.w1(32'h3a35432e),
	.w2(32'h3962948d),
	.w3(32'h3b2d8768),
	.w4(32'h3bf90765),
	.w5(32'h3c72d785),
	.w6(32'hbc20c352),
	.w7(32'h3bb0fe60),
	.w8(32'h3c061304),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f06dd),
	.w1(32'h3d02dbad),
	.w2(32'hbb0e1fa7),
	.w3(32'h3923bc6a),
	.w4(32'h3ca4eb0c),
	.w5(32'hbb76096a),
	.w6(32'h3cc3f626),
	.w7(32'h3c125ec8),
	.w8(32'hbc692353),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd21916d),
	.w1(32'hbaa23df1),
	.w2(32'hbc161f47),
	.w3(32'hbccfb2a4),
	.w4(32'hbb804e1a),
	.w5(32'hbb8c7f33),
	.w6(32'h3b909ee9),
	.w7(32'hbb9825f7),
	.w8(32'hbc7294b9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6d840),
	.w1(32'hbc4765e5),
	.w2(32'hbb94e13f),
	.w3(32'hbb660766),
	.w4(32'hbbdfb168),
	.w5(32'hba8ca561),
	.w6(32'hbb36c239),
	.w7(32'hbaa70af4),
	.w8(32'h3b817ba2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f82b0),
	.w1(32'h3ba136b8),
	.w2(32'h3be33b7f),
	.w3(32'h3c5276f7),
	.w4(32'h3c1791be),
	.w5(32'h3c19dde2),
	.w6(32'h3c02a69f),
	.w7(32'h3ad80451),
	.w8(32'hbc062c22),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae2721),
	.w1(32'h3d126450),
	.w2(32'hbbb4c087),
	.w3(32'h3b014ca8),
	.w4(32'h3ccf6fb6),
	.w5(32'hbbb820b7),
	.w6(32'h3d01b973),
	.w7(32'h3c28b3b1),
	.w8(32'hbc44a153),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2eefb3),
	.w1(32'hbbbd01b1),
	.w2(32'hbb427550),
	.w3(32'hbd022f66),
	.w4(32'hbc273956),
	.w5(32'hbb00e809),
	.w6(32'hbb3b4bba),
	.w7(32'h3bf1b72f),
	.w8(32'h3b366d4d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9b0a6),
	.w1(32'h3cbe97bb),
	.w2(32'h3c66de32),
	.w3(32'hba40c2eb),
	.w4(32'h3caf687a),
	.w5(32'h3c93e942),
	.w6(32'h38a46ac8),
	.w7(32'h3bce653e),
	.w8(32'h3be25b99),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e9086),
	.w1(32'hbae4bf4a),
	.w2(32'h3b802648),
	.w3(32'h3af1c0fe),
	.w4(32'hbbb81aca),
	.w5(32'hbb194b7e),
	.w6(32'hbbdc2b4a),
	.w7(32'hbb373482),
	.w8(32'h3bdd4814),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ad45),
	.w1(32'hbaf4dec4),
	.w2(32'h3b0210aa),
	.w3(32'hbb284baa),
	.w4(32'hbb84fa0e),
	.w5(32'hbba0aa33),
	.w6(32'h3ba451ef),
	.w7(32'h3c03d10d),
	.w8(32'h3b4af2d0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c87de),
	.w1(32'hbb3497e2),
	.w2(32'h3bbf7f45),
	.w3(32'hbb3e474f),
	.w4(32'h3a257a6e),
	.w5(32'h3b531ede),
	.w6(32'hba15b80a),
	.w7(32'h3ac660c1),
	.w8(32'hb9d866d5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc45ea1),
	.w1(32'hbcfd930a),
	.w2(32'h3b2fe1e9),
	.w3(32'hbb32959d),
	.w4(32'hbc865099),
	.w5(32'h3bb87235),
	.w6(32'hbc9044c6),
	.w7(32'hbb3cb35a),
	.w8(32'h3c9a69df),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1de459),
	.w1(32'h3bb9914f),
	.w2(32'h3b837872),
	.w3(32'h3cddd352),
	.w4(32'h3a281b6b),
	.w5(32'h3bd8729b),
	.w6(32'h3ba6ce71),
	.w7(32'h3be7c3c4),
	.w8(32'h3c8ce427),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd10775),
	.w1(32'h3b2cc7f2),
	.w2(32'h3b687904),
	.w3(32'h3bfdea0b),
	.w4(32'hb9b56753),
	.w5(32'h3b1de4a6),
	.w6(32'hb9ddf996),
	.w7(32'h3b5cb24e),
	.w8(32'h3b42ecd2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15011c),
	.w1(32'h3c4f4fee),
	.w2(32'h3c56d86f),
	.w3(32'h3b37e0fd),
	.w4(32'h3bc55a0c),
	.w5(32'h39e95612),
	.w6(32'h3c0d2265),
	.w7(32'h3c201ef6),
	.w8(32'h3c0afc45),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c0596),
	.w1(32'h3cd3973b),
	.w2(32'h3d0a69d9),
	.w3(32'hbc2b6e2c),
	.w4(32'h3c4b3018),
	.w5(32'h3c165c62),
	.w6(32'hbc9b04b2),
	.w7(32'hbb8c0837),
	.w8(32'hbbfc00e7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51e74e),
	.w1(32'hbc9a2cab),
	.w2(32'h3adef099),
	.w3(32'h3b0ca6e6),
	.w4(32'hbc187fb2),
	.w5(32'hbace4e6a),
	.w6(32'h3a363556),
	.w7(32'h3c3e3b37),
	.w8(32'h3c89a1e5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01a9f6),
	.w1(32'hbbcaf06e),
	.w2(32'hbbcec279),
	.w3(32'h3c8f9f3a),
	.w4(32'hbc3ef13b),
	.w5(32'hbb1ea09e),
	.w6(32'hba2ed7b8),
	.w7(32'hbc4c6fb0),
	.w8(32'hbc5a7cac),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e2637),
	.w1(32'hbbfc7b15),
	.w2(32'hbc21a21c),
	.w3(32'h396af64d),
	.w4(32'hbac2b8e5),
	.w5(32'hbbc38188),
	.w6(32'h39bacd02),
	.w7(32'hbc2294ea),
	.w8(32'hbbce2563),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4012f),
	.w1(32'h3c8131ad),
	.w2(32'h3ce708cd),
	.w3(32'hbb9339ce),
	.w4(32'h3c5fc1a0),
	.w5(32'h3ccd847b),
	.w6(32'hbca82360),
	.w7(32'h3c015fc0),
	.w8(32'h3c2bc2c2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9dec6),
	.w1(32'hbbddcb24),
	.w2(32'hbc2a5e06),
	.w3(32'hba256a11),
	.w4(32'hbc14145e),
	.w5(32'hbc00fc20),
	.w6(32'hbbaee37a),
	.w7(32'hbbf9cf1a),
	.w8(32'hbbe19a8f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe45399),
	.w1(32'hba75e117),
	.w2(32'h3b4ac69a),
	.w3(32'hbba5864d),
	.w4(32'h3b09a4dd),
	.w5(32'h3b8b407d),
	.w6(32'hbb2e3e7d),
	.w7(32'h3b54347e),
	.w8(32'h3b632a0e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee0e27),
	.w1(32'hbc35f323),
	.w2(32'hbbdd5102),
	.w3(32'hbaea3668),
	.w4(32'h3bec22f7),
	.w5(32'hbbb7c65c),
	.w6(32'hbcc294c1),
	.w7(32'hbc921148),
	.w8(32'hbbd44c2a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a095c),
	.w1(32'hbc0aba1f),
	.w2(32'hbc657e22),
	.w3(32'hbc183ff3),
	.w4(32'hbb8e1cbc),
	.w5(32'hbbaa3305),
	.w6(32'hbc5767d6),
	.w7(32'hbc1ef649),
	.w8(32'hbc08433d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd51c933),
	.w1(32'h3d0960a3),
	.w2(32'h3d17c2d2),
	.w3(32'h3d07f6d5),
	.w4(32'h3cad38a8),
	.w5(32'h3d12bea4),
	.w6(32'hbdaf5061),
	.w7(32'hbd7987bf),
	.w8(32'hbda2cdaf),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fed2a),
	.w1(32'h3c986c41),
	.w2(32'h3c222083),
	.w3(32'h3ac0fbd6),
	.w4(32'h3c4f5d26),
	.w5(32'h3b3d5331),
	.w6(32'h3c4a1b19),
	.w7(32'h3c0a1096),
	.w8(32'h3b022aa8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c4b5),
	.w1(32'hbb15e6be),
	.w2(32'hbb2197fa),
	.w3(32'hbb3f6bfc),
	.w4(32'hbc0372c7),
	.w5(32'hbc251965),
	.w6(32'hba073921),
	.w7(32'hbac2a6d9),
	.w8(32'h3b55385e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceb97a),
	.w1(32'hba2a4bce),
	.w2(32'hba261923),
	.w3(32'hbbf19e93),
	.w4(32'hbac0cf4c),
	.w5(32'hbab23503),
	.w6(32'h3a895477),
	.w7(32'hbb84d2a6),
	.w8(32'hbb3214d4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a3439),
	.w1(32'h3b3a0e86),
	.w2(32'h3b1c5ddc),
	.w3(32'hbb40aff2),
	.w4(32'h3b37c99e),
	.w5(32'hbb724d33),
	.w6(32'h3c1c32f7),
	.w7(32'h3abc3095),
	.w8(32'h3a7bdc82),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6061f8),
	.w1(32'h3b533a86),
	.w2(32'hbb0db6ee),
	.w3(32'hbb87e02d),
	.w4(32'hbbc88335),
	.w5(32'hbab1cb18),
	.w6(32'hbb0ed9c2),
	.w7(32'hbacbef16),
	.w8(32'hbb0c9680),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaea060),
	.w1(32'hbc28a319),
	.w2(32'hbc5ae09a),
	.w3(32'hbb4a6baf),
	.w4(32'hbc1c38fa),
	.w5(32'hbc2f392d),
	.w6(32'hbbc98eda),
	.w7(32'hbc3b4b92),
	.w8(32'hbbcaf2c6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a2291),
	.w1(32'hbbb7842d),
	.w2(32'hbbc65614),
	.w3(32'hbc875fc6),
	.w4(32'hbbb0bd71),
	.w5(32'hbbe38941),
	.w6(32'h3bfdd488),
	.w7(32'h3ba1491d),
	.w8(32'h3ba480d3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceacad),
	.w1(32'h3a012401),
	.w2(32'h3ba9e2b1),
	.w3(32'h3aa2de6b),
	.w4(32'hba0c3c2b),
	.w5(32'hbb60a0b9),
	.w6(32'hbbb58c3f),
	.w7(32'hbb011798),
	.w8(32'hbbbc6174),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0b22e),
	.w1(32'h3af06c74),
	.w2(32'h3b03b156),
	.w3(32'hbbb05ca8),
	.w4(32'h3b45c52e),
	.w5(32'h3ae9f432),
	.w6(32'h3abe0c50),
	.w7(32'h3af4bc08),
	.w8(32'h3aeba885),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8dea1),
	.w1(32'hbb1d6818),
	.w2(32'h3c1213a4),
	.w3(32'h3aab48bb),
	.w4(32'h3ae7fd74),
	.w5(32'h3c1a7052),
	.w6(32'hba946370),
	.w7(32'h3b986845),
	.w8(32'h3c59b50d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57e470),
	.w1(32'hba8ee680),
	.w2(32'h399624dc),
	.w3(32'h3c4fc988),
	.w4(32'hba87a21c),
	.w5(32'hbba1f466),
	.w6(32'hbb47365e),
	.w7(32'hbba9df98),
	.w8(32'hbb90dbf8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa45ffa),
	.w1(32'hbc05a116),
	.w2(32'hbc4ac473),
	.w3(32'h3a0ea7a6),
	.w4(32'hbc099d36),
	.w5(32'hbc1debb6),
	.w6(32'hbc1d0293),
	.w7(32'hbc4c1d5c),
	.w8(32'hbb9edb0d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56a78d),
	.w1(32'h3b623e5f),
	.w2(32'hb9530c7a),
	.w3(32'hbbddf54d),
	.w4(32'h3c0fd90a),
	.w5(32'h3b493624),
	.w6(32'hbc7b62fe),
	.w7(32'hbaf17a27),
	.w8(32'h3c581e4c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375a3f),
	.w1(32'h3c1fcd63),
	.w2(32'h3c49f3c1),
	.w3(32'hbb2f7884),
	.w4(32'h3adc91e7),
	.w5(32'h3bf6943d),
	.w6(32'h3b9f5160),
	.w7(32'h3bac1ed2),
	.w8(32'h3c008ab8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10e5b9),
	.w1(32'h3bd9ee48),
	.w2(32'h3be8440b),
	.w3(32'h3bc8e9b8),
	.w4(32'h3c1d2a2f),
	.w5(32'h3c23468a),
	.w6(32'h3c041f32),
	.w7(32'h3b30b5aa),
	.w8(32'h3b0ac18d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff58e6),
	.w1(32'h3b1b00ba),
	.w2(32'h383f46b6),
	.w3(32'h3aa363b1),
	.w4(32'h3b5a28fc),
	.w5(32'hbb896ad1),
	.w6(32'hbae28767),
	.w7(32'hbb5db73a),
	.w8(32'h3b0c262b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe45881),
	.w1(32'h3bb3cc21),
	.w2(32'hba6b4b3e),
	.w3(32'hbb3ef8d9),
	.w4(32'h3a43cfac),
	.w5(32'h39f9b736),
	.w6(32'hbc213fe1),
	.w7(32'hbbf80358),
	.w8(32'hbbe3420d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea19cf),
	.w1(32'hbcf005ab),
	.w2(32'hbc6e905d),
	.w3(32'hbc122e8f),
	.w4(32'hbc997bbf),
	.w5(32'hbbfa26a8),
	.w6(32'hbc863aa1),
	.w7(32'hbc4af868),
	.w8(32'h3b7e73aa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ebaa6),
	.w1(32'h3b4711da),
	.w2(32'hb9981618),
	.w3(32'h3c1c38b6),
	.w4(32'h3ba07ab4),
	.w5(32'h3b2830ca),
	.w6(32'h3c176f7e),
	.w7(32'h3b5f8ec8),
	.w8(32'h3bf2fa5d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38960),
	.w1(32'hbbe5e791),
	.w2(32'h3b466f88),
	.w3(32'h3ae7c4c5),
	.w4(32'hbab6f1ce),
	.w5(32'hba3132c4),
	.w6(32'hbc62e9e3),
	.w7(32'hbc26bccc),
	.w8(32'hbbfb79fd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4470b4),
	.w1(32'hbab52980),
	.w2(32'hbb35e0cd),
	.w3(32'h3b80e96f),
	.w4(32'h3b8c89ae),
	.w5(32'h3b64a11e),
	.w6(32'hb9d54de2),
	.w7(32'h3a5915a1),
	.w8(32'hbac671f6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf721d),
	.w1(32'h3bddf918),
	.w2(32'h3c220ede),
	.w3(32'hbaf2acac),
	.w4(32'h3c5d5553),
	.w5(32'h3c363cec),
	.w6(32'hbbaa8401),
	.w7(32'hb9cb70f4),
	.w8(32'h3c2ca46b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb114f14),
	.w1(32'hbc1c2bb1),
	.w2(32'hbb8b33db),
	.w3(32'hbabf09c7),
	.w4(32'hbc2b291f),
	.w5(32'hbb678c78),
	.w6(32'hbb754fba),
	.w7(32'hbc21d8d1),
	.w8(32'hb9ff49ea),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b3d7a),
	.w1(32'h3c3f9fd2),
	.w2(32'h3b839d60),
	.w3(32'h3c37628f),
	.w4(32'h3caeb5cf),
	.w5(32'h3c617722),
	.w6(32'hbcd14c61),
	.w7(32'hbbf84fbf),
	.w8(32'hbc6ddba5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5e9f3),
	.w1(32'hba92edf1),
	.w2(32'hbc12eb64),
	.w3(32'h3b838f8e),
	.w4(32'h3b0b5d16),
	.w5(32'hbb8a6e5f),
	.w6(32'hbc2f2b45),
	.w7(32'hbbdf1ca4),
	.w8(32'hbba1af55),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc396b72),
	.w1(32'h3ab6f6e4),
	.w2(32'h3c8a6d77),
	.w3(32'hbbf83876),
	.w4(32'hbb1efa6b),
	.w5(32'h3b40c27c),
	.w6(32'h3bcb4ec0),
	.w7(32'h3c6c9a9f),
	.w8(32'h3bf9dbaa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b370ec3),
	.w1(32'h3a938420),
	.w2(32'h3c22bffa),
	.w3(32'hbba55a51),
	.w4(32'hbb74b20b),
	.w5(32'h3a320c11),
	.w6(32'hbad24c6d),
	.w7(32'h3c0b1e0a),
	.w8(32'hbac73881),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce66ada),
	.w1(32'hbc68012f),
	.w2(32'hba891a34),
	.w3(32'hbc891b4e),
	.w4(32'hbca2cd59),
	.w5(32'hbc88aa7f),
	.w6(32'hbc9e6b22),
	.w7(32'hbc27087d),
	.w8(32'hbbb6ceb0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21c1fd),
	.w1(32'hbb5d5ecf),
	.w2(32'h3c7437c4),
	.w3(32'hbc4b1c91),
	.w4(32'hbb92a7d1),
	.w5(32'h3c3bb492),
	.w6(32'h3b2d757e),
	.w7(32'h3b583dbb),
	.w8(32'h3ba8a45d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c442157),
	.w1(32'h3bf2d01f),
	.w2(32'h3bed4939),
	.w3(32'h3c12e30e),
	.w4(32'h3b9848f8),
	.w5(32'h3c10da18),
	.w6(32'hbb4c9c66),
	.w7(32'h3b82bd1e),
	.w8(32'hbb289acb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a091),
	.w1(32'hbbb65dcd),
	.w2(32'hbb039744),
	.w3(32'hb9b1e568),
	.w4(32'hbb1d191c),
	.w5(32'h3b724db4),
	.w6(32'hbc5466fc),
	.w7(32'hbc46ff48),
	.w8(32'hbba0a64e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a445022),
	.w1(32'hbc100b81),
	.w2(32'hbc128544),
	.w3(32'h3b84bed8),
	.w4(32'h3b5a9db1),
	.w5(32'h3b21f32f),
	.w6(32'hbc872f3f),
	.w7(32'hbc532f61),
	.w8(32'hbb6ad801),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0a2f6),
	.w1(32'hbb6202c8),
	.w2(32'hbb31773a),
	.w3(32'hbbe7bb4d),
	.w4(32'h3b57f644),
	.w5(32'h3a1b7bfc),
	.w6(32'hbb3a1784),
	.w7(32'hbb3f2091),
	.w8(32'hbb5e5886),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c194),
	.w1(32'h3ba4f859),
	.w2(32'hbb50ab43),
	.w3(32'hbadf4b42),
	.w4(32'h3b8e7e6b),
	.w5(32'hbb4405ea),
	.w6(32'h3b719a11),
	.w7(32'h3aa2122e),
	.w8(32'h3a95c525),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ca963),
	.w1(32'h3c07bb91),
	.w2(32'hb89524d4),
	.w3(32'hbb322d89),
	.w4(32'hba5958ee),
	.w5(32'hbc0164bf),
	.w6(32'hbbd5177f),
	.w7(32'hbb8e26c7),
	.w8(32'hba02d97f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a6d13),
	.w1(32'hb9f379e3),
	.w2(32'hb8cf47e6),
	.w3(32'hbbb94bcf),
	.w4(32'h3a421314),
	.w5(32'h3a390fc3),
	.w6(32'h3b44e115),
	.w7(32'h3b8eac29),
	.w8(32'h3c000705),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0867e),
	.w1(32'hbbfeb362),
	.w2(32'h3bd1f28b),
	.w3(32'h3b6fd702),
	.w4(32'hbb9e7c64),
	.w5(32'h3bcc5987),
	.w6(32'hbbd30f68),
	.w7(32'h3afe640c),
	.w8(32'h3c49deda),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c944a75),
	.w1(32'hbbfcf6e6),
	.w2(32'hbc233bb0),
	.w3(32'h3c744ef6),
	.w4(32'hbbe5cc56),
	.w5(32'hbc42e5f0),
	.w6(32'hbb79a7b0),
	.w7(32'hbc0c2ecd),
	.w8(32'hbc3ffcf8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28de4b),
	.w1(32'hbbcbbd3e),
	.w2(32'hbc711f9e),
	.w3(32'hbbf6daf0),
	.w4(32'hbbcaa11e),
	.w5(32'hbc2f5d04),
	.w6(32'hbb9ab95e),
	.w7(32'hbc1be7ba),
	.w8(32'hbc20c01d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91967f),
	.w1(32'hbbb50dea),
	.w2(32'hba576716),
	.w3(32'hbc431028),
	.w4(32'hbb803fd0),
	.w5(32'hbbd80641),
	.w6(32'hbb84f6e9),
	.w7(32'hbbd579af),
	.w8(32'hbb3e1973),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93239f),
	.w1(32'hbbb3ef64),
	.w2(32'hbc0aed1f),
	.w3(32'h3bc0a610),
	.w4(32'hbb593770),
	.w5(32'hbbf8e9b2),
	.w6(32'hbb9a00a0),
	.w7(32'hbc24c5d1),
	.w8(32'hbbb295e8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb366bc),
	.w1(32'h3b6c351c),
	.w2(32'h3c3f831c),
	.w3(32'h3b50300f),
	.w4(32'h3ca3b48e),
	.w5(32'h3cc05c75),
	.w6(32'hbc82796d),
	.w7(32'hbc4ff6a7),
	.w8(32'hbc0b57a5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9cbb7),
	.w1(32'h3ac4121d),
	.w2(32'hbc094723),
	.w3(32'h3b6d89b3),
	.w4(32'h3b64b2c0),
	.w5(32'hbbebb3e8),
	.w6(32'h3ba56eb7),
	.w7(32'hbbb425cb),
	.w8(32'hbb913281),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39d1b1),
	.w1(32'h3a8c1658),
	.w2(32'h3b9b5d05),
	.w3(32'hbbd4d43a),
	.w4(32'h3bb4b0ff),
	.w5(32'h3ba61daa),
	.w6(32'h3b9a79c2),
	.w7(32'h3bc095ef),
	.w8(32'h39b695c9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1a001),
	.w1(32'hbbb25f6b),
	.w2(32'hbbf8e302),
	.w3(32'h3b62121f),
	.w4(32'hbb6aab30),
	.w5(32'hbb30d84e),
	.w6(32'h3b840a9a),
	.w7(32'h37fd7f21),
	.w8(32'h3ab9a47e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0110aa),
	.w1(32'hbaa826b3),
	.w2(32'h3bc70161),
	.w3(32'hbb2b9a7f),
	.w4(32'hbb0fafe8),
	.w5(32'h3b394ace),
	.w6(32'h3b6a2b72),
	.w7(32'h3be90289),
	.w8(32'h3bfd249e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ca2aa),
	.w1(32'h3c02e7b4),
	.w2(32'h3c348768),
	.w3(32'h3af7161e),
	.w4(32'h3bde6aea),
	.w5(32'h3c088bdc),
	.w6(32'h3b1059b2),
	.w7(32'h3b865c3e),
	.w8(32'h3a17a250),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b529a16),
	.w1(32'h3c30bc02),
	.w2(32'h3c1774f7),
	.w3(32'hbab39752),
	.w4(32'h3b6e6a56),
	.w5(32'h3be3d3b4),
	.w6(32'h3aa3a9f8),
	.w7(32'h3b1be64d),
	.w8(32'hbae73ad3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f979),
	.w1(32'h3b78c9bf),
	.w2(32'h3c1b4e28),
	.w3(32'h3b8a200b),
	.w4(32'h3b0f9f8f),
	.w5(32'h3b9d34e9),
	.w6(32'h3bc7b619),
	.w7(32'h3bb5ad88),
	.w8(32'h3a227284),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac85b28),
	.w1(32'h3c9d4b17),
	.w2(32'h3cd77e7b),
	.w3(32'hb944d18d),
	.w4(32'h3c89e44d),
	.w5(32'h3ca0d2c5),
	.w6(32'hb9e9b6f6),
	.w7(32'h3b8b5f4d),
	.w8(32'h3b70c306),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae551f),
	.w1(32'hbb12d7a4),
	.w2(32'h3c143d74),
	.w3(32'h39ed43a2),
	.w4(32'hba8f3f15),
	.w5(32'h3b7b06ee),
	.w6(32'hbab55cc2),
	.w7(32'h3b106203),
	.w8(32'h3ad8f67c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb053901),
	.w1(32'hbb87aa5d),
	.w2(32'hbc0b074d),
	.w3(32'h3a9ae449),
	.w4(32'hbb20f554),
	.w5(32'hbb838492),
	.w6(32'hbaab1ed2),
	.w7(32'h3b169eee),
	.w8(32'hbb3765c9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79cc50),
	.w1(32'hbc0454a2),
	.w2(32'hbac315a2),
	.w3(32'h3a71c209),
	.w4(32'hbb9813ff),
	.w5(32'hbb049bab),
	.w6(32'hbb234c6a),
	.w7(32'hba191616),
	.w8(32'h3a567ca9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13b855),
	.w1(32'hbb1dda99),
	.w2(32'h3b07850b),
	.w3(32'hbb80b342),
	.w4(32'h3b81f0b7),
	.w5(32'hb91577e8),
	.w6(32'hbbe0fe0c),
	.w7(32'hbbe315d7),
	.w8(32'hbbb07938),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12893c),
	.w1(32'h3c1e6e32),
	.w2(32'h3c874842),
	.w3(32'h3a0536c9),
	.w4(32'h3c0a9dd1),
	.w5(32'h3bc3c26b),
	.w6(32'hbacc0e93),
	.w7(32'h3bcec73c),
	.w8(32'h3ac8cb6c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85844a),
	.w1(32'h3b9291ec),
	.w2(32'h3c86b5ac),
	.w3(32'hbb733a72),
	.w4(32'h3c495d0c),
	.w5(32'h3c98e485),
	.w6(32'hbc42aa00),
	.w7(32'h3c48504a),
	.w8(32'h3c40d3a7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd041b1),
	.w1(32'h3bdc1e1d),
	.w2(32'h3c6e7a5d),
	.w3(32'hbb1784c7),
	.w4(32'h3c331f9f),
	.w5(32'h3c6fb93e),
	.w6(32'hbc7d6841),
	.w7(32'hbb1e673b),
	.w8(32'hbada448c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cacd0),
	.w1(32'h3be9cf3d),
	.w2(32'h3aed1536),
	.w3(32'h3b05a2ba),
	.w4(32'h3b5cff4a),
	.w5(32'h3b7da885),
	.w6(32'hbace865d),
	.w7(32'h3bbeaf3c),
	.w8(32'h3bb94d23),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3642b1),
	.w1(32'h3aad6235),
	.w2(32'h3afa6eab),
	.w3(32'h3916edd5),
	.w4(32'h39bf1372),
	.w5(32'h3af92189),
	.w6(32'h3b404b63),
	.w7(32'h3b61d4f1),
	.w8(32'h3afbbe10),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3b94),
	.w1(32'h3b8d6709),
	.w2(32'hb9c03342),
	.w3(32'h3914d31f),
	.w4(32'h3bd32e80),
	.w5(32'h3b08750b),
	.w6(32'h3b80dcaa),
	.w7(32'h3b9efb58),
	.w8(32'h3bc44289),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05527b),
	.w1(32'hbbafef9e),
	.w2(32'hbb2d7fde),
	.w3(32'h39e57b47),
	.w4(32'hbb578c7e),
	.w5(32'hbabeabef),
	.w6(32'h3a07f31b),
	.w7(32'h3a9c5871),
	.w8(32'hba015ee2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb74a75),
	.w1(32'hbbd06c94),
	.w2(32'h3b0dec3e),
	.w3(32'hbb0fe8aa),
	.w4(32'hbae8171d),
	.w5(32'h3be91de5),
	.w6(32'hbbae9cbc),
	.w7(32'hba413e5c),
	.w8(32'hba23cbf0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43b0ce),
	.w1(32'h380ce995),
	.w2(32'h3b8a6766),
	.w3(32'hb98f666d),
	.w4(32'h388799c2),
	.w5(32'hb946a594),
	.w6(32'hbb82d819),
	.w7(32'hbaae7f4d),
	.w8(32'hbb397211),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fd77a),
	.w1(32'hbb9badc2),
	.w2(32'hbba198e6),
	.w3(32'h3a149c5f),
	.w4(32'hbbe148d1),
	.w5(32'hbc01fe53),
	.w6(32'hbb77ca9f),
	.w7(32'h3943ec74),
	.w8(32'hba0482a9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b3f22),
	.w1(32'h3c19521a),
	.w2(32'hbbbbf6a7),
	.w3(32'h3aa13a46),
	.w4(32'h3c28c3f4),
	.w5(32'hb91577e6),
	.w6(32'h3c1b966a),
	.w7(32'h3b9b6fb3),
	.w8(32'hbb765fde),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32776e),
	.w1(32'h3c82adf4),
	.w2(32'h3b4df2a6),
	.w3(32'hbc426974),
	.w4(32'h3c1c53d0),
	.w5(32'hba263ca6),
	.w6(32'h3bc83b1b),
	.w7(32'h3ad7efd6),
	.w8(32'hbbafdc13),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83159e),
	.w1(32'h3c2c5818),
	.w2(32'h3c4105aa),
	.w3(32'hbc40ef86),
	.w4(32'h3c144772),
	.w5(32'h3bc0aa89),
	.w6(32'h3c817491),
	.w7(32'h3c31a44a),
	.w8(32'h3c049ed5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b865be1),
	.w1(32'hba4e8bce),
	.w2(32'h3b9591fb),
	.w3(32'hbbe7e02e),
	.w4(32'hbb9bb520),
	.w5(32'hbaf7337a),
	.w6(32'hb65119ec),
	.w7(32'h3b587c49),
	.w8(32'h3adfca64),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b958dc5),
	.w1(32'h3c8ac75c),
	.w2(32'h3c2efbc5),
	.w3(32'hbb2f0107),
	.w4(32'h3c5736a6),
	.w5(32'h3bcc040b),
	.w6(32'h3a3e4035),
	.w7(32'h3b9b242a),
	.w8(32'hb5a330f2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd160d),
	.w1(32'hb97cc3f4),
	.w2(32'hb716aa71),
	.w3(32'h3b75c69b),
	.w4(32'hbb2cca7d),
	.w5(32'hbb42710f),
	.w6(32'h3b3fb283),
	.w7(32'hbb82c3ff),
	.w8(32'hbb8473dd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3623f7),
	.w1(32'h3b20b93c),
	.w2(32'h3b5cca43),
	.w3(32'hbb1b6454),
	.w4(32'h3aa3b51a),
	.w5(32'h3a85eb1f),
	.w6(32'h3ba6c445),
	.w7(32'h39b78ac8),
	.w8(32'h3bc250bc),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b05e7),
	.w1(32'h3b214b2a),
	.w2(32'h3b8907d7),
	.w3(32'h3bf059b5),
	.w4(32'hbb237368),
	.w5(32'h3929c69d),
	.w6(32'hb9e12ce3),
	.w7(32'hba18e95e),
	.w8(32'h3a9b2564),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5050e7),
	.w1(32'h3b5d2e38),
	.w2(32'h3af5412a),
	.w3(32'h3a37f218),
	.w4(32'h3b4dc127),
	.w5(32'h3ada933b),
	.w6(32'h3b97d8d8),
	.w7(32'h3a792cd5),
	.w8(32'hbbf475d4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb411ad8),
	.w1(32'h3ac0e7c8),
	.w2(32'hbbbd9170),
	.w3(32'hb8fae2f0),
	.w4(32'hbac0c38e),
	.w5(32'h3b725584),
	.w6(32'h3a60eb8c),
	.w7(32'h3b4aea83),
	.w8(32'hba867296),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba56540),
	.w1(32'hba88fceb),
	.w2(32'hb95e60ad),
	.w3(32'hbbcd519b),
	.w4(32'hbb911a0c),
	.w5(32'hbb639675),
	.w6(32'hb9a97c28),
	.w7(32'hbb2be219),
	.w8(32'hbb9762a8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab297ff),
	.w1(32'hbb99c48d),
	.w2(32'hba2b2f29),
	.w3(32'hbb3617c9),
	.w4(32'h3b0b33f7),
	.w5(32'h3a53ea20),
	.w6(32'hbb14e34d),
	.w7(32'h3bc44d8e),
	.w8(32'hb9aba3eb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71f635),
	.w1(32'h3b98e3d4),
	.w2(32'h3c1d2179),
	.w3(32'hbb014e07),
	.w4(32'h3a612bfd),
	.w5(32'h3b269ee1),
	.w6(32'hbacd63ed),
	.w7(32'h3c472b88),
	.w8(32'h3c1a4c8c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd4249),
	.w1(32'hbcd9833c),
	.w2(32'hbac2ea42),
	.w3(32'h3bf2b291),
	.w4(32'hbbc98ec9),
	.w5(32'h3be2303f),
	.w6(32'hbce80fbd),
	.w7(32'hbc786bc1),
	.w8(32'h3c361d47),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8db98),
	.w1(32'h3a498d2e),
	.w2(32'h3b73414d),
	.w3(32'h3cb092d3),
	.w4(32'h3b477c06),
	.w5(32'h3b97232d),
	.w6(32'h3b02b5ae),
	.w7(32'h3ad45fc8),
	.w8(32'h3aa312db),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d027a),
	.w1(32'h3af40995),
	.w2(32'h3bc85475),
	.w3(32'h3b2d738c),
	.w4(32'h3b97e0ce),
	.w5(32'h3baf856f),
	.w6(32'h3b5b36e6),
	.w7(32'h3b9808aa),
	.w8(32'h3b09bc91),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae2e1c),
	.w1(32'hbb456d1d),
	.w2(32'hbc1d0046),
	.w3(32'h3b49f918),
	.w4(32'hbaf8c795),
	.w5(32'hbbec8d6e),
	.w6(32'h3af4f6a2),
	.w7(32'hbb4c46da),
	.w8(32'hbac51806),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed86d0),
	.w1(32'h3c541b56),
	.w2(32'h39d76124),
	.w3(32'hbbe946b5),
	.w4(32'h3c0d956f),
	.w5(32'h396c3599),
	.w6(32'h3b67a8ee),
	.w7(32'h3925f534),
	.w8(32'hbbecec61),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc919ef3),
	.w1(32'h3a38238e),
	.w2(32'hb8d3f969),
	.w3(32'hbc80d190),
	.w4(32'hbbd99e62),
	.w5(32'hbb8d3a97),
	.w6(32'hba8ff19c),
	.w7(32'hbbc8f721),
	.w8(32'hbc282192),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae2262),
	.w1(32'hbb0dda12),
	.w2(32'hbb82299b),
	.w3(32'hbbaf70dc),
	.w4(32'hbb945c66),
	.w5(32'hbbbf1be1),
	.w6(32'h37c81ec2),
	.w7(32'h3aae31fa),
	.w8(32'h3b8f50b9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc9547),
	.w1(32'hbb654572),
	.w2(32'hba079a0c),
	.w3(32'h3bcbbf00),
	.w4(32'hbb10d3bc),
	.w5(32'hbba7b1e0),
	.w6(32'h3b23d1a7),
	.w7(32'h3b98336e),
	.w8(32'h3ac9fefc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc047f61),
	.w1(32'hbbc02b18),
	.w2(32'hbbc66bbe),
	.w3(32'hbbbf91eb),
	.w4(32'hba72edd7),
	.w5(32'hbbd60ea4),
	.w6(32'hbbb3eaa4),
	.w7(32'hbba2ad6d),
	.w8(32'hbb888095),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdadb74),
	.w1(32'hbb2df988),
	.w2(32'h3af25f54),
	.w3(32'hbc300248),
	.w4(32'hbb14e69c),
	.w5(32'h3b8307e2),
	.w6(32'hbab76bbb),
	.w7(32'h3a903036),
	.w8(32'h3b235fe1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28b68c),
	.w1(32'h3b750cd7),
	.w2(32'h3aa831f3),
	.w3(32'h3b2b74e2),
	.w4(32'h3b037300),
	.w5(32'h3a75eb18),
	.w6(32'hbb38d1f6),
	.w7(32'hbb00c620),
	.w8(32'hbb4b4bd5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba36ece),
	.w1(32'h3bdc9d1f),
	.w2(32'h3b850370),
	.w3(32'hbb10a0df),
	.w4(32'h3bb17e6b),
	.w5(32'h3b777f34),
	.w6(32'h3b8a254a),
	.w7(32'h3b0d57b0),
	.w8(32'h3b9118ea),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca34a),
	.w1(32'h3b757b2f),
	.w2(32'h3a84bdcc),
	.w3(32'h3b9531c9),
	.w4(32'h3bc128ce),
	.w5(32'h3b2400e5),
	.w6(32'hbc28fe76),
	.w7(32'hbb0f9e4b),
	.w8(32'hbb700a66),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb200ac4),
	.w1(32'hbbe2a6d7),
	.w2(32'hbbae70fb),
	.w3(32'hbb291f2a),
	.w4(32'h394ee48d),
	.w5(32'hbb486c38),
	.w6(32'hbc14b48e),
	.w7(32'hbc03ca65),
	.w8(32'hbbce6c2c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14896f),
	.w1(32'h3b1cb82b),
	.w2(32'h3c19f231),
	.w3(32'hbc2cb5f4),
	.w4(32'h3b120451),
	.w5(32'h3b8edbe6),
	.w6(32'h3a81581d),
	.w7(32'h3b75549c),
	.w8(32'h3a029026),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97d308),
	.w1(32'hbc1de927),
	.w2(32'hbc00b32a),
	.w3(32'hbbe904d0),
	.w4(32'hb9ee7d42),
	.w5(32'hbbf9d9fe),
	.w6(32'hbb62b2de),
	.w7(32'h3a049198),
	.w8(32'hbaca7588),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e5f69),
	.w1(32'h3b5eb914),
	.w2(32'h3bf91b70),
	.w3(32'hbc0f5466),
	.w4(32'h3bafec1f),
	.w5(32'h3b8bd1cd),
	.w6(32'h3b9e4a63),
	.w7(32'h3b848d7f),
	.w8(32'h3c192e15),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07e629),
	.w1(32'h3c7759aa),
	.w2(32'hbbb4d99b),
	.w3(32'h3b978747),
	.w4(32'h3c281b22),
	.w5(32'hbb966fee),
	.w6(32'h3c272dd7),
	.w7(32'h3ac51210),
	.w8(32'hbc1155f3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb9905),
	.w1(32'h3b382704),
	.w2(32'hbbbc8f2a),
	.w3(32'hbc7b013f),
	.w4(32'h3a8f6602),
	.w5(32'hbafd32ae),
	.w6(32'hb833e84b),
	.w7(32'hbb9e327a),
	.w8(32'hbbe44569),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfbebe),
	.w1(32'h3a1c5fe0),
	.w2(32'h3a20ff3c),
	.w3(32'hbb99ecd9),
	.w4(32'hb9a4c3af),
	.w5(32'h3bae91a6),
	.w6(32'hb8934310),
	.w7(32'h3a838563),
	.w8(32'hbb8210de),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac477ea),
	.w1(32'hbc2f4f53),
	.w2(32'hbb0a33a4),
	.w3(32'hba967deb),
	.w4(32'h3acdd6b5),
	.w5(32'hbb371aeb),
	.w6(32'hbaf07756),
	.w7(32'hbbb9632e),
	.w8(32'hbbfbfa4d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ae0c2),
	.w1(32'hb981b91e),
	.w2(32'hbaf1e671),
	.w3(32'hbbc49532),
	.w4(32'hbb42c659),
	.w5(32'hbb923654),
	.w6(32'h394fea75),
	.w7(32'hbb0a5ea3),
	.w8(32'h392dbc24),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafe621),
	.w1(32'hbbe5b499),
	.w2(32'hbce6c4ee),
	.w3(32'hbbb5c80b),
	.w4(32'hbb06de93),
	.w5(32'hbc873b95),
	.w6(32'h3ba76bf6),
	.w7(32'hbc0edf0b),
	.w8(32'h3b628df2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule