module layer_10_featuremap_47(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42b25d),
	.w1(32'h3c2e6dc0),
	.w2(32'hbc20a0ff),
	.w3(32'h3c851c3b),
	.w4(32'h3c8a9df0),
	.w5(32'hbbb12f67),
	.w6(32'h3c37386f),
	.w7(32'h3c1a3611),
	.w8(32'h3b2f9379),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3029a),
	.w1(32'h3c1e347a),
	.w2(32'hba0c2a3e),
	.w3(32'hbaaf6ccf),
	.w4(32'hbbcd3f28),
	.w5(32'h3baa4d91),
	.w6(32'h3bda396e),
	.w7(32'hbc9a95ce),
	.w8(32'hbb78101a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c5377),
	.w1(32'h3bf947cb),
	.w2(32'hbb6f8d9f),
	.w3(32'h3b674533),
	.w4(32'h3b94be01),
	.w5(32'hbbdc59ca),
	.w6(32'h3b266f1e),
	.w7(32'hbb12df14),
	.w8(32'h3a81b165),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6dcbb),
	.w1(32'h3c12cf61),
	.w2(32'h3ba60a1b),
	.w3(32'hbbdda3e1),
	.w4(32'hbbaf2eec),
	.w5(32'h3c853c4e),
	.w6(32'h3a4a8851),
	.w7(32'hbb84e318),
	.w8(32'h3917590b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce91fa),
	.w1(32'hbbaf1e53),
	.w2(32'hbafe3e8b),
	.w3(32'h3be73e80),
	.w4(32'h3b17aea9),
	.w5(32'h3acf8cb1),
	.w6(32'hba5c2315),
	.w7(32'h3b8203db),
	.w8(32'h3bad291a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5207a6),
	.w1(32'h3b57bb35),
	.w2(32'hbab8e5e7),
	.w3(32'h3a84e8d0),
	.w4(32'h3be5c84e),
	.w5(32'hbb86c54c),
	.w6(32'hb9b51078),
	.w7(32'h3ac11c27),
	.w8(32'hba9a111f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb6a18),
	.w1(32'h38537920),
	.w2(32'h3b7d5c0f),
	.w3(32'hbbe9f8f6),
	.w4(32'h3b868110),
	.w5(32'hb9f73696),
	.w6(32'hbbdd1cc3),
	.w7(32'h3c13a19d),
	.w8(32'h3bf8a1ae),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab592a),
	.w1(32'hbb688f35),
	.w2(32'hbb304e2d),
	.w3(32'hbc2ab671),
	.w4(32'hbc149564),
	.w5(32'hbc54862d),
	.w6(32'hbc0b42da),
	.w7(32'h3c44fbe2),
	.w8(32'hbc46f6ba),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c721731),
	.w1(32'h3c27446c),
	.w2(32'h3b83c329),
	.w3(32'h3c43f31b),
	.w4(32'h3c029b51),
	.w5(32'h3c1c9061),
	.w6(32'h3bcd20c8),
	.w7(32'h3b828318),
	.w8(32'h3bfee3d2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8e3d6),
	.w1(32'hbc175637),
	.w2(32'h3bd738bd),
	.w3(32'h3c9a4055),
	.w4(32'hbaef53b5),
	.w5(32'h39b02062),
	.w6(32'h3c92127b),
	.w7(32'h3bc7b990),
	.w8(32'hbad07b34),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12ae6d),
	.w1(32'h3b08fc5f),
	.w2(32'h3bc935e3),
	.w3(32'h3a3c52bc),
	.w4(32'h3b147145),
	.w5(32'h3b218b39),
	.w6(32'h39097618),
	.w7(32'h3ae93e97),
	.w8(32'h3b882c73),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c1ab6),
	.w1(32'hbc080498),
	.w2(32'h3c13f9b7),
	.w3(32'hbb80e063),
	.w4(32'h3c396317),
	.w5(32'h3b29479a),
	.w6(32'hbbc75594),
	.w7(32'h3c290a08),
	.w8(32'h3c548716),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eede6),
	.w1(32'hbc68cf8e),
	.w2(32'hbabd57cf),
	.w3(32'hbbbf4f8e),
	.w4(32'hbc396ef4),
	.w5(32'h3accdcaa),
	.w6(32'hbbedad1f),
	.w7(32'hbb8c25ca),
	.w8(32'h3b170bd6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b7c98),
	.w1(32'h3be2899c),
	.w2(32'hb88f60d5),
	.w3(32'h3c083ffe),
	.w4(32'h3b89abd2),
	.w5(32'hbc0895db),
	.w6(32'h3bc7b9ca),
	.w7(32'h3ba724f8),
	.w8(32'hbc151283),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82037d),
	.w1(32'hb8e55acc),
	.w2(32'hbc1d2629),
	.w3(32'h3b0d01bd),
	.w4(32'hbc171d27),
	.w5(32'hbc86c1f4),
	.w6(32'h3b889be1),
	.w7(32'hbc1784ed),
	.w8(32'hbc2275eb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8aa79),
	.w1(32'hbc1269ab),
	.w2(32'h3b1733a1),
	.w3(32'hbcc7604e),
	.w4(32'hbd0176d2),
	.w5(32'hbc09a6e1),
	.w6(32'hbc33e070),
	.w7(32'hbcdfa2ed),
	.w8(32'hbc820f5c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe63d1),
	.w1(32'h3aa5c0c9),
	.w2(32'h3c0afe4c),
	.w3(32'h39e3f100),
	.w4(32'h3a754121),
	.w5(32'h3c655704),
	.w6(32'hba5ac2f3),
	.w7(32'h3a86f332),
	.w8(32'h3ca90a89),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c9fc),
	.w1(32'hbc7342f3),
	.w2(32'hbc3f2e78),
	.w3(32'h3c4418d3),
	.w4(32'hbac42fc0),
	.w5(32'hbb96cc35),
	.w6(32'h3c8adefb),
	.w7(32'h3ce35691),
	.w8(32'hbb5b6ed0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda87d0),
	.w1(32'hbc4045be),
	.w2(32'hbca4f9b0),
	.w3(32'hbb5e07a3),
	.w4(32'hbb832553),
	.w5(32'hbce5e6fd),
	.w6(32'h3ae7d850),
	.w7(32'h3c2d0843),
	.w8(32'hbc4d53ca),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc457cab),
	.w1(32'h3b99192b),
	.w2(32'hba7d311f),
	.w3(32'hbcd75e12),
	.w4(32'hbc09e9b2),
	.w5(32'h38975b85),
	.w6(32'hbc88633d),
	.w7(32'hbc7f0ca7),
	.w8(32'h3970059d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a0e28),
	.w1(32'hbaf498cb),
	.w2(32'h39d239ca),
	.w3(32'hbb21f9c8),
	.w4(32'hbb4e0be0),
	.w5(32'hbb667dd4),
	.w6(32'h3a41381d),
	.w7(32'h37932751),
	.w8(32'h3bc0a170),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e8771),
	.w1(32'h3bfbe5ee),
	.w2(32'hbb89d76e),
	.w3(32'hbbd142a8),
	.w4(32'hbb7b15f1),
	.w5(32'hbbeee6de),
	.w6(32'h3b7f75ea),
	.w7(32'hbba62882),
	.w8(32'hbb944c81),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85223d),
	.w1(32'hbc6db7cc),
	.w2(32'hbba1760e),
	.w3(32'hbb87192d),
	.w4(32'h38f41f05),
	.w5(32'h3a1ee4e3),
	.w6(32'h3ba3aaa7),
	.w7(32'h3c35c61b),
	.w8(32'h3bb9fc57),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ef493),
	.w1(32'hba9a3c28),
	.w2(32'h3c32e2c0),
	.w3(32'hbbcb610a),
	.w4(32'hbb9400b1),
	.w5(32'h3c425649),
	.w6(32'hbbb00518),
	.w7(32'hbba2e549),
	.w8(32'h3bca9242),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7217a9),
	.w1(32'h3bb14ae0),
	.w2(32'h3c0af3c9),
	.w3(32'h3c2572f4),
	.w4(32'hbb3d2ddc),
	.w5(32'h3c0f7134),
	.w6(32'h3c6e7488),
	.w7(32'hbbbf6102),
	.w8(32'hbb0fe683),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd9c04),
	.w1(32'hb956fb1f),
	.w2(32'h3a5b3c45),
	.w3(32'h3bcc5268),
	.w4(32'hbb76e896),
	.w5(32'hba5864fd),
	.w6(32'h3b09de17),
	.w7(32'h3ba85244),
	.w8(32'hba423d6d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5e73f),
	.w1(32'h3b196341),
	.w2(32'h39b44552),
	.w3(32'hbbc4bead),
	.w4(32'hbbb54f9f),
	.w5(32'h3a0e44df),
	.w6(32'hbb4384a9),
	.w7(32'hbb63da6c),
	.w8(32'hb8bb3013),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cf26e),
	.w1(32'h3b26fab0),
	.w2(32'hbc2799a5),
	.w3(32'h3bcce094),
	.w4(32'hbbe9250c),
	.w5(32'hbb5ba491),
	.w6(32'h3b187aff),
	.w7(32'hbbfcf6cd),
	.w8(32'hbcbdfb4b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b2536),
	.w1(32'h3bbaabf7),
	.w2(32'hbb26e29e),
	.w3(32'h3c0be98f),
	.w4(32'h3c2e9e2f),
	.w5(32'hbc05432f),
	.w6(32'h390e10c3),
	.w7(32'hbb0d4f35),
	.w8(32'hbb67d361),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0fe13),
	.w1(32'h3b8337ef),
	.w2(32'h3bc68121),
	.w3(32'h3b64e0aa),
	.w4(32'hbbee7e30),
	.w5(32'h3b9e0cfc),
	.w6(32'h3c61a2e6),
	.w7(32'hbc423f27),
	.w8(32'hbc0c0761),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ece60),
	.w1(32'hbb96f1d4),
	.w2(32'h3a4659bc),
	.w3(32'h3b85a463),
	.w4(32'h3b34040a),
	.w5(32'hbce22b3f),
	.w6(32'hbb2b7db6),
	.w7(32'hbad36cfa),
	.w8(32'h3ca97c5f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1956c),
	.w1(32'hbc0bd824),
	.w2(32'hbbe43f89),
	.w3(32'hbcd0e80b),
	.w4(32'hbcdf60c0),
	.w5(32'hbc1ee0eb),
	.w6(32'h3c6d709d),
	.w7(32'h3bf1c122),
	.w8(32'h3c0c8c12),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d04da),
	.w1(32'hbc1b3289),
	.w2(32'h3aea5166),
	.w3(32'hbbcc4aa2),
	.w4(32'hbbc3c76e),
	.w5(32'h39701300),
	.w6(32'hbba8e576),
	.w7(32'hbb71a23f),
	.w8(32'hb9fc09b7),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75953c),
	.w1(32'h3bb22380),
	.w2(32'h3990f980),
	.w3(32'h3bc2be12),
	.w4(32'h3ba64029),
	.w5(32'h3be0580c),
	.w6(32'h3b729fc3),
	.w7(32'h3ad24c4b),
	.w8(32'hbacbda0b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fe5d0),
	.w1(32'hbbe3d403),
	.w2(32'h3a02b4e3),
	.w3(32'h3add8e0a),
	.w4(32'hbb2f4da9),
	.w5(32'hba151768),
	.w6(32'hbbee5b20),
	.w7(32'hbc570ea4),
	.w8(32'h3a1d5bac),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfca241),
	.w1(32'hbb22eda2),
	.w2(32'h3bee7205),
	.w3(32'hbbd7ab4b),
	.w4(32'h387f1c4e),
	.w5(32'hbcb2c2ef),
	.w6(32'hbbc644f3),
	.w7(32'h3a213b52),
	.w8(32'h3bf52ef7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d3589),
	.w1(32'hbd01bc7b),
	.w2(32'h3c6078ea),
	.w3(32'hbc8d40f1),
	.w4(32'hbcda1d79),
	.w5(32'h3c95905e),
	.w6(32'h39a3a9c2),
	.w7(32'hbb407d37),
	.w8(32'h3cbe3a29),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceade35),
	.w1(32'h3c98abce),
	.w2(32'hbbfb75d7),
	.w3(32'h3cc406e9),
	.w4(32'h3c2b27cb),
	.w5(32'h3c9559df),
	.w6(32'h3cefbbc8),
	.w7(32'h3b242c07),
	.w8(32'hbc086131),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2b593),
	.w1(32'h3ce2fc7c),
	.w2(32'h3caefe80),
	.w3(32'h3cc08473),
	.w4(32'h3cc4581e),
	.w5(32'h3bbf69ad),
	.w6(32'h3c54dcf1),
	.w7(32'h3b6a6a5d),
	.w8(32'h3c17a550),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4cbb3),
	.w1(32'h3ba64f4e),
	.w2(32'hbb867419),
	.w3(32'h3c4c5636),
	.w4(32'hb91fd4a0),
	.w5(32'hbafe66f7),
	.w6(32'h3af3d441),
	.w7(32'h3b88ac88),
	.w8(32'h399fb827),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2bdfa),
	.w1(32'hbb302172),
	.w2(32'hbbaebdb0),
	.w3(32'hbb1c8bc8),
	.w4(32'h3ba0b050),
	.w5(32'h3b85fa8f),
	.w6(32'h3c2d3158),
	.w7(32'h3c8caf91),
	.w8(32'hbbc343d5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd922af),
	.w1(32'h3b8ddf85),
	.w2(32'hbbb5e691),
	.w3(32'h3be5e93f),
	.w4(32'h3c000b2e),
	.w5(32'hbc5427d0),
	.w6(32'hbbae68e6),
	.w7(32'hbaf70ef0),
	.w8(32'h3c0046e9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21ee9e),
	.w1(32'hb986a975),
	.w2(32'hba925410),
	.w3(32'hbc7591ef),
	.w4(32'hbc373d3a),
	.w5(32'h3a94b637),
	.w6(32'h3c95dfcc),
	.w7(32'h3bcd8d17),
	.w8(32'h3868fee0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9ca06),
	.w1(32'hbbaa27b4),
	.w2(32'h3b127c55),
	.w3(32'hbb54a9c7),
	.w4(32'hbc1028a0),
	.w5(32'hbc7c1117),
	.w6(32'hbaa49ff4),
	.w7(32'h39d2365b),
	.w8(32'hbb192d41),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfa31f),
	.w1(32'h3ba86a0c),
	.w2(32'h3cae58d2),
	.w3(32'hbc8f0bf8),
	.w4(32'hbcc9a131),
	.w5(32'hbbfd2058),
	.w6(32'hbbae5ec5),
	.w7(32'hbc8fc00d),
	.w8(32'h3b8ffba1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15761e),
	.w1(32'h3be98143),
	.w2(32'h3c179edf),
	.w3(32'hbccebea7),
	.w4(32'hbc911dc5),
	.w5(32'h3c1debcc),
	.w6(32'hbb4013de),
	.w7(32'hbbf9664a),
	.w8(32'hbb05deb8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad34a0),
	.w1(32'hbc5bf071),
	.w2(32'h3988d23d),
	.w3(32'h3bd105da),
	.w4(32'h3b3eb6ac),
	.w5(32'h3c27e260),
	.w6(32'hbc2977d7),
	.w7(32'hba9f245a),
	.w8(32'hb9c74015),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc814c6),
	.w1(32'hbcc38fcb),
	.w2(32'hbc0dccd0),
	.w3(32'hbc873ec9),
	.w4(32'hbc365d7f),
	.w5(32'hbc37422a),
	.w6(32'hbca11eca),
	.w7(32'h3ac87456),
	.w8(32'h3bf9ad75),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9804bb3),
	.w1(32'h39ad9ed6),
	.w2(32'hbb456816),
	.w3(32'hbb447801),
	.w4(32'hbb7a08f5),
	.w5(32'h3a9e8f8e),
	.w6(32'hbad9aea9),
	.w7(32'hbb418422),
	.w8(32'h3cd3400a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ad88c),
	.w1(32'hb99c54ad),
	.w2(32'hbb0716e9),
	.w3(32'hbbe873c4),
	.w4(32'h3b6fc7ed),
	.w5(32'h3cc2cef7),
	.w6(32'h3d14f4f7),
	.w7(32'h3cc6cc3a),
	.w8(32'hbb7eaa1a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b351f55),
	.w1(32'h3ba41f2a),
	.w2(32'h3a3b3682),
	.w3(32'h3cc6d0e9),
	.w4(32'h3c4e3e26),
	.w5(32'h3b349ba0),
	.w6(32'hbc1be42c),
	.w7(32'hbbc1dbc6),
	.w8(32'hbb10cf18),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82fddc),
	.w1(32'hba9c3274),
	.w2(32'hbbb5518a),
	.w3(32'hbb479cf9),
	.w4(32'hbc0ba929),
	.w5(32'h3c4244cd),
	.w6(32'hbc21481e),
	.w7(32'hbca41900),
	.w8(32'hbb8943cc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1559f),
	.w1(32'h3bcaca0f),
	.w2(32'h3b8849a1),
	.w3(32'h3cbfccf1),
	.w4(32'h3c911eab),
	.w5(32'hbc81fc7a),
	.w6(32'hbc820a92),
	.w7(32'hbc2e4eb5),
	.w8(32'h3c0fd0ff),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e5c43),
	.w1(32'hbc8d9a4c),
	.w2(32'hbb3f44f6),
	.w3(32'hbcef3d30),
	.w4(32'hbcdaf023),
	.w5(32'hbc8274d7),
	.w6(32'h3b4522c7),
	.w7(32'h3c3bbd6a),
	.w8(32'h3c955274),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef19c5),
	.w1(32'hbb1a5c8d),
	.w2(32'hbc0eb0ba),
	.w3(32'hbc9ec4d1),
	.w4(32'hbc5d2a1c),
	.w5(32'h3bd2a8c9),
	.w6(32'h3ca90d2b),
	.w7(32'h3c95fbc2),
	.w8(32'h3c1ea733),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb764d),
	.w1(32'hbbc4216f),
	.w2(32'hbabf0231),
	.w3(32'h3c60e4e1),
	.w4(32'h3c426dc6),
	.w5(32'hbbe5270c),
	.w6(32'h3c47653b),
	.w7(32'h3c30ec73),
	.w8(32'hbc644e98),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1d068),
	.w1(32'hbbe64772),
	.w2(32'hbb701979),
	.w3(32'h3bd24976),
	.w4(32'h3bb6d4b2),
	.w5(32'h3b7bf778),
	.w6(32'hbbeafcda),
	.w7(32'h3ad538fe),
	.w8(32'h3b636d83),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936a29f),
	.w1(32'h378bf383),
	.w2(32'hba73557d),
	.w3(32'h3b2745e7),
	.w4(32'h3b50d673),
	.w5(32'hb8fe08a6),
	.w6(32'h3b714ee7),
	.w7(32'h3a7339d7),
	.w8(32'h3b30ae85),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f750b),
	.w1(32'h3a6e1cdd),
	.w2(32'hba995fbb),
	.w3(32'h390ad634),
	.w4(32'h3ba4f6a4),
	.w5(32'hbbb25960),
	.w6(32'h3c05cf6c),
	.w7(32'h3c689f58),
	.w8(32'h3c072f48),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98b34c),
	.w1(32'h3b8bb514),
	.w2(32'hbc0453fe),
	.w3(32'hbbe0dfed),
	.w4(32'hbbe16907),
	.w5(32'h3c24f901),
	.w6(32'h3c02ec46),
	.w7(32'h3bc4ebec),
	.w8(32'hbb9f43bd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc979bd1),
	.w1(32'hbc467f13),
	.w2(32'hbc61232c),
	.w3(32'hb9e1bf5d),
	.w4(32'hbbb1fb73),
	.w5(32'hba4dcb00),
	.w6(32'hb97f417c),
	.w7(32'hbb01c46a),
	.w8(32'hbc41df08),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9bfcc),
	.w1(32'hbb8da492),
	.w2(32'hbbeab242),
	.w3(32'h3bc5fab2),
	.w4(32'hbb946635),
	.w5(32'h398bbb05),
	.w6(32'hbb0f2b7d),
	.w7(32'hbb9ec4a3),
	.w8(32'hbcbbee62),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c8a1e),
	.w1(32'h3bcd1a94),
	.w2(32'h3aeef8be),
	.w3(32'h3aa21f33),
	.w4(32'h3c6cf132),
	.w5(32'hbb184006),
	.w6(32'hbcc505d3),
	.w7(32'hbca24f39),
	.w8(32'h3b73bc30),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab648ba),
	.w1(32'hbb0816ec),
	.w2(32'hbaa35ab9),
	.w3(32'hbbd140a9),
	.w4(32'hbc043003),
	.w5(32'hbc496352),
	.w6(32'h3c1cb224),
	.w7(32'h3b70983b),
	.w8(32'hba7b33f2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc722d),
	.w1(32'hbb1012b2),
	.w2(32'h39c54eea),
	.w3(32'hbc48906b),
	.w4(32'hbc30e742),
	.w5(32'h3ae3226b),
	.w6(32'h3b53084b),
	.w7(32'h3c696c21),
	.w8(32'h3b4d3c54),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab562f6),
	.w1(32'hbaabd2f2),
	.w2(32'hbae88dad),
	.w3(32'h3895845a),
	.w4(32'hba4ecd17),
	.w5(32'h3b4b4949),
	.w6(32'h3b13bfa2),
	.w7(32'hb7d03d14),
	.w8(32'hbbaa7aee),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca58daf),
	.w1(32'hbcae986d),
	.w2(32'hbc83cb46),
	.w3(32'h3b51ff46),
	.w4(32'hbc3c1ae1),
	.w5(32'hbc28a688),
	.w6(32'hbb6fa7c7),
	.w7(32'hba736831),
	.w8(32'hbcd23f40),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a13eb),
	.w1(32'hbc640697),
	.w2(32'h3bf697d7),
	.w3(32'hbc12cbc0),
	.w4(32'hbbeee3be),
	.w5(32'h3bf53bf8),
	.w6(32'hbc995b33),
	.w7(32'h3ae4cc1d),
	.w8(32'hbc92002b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a977c),
	.w1(32'hbc293b6e),
	.w2(32'hbc4f19da),
	.w3(32'h3c7def20),
	.w4(32'h3bb24f94),
	.w5(32'hbc1f1f66),
	.w6(32'hbcab4e06),
	.w7(32'hbcb35af0),
	.w8(32'hbc427530),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1c9b0),
	.w1(32'hbb8c2669),
	.w2(32'h3c308a44),
	.w3(32'h3a480d29),
	.w4(32'hbc24e63b),
	.w5(32'h3c6c6f42),
	.w6(32'h3be71179),
	.w7(32'hbcda0caf),
	.w8(32'hbb174d2c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5219c),
	.w1(32'hbb3366ad),
	.w2(32'hbac52de0),
	.w3(32'h3ba70655),
	.w4(32'h3b4027e7),
	.w5(32'hba647bbc),
	.w6(32'h3be075aa),
	.w7(32'h3b57c0a4),
	.w8(32'h3ba8e602),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2e9a9),
	.w1(32'h3a794aff),
	.w2(32'h399cd676),
	.w3(32'hba142ae4),
	.w4(32'h3bf18ecc),
	.w5(32'h3c211d76),
	.w6(32'hbb8f5b7c),
	.w7(32'h3a13b10a),
	.w8(32'h39adf15c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc016ddd),
	.w1(32'hbc431995),
	.w2(32'h3aebb6cc),
	.w3(32'h3bfd643e),
	.w4(32'hba493b30),
	.w5(32'hbcf7ede0),
	.w6(32'hbbdd0d36),
	.w7(32'h3be9f1cc),
	.w8(32'h3c481994),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f03e),
	.w1(32'h3af41e32),
	.w2(32'hbb9a2cbb),
	.w3(32'hbcc1924f),
	.w4(32'hbce1d106),
	.w5(32'hbb89f4ff),
	.w6(32'h3c8ec908),
	.w7(32'h3c12002e),
	.w8(32'hbbfb9d1d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8555fc),
	.w1(32'hbbc3b27f),
	.w2(32'hbb85c799),
	.w3(32'h388650ee),
	.w4(32'hbb0503ca),
	.w5(32'hbb855207),
	.w6(32'hbbed223c),
	.w7(32'hbc0b03a6),
	.w8(32'hbbafd129),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6adb31),
	.w1(32'hbc53121e),
	.w2(32'h3be2827f),
	.w3(32'hbc554cab),
	.w4(32'hbc49d2e3),
	.w5(32'hbba2ea7f),
	.w6(32'hbc5cd396),
	.w7(32'hbbd47cc0),
	.w8(32'hbc8bc48b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc542c1),
	.w1(32'hbc329170),
	.w2(32'hbc1a9ea4),
	.w3(32'hbb2f1a5e),
	.w4(32'hbbd9dcc2),
	.w5(32'hbc9c1100),
	.w6(32'hbd3ea599),
	.w7(32'hbc97880a),
	.w8(32'hbb45b331),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b542371),
	.w1(32'h3b788a36),
	.w2(32'hba47d7bf),
	.w3(32'hbbe9c6e9),
	.w4(32'hbc9f5a73),
	.w5(32'hbbbe30d3),
	.w6(32'hbc32154e),
	.w7(32'hbcabf785),
	.w8(32'hbbe03147),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49f057),
	.w1(32'hbc669628),
	.w2(32'hba093654),
	.w3(32'hbb8283b1),
	.w4(32'hbbacb4f3),
	.w5(32'hba1d6204),
	.w6(32'hbc4886d8),
	.w7(32'hbbf037df),
	.w8(32'hbbb79557),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27fe0f),
	.w1(32'hbc200c5e),
	.w2(32'h3b199d8a),
	.w3(32'h3ba1bf84),
	.w4(32'h3ac6a3be),
	.w5(32'h3b9111c2),
	.w6(32'h3bd3a965),
	.w7(32'h3b4b3e6d),
	.w8(32'hbbc10866),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1837c),
	.w1(32'hbbaa41d5),
	.w2(32'h3b267e12),
	.w3(32'h3aea2931),
	.w4(32'hbb2a6508),
	.w5(32'h3bfa5672),
	.w6(32'hbbd495ba),
	.w7(32'hbc52f2f6),
	.w8(32'hbc094ccc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b41c2),
	.w1(32'hbc5c449c),
	.w2(32'h3bf2237b),
	.w3(32'h395f0cff),
	.w4(32'hbb87b319),
	.w5(32'h3bb1967c),
	.w6(32'hbbffa74c),
	.w7(32'hbb25d813),
	.w8(32'h3b4e41a5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef1017),
	.w1(32'hbb8f3856),
	.w2(32'hbbbe3954),
	.w3(32'h3bd19316),
	.w4(32'hbb6db506),
	.w5(32'h3b555c92),
	.w6(32'hbbfc6048),
	.w7(32'hbb2585c4),
	.w8(32'hbc0d295c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd825),
	.w1(32'hbb65fb4e),
	.w2(32'h3a6679c5),
	.w3(32'h3b872048),
	.w4(32'h3b961123),
	.w5(32'h3c46c21d),
	.w6(32'hbc98a9de),
	.w7(32'hbc067da1),
	.w8(32'hbc284317),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7d415),
	.w1(32'hbc11c605),
	.w2(32'hbc33b20e),
	.w3(32'h3c4e82d6),
	.w4(32'h3c86b8f8),
	.w5(32'h3b784612),
	.w6(32'hbbbeb589),
	.w7(32'hbb661521),
	.w8(32'hbbb055c2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb069316),
	.w1(32'hb9e55303),
	.w2(32'hbbb9c3a5),
	.w3(32'hbb6c16d2),
	.w4(32'h3b545c9d),
	.w5(32'hba9de4f5),
	.w6(32'hbc025dad),
	.w7(32'hbb8f5168),
	.w8(32'hbab50ce7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82b0e6),
	.w1(32'h3bdd4671),
	.w2(32'h3c38ed85),
	.w3(32'hba8893b3),
	.w4(32'h3b547940),
	.w5(32'h3c123de9),
	.w6(32'h3b19e89a),
	.w7(32'hbbda38ed),
	.w8(32'h3ac3565f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2a57a),
	.w1(32'h3a9828ed),
	.w2(32'hbbd49f60),
	.w3(32'h3b82b671),
	.w4(32'h3b7cd9a7),
	.w5(32'h3c6d48bc),
	.w6(32'hbac478d9),
	.w7(32'hbacd9c6d),
	.w8(32'hbb2e3791),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3e7f3),
	.w1(32'hbb30d413),
	.w2(32'h3be48c8e),
	.w3(32'h3bfba483),
	.w4(32'h3c77f5eb),
	.w5(32'h3c34d80d),
	.w6(32'hbb8646d0),
	.w7(32'hbc7e32ee),
	.w8(32'h3c1a0c75),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac07a64),
	.w1(32'h3ad9950d),
	.w2(32'h3b884b96),
	.w3(32'h3c170e46),
	.w4(32'h3c1f4ed3),
	.w5(32'hbbdbb804),
	.w6(32'h3bb40da4),
	.w7(32'h3cb9621d),
	.w8(32'h3af34eba),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c870cc1),
	.w1(32'h3c032a8e),
	.w2(32'h3ab636c3),
	.w3(32'h3bb8e6e9),
	.w4(32'h3b3639f7),
	.w5(32'h3ab5b153),
	.w6(32'h3b81aa63),
	.w7(32'hbb84d761),
	.w8(32'h3c4a9eb5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1bff5f),
	.w1(32'hbc5e57ad),
	.w2(32'h3ba138ee),
	.w3(32'hbcac20a0),
	.w4(32'hbba720d2),
	.w5(32'h3c0e234b),
	.w6(32'h3c5c9f36),
	.w7(32'h3c444e14),
	.w8(32'h3b685b2b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ff7f9),
	.w1(32'hba8ef8a7),
	.w2(32'h3bc6de2e),
	.w3(32'h3babceaf),
	.w4(32'h3b5cda4c),
	.w5(32'h3bc60b07),
	.w6(32'h3a98997e),
	.w7(32'h3b63c47d),
	.w8(32'hba4c2bb3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad567c7),
	.w1(32'h3b83a9e1),
	.w2(32'hbc387d95),
	.w3(32'h3c3e3201),
	.w4(32'h3bc93deb),
	.w5(32'hba990522),
	.w6(32'h3c404dbe),
	.w7(32'h3c3c5933),
	.w8(32'hbcb0a450),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3be63e),
	.w1(32'h3c2726e5),
	.w2(32'h3c01785c),
	.w3(32'h3c3a9bc0),
	.w4(32'h3bc908a4),
	.w5(32'hbc13d53c),
	.w6(32'hbc966786),
	.w7(32'hbc4442cc),
	.w8(32'h3ced78c0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf0b16),
	.w1(32'h3ad0f2e3),
	.w2(32'hbc08e8dc),
	.w3(32'hbc389a24),
	.w4(32'hbc0c8ad4),
	.w5(32'hbaa58452),
	.w6(32'h3d47eb01),
	.w7(32'h3cf14fdd),
	.w8(32'hbc3ea1d7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcafaa),
	.w1(32'hbc0f67f8),
	.w2(32'h3bde74a9),
	.w3(32'hbab0f456),
	.w4(32'hbb4b962d),
	.w5(32'h3a8ee4e8),
	.w6(32'hbc65d5e3),
	.w7(32'hbc00b9cf),
	.w8(32'hbc4fad35),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcea68),
	.w1(32'hbbbedacd),
	.w2(32'h3b84d273),
	.w3(32'h3a6379c0),
	.w4(32'h3c0344e5),
	.w5(32'hbc01a9f2),
	.w6(32'hbcd10a2a),
	.w7(32'hbc6f2b19),
	.w8(32'h3c56315d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd14698b),
	.w1(32'hbcaeed17),
	.w2(32'h3bd4b33d),
	.w3(32'hbc95463e),
	.w4(32'hbcc4a260),
	.w5(32'h3c977962),
	.w6(32'h3aaede2a),
	.w7(32'h3b83bb58),
	.w8(32'h3b843da7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65bf1a),
	.w1(32'hbccaa3ff),
	.w2(32'hbc7959fb),
	.w3(32'hbc5343bf),
	.w4(32'hbbdea9d4),
	.w5(32'hbc9fb3a1),
	.w6(32'hbcf92754),
	.w7(32'hbcffd459),
	.w8(32'h3d3ff97e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf5acc4),
	.w1(32'h3c6ad2ec),
	.w2(32'h3b652382),
	.w3(32'h3c97e1ba),
	.w4(32'hbbacc7bd),
	.w5(32'hbc9fcece),
	.w6(32'h3d8d8169),
	.w7(32'h3d1d4846),
	.w8(32'h3cde4050),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde4ac6),
	.w1(32'hbc2eedf1),
	.w2(32'h3c8d4b6f),
	.w3(32'hbca64a18),
	.w4(32'hbcaf1e15),
	.w5(32'h3ca8e3fa),
	.w6(32'h3d393106),
	.w7(32'h3d0b506e),
	.w8(32'h3b153e23),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb137f9),
	.w1(32'hbc9f1989),
	.w2(32'h3c06f2e1),
	.w3(32'h3bded5f5),
	.w4(32'h3c8279d1),
	.w5(32'h3c36c19a),
	.w6(32'h39ec7355),
	.w7(32'h3c4dba72),
	.w8(32'h3c5f0d59),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e67d),
	.w1(32'hbb17693a),
	.w2(32'hbb00e756),
	.w3(32'h39c820ba),
	.w4(32'hbaff072b),
	.w5(32'h3c27bcec),
	.w6(32'h3a8cffe3),
	.w7(32'hbb16ba11),
	.w8(32'hbc402b99),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd5b66a),
	.w1(32'hbcdde84f),
	.w2(32'hbcb8c6a1),
	.w3(32'hbba50b69),
	.w4(32'hbc4e7b2e),
	.w5(32'hbbcce712),
	.w6(32'hbc8ec164),
	.w7(32'hbce98644),
	.w8(32'h3bc0c519),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30fdde),
	.w1(32'hbc065d72),
	.w2(32'hbbfe640e),
	.w3(32'hbbdabfa5),
	.w4(32'hbb4a7bed),
	.w5(32'hbb0c8d6b),
	.w6(32'hbbe6c175),
	.w7(32'hbc279db7),
	.w8(32'h3c0f85ca),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30f6cf),
	.w1(32'h3ad184f7),
	.w2(32'hbb8a4464),
	.w3(32'hba9e9ef7),
	.w4(32'h3a97013f),
	.w5(32'hbc042ef8),
	.w6(32'hbb14c459),
	.w7(32'hba55d382),
	.w8(32'h3a9f890a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6c0e),
	.w1(32'h3b42cc66),
	.w2(32'hbb284eba),
	.w3(32'hbc0b6e9c),
	.w4(32'hbb66a839),
	.w5(32'h3c2208c7),
	.w6(32'h3b209a84),
	.w7(32'hbb83752d),
	.w8(32'hbc0b9f05),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f5f0d),
	.w1(32'hbb06ebee),
	.w2(32'h3a731cbc),
	.w3(32'h3c88d74c),
	.w4(32'h3b132f65),
	.w5(32'hbc93efb5),
	.w6(32'hbac8e419),
	.w7(32'h3bf84aba),
	.w8(32'h3ce71580),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35b768),
	.w1(32'h3b98c572),
	.w2(32'h3c450b52),
	.w3(32'hbc4af946),
	.w4(32'hbc74c7cc),
	.w5(32'h3c1018f6),
	.w6(32'h3d07c830),
	.w7(32'h3cc37307),
	.w8(32'hbc13612d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dee62),
	.w1(32'h3c4f67be),
	.w2(32'hbbc3b16d),
	.w3(32'hbb8b885c),
	.w4(32'h3bcb23fe),
	.w5(32'h3c49a54f),
	.w6(32'hbc458d61),
	.w7(32'hbcca4e29),
	.w8(32'hbbd24802),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19173f),
	.w1(32'hbbb7197e),
	.w2(32'hbb873279),
	.w3(32'h3bab28b4),
	.w4(32'hb9b524ad),
	.w5(32'h3b1a8514),
	.w6(32'hba35def9),
	.w7(32'hbb318818),
	.w8(32'hb986559a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc737241),
	.w1(32'hbc09b236),
	.w2(32'h3c050dec),
	.w3(32'hbb7d3c0b),
	.w4(32'hbbd68b6c),
	.w5(32'hbc8df4f9),
	.w6(32'hbb46d3b8),
	.w7(32'hbbc520ee),
	.w8(32'h3c51fce4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe7df1),
	.w1(32'hbc062b59),
	.w2(32'hbc2f18b5),
	.w3(32'hbcb63445),
	.w4(32'hbcfe6c81),
	.w5(32'hbc1ef7e2),
	.w6(32'h3c45d91c),
	.w7(32'hbaa9403a),
	.w8(32'h3a572288),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf27163),
	.w1(32'hba157b3a),
	.w2(32'h3b924e00),
	.w3(32'hbbdc58e5),
	.w4(32'hbb897125),
	.w5(32'h3b7c441f),
	.w6(32'h3c60ab0d),
	.w7(32'h3c35fa44),
	.w8(32'h3a2b4939),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1b1b1),
	.w1(32'h3b60149a),
	.w2(32'h3a361233),
	.w3(32'hbaba91b3),
	.w4(32'h3af0c6b0),
	.w5(32'hbb63fe83),
	.w6(32'hb9b44581),
	.w7(32'hbb39c819),
	.w8(32'hbbe33ce2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac749bb),
	.w1(32'hba051030),
	.w2(32'hbb47cb47),
	.w3(32'h39228067),
	.w4(32'h3b15f404),
	.w5(32'hbbb0b340),
	.w6(32'hbb7a2c00),
	.w7(32'hbb2d290c),
	.w8(32'hb9f72d0b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57c149),
	.w1(32'h3abbf8a4),
	.w2(32'hbbac7ef3),
	.w3(32'hbb349082),
	.w4(32'hbae43f33),
	.w5(32'hbcf1390d),
	.w6(32'h3bb57ff4),
	.w7(32'h3ac66391),
	.w8(32'h3bbcb02b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23dfdc),
	.w1(32'hbc1d3c34),
	.w2(32'hbb8e54fe),
	.w3(32'hbca874a9),
	.w4(32'hbc9ac8f7),
	.w5(32'hbc1d7549),
	.w6(32'h3b992791),
	.w7(32'h3b877f2f),
	.w8(32'h3cc8d42c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2890f9),
	.w1(32'hbc1b7ebd),
	.w2(32'h3c3c8f76),
	.w3(32'hbbd4ff99),
	.w4(32'hbc4ca148),
	.w5(32'h3b1c505a),
	.w6(32'h3d1c2562),
	.w7(32'h3cc27c2b),
	.w8(32'hbb81abdc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab036ff),
	.w1(32'h3b201947),
	.w2(32'h39ecf436),
	.w3(32'hb9c35c43),
	.w4(32'h3c06271c),
	.w5(32'h3b67f7ea),
	.w6(32'hbcd96bbf),
	.w7(32'hbceee9fb),
	.w8(32'hbab75118),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf61896),
	.w1(32'hbc1e91cc),
	.w2(32'h3a9e4af0),
	.w3(32'h3a125cfd),
	.w4(32'hb895b5cd),
	.w5(32'h3a11326b),
	.w6(32'hbb9da26b),
	.w7(32'hba61bdb7),
	.w8(32'h3b02ac4c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc29f8),
	.w1(32'h3bf0ed34),
	.w2(32'h397e3b53),
	.w3(32'h3c041dde),
	.w4(32'hbb0b21a1),
	.w5(32'h386209f8),
	.w6(32'h3c3f0333),
	.w7(32'hbc00e9ad),
	.w8(32'hbc1ceaed),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef8604),
	.w1(32'hbb58093b),
	.w2(32'hbb47ccc4),
	.w3(32'h3af835f9),
	.w4(32'h3a82d422),
	.w5(32'hba08127f),
	.w6(32'hbc090de7),
	.w7(32'hbc999d42),
	.w8(32'hbb24a234),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a4d16),
	.w1(32'h3aa3fafa),
	.w2(32'hba714ccf),
	.w3(32'h3b74ba9e),
	.w4(32'h3b35e945),
	.w5(32'h3c29e9e5),
	.w6(32'hb9dc6cb7),
	.w7(32'hbb88de08),
	.w8(32'hb98c53e6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28c3b3),
	.w1(32'hba424762),
	.w2(32'hbc06289a),
	.w3(32'hbaf6bb95),
	.w4(32'hba2d046d),
	.w5(32'h3ba50910),
	.w6(32'hbb86eb24),
	.w7(32'hbc143785),
	.w8(32'hbad74863),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a111d),
	.w1(32'hbc1735cc),
	.w2(32'hbb78c86b),
	.w3(32'h3ae82d6b),
	.w4(32'hbb17716e),
	.w5(32'hbb1b6ff5),
	.w6(32'hbb81efaf),
	.w7(32'h3b4661fb),
	.w8(32'hbb0ec5c9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc57cab),
	.w1(32'hbc384973),
	.w2(32'h3bd3d3a8),
	.w3(32'hbc97a8c2),
	.w4(32'hbbce97cc),
	.w5(32'hbba7b296),
	.w6(32'hbc76fea8),
	.w7(32'hbaa191cb),
	.w8(32'h3c1ea884),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fa37a),
	.w1(32'hbc4699e3),
	.w2(32'h3a8cb6d9),
	.w3(32'hbbaa9b85),
	.w4(32'hbc3cf73b),
	.w5(32'h39e40fc6),
	.w6(32'h3b376167),
	.w7(32'h3b81e973),
	.w8(32'h3c1c3ee6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb154c00),
	.w1(32'hbb6888f1),
	.w2(32'hbb2d049d),
	.w3(32'hbba9c69f),
	.w4(32'hbc18c085),
	.w5(32'hbc44a4b2),
	.w6(32'h3c96b1fd),
	.w7(32'h3cd90439),
	.w8(32'h3c65f615),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1709c5),
	.w1(32'hbbf613ab),
	.w2(32'h3ac32ebc),
	.w3(32'hbb85a5b2),
	.w4(32'hbbb2a050),
	.w5(32'hbc1ca2d2),
	.w6(32'h3c753b65),
	.w7(32'h3c516d5d),
	.w8(32'hbad4432b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babfa7b),
	.w1(32'h3acbf504),
	.w2(32'hbb7021b0),
	.w3(32'hbc17744d),
	.w4(32'hbb905ff9),
	.w5(32'hbb5391f9),
	.w6(32'h39f8affd),
	.w7(32'hbc84ea4e),
	.w8(32'hbaafefe6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97388e),
	.w1(32'hbc132890),
	.w2(32'hbc6874ee),
	.w3(32'hbc6674b5),
	.w4(32'hbc1e662a),
	.w5(32'hbc123f10),
	.w6(32'hbc094153),
	.w7(32'hbb4f6457),
	.w8(32'hbb68e4ea),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a6fbc),
	.w1(32'hbb447f27),
	.w2(32'h3bad16fb),
	.w3(32'hb97c60ad),
	.w4(32'hbc0f38d4),
	.w5(32'h3b9963bc),
	.w6(32'h3c33d64b),
	.w7(32'h3be78f9a),
	.w8(32'hbbe8bd8c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc945020),
	.w1(32'hbcb5680b),
	.w2(32'hbb3884a7),
	.w3(32'hbc03b2af),
	.w4(32'hbc17b49f),
	.w5(32'hbc548818),
	.w6(32'hbc261dcd),
	.w7(32'hbb951282),
	.w8(32'h3bbe26e6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc30e00),
	.w1(32'h3b4c2de0),
	.w2(32'h3ab2290c),
	.w3(32'hbbbf596c),
	.w4(32'hbc074280),
	.w5(32'hbbf8656d),
	.w6(32'h3c83ece1),
	.w7(32'h3af5339f),
	.w8(32'h3bb6f0d7),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a2780),
	.w1(32'hbb8f50c6),
	.w2(32'hba612866),
	.w3(32'hbc7f460a),
	.w4(32'hbc0d2278),
	.w5(32'hbb85200a),
	.w6(32'h3a4b9cd4),
	.w7(32'hbc0686d8),
	.w8(32'h3b999eaf),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58303c),
	.w1(32'hbb7b8e68),
	.w2(32'h3bbd08af),
	.w3(32'hbbebd0c3),
	.w4(32'h3b6e9e08),
	.w5(32'h3bef7f6e),
	.w6(32'h3c095721),
	.w7(32'h3c9d8719),
	.w8(32'h3c0d8f65),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe6469),
	.w1(32'h39fe9667),
	.w2(32'h3aa7acb4),
	.w3(32'h3b1331e1),
	.w4(32'h3b2627f9),
	.w5(32'hbc1fa236),
	.w6(32'hba60f356),
	.w7(32'hbbc14bdb),
	.w8(32'h3bcb9649),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc708832),
	.w1(32'hbc2dad8a),
	.w2(32'h3b812ec3),
	.w3(32'hbc1ded62),
	.w4(32'hbbb233bb),
	.w5(32'hbb62807b),
	.w6(32'h3c274a72),
	.w7(32'hbb9799db),
	.w8(32'hbb97d495),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d8434),
	.w1(32'h3ab70bb1),
	.w2(32'h3bfcd2c2),
	.w3(32'hbb0e96b8),
	.w4(32'hbb1942f9),
	.w5(32'hb89960b9),
	.w6(32'h3a947a35),
	.w7(32'hbb058275),
	.w8(32'hbc370939),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92f138),
	.w1(32'h3c8f2bbd),
	.w2(32'hba2fc6f4),
	.w3(32'h3c9aad22),
	.w4(32'h3b26623d),
	.w5(32'h3bb793c3),
	.w6(32'h3c40dd9e),
	.w7(32'hbbda9184),
	.w8(32'h3c97352e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4750e9),
	.w1(32'h3a139669),
	.w2(32'h39a320ca),
	.w3(32'h3b921edf),
	.w4(32'h3af78df7),
	.w5(32'h3a80f77a),
	.w6(32'h3cbdce94),
	.w7(32'h3ce1d640),
	.w8(32'h3bc44cb1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39620367),
	.w1(32'hb9b15c98),
	.w2(32'hbb0cd940),
	.w3(32'hbb3be16d),
	.w4(32'hbb8d4467),
	.w5(32'h3a278dfb),
	.w6(32'h3beda1b3),
	.w7(32'h3b1a9161),
	.w8(32'hbb925cbd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf107a9),
	.w1(32'hbb32e16d),
	.w2(32'hb98dad67),
	.w3(32'h3ad29685),
	.w4(32'h3913b9a6),
	.w5(32'hbb961b4b),
	.w6(32'hbad9b585),
	.w7(32'hbb302edd),
	.w8(32'h3c15021b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc09906),
	.w1(32'hbbf90bdb),
	.w2(32'hb9aaace4),
	.w3(32'hbb9dab3c),
	.w4(32'hbc3b57bd),
	.w5(32'hb9977aef),
	.w6(32'h3c1dd899),
	.w7(32'h3b626a59),
	.w8(32'hbc128023),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47d6cc),
	.w1(32'h3bb7e624),
	.w2(32'h3be5f0c1),
	.w3(32'h3ae0b4bb),
	.w4(32'hba1eeee9),
	.w5(32'hbaac69b2),
	.w6(32'h3b461c58),
	.w7(32'hbc03d681),
	.w8(32'h38fe4364),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71a1dc),
	.w1(32'hbbed0516),
	.w2(32'hbb1ee85d),
	.w3(32'hbcb135f0),
	.w4(32'hbbdaa101),
	.w5(32'hbba2e44a),
	.w6(32'hbc0f79d9),
	.w7(32'h3b103949),
	.w8(32'hbc0a51be),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acee305),
	.w1(32'hbab38268),
	.w2(32'h3bf82de1),
	.w3(32'h3a80bbef),
	.w4(32'hbba38dd7),
	.w5(32'h3c73f7be),
	.w6(32'h39d85dba),
	.w7(32'hb96fac44),
	.w8(32'hbc2576a2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff563e),
	.w1(32'h3b3f8c52),
	.w2(32'h3bb96a2a),
	.w3(32'h3c7e0024),
	.w4(32'h3cae17f5),
	.w5(32'hbb05d553),
	.w6(32'hbccea6f1),
	.w7(32'hbc86adae),
	.w8(32'hbb77e905),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2daf38),
	.w1(32'hba90952a),
	.w2(32'h3c0be5c7),
	.w3(32'h3ad76edc),
	.w4(32'h3a2405c2),
	.w5(32'h3bc6a38f),
	.w6(32'hbba2d3f4),
	.w7(32'hbbe50997),
	.w8(32'h3b0d2f9c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40b732),
	.w1(32'hbc3e7f60),
	.w2(32'hbba9e962),
	.w3(32'hba9f2c81),
	.w4(32'hbb23a090),
	.w5(32'hbaef1667),
	.w6(32'h3a9ec54d),
	.w7(32'h3baa59a5),
	.w8(32'hbbfe6b6b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee65a1),
	.w1(32'hbaef2928),
	.w2(32'hbc1341bf),
	.w3(32'hbbeb5d4a),
	.w4(32'hbca5804e),
	.w5(32'h3cbc4025),
	.w6(32'hbbb53fd2),
	.w7(32'hbc8385ef),
	.w8(32'hbc31a595),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6c77e),
	.w1(32'h3c4a25ed),
	.w2(32'h3c169c17),
	.w3(32'h3c04b29b),
	.w4(32'h3b19dc19),
	.w5(32'h3be14dd4),
	.w6(32'h3c663ecb),
	.w7(32'h3c9bad07),
	.w8(32'hbc9a3989),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82281a),
	.w1(32'h3c728879),
	.w2(32'h3af8013e),
	.w3(32'h3bbe46d9),
	.w4(32'h3b296bf0),
	.w5(32'h3a8eaf0f),
	.w6(32'hbca4c30c),
	.w7(32'hbd01d851),
	.w8(32'h3a560ea5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e036b),
	.w1(32'h3acb01e7),
	.w2(32'hbbcdfc85),
	.w3(32'h3b852cf5),
	.w4(32'h3a1eadd5),
	.w5(32'hbc7c80cf),
	.w6(32'h3be6e1d3),
	.w7(32'h3a5e0b6b),
	.w8(32'hbbc80d43),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc160f10),
	.w1(32'h3ba0e29a),
	.w2(32'h3bf4d216),
	.w3(32'hbc949578),
	.w4(32'hbbc79c76),
	.w5(32'h3b360488),
	.w6(32'hbbc1528e),
	.w7(32'hbb55072b),
	.w8(32'h3b90edcb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd78bf8),
	.w1(32'h3b51ac81),
	.w2(32'hbb8beb19),
	.w3(32'hbbcd582e),
	.w4(32'hbc15a6bb),
	.w5(32'hbbaa3227),
	.w6(32'hbb24557d),
	.w7(32'hbc0a2d4d),
	.w8(32'hbb47f733),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab21c4),
	.w1(32'hbb1ef09b),
	.w2(32'h3aa2c4f0),
	.w3(32'hbb5cc219),
	.w4(32'hbb02399d),
	.w5(32'h3ba4ea77),
	.w6(32'hbb211df4),
	.w7(32'h3a2c8d8c),
	.w8(32'hba62fadf),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac391db),
	.w1(32'hbbbb9c31),
	.w2(32'hbbd13637),
	.w3(32'h3b514a47),
	.w4(32'hbb90b5c7),
	.w5(32'h3bb78c6d),
	.w6(32'hbad2db37),
	.w7(32'hbbc66e0b),
	.w8(32'h3bdab649),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc528d61),
	.w1(32'hbc04703f),
	.w2(32'h3ab6c0b4),
	.w3(32'hbc0dd664),
	.w4(32'hbad1a052),
	.w5(32'hbb89a812),
	.w6(32'hbb64ec3c),
	.w7(32'hbbab527a),
	.w8(32'h3bad0432),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08a79e),
	.w1(32'h3b012dfe),
	.w2(32'h3b57963b),
	.w3(32'h3a14e49b),
	.w4(32'h3b108465),
	.w5(32'h3c84648d),
	.w6(32'h3b047da5),
	.w7(32'h3b7197ef),
	.w8(32'h3c84444f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d059a),
	.w1(32'h3ba5b0c2),
	.w2(32'hbac743b8),
	.w3(32'h3c825316),
	.w4(32'h3bad8ce8),
	.w5(32'hbb8e7cd6),
	.w6(32'h3c7acccb),
	.w7(32'hbb8df757),
	.w8(32'hbb96d8d0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb15e88),
	.w1(32'hbbb2fe42),
	.w2(32'hbb70ab2f),
	.w3(32'hbbeffd83),
	.w4(32'hbbd80608),
	.w5(32'hbbd733be),
	.w6(32'hbbd74482),
	.w7(32'hbbd6aa0a),
	.w8(32'hbc09ebd8),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaac868),
	.w1(32'hbc6f2108),
	.w2(32'hbc8689ea),
	.w3(32'hbca272f3),
	.w4(32'hbc8e9d0f),
	.w5(32'hbcb10f14),
	.w6(32'hbcc0e217),
	.w7(32'hbca4b8d7),
	.w8(32'hbbebe206),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc042d74),
	.w1(32'hbb31f9b6),
	.w2(32'h3bfa2232),
	.w3(32'hbbc716ae),
	.w4(32'hbb628eb0),
	.w5(32'h3b8d4e12),
	.w6(32'h39a8fc22),
	.w7(32'hb9c5167d),
	.w8(32'hbbbf09e0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec4a33),
	.w1(32'hbc8dd763),
	.w2(32'hbba7c17e),
	.w3(32'hbc372488),
	.w4(32'hbcb0ca1d),
	.w5(32'hbb51eb1b),
	.w6(32'hbc7ffde0),
	.w7(32'hbc57b7db),
	.w8(32'hbba7176f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fbd42),
	.w1(32'hbafd6d29),
	.w2(32'h3bce8d35),
	.w3(32'hba7a585f),
	.w4(32'h3b5e4de4),
	.w5(32'h3bd712ca),
	.w6(32'h3c2dd737),
	.w7(32'h3b9862e0),
	.w8(32'h39a10716),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf3f9d),
	.w1(32'hbbabb7d8),
	.w2(32'h3c32a619),
	.w3(32'hbbd62da1),
	.w4(32'hba9c6349),
	.w5(32'h3c13de0f),
	.w6(32'hbc7f4c4f),
	.w7(32'hbb9bca5d),
	.w8(32'h3c865457),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3af1f9),
	.w1(32'h3b85ba54),
	.w2(32'h3c136b3e),
	.w3(32'hba169cfa),
	.w4(32'hbbdb6203),
	.w5(32'h3bbcc346),
	.w6(32'hbbdadd0c),
	.w7(32'hbc2ce0f9),
	.w8(32'h3b85c8c4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be541f6),
	.w1(32'h3b9ef419),
	.w2(32'h3bf47e86),
	.w3(32'h3bae6ec1),
	.w4(32'hbb91f782),
	.w5(32'h3b9683e6),
	.w6(32'h3b281b1d),
	.w7(32'hbbe9ee9e),
	.w8(32'h3b3a0619),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae95a06),
	.w1(32'h3b08021c),
	.w2(32'h3c142fa5),
	.w3(32'h3b35bed4),
	.w4(32'hb914a015),
	.w5(32'h3c8739e5),
	.w6(32'h3b36c1ef),
	.w7(32'h393c8410),
	.w8(32'h3c6db97d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8da110),
	.w1(32'h3b834777),
	.w2(32'hbc0f4f48),
	.w3(32'h3c727d55),
	.w4(32'h3b1c5790),
	.w5(32'hbc88541d),
	.w6(32'h3c90edbe),
	.w7(32'hb8768995),
	.w8(32'hbc8b1136),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08d93f),
	.w1(32'h3aa4674a),
	.w2(32'hbb96a102),
	.w3(32'hbbf9b665),
	.w4(32'h3b3b69a9),
	.w5(32'hbbe60b85),
	.w6(32'h3bbf6920),
	.w7(32'h3bcd47fb),
	.w8(32'h3b328346),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc703d7d),
	.w1(32'hbc4c6236),
	.w2(32'h3c6d0354),
	.w3(32'hbc28ca82),
	.w4(32'hbc735eb2),
	.w5(32'h3cd32e4a),
	.w6(32'hbc3f6daf),
	.w7(32'hbbe07b21),
	.w8(32'h3c69d31e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bad11),
	.w1(32'h3c1e71da),
	.w2(32'hbaf12756),
	.w3(32'h3cb9b38f),
	.w4(32'h3be453d8),
	.w5(32'hbb666fe3),
	.w6(32'h3b468be1),
	.w7(32'hbbb767da),
	.w8(32'hbb2b7f12),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d959),
	.w1(32'h3b57ea39),
	.w2(32'h3a5a51fe),
	.w3(32'h3a6fbd16),
	.w4(32'h3988ab2c),
	.w5(32'h3adcaeca),
	.w6(32'h3bc49cdb),
	.w7(32'h3b27c163),
	.w8(32'h3b27ec85),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5adf12),
	.w1(32'h3bbf6ea2),
	.w2(32'hbb03b24f),
	.w3(32'h3bc747bb),
	.w4(32'h3be2de17),
	.w5(32'h3a93b6c5),
	.w6(32'h3c01774f),
	.w7(32'h3bbf3505),
	.w8(32'hba744fb8),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ab5c1),
	.w1(32'hbac1f7ed),
	.w2(32'h3c282551),
	.w3(32'hba9cf6e5),
	.w4(32'hbb13ae58),
	.w5(32'h3c5b5843),
	.w6(32'hbb9e92f7),
	.w7(32'hbb32a580),
	.w8(32'h3996ec7f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3e346),
	.w1(32'hbbe05d20),
	.w2(32'hbc2f72a4),
	.w3(32'hba152481),
	.w4(32'hbc2e81ca),
	.w5(32'hbaf045e6),
	.w6(32'hbc0c1926),
	.w7(32'hbc2317a3),
	.w8(32'h3b8042bd),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc134aab),
	.w1(32'h37531404),
	.w2(32'h3bc1f3a0),
	.w3(32'hb90e2d11),
	.w4(32'hbc1b3a8d),
	.w5(32'h3b7278f9),
	.w6(32'h3bfa8fe5),
	.w7(32'hb982ac18),
	.w8(32'hbb81833a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde4d01),
	.w1(32'hbb89d678),
	.w2(32'hbb0cdd30),
	.w3(32'h3bed732b),
	.w4(32'hbaecd11b),
	.w5(32'hbc38287b),
	.w6(32'h38449d5b),
	.w7(32'hbb9b1e4c),
	.w8(32'hbb7a289f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb905268),
	.w1(32'h3c186b88),
	.w2(32'h38eefb42),
	.w3(32'hbbc316d3),
	.w4(32'h3aca98a8),
	.w5(32'h3cb61c3f),
	.w6(32'hbbf224c8),
	.w7(32'hbb80efb3),
	.w8(32'h3c3b10e5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a74d0),
	.w1(32'hb9190fdc),
	.w2(32'hbaf05357),
	.w3(32'h3cab11a7),
	.w4(32'h3c7832bc),
	.w5(32'h3a3ec874),
	.w6(32'h3c993ec9),
	.w7(32'h3c3039f6),
	.w8(32'hbc15f7e7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2b522),
	.w1(32'hba5742dd),
	.w2(32'h3bd601bf),
	.w3(32'h3be2a124),
	.w4(32'h3c07f3a2),
	.w5(32'h3beb1fdd),
	.w6(32'hbb265a48),
	.w7(32'hbc007497),
	.w8(32'h3bd4466d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29d9c8),
	.w1(32'hbb55f120),
	.w2(32'h3bbe8c78),
	.w3(32'hbc1d51de),
	.w4(32'hbb320cbb),
	.w5(32'h3b1b47fc),
	.w6(32'hbbd8d763),
	.w7(32'h3bb7fc3d),
	.w8(32'h3c4847f6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba835d3f),
	.w1(32'hbbf9146d),
	.w2(32'h3b64ff07),
	.w3(32'hbb49247e),
	.w4(32'hbc2a5f9c),
	.w5(32'h3a8d0da0),
	.w6(32'hb9a1068b),
	.w7(32'hbbeb28f8),
	.w8(32'hbbbcd9c1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcef7162),
	.w1(32'hbcda372f),
	.w2(32'hbc5304b8),
	.w3(32'hbcb49fcc),
	.w4(32'hbcc0f78e),
	.w5(32'hbc27562f),
	.w6(32'hbcd7b074),
	.w7(32'hbca75706),
	.w8(32'hbbf55e23),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02ed96),
	.w1(32'h3c882b06),
	.w2(32'h3ba4dbd3),
	.w3(32'h3c2dab33),
	.w4(32'h3b0f44c3),
	.w5(32'h3c5c8951),
	.w6(32'h3c775ea8),
	.w7(32'h3baa188c),
	.w8(32'hbc519182),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a0a9),
	.w1(32'hbc1bf096),
	.w2(32'h3bb7c821),
	.w3(32'hbad31c47),
	.w4(32'hbaa6349a),
	.w5(32'h3ae609d8),
	.w6(32'h3bce5d0a),
	.w7(32'h3abe7bf8),
	.w8(32'h3bba6b1c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9a5a4),
	.w1(32'hb9a8e72c),
	.w2(32'hbc005f43),
	.w3(32'h39282a67),
	.w4(32'hbacaa9e6),
	.w5(32'hbc841ddb),
	.w6(32'hbb9e3089),
	.w7(32'hbb99a06b),
	.w8(32'hba023716),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383efc3f),
	.w1(32'h3b6a982b),
	.w2(32'h3c1e4368),
	.w3(32'hbbb9cac8),
	.w4(32'h3a029ec2),
	.w5(32'hb9e16969),
	.w6(32'h3b72ba9b),
	.w7(32'h385e1a85),
	.w8(32'h3bf91c87),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0872b5),
	.w1(32'h3a715e49),
	.w2(32'hbbecfd52),
	.w3(32'h3bd14d57),
	.w4(32'hbbd55820),
	.w5(32'hbbaa0fce),
	.w6(32'h3a1261fb),
	.w7(32'hbaf292be),
	.w8(32'h3afb9416),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72407f),
	.w1(32'hbb1b83d4),
	.w2(32'h3b367910),
	.w3(32'hbbd32371),
	.w4(32'h3b7dfe24),
	.w5(32'h39fbf300),
	.w6(32'hbb6deac3),
	.w7(32'h3be7bb71),
	.w8(32'h3b6a8037),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384764b9),
	.w1(32'hbb2d8ee7),
	.w2(32'hb9163d5e),
	.w3(32'h3ab8469f),
	.w4(32'h3a83c445),
	.w5(32'h3b36b11e),
	.w6(32'h3ae4de4c),
	.w7(32'h3b0a240b),
	.w8(32'h3a8520a0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdabd6d),
	.w1(32'hbaf19809),
	.w2(32'h3c88bd54),
	.w3(32'hbb82db90),
	.w4(32'hbbf7423c),
	.w5(32'h3bbc15d2),
	.w6(32'hbb88b598),
	.w7(32'hbc35f92b),
	.w8(32'hbada40e2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dd3c6),
	.w1(32'hba146460),
	.w2(32'hbacf1e86),
	.w3(32'hbad1f156),
	.w4(32'hbb1df856),
	.w5(32'hbab22796),
	.w6(32'hbb24e0a9),
	.w7(32'hbadd7f1c),
	.w8(32'hbb206085),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40f025),
	.w1(32'hbc4eed0c),
	.w2(32'h3bd6b91e),
	.w3(32'hbc2dbec4),
	.w4(32'hbc2fe7bf),
	.w5(32'h3c081032),
	.w6(32'hbbbd1edc),
	.w7(32'hbb671195),
	.w8(32'h3ac12ce2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb9954),
	.w1(32'hba0575b1),
	.w2(32'hbc0f9c89),
	.w3(32'h3b9dfcec),
	.w4(32'hbb071164),
	.w5(32'hbb9d9568),
	.w6(32'hbc1dcb25),
	.w7(32'hbc76c828),
	.w8(32'hbae4e941),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd81a9e),
	.w1(32'hbc0c97e8),
	.w2(32'h3b82a157),
	.w3(32'hbbc70631),
	.w4(32'hbc1d42e8),
	.w5(32'h3b90a750),
	.w6(32'hbb2b51ad),
	.w7(32'hbbb2aabb),
	.w8(32'h3bbd0292),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad96950),
	.w1(32'hbb488daa),
	.w2(32'hbc056baa),
	.w3(32'h3bbc7734),
	.w4(32'hba73ffa9),
	.w5(32'hbc0c2252),
	.w6(32'h3b5562f7),
	.w7(32'h3ba6d205),
	.w8(32'hbae3f075),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf2bae),
	.w1(32'hbbb6640e),
	.w2(32'h3ae4a79e),
	.w3(32'hba4eef2d),
	.w4(32'hbba01ac5),
	.w5(32'hbb5a8cba),
	.w6(32'h3b993e62),
	.w7(32'hbbcc611c),
	.w8(32'h3b23f1f7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000778),
	.w1(32'hbb2c5c72),
	.w2(32'hbadf891a),
	.w3(32'hbc598438),
	.w4(32'hbc5b60d0),
	.w5(32'hbbef3626),
	.w6(32'hbbbbe1b3),
	.w7(32'hbc03501d),
	.w8(32'hbbce41c4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b97d4),
	.w1(32'hbb36eace),
	.w2(32'h3c44bf61),
	.w3(32'hbafdaa98),
	.w4(32'hbc603856),
	.w5(32'h3c19d9be),
	.w6(32'hbb91fa65),
	.w7(32'hbca91492),
	.w8(32'h3b92bf04),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac67f4),
	.w1(32'hb9ac2ddf),
	.w2(32'h3b9398c6),
	.w3(32'h3b94c279),
	.w4(32'h3a9e94bb),
	.w5(32'h3bc4ad3f),
	.w6(32'h3c2855fe),
	.w7(32'h3b880dc6),
	.w8(32'h3b2aed34),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcdbbf),
	.w1(32'hba9c9976),
	.w2(32'h38ce6a1c),
	.w3(32'h3bf51856),
	.w4(32'h3c0d229c),
	.w5(32'h3bda99ab),
	.w6(32'hbb290367),
	.w7(32'hba18e8ad),
	.w8(32'h3b3f9b19),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18260f),
	.w1(32'h3bc05e67),
	.w2(32'h3be452ec),
	.w3(32'h3c1fd6df),
	.w4(32'hba5907a2),
	.w5(32'h3bbb7b4b),
	.w6(32'h3c80e20f),
	.w7(32'hbb393c41),
	.w8(32'h3a8f2ffd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b0d5c),
	.w1(32'hbbb4d04c),
	.w2(32'h3bba2a6c),
	.w3(32'hbb74df92),
	.w4(32'hbc1d0ac3),
	.w5(32'h3c2140b3),
	.w6(32'hbb91b20b),
	.w7(32'hbb438e7b),
	.w8(32'h3b698344),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a546016),
	.w1(32'hbbda3a89),
	.w2(32'hb98bedcd),
	.w3(32'h3bbef4b8),
	.w4(32'hbb79bf34),
	.w5(32'hbaed1ed7),
	.w6(32'hbb8e26bb),
	.w7(32'hbc385a7d),
	.w8(32'h38ae1917),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9478a66),
	.w1(32'hba577cf8),
	.w2(32'hbb64b31b),
	.w3(32'hbb44ee42),
	.w4(32'hbb29fd47),
	.w5(32'hbbbd92bb),
	.w6(32'hbb44fc8b),
	.w7(32'hbb274daa),
	.w8(32'hbbefdd21),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b6c78),
	.w1(32'hbb98e99f),
	.w2(32'hbb1cf09b),
	.w3(32'hbc821440),
	.w4(32'hbbcff706),
	.w5(32'hbc4fe96d),
	.w6(32'hbc317fe4),
	.w7(32'hb9f31a6b),
	.w8(32'hbba66c6e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc147437),
	.w1(32'hbb8dcb67),
	.w2(32'h3ca6c9cb),
	.w3(32'hbc97e751),
	.w4(32'h39f7156e),
	.w5(32'h3cc7100a),
	.w6(32'hbbe6c736),
	.w7(32'h3b154940),
	.w8(32'h3ca22eb0),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb478dda),
	.w1(32'hbb6b0843),
	.w2(32'hbc02d1d3),
	.w3(32'hbbea21aa),
	.w4(32'h3ba7e8b4),
	.w5(32'h3ba138b8),
	.w6(32'hbacafebc),
	.w7(32'hb8a62abc),
	.w8(32'h3c24f2a8),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907afc8),
	.w1(32'h3af2200a),
	.w2(32'h3b32ba34),
	.w3(32'hbb475e76),
	.w4(32'h3a272ea5),
	.w5(32'hbb3d32b0),
	.w6(32'h3b756846),
	.w7(32'hbaf3e649),
	.w8(32'hba78ef11),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1cc657),
	.w1(32'hbc2b97c7),
	.w2(32'hbb027569),
	.w3(32'hbc794126),
	.w4(32'hbb0962be),
	.w5(32'h3b0eb4ca),
	.w6(32'h3b88efbb),
	.w7(32'h3ba0e2e6),
	.w8(32'hbbc876e5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a7cb),
	.w1(32'hbb692d7b),
	.w2(32'hba3ea8e7),
	.w3(32'hbb52cd10),
	.w4(32'hbbb4b409),
	.w5(32'h3bca2f36),
	.w6(32'hbb8d043e),
	.w7(32'hbb972d3e),
	.w8(32'hbb9bd2d7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1734bf),
	.w1(32'hbb0c74f7),
	.w2(32'h3b181b88),
	.w3(32'hbb38ae67),
	.w4(32'h3a8e8576),
	.w5(32'h3c0521c6),
	.w6(32'hba2d0101),
	.w7(32'h3baf33fe),
	.w8(32'h3bba9cbb),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2e90e),
	.w1(32'hbc864307),
	.w2(32'h3c6ee60a),
	.w3(32'hbba38cda),
	.w4(32'h3baaeba5),
	.w5(32'h3ca14b39),
	.w6(32'hbc0397d7),
	.w7(32'hb9fcd067),
	.w8(32'h3d0c8d6d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27ebe6),
	.w1(32'hbc96eeec),
	.w2(32'hbc0db0da),
	.w3(32'h3bd24599),
	.w4(32'hbb184cbd),
	.w5(32'hbbc92b58),
	.w6(32'h3c2114d4),
	.w7(32'h3c25063c),
	.w8(32'h3b0dfc7c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd452a7),
	.w1(32'h3b98bc95),
	.w2(32'hbbb3db82),
	.w3(32'h3b9a34e4),
	.w4(32'h3c8bda3f),
	.w5(32'hbabf73a1),
	.w6(32'h3c159d14),
	.w7(32'h3cb2b0f0),
	.w8(32'h3bef4a8c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fbcd1),
	.w1(32'h3b574a51),
	.w2(32'h3bf59239),
	.w3(32'h3bbb0550),
	.w4(32'hbb0fd46c),
	.w5(32'h3b9fff66),
	.w6(32'h3be3c156),
	.w7(32'hbba6f541),
	.w8(32'hbb678039),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bf4a3),
	.w1(32'h3c072776),
	.w2(32'h3c9616e0),
	.w3(32'h3b849e41),
	.w4(32'hbb8c83ad),
	.w5(32'h3c1fd6d1),
	.w6(32'h3b8c2624),
	.w7(32'hbbd4a2a8),
	.w8(32'h3ba1faae),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b318032),
	.w1(32'h3a496452),
	.w2(32'h3b784a0a),
	.w3(32'h3bb66cb6),
	.w4(32'h3a513b0f),
	.w5(32'h3c043e52),
	.w6(32'hbba990d6),
	.w7(32'h3b2582d2),
	.w8(32'h3b855bc4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad09192),
	.w1(32'h3b59b572),
	.w2(32'h3badc8d4),
	.w3(32'h3c61f3a6),
	.w4(32'h3c2986e2),
	.w5(32'h3b024d34),
	.w6(32'h3c748487),
	.w7(32'h3bbbf119),
	.w8(32'h3b02268b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb2768),
	.w1(32'h3bfc5597),
	.w2(32'h3c2bab1a),
	.w3(32'hbc14ae2f),
	.w4(32'h3b4da91a),
	.w5(32'h3bce700f),
	.w6(32'hbbc68fc6),
	.w7(32'h3be7b74c),
	.w8(32'h3c7b3719),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6913e3),
	.w1(32'h3b8dba53),
	.w2(32'hbbc859b0),
	.w3(32'h3b84be8e),
	.w4(32'h3ab8e51c),
	.w5(32'hba8db996),
	.w6(32'hb9c39295),
	.w7(32'hbc153878),
	.w8(32'h3c0e6f05),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87b9bcd),
	.w1(32'h3b0977c8),
	.w2(32'h3c87458c),
	.w3(32'h3c2ae7a3),
	.w4(32'h3aeb5a96),
	.w5(32'h3c696e78),
	.w6(32'h3bc43bf0),
	.w7(32'hbad8249d),
	.w8(32'h3c258c54),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d70eb),
	.w1(32'h3c59c326),
	.w2(32'hbb2ad12b),
	.w3(32'h3cab4043),
	.w4(32'h3c94e440),
	.w5(32'h3b17e2a2),
	.w6(32'h3c804c21),
	.w7(32'h3c54566a),
	.w8(32'hbac8f162),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe0c33),
	.w1(32'h3b0471f5),
	.w2(32'h3be579ec),
	.w3(32'h3c20c8a6),
	.w4(32'h3a564bea),
	.w5(32'h3bee107e),
	.w6(32'h3b6d445d),
	.w7(32'h3b753657),
	.w8(32'h3ba58443),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99ecd0),
	.w1(32'hbb7f8e18),
	.w2(32'hbba32949),
	.w3(32'h3c2432c7),
	.w4(32'hbb134d64),
	.w5(32'h3a9eafb2),
	.w6(32'h3baf74a6),
	.w7(32'hba595561),
	.w8(32'h3bcee4cb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdabeeb),
	.w1(32'hbc975ed4),
	.w2(32'h3bad0ab9),
	.w3(32'hbc61b910),
	.w4(32'h3a8d9a82),
	.w5(32'h3ca122ec),
	.w6(32'hbc4ce6c2),
	.w7(32'h3bc78953),
	.w8(32'h3ceba981),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba75a67),
	.w1(32'hb9ebe555),
	.w2(32'h39b635b6),
	.w3(32'h3c45dfc8),
	.w4(32'h3c490ddd),
	.w5(32'h3c317ce3),
	.w6(32'h3c06b7e1),
	.w7(32'h3b4902eb),
	.w8(32'h3b2200e7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36ee96),
	.w1(32'h3baa7816),
	.w2(32'hbb6359ca),
	.w3(32'h3c6d22e2),
	.w4(32'hbb4985a8),
	.w5(32'hb9e7d080),
	.w6(32'h3bf31ed2),
	.w7(32'hbb94d765),
	.w8(32'h3b71a173),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f388c),
	.w1(32'hbc05cf2a),
	.w2(32'hbbb03923),
	.w3(32'hbc617650),
	.w4(32'hbbd32b38),
	.w5(32'hbbc9129f),
	.w6(32'hbc107ff2),
	.w7(32'hbb42ce0c),
	.w8(32'h3a7ea5b3),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe478e9),
	.w1(32'hbb80fb6a),
	.w2(32'h3c275bcc),
	.w3(32'hbc30ea39),
	.w4(32'hbbb5f5cf),
	.w5(32'h3b140f4e),
	.w6(32'hbc348409),
	.w7(32'hbc2b7231),
	.w8(32'hbb461c44),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0157b1),
	.w1(32'h3b3cf3fa),
	.w2(32'h3ab8487f),
	.w3(32'hbb602951),
	.w4(32'hbbd22f67),
	.w5(32'h3b962e37),
	.w6(32'hbc292111),
	.w7(32'hbc6bc7ef),
	.w8(32'h3bc3b9c8),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f94a2),
	.w1(32'hbb9a90ed),
	.w2(32'hbc1000de),
	.w3(32'hbb6be8e1),
	.w4(32'h3ad7acdf),
	.w5(32'hbb9bcc52),
	.w6(32'h3bad6333),
	.w7(32'hbb69aa02),
	.w8(32'hbb848b31),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eb1d5e),
	.w1(32'h3a5a7756),
	.w2(32'h3bf9e772),
	.w3(32'h3b589e36),
	.w4(32'h3bcff975),
	.w5(32'hba4fc5c4),
	.w6(32'hba25ce4b),
	.w7(32'hb9ed6d1b),
	.w8(32'h3c096d30),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beac154),
	.w1(32'h3c337100),
	.w2(32'hbbf5e23f),
	.w3(32'h3bfa9cb9),
	.w4(32'h3b099f60),
	.w5(32'h3b8bb31d),
	.w6(32'h3b359cad),
	.w7(32'h3acede9d),
	.w8(32'h3b1d0cb4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc010446),
	.w1(32'hbc255872),
	.w2(32'hb94dea90),
	.w3(32'hbb94711d),
	.w4(32'hbc75e5b5),
	.w5(32'h3aa6f53b),
	.w6(32'h399577f2),
	.w7(32'hbc118ec3),
	.w8(32'hbaa30ef4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76be4dd),
	.w1(32'h3a23dcf4),
	.w2(32'h3babaf9b),
	.w3(32'hb91781fb),
	.w4(32'hba056511),
	.w5(32'h3aab688a),
	.w6(32'h3a868506),
	.w7(32'h3be32768),
	.w8(32'h3c21955f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1444f5),
	.w1(32'hbbcf42cb),
	.w2(32'h3bb75d0d),
	.w3(32'hbb00f445),
	.w4(32'hbc3b1285),
	.w5(32'h3bb988d1),
	.w6(32'h3b0dfa68),
	.w7(32'hbb8ee0f8),
	.w8(32'h3c295cf4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c294bca),
	.w1(32'h3bdd36ed),
	.w2(32'hbb57914b),
	.w3(32'h3c1c699c),
	.w4(32'h3bac49f3),
	.w5(32'hbc232aae),
	.w6(32'h3c1d2c93),
	.w7(32'h3b371440),
	.w8(32'hbc133d2b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aa7be),
	.w1(32'hbb3ac8a8),
	.w2(32'hbbac050d),
	.w3(32'hbc529e8e),
	.w4(32'hbc375b0d),
	.w5(32'hbb3eefae),
	.w6(32'hbc540363),
	.w7(32'hbc084268),
	.w8(32'hbb9ead95),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81ed48),
	.w1(32'hbc3039d2),
	.w2(32'hb959b334),
	.w3(32'hb9e93e8e),
	.w4(32'hbbb13732),
	.w5(32'hbb940587),
	.w6(32'hbb4662cc),
	.w7(32'hbbdbd933),
	.w8(32'hbb9b03a3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba869823),
	.w1(32'hbabf67ae),
	.w2(32'hbb1ebc8d),
	.w3(32'hbc13f7c7),
	.w4(32'hbc14131f),
	.w5(32'h3bae248f),
	.w6(32'hbc294c18),
	.w7(32'hbc349691),
	.w8(32'hba6f93c8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08e5e3),
	.w1(32'hbc512223),
	.w2(32'h3bd23fc9),
	.w3(32'h3b914220),
	.w4(32'hbba62f76),
	.w5(32'hbbfeb774),
	.w6(32'hbabd35cf),
	.w7(32'hba6fe911),
	.w8(32'hbbd28497),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0976),
	.w1(32'hbb272453),
	.w2(32'h3ba63c40),
	.w3(32'hbaefa869),
	.w4(32'hbbd1c86c),
	.w5(32'hba685abe),
	.w6(32'h3953e06c),
	.w7(32'hbb06eb7a),
	.w8(32'h3a9eb579),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9415c7b),
	.w1(32'hbb6c5e90),
	.w2(32'h39b85517),
	.w3(32'hbb72ffd8),
	.w4(32'hbbbeb205),
	.w5(32'h3a12e770),
	.w6(32'hbbb2b93a),
	.w7(32'hbc24a34b),
	.w8(32'h396af907),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6066c9),
	.w1(32'hbb672cf3),
	.w2(32'hbb701c6c),
	.w3(32'hba9dba5c),
	.w4(32'hbbc1072e),
	.w5(32'hbbcec8ca),
	.w6(32'hba020351),
	.w7(32'hbbfafe69),
	.w8(32'hbbb6a817),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cd456),
	.w1(32'hbb9152bb),
	.w2(32'h3b6ca009),
	.w3(32'hbb847118),
	.w4(32'hbbe56870),
	.w5(32'hba13728c),
	.w6(32'hbbfa39a8),
	.w7(32'hbc064621),
	.w8(32'h3c0f5a4a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf1ff2),
	.w1(32'hbb121082),
	.w2(32'hbc2c9406),
	.w3(32'hbbf09d52),
	.w4(32'hbb04344c),
	.w5(32'hbc66aea7),
	.w6(32'h3bfe86b1),
	.w7(32'h3bda4535),
	.w8(32'hbc1025dc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42fb6c),
	.w1(32'hbbcc3edf),
	.w2(32'hbc2d3cbf),
	.w3(32'hbc92ecb0),
	.w4(32'hbc36211c),
	.w5(32'h3af3a19c),
	.w6(32'hbc48d176),
	.w7(32'hbbfd17c1),
	.w8(32'hbacb1bc5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39176c),
	.w1(32'hbc7bc0f0),
	.w2(32'hbc8d87c0),
	.w3(32'h3bcee94a),
	.w4(32'hbc3ec808),
	.w5(32'hbca130c9),
	.w6(32'h3c8b749a),
	.w7(32'h3be07eca),
	.w8(32'hbccec457),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fcefa),
	.w1(32'h3b95e975),
	.w2(32'hba159804),
	.w3(32'hbad4ed7d),
	.w4(32'h3b558293),
	.w5(32'h3a76c775),
	.w6(32'hbbdf4917),
	.w7(32'h3b908bf8),
	.w8(32'h3b394b83),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf8dc0),
	.w1(32'h3ab06c7d),
	.w2(32'h3c8a64ad),
	.w3(32'h3bfcb995),
	.w4(32'h3b8d1d91),
	.w5(32'h3c0078ec),
	.w6(32'h3be2dbfa),
	.w7(32'h3c084f7d),
	.w8(32'h3a32d50b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule