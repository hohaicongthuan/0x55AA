module layer_10_featuremap_115(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4cd0edf),
	.w1(32'hb48716bc),
	.w2(32'h36ba06c4),
	.w3(32'h3666c107),
	.w4(32'hb6cc4eb2),
	.w5(32'h36725d56),
	.w6(32'h3684e866),
	.w7(32'h36d47de4),
	.w8(32'h36fd6b9f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ed390),
	.w1(32'h3986088b),
	.w2(32'hb80535b0),
	.w3(32'h39641d65),
	.w4(32'h3a07571c),
	.w5(32'h37b8fa38),
	.w6(32'h393176cb),
	.w7(32'h3a294ddd),
	.w8(32'h392ca6da),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69f40c6),
	.w1(32'hb6abf4ed),
	.w2(32'hb640bfef),
	.w3(32'hb698649b),
	.w4(32'hb43ba9bb),
	.w5(32'h36483548),
	.w6(32'hb6cd2692),
	.w7(32'hb5d54c91),
	.w8(32'hb68457a4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87931e8),
	.w1(32'hb9f70305),
	.w2(32'hb9e2765d),
	.w3(32'h3982803a),
	.w4(32'h39173770),
	.w5(32'hb799d3b3),
	.w6(32'h395121e4),
	.w7(32'h39484ade),
	.w8(32'hb86f4ed5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb784b327),
	.w1(32'hb6b86da6),
	.w2(32'hb738b3fa),
	.w3(32'hb76ce8d8),
	.w4(32'hb717f343),
	.w5(32'hb755c0c9),
	.w6(32'hb71f6122),
	.w7(32'hb7038818),
	.w8(32'hb6f41bcd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb570b7de),
	.w1(32'h3563dfbf),
	.w2(32'hb61cb975),
	.w3(32'hb6d3a79b),
	.w4(32'h3572e815),
	.w5(32'h358fc6c1),
	.w6(32'h36fa4dbb),
	.w7(32'h369ad6db),
	.w8(32'h35feca30),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1001b2),
	.w1(32'hba0debca),
	.w2(32'h38d88683),
	.w3(32'h39eab04c),
	.w4(32'h39f11550),
	.w5(32'h3ab35a39),
	.w6(32'h3a5fc9fc),
	.w7(32'hba661bcc),
	.w8(32'h39308f6c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f5a176),
	.w1(32'hbb0d3f64),
	.w2(32'h3a9bd8d1),
	.w3(32'h3b03aca5),
	.w4(32'h3b72999f),
	.w5(32'h3aebf02c),
	.w6(32'hbaa0ce77),
	.w7(32'h3aba2152),
	.w8(32'hb775c9a9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3851f3e5),
	.w1(32'hb7de9be4),
	.w2(32'h390b0181),
	.w3(32'h3656b30e),
	.w4(32'hb82b0ecd),
	.w5(32'h38b6a751),
	.w6(32'h3715e592),
	.w7(32'hb82eb6ea),
	.w8(32'h3626f620),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaa746),
	.w1(32'hba4486a8),
	.w2(32'h3a611f83),
	.w3(32'hba2fac9f),
	.w4(32'h38de9b2b),
	.w5(32'hb8710fb0),
	.w6(32'h3a4733eb),
	.w7(32'h39acada4),
	.w8(32'h3760365a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88dfa7a),
	.w1(32'hb893bd1f),
	.w2(32'hb94a577c),
	.w3(32'h36decd8f),
	.w4(32'hb9006a64),
	.w5(32'hb95bc7c7),
	.w6(32'h3808ca53),
	.w7(32'hb7e5acd9),
	.w8(32'hb90e7edc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d736e),
	.w1(32'hbb7a7098),
	.w2(32'hbb10677b),
	.w3(32'hbac21d24),
	.w4(32'hbab2c7e3),
	.w5(32'hbac68f90),
	.w6(32'h3a1542c6),
	.w7(32'hba661bc3),
	.w8(32'hb98eaa5b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb177b06),
	.w1(32'hba23367f),
	.w2(32'h3a426158),
	.w3(32'hba42fb4e),
	.w4(32'hb8ceb786),
	.w5(32'h389691c0),
	.w6(32'h395b0973),
	.w7(32'hb972d4c6),
	.w8(32'h391adc32),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3bd85),
	.w1(32'hba1c7ba6),
	.w2(32'h39fe1b57),
	.w3(32'hba3ebe62),
	.w4(32'h3935b32f),
	.w5(32'h3aa7d250),
	.w6(32'hba37489e),
	.w7(32'h3985dcbe),
	.w8(32'h3a7201a6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2581db),
	.w1(32'h3a20dd78),
	.w2(32'h3955fc2f),
	.w3(32'hb8872067),
	.w4(32'hb85681fb),
	.w5(32'hb9e16f80),
	.w6(32'hb68bfbca),
	.w7(32'h395b5913),
	.w8(32'hb90b23ce),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc50be),
	.w1(32'h3998b8dd),
	.w2(32'h3a6b54f0),
	.w3(32'hba31e747),
	.w4(32'h3a81bfbc),
	.w5(32'h3afa9841),
	.w6(32'h3a899b31),
	.w7(32'h3b0b01cb),
	.w8(32'h3acaa917),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce11b2),
	.w1(32'hb8a67c35),
	.w2(32'hb8413c8a),
	.w3(32'hb904d9c7),
	.w4(32'hb94a604f),
	.w5(32'hb8be4160),
	.w6(32'hb7bfab0f),
	.w7(32'hb9173772),
	.w8(32'hb8c8de26),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e82c),
	.w1(32'hb9b8d538),
	.w2(32'h3a7ef94a),
	.w3(32'h3a74e0c9),
	.w4(32'h3a046a45),
	.w5(32'h3a983124),
	.w6(32'h3af18323),
	.w7(32'h3aab0199),
	.w8(32'h3afbb510),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede648),
	.w1(32'hb9809c5d),
	.w2(32'h39c7c9cc),
	.w3(32'h38fa6334),
	.w4(32'h394e84a1),
	.w5(32'h39831cfa),
	.w6(32'h3a3da0c3),
	.w7(32'h39508a1b),
	.w8(32'h3a00324c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37acf180),
	.w1(32'hb7f2b2ff),
	.w2(32'hb7a85f1c),
	.w3(32'hb6ee77e7),
	.w4(32'hb81504bf),
	.w5(32'hb7ecb8bd),
	.w6(32'hb6604cd7),
	.w7(32'hb77caa96),
	.w8(32'hb7f70bfb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb800aaf5),
	.w1(32'hb7d4bd4d),
	.w2(32'h372347b6),
	.w3(32'hb749f68e),
	.w4(32'hb6db6b8c),
	.w5(32'h378213c5),
	.w6(32'hb7b49953),
	.w7(32'h3707df5f),
	.w8(32'h372a9bc1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9914b),
	.w1(32'h398bb87d),
	.w2(32'hb921cc70),
	.w3(32'hb56c3b8c),
	.w4(32'h381ffcdd),
	.w5(32'hb8c97dd6),
	.w6(32'h36f16267),
	.w7(32'h3935f287),
	.w8(32'hb897b9c8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31585c),
	.w1(32'h3b167534),
	.w2(32'h3b2b5c5e),
	.w3(32'hbaf08d5d),
	.w4(32'h3b2e8444),
	.w5(32'h3b11f503),
	.w6(32'h3afd0537),
	.w7(32'h397db327),
	.w8(32'h3a5d8a54),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a031c15),
	.w1(32'h39cdb7bd),
	.w2(32'h3a45cc26),
	.w3(32'hb644006c),
	.w4(32'h37adf97b),
	.w5(32'h398f93f2),
	.w6(32'hb866322e),
	.w7(32'hb91cf779),
	.w8(32'hb8ed4a77),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b4814),
	.w1(32'h3a36f2ef),
	.w2(32'h391c72ad),
	.w3(32'hb99642c0),
	.w4(32'h3a06a7d6),
	.w5(32'hb986151f),
	.w6(32'hba74b66d),
	.w7(32'h3984c203),
	.w8(32'hb9a81198),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895cfab),
	.w1(32'hb81cfb87),
	.w2(32'hb82f0b42),
	.w3(32'h38ca2e7d),
	.w4(32'hb75f92d1),
	.w5(32'hb80074a6),
	.w6(32'h37804061),
	.w7(32'h3551a331),
	.w8(32'hb7624b56),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7388450),
	.w1(32'hb7636b3e),
	.w2(32'hb8109dc1),
	.w3(32'hb7b8ac42),
	.w4(32'hb7ab18f7),
	.w5(32'hb80eaec5),
	.w6(32'hb6f72b3c),
	.w7(32'h36aa7742),
	.w8(32'hb78552b2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68d5b7),
	.w1(32'h3af57b86),
	.w2(32'h3b0b72b4),
	.w3(32'hb9abab3f),
	.w4(32'h3aaf407e),
	.w5(32'h393819d0),
	.w6(32'hba01d85d),
	.w7(32'h39062548),
	.w8(32'h38e682c1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93eeab6),
	.w1(32'hb8e3e591),
	.w2(32'hb97160e9),
	.w3(32'hb928530b),
	.w4(32'hb9599114),
	.w5(32'hb9c8e967),
	.w6(32'hb963ff1a),
	.w7(32'hb99ad252),
	.w8(32'hb9c501e6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a7020),
	.w1(32'h3ab02841),
	.w2(32'h3a329335),
	.w3(32'hba982575),
	.w4(32'h3995b0ee),
	.w5(32'h39c947db),
	.w6(32'hbb21268f),
	.w7(32'h3958b75f),
	.w8(32'hb8951c58),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a2a816),
	.w1(32'hb73f82ac),
	.w2(32'hb79d9bba),
	.w3(32'hb6f3a5fb),
	.w4(32'hb76f1824),
	.w5(32'hb79fd496),
	.w6(32'hb5278a83),
	.w7(32'hb6d43cd9),
	.w8(32'hb6e07a9d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ccc697),
	.w1(32'hb78ff484),
	.w2(32'hb849e226),
	.w3(32'h384e5de4),
	.w4(32'hb764f058),
	.w5(32'hb8b4a637),
	.w6(32'h3826c65f),
	.w7(32'hb7a93660),
	.w8(32'hb88cab2a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba965a5a),
	.w1(32'hba1de4cd),
	.w2(32'hb88754a4),
	.w3(32'hb9f21860),
	.w4(32'hb90d805f),
	.w5(32'hb87996e2),
	.w6(32'h390aa676),
	.w7(32'h38e15903),
	.w8(32'h3990eae1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fa4aa),
	.w1(32'h399532a4),
	.w2(32'h39ce9b39),
	.w3(32'h39a19ca6),
	.w4(32'h3a21cfa2),
	.w5(32'h39d7aacf),
	.w6(32'hb8bd5358),
	.w7(32'h39fb6815),
	.w8(32'h39c7aa9e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82af51),
	.w1(32'hba49e5a1),
	.w2(32'hb99e3f62),
	.w3(32'hb8e5b836),
	.w4(32'h389e1b11),
	.w5(32'h35890d31),
	.w6(32'h38ead259),
	.w7(32'h388b7eba),
	.w8(32'h3945c6db),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa56ad4),
	.w1(32'hb955f595),
	.w2(32'h386a58b9),
	.w3(32'h39ac6c6d),
	.w4(32'h3a45aa34),
	.w5(32'h3a29238e),
	.w6(32'h3800b658),
	.w7(32'hb8fb6412),
	.w8(32'h3982af51),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0966b),
	.w1(32'hbb7837a0),
	.w2(32'hbaefe755),
	.w3(32'hbafdef07),
	.w4(32'h3a6a80a4),
	.w5(32'hbb8a0568),
	.w6(32'hba7717fa),
	.w7(32'h39709098),
	.w8(32'hbad8b49d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11eddf),
	.w1(32'h3b541776),
	.w2(32'h3a02f0d0),
	.w3(32'hba55143e),
	.w4(32'hb948b410),
	.w5(32'hbad5a768),
	.w6(32'hbabe1b49),
	.w7(32'hb8d6a8bb),
	.w8(32'hba9850c1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbc0f9),
	.w1(32'h3b68649d),
	.w2(32'h3b2bdac3),
	.w3(32'hbab96f50),
	.w4(32'h3860e52a),
	.w5(32'h3838b388),
	.w6(32'hba95a293),
	.w7(32'h3a1af626),
	.w8(32'hb979dd84),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c69565),
	.w1(32'h390b2a15),
	.w2(32'hb9b0da00),
	.w3(32'hb8374c95),
	.w4(32'hb88b435c),
	.w5(32'hb9ffda38),
	.w6(32'h37b87237),
	.w7(32'h39234cfd),
	.w8(32'hb8f77a47),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927500d),
	.w1(32'h38839690),
	.w2(32'h37ac7b3e),
	.w3(32'h3917a438),
	.w4(32'h38448c8f),
	.w5(32'h375038ab),
	.w6(32'h37de20db),
	.w7(32'hb727609c),
	.w8(32'hb814486d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c8b030),
	.w1(32'h36b0633a),
	.w2(32'hb7bbd98a),
	.w3(32'hb793b56a),
	.w4(32'hb821553d),
	.w5(32'hb81687e7),
	.w6(32'hb859d98c),
	.w7(32'hb78fec53),
	.w8(32'hb88f9af7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f303ef),
	.w1(32'hb7a7c4eb),
	.w2(32'hb952de35),
	.w3(32'h38da2589),
	.w4(32'h379f59c4),
	.w5(32'hb95754c6),
	.w6(32'h38d2bf09),
	.w7(32'hb8280f1a),
	.w8(32'hb96a52b3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa44995),
	.w1(32'h39a65bbc),
	.w2(32'h3b21ff31),
	.w3(32'hba1d48aa),
	.w4(32'hba1e6971),
	.w5(32'h3a046fa3),
	.w6(32'h3ac0732b),
	.w7(32'hb73c4703),
	.w8(32'h36c1ec56),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdeca4),
	.w1(32'h3a68aeee),
	.w2(32'h3a02bd52),
	.w3(32'hb96f6fc6),
	.w4(32'hb9d9ee1f),
	.w5(32'hb9db03c0),
	.w6(32'hb9e4a9f9),
	.w7(32'hb9c4e8a2),
	.w8(32'hba2c60c1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e2a97),
	.w1(32'h3aafa1ec),
	.w2(32'h3813ebd8),
	.w3(32'hb889bef5),
	.w4(32'h382aeb24),
	.w5(32'h3927d9a4),
	.w6(32'h392fc217),
	.w7(32'h380b9ef0),
	.w8(32'h38eac4e6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03f81e),
	.w1(32'h391af923),
	.w2(32'h39ebfc1b),
	.w3(32'hb9cb0551),
	.w4(32'hb79f8bc5),
	.w5(32'hb5bba894),
	.w6(32'hb9bae99e),
	.w7(32'h38e7bfe4),
	.w8(32'hb98f995a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cb19c),
	.w1(32'hbaf04437),
	.w2(32'hb8238387),
	.w3(32'hba874619),
	.w4(32'hb6d58b23),
	.w5(32'h39faa0e0),
	.w6(32'h3ad06701),
	.w7(32'h3a27f4dd),
	.w8(32'h3a8a825f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c84473),
	.w1(32'h38b9c104),
	.w2(32'h38c1ec23),
	.w3(32'hb854887f),
	.w4(32'hb84873de),
	.w5(32'h378f8eb7),
	.w6(32'hb80ea8c4),
	.w7(32'h37b47962),
	.w8(32'h35f53d18),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b87b0),
	.w1(32'h38ac8e7a),
	.w2(32'h397fe72d),
	.w3(32'hb7491c7d),
	.w4(32'h38fd2090),
	.w5(32'h398d0d53),
	.w6(32'hb90fdf34),
	.w7(32'hb8d4668f),
	.w8(32'hb7c22944),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87898df),
	.w1(32'hb88e10a2),
	.w2(32'h38be0fb8),
	.w3(32'hb934b464),
	.w4(32'hb893de4f),
	.w5(32'h38d0db30),
	.w6(32'hb987b364),
	.w7(32'hb96734b4),
	.w8(32'hb79f0cb1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c9d71),
	.w1(32'h3ac60cb1),
	.w2(32'h3a2bb3a9),
	.w3(32'h39eed780),
	.w4(32'h3a753ed3),
	.w5(32'h39a9daf2),
	.w6(32'h38db9215),
	.w7(32'hb992c576),
	.w8(32'hba024cf4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd5983),
	.w1(32'hb91dd296),
	.w2(32'h398d1645),
	.w3(32'h39563c60),
	.w4(32'h3a256b5b),
	.w5(32'h39c59f5b),
	.w6(32'h38a0f231),
	.w7(32'h39cafb14),
	.w8(32'h39dc04a9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8910e2),
	.w1(32'hbad6f696),
	.w2(32'h38a62753),
	.w3(32'hbac95d8e),
	.w4(32'hb92bcf9e),
	.w5(32'h39e33426),
	.w6(32'h3ae2837c),
	.w7(32'h3a9ca2c1),
	.w8(32'h3ad9410a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922cb7c),
	.w1(32'h39e96d6a),
	.w2(32'h39b619fd),
	.w3(32'h3a182614),
	.w4(32'h398874ec),
	.w5(32'h39b6324c),
	.w6(32'hb980797b),
	.w7(32'h38237cf1),
	.w8(32'h38cdee44),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de2625),
	.w1(32'h3888a19e),
	.w2(32'h37fda1c7),
	.w3(32'hb7c4a7fc),
	.w4(32'h37ca2390),
	.w5(32'hb8185184),
	.w6(32'hb8abe73d),
	.w7(32'hb68ac165),
	.w8(32'hb82dc6de),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378571e2),
	.w1(32'h356f35ad),
	.w2(32'h3660a7a9),
	.w3(32'hb504fb62),
	.w4(32'hb5abbe94),
	.w5(32'h35c41258),
	.w6(32'h3598648c),
	.w7(32'h374223d5),
	.w8(32'h37448537),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a9d522),
	.w1(32'h38be36b2),
	.w2(32'hb7bde565),
	.w3(32'h37c4bb85),
	.w4(32'hb90e4a55),
	.w5(32'hb8864dbd),
	.w6(32'hb7d3dd2c),
	.w7(32'hb858f096),
	.w8(32'h37081f88),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88da25a),
	.w1(32'hb89cb75c),
	.w2(32'hb9693582),
	.w3(32'hb90455ea),
	.w4(32'hb8e39445),
	.w5(32'hb92cfa5a),
	.w6(32'hb84ba38f),
	.w7(32'hb81cc6c0),
	.w8(32'hb822449b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3e359),
	.w1(32'hb97f92fa),
	.w2(32'hb925380d),
	.w3(32'h38e05947),
	.w4(32'h388eb489),
	.w5(32'h3817bbf9),
	.w6(32'h38d5fc38),
	.w7(32'h37ab5520),
	.w8(32'h38a21536),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7cd9),
	.w1(32'hb9889ba9),
	.w2(32'h3a15ee7c),
	.w3(32'h396a5e81),
	.w4(32'h39d2df5c),
	.w5(32'h3a1b34ec),
	.w6(32'h3a3a58f2),
	.w7(32'h39d39339),
	.w8(32'h3a2c3b00),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f012d),
	.w1(32'h3a951e66),
	.w2(32'h3aaf2d05),
	.w3(32'h3a36c863),
	.w4(32'h3a3967a5),
	.w5(32'h3a826919),
	.w6(32'hb7e92341),
	.w7(32'h3975d432),
	.w8(32'h39aa4734),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382bf2be),
	.w1(32'hb66a0eda),
	.w2(32'h37793a60),
	.w3(32'h3791835c),
	.w4(32'hb7b779a7),
	.w5(32'hb6b7ae7c),
	.w6(32'hb5fa65b2),
	.w7(32'hb7dd4130),
	.w8(32'hb85d209f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ccd62f),
	.w1(32'h367c722b),
	.w2(32'hb665f2a6),
	.w3(32'hb7be1c46),
	.w4(32'h365f96a9),
	.w5(32'hb6098e8f),
	.w6(32'h369f953e),
	.w7(32'h360e22ba),
	.w8(32'hb6f3f9ff),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e52cf7),
	.w1(32'hb7675329),
	.w2(32'hb84e2274),
	.w3(32'h341220ca),
	.w4(32'hb6c76525),
	.w5(32'hb857cf0a),
	.w6(32'h3722f153),
	.w7(32'hb7401136),
	.w8(32'hb7f70055),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6aac429),
	.w1(32'hb7708e98),
	.w2(32'hb7ed6ac3),
	.w3(32'h350a3d6a),
	.w4(32'hb69eef76),
	.w5(32'hb786da04),
	.w6(32'h3523a753),
	.w7(32'h3568a2be),
	.w8(32'hb6f364ae),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03cfd1),
	.w1(32'hbba27d79),
	.w2(32'hb8f3a645),
	.w3(32'hbb3e96b5),
	.w4(32'hba8cb084),
	.w5(32'hb92846d0),
	.w6(32'h3b05c466),
	.w7(32'h3b35f68a),
	.w8(32'h3b4d8c79),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b055a),
	.w1(32'hba9ffe33),
	.w2(32'hba09eaff),
	.w3(32'h3b0ada55),
	.w4(32'h3b1fd00d),
	.w5(32'h3b0f3388),
	.w6(32'hba705e34),
	.w7(32'h3a88ceac),
	.w8(32'h3b2e3a66),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47aeb2),
	.w1(32'h3a96ae4c),
	.w2(32'h3b032892),
	.w3(32'h3aaa44e9),
	.w4(32'h3a91fadb),
	.w5(32'h3ac96140),
	.w6(32'hb72a1e2c),
	.w7(32'h3a210a34),
	.w8(32'h3a6ab8df),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa6929),
	.w1(32'h3ad9df84),
	.w2(32'h3929bec4),
	.w3(32'hba756590),
	.w4(32'hb93de352),
	.w5(32'hbaa2241a),
	.w6(32'hba986e40),
	.w7(32'hb854134d),
	.w8(32'hba74777a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36030b7f),
	.w1(32'hb7aa2b3f),
	.w2(32'hb7a618a2),
	.w3(32'hb682b2da),
	.w4(32'hb74fefce),
	.w5(32'hb735dfc3),
	.w6(32'hb717d45e),
	.w7(32'hb67cd75e),
	.w8(32'hb6c897e1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5cc813f),
	.w1(32'hb55c55c6),
	.w2(32'hb790a26c),
	.w3(32'hb70de831),
	.w4(32'h363b77e1),
	.w5(32'hb6ff09c6),
	.w6(32'hb5b079fc),
	.w7(32'h36b17422),
	.w8(32'hb6f102f6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72c82c6),
	.w1(32'hb7269b05),
	.w2(32'hb8067fd0),
	.w3(32'hb39619f9),
	.w4(32'hb6fd93c3),
	.w5(32'hb782c964),
	.w6(32'h35b8ddf9),
	.w7(32'hb699b1a5),
	.w8(32'hb6bda665),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba342296),
	.w1(32'hba0005f9),
	.w2(32'hb8d8d214),
	.w3(32'h395c1cc6),
	.w4(32'hb857005b),
	.w5(32'h3692e27e),
	.w6(32'h39d3dea4),
	.w7(32'h39950356),
	.w8(32'h399ae049),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368dcbc9),
	.w1(32'h37bf1115),
	.w2(32'h376bc434),
	.w3(32'hb7b0bcd5),
	.w4(32'h36df98ce),
	.w5(32'h37707061),
	.w6(32'hb7bd545a),
	.w7(32'hb534073a),
	.w8(32'hb75e7f9e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03b869),
	.w1(32'hbaa15701),
	.w2(32'h39c74938),
	.w3(32'hbad09b64),
	.w4(32'h39b008d0),
	.w5(32'hba1101d1),
	.w6(32'h3a08a75d),
	.w7(32'h3a46ab48),
	.w8(32'h399772dc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ec2c0),
	.w1(32'hbaf75a1a),
	.w2(32'hb90632cc),
	.w3(32'h38c43998),
	.w4(32'h3abc69e6),
	.w5(32'h3a5d9ed4),
	.w6(32'h3a556cf7),
	.w7(32'h3afbf8da),
	.w8(32'h3ab5fbbc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90d50e),
	.w1(32'h3a3660f7),
	.w2(32'h395a42d4),
	.w3(32'hb9b56515),
	.w4(32'hb98fbbee),
	.w5(32'hba0378f6),
	.w6(32'hb9b57fbb),
	.w7(32'hb98cc911),
	.w8(32'hba358008),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba488a4e),
	.w1(32'hb9648649),
	.w2(32'h3a530294),
	.w3(32'hb9f554b1),
	.w4(32'h378ec3c6),
	.w5(32'h3a24b581),
	.w6(32'hb98a28ec),
	.w7(32'h39c6cee2),
	.w8(32'h3a2b29dc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f60bc),
	.w1(32'hbb449d97),
	.w2(32'hbaabb485),
	.w3(32'hbad945b0),
	.w4(32'h391c60f8),
	.w5(32'hba33f715),
	.w6(32'h3a4edef2),
	.w7(32'h3a62cf00),
	.w8(32'h3a59f2a4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e7cbd),
	.w1(32'h3a112e3a),
	.w2(32'h3a2f92e1),
	.w3(32'hb9c94c54),
	.w4(32'hb9a03405),
	.w5(32'hb87e8bc3),
	.w6(32'hba175eff),
	.w7(32'hb8bde2d6),
	.w8(32'hb9a692c2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc8e51),
	.w1(32'hba074e6d),
	.w2(32'h39682012),
	.w3(32'hb9fb1dc3),
	.w4(32'h36d3f004),
	.w5(32'h38bffd15),
	.w6(32'h398af434),
	.w7(32'h381c9cc7),
	.w8(32'h394fb2c7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6abe251),
	.w1(32'h3537948c),
	.w2(32'h363f52d2),
	.w3(32'h361bc3b8),
	.w4(32'h35aff47a),
	.w5(32'h370ebac6),
	.w6(32'hb6199b18),
	.w7(32'h3568ca87),
	.w8(32'hb5838c02),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369c8e9f),
	.w1(32'h3716e89c),
	.w2(32'h378e5223),
	.w3(32'h365cbc31),
	.w4(32'h374addd1),
	.w5(32'h37b362c3),
	.w6(32'h37422bd2),
	.w7(32'h374c291a),
	.w8(32'h377e2881),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67d3982),
	.w1(32'hb4de4133),
	.w2(32'h373a07ba),
	.w3(32'hb5dbb66d),
	.w4(32'hb7879038),
	.w5(32'hb5af2d1b),
	.w6(32'hb77e371e),
	.w7(32'hb6223097),
	.w8(32'hb6b3cf74),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e6fd5),
	.w1(32'h3982c75d),
	.w2(32'h38121d98),
	.w3(32'h370a93a1),
	.w4(32'h381d5213),
	.w5(32'hb7f4d054),
	.w6(32'hb883bd05),
	.w7(32'hb7548e61),
	.w8(32'hb78de0e1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb636f),
	.w1(32'h3921d1b5),
	.w2(32'hb5f52a92),
	.w3(32'h38879ce0),
	.w4(32'hb962eeed),
	.w5(32'hb9f21a74),
	.w6(32'hb74a1d4a),
	.w7(32'h394f38a8),
	.w8(32'hba03e3cf),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d5cf32),
	.w1(32'hb90cfe44),
	.w2(32'hb944bbcb),
	.w3(32'hb7c7f62a),
	.w4(32'hb8725eac),
	.w5(32'hb8e5478e),
	.w6(32'h33fd14b6),
	.w7(32'hb791e4a5),
	.w8(32'hb8549dc8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a29a7),
	.w1(32'h3903ede3),
	.w2(32'hba1a36ce),
	.w3(32'h3a3d7581),
	.w4(32'h3a403198),
	.w5(32'h384c1b5e),
	.w6(32'h3a36a1fa),
	.w7(32'h3aa2a0e7),
	.w8(32'h3a25efb8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21d2f4),
	.w1(32'hb8ac4832),
	.w2(32'h3a2919b4),
	.w3(32'hb9333e35),
	.w4(32'h3a950034),
	.w5(32'h3a079d92),
	.w6(32'h3a383acc),
	.w7(32'h3a9dbede),
	.w8(32'h3a9ccd1f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59ebe5),
	.w1(32'h3ad98d52),
	.w2(32'h3a6c39fc),
	.w3(32'hba2c72b9),
	.w4(32'h3945c919),
	.w5(32'hb9458cb0),
	.w6(32'hb949bb4f),
	.w7(32'hb8307630),
	.w8(32'hb9bf419d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1039f),
	.w1(32'hbb062adb),
	.w2(32'hb9df1002),
	.w3(32'hbb06a801),
	.w4(32'hbac98f6b),
	.w5(32'hba79e470),
	.w6(32'h3ae6ad47),
	.w7(32'h3a552d34),
	.w8(32'h39aba4c4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abec77a),
	.w1(32'h3abd0e66),
	.w2(32'h3a22404c),
	.w3(32'hb69688cf),
	.w4(32'h39a432d5),
	.w5(32'hb9fef8c6),
	.w6(32'hb9065fc9),
	.w7(32'hba4e6286),
	.w8(32'hba22827b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fe67e),
	.w1(32'hbaf4af00),
	.w2(32'h3a029530),
	.w3(32'hba8853f8),
	.w4(32'h392cbad1),
	.w5(32'h3a944082),
	.w6(32'hb9e37d77),
	.w7(32'h3ade62d1),
	.w8(32'h3af6e952),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac31fee),
	.w1(32'hb9b8c114),
	.w2(32'h39b1dbae),
	.w3(32'hb98f41a6),
	.w4(32'hb91192fb),
	.w5(32'h391addc1),
	.w6(32'hb9b7c6ae),
	.w7(32'h3a109493),
	.w8(32'h3a368267),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37817796),
	.w1(32'h3a9bc941),
	.w2(32'h39160216),
	.w3(32'hba100c41),
	.w4(32'h3993eb64),
	.w5(32'hb9c1549a),
	.w6(32'hba373e35),
	.w7(32'h3967c310),
	.w8(32'hb8a9b874),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9f684),
	.w1(32'hb8b9aada),
	.w2(32'h39269e14),
	.w3(32'hb9984889),
	.w4(32'h38ccc6f0),
	.w5(32'h3985ee79),
	.w6(32'hb9017ea3),
	.w7(32'hb7960925),
	.w8(32'hb8176127),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9ea83),
	.w1(32'hb9dff9cf),
	.w2(32'h3a7ca778),
	.w3(32'hb89a10c4),
	.w4(32'h39e8b0fb),
	.w5(32'h3a6e7aa1),
	.w6(32'h3a08bb37),
	.w7(32'h394a333a),
	.w8(32'h3a601ec2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4ea2),
	.w1(32'hbb2eec4a),
	.w2(32'hb940ed3d),
	.w3(32'hbb497707),
	.w4(32'hbac1d0c5),
	.w5(32'hbae113ae),
	.w6(32'h3a0010f8),
	.w7(32'hb999548e),
	.w8(32'hba90d3f1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390099ce),
	.w1(32'hba925120),
	.w2(32'hba62268c),
	.w3(32'hb9208c40),
	.w4(32'h3b247bd7),
	.w5(32'h39b9d2e8),
	.w6(32'hb9c903aa),
	.w7(32'hba7747af),
	.w8(32'h39cb5cc3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e1cbd),
	.w1(32'h3ac17ba9),
	.w2(32'hba0b5a9f),
	.w3(32'h36e21a4e),
	.w4(32'h391de8ae),
	.w5(32'hbac992a8),
	.w6(32'hb8d3a61d),
	.w7(32'h3982d914),
	.w8(32'hba825a6b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa03657),
	.w1(32'h3a671047),
	.w2(32'h39cc9835),
	.w3(32'h39ae8b93),
	.w4(32'h396a7f11),
	.w5(32'hb84a26cd),
	.w6(32'hb973fc7e),
	.w7(32'h3908399b),
	.w8(32'hb97b92db),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995055),
	.w1(32'hbb4d4183),
	.w2(32'hba93ffd2),
	.w3(32'hbaca75d2),
	.w4(32'hba8bdc5d),
	.w5(32'hbab76f7a),
	.w6(32'h3a203e00),
	.w7(32'hb96a1cc9),
	.w8(32'h38a247c0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ac84e),
	.w1(32'h3998ffd0),
	.w2(32'h39b4f11f),
	.w3(32'hb9d66f4c),
	.w4(32'h392c99f6),
	.w5(32'h3a0ae4cf),
	.w6(32'hb9ba7813),
	.w7(32'hb7570a60),
	.w8(32'h39952c09),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44be06),
	.w1(32'hbb92baae),
	.w2(32'h3a8abd50),
	.w3(32'hbb2971d8),
	.w4(32'h3a89080e),
	.w5(32'hba8530a6),
	.w6(32'h39cb27dc),
	.w7(32'h3aadfe13),
	.w8(32'hbac7a168),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991f444),
	.w1(32'hbb03c5a2),
	.w2(32'h3a80d19d),
	.w3(32'h3923ada1),
	.w4(32'hbac2df2e),
	.w5(32'hb8f6e23a),
	.w6(32'h398cfd32),
	.w7(32'hba7e546a),
	.w8(32'hba8821c9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a216ce),
	.w1(32'hb68b41fa),
	.w2(32'hb67ace8b),
	.w3(32'hb92c2e39),
	.w4(32'hb88a9ddc),
	.w5(32'hb805ad96),
	.w6(32'hb890ffc6),
	.w7(32'h36cf17d6),
	.w8(32'h3752225a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29b57b),
	.w1(32'h39daa7ed),
	.w2(32'hb8c5ecb5),
	.w3(32'hb986d1bc),
	.w4(32'h39cd2aa9),
	.w5(32'h388d689c),
	.w6(32'h39585f29),
	.w7(32'h39cf6f83),
	.w8(32'h38846114),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99a285),
	.w1(32'hba1b4af2),
	.w2(32'h3998f666),
	.w3(32'hba328395),
	.w4(32'hb9349741),
	.w5(32'h397eb24d),
	.w6(32'h38c9a3d7),
	.w7(32'h388a04b4),
	.w8(32'h3987afc7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a087852),
	.w1(32'h39c4b882),
	.w2(32'h39e0881c),
	.w3(32'hba38195d),
	.w4(32'hba11310e),
	.w5(32'hb9e96887),
	.w6(32'hba2bbcfe),
	.w7(32'hba234e82),
	.w8(32'hba6b072d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8084e1),
	.w1(32'h3ad08e36),
	.w2(32'h3a8a07ad),
	.w3(32'hba72e8ab),
	.w4(32'hb8a5cc19),
	.w5(32'hb99c3972),
	.w6(32'h39f444eb),
	.w7(32'h390b83be),
	.w8(32'hb9cc8c08),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a670aa6),
	.w1(32'h39da3d50),
	.w2(32'h38f342f7),
	.w3(32'h38588db5),
	.w4(32'h39cec0ac),
	.w5(32'hb8550a7e),
	.w6(32'hb969d7d3),
	.w7(32'h397d018d),
	.w8(32'h3911761b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d0ef),
	.w1(32'hbb0ff92b),
	.w2(32'hbb1952f7),
	.w3(32'h3ab66a3a),
	.w4(32'h3a847915),
	.w5(32'h3878f1ba),
	.w6(32'h3a52f128),
	.w7(32'h3a8c01f6),
	.w8(32'h392594c5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd2694),
	.w1(32'hb933ae91),
	.w2(32'h3a6c82cf),
	.w3(32'hb9e55730),
	.w4(32'h39ee86c4),
	.w5(32'h3ad1a7f8),
	.w6(32'h3a9c6cbf),
	.w7(32'h3abc0cf8),
	.w8(32'h3ac1c413),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a181854),
	.w1(32'h39e0adab),
	.w2(32'h39655692),
	.w3(32'hb72c38a7),
	.w4(32'hb9262c1c),
	.w5(32'hb7ca63a9),
	.w6(32'hb91428be),
	.w7(32'hb9828b05),
	.w8(32'hb990391d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3616c6c7),
	.w1(32'h36a04db7),
	.w2(32'h36451f88),
	.w3(32'h369146ba),
	.w4(32'h36c78584),
	.w5(32'h3653360b),
	.w6(32'h37a48672),
	.w7(32'h36e6325e),
	.w8(32'h379ce775),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39005cd8),
	.w1(32'h38d0a7fa),
	.w2(32'h38afc40a),
	.w3(32'h3874bbee),
	.w4(32'h3934d9cb),
	.w5(32'h394760a4),
	.w6(32'h38da6df5),
	.w7(32'h39ec26f7),
	.w8(32'h39aed5d4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35635594),
	.w1(32'h353ace32),
	.w2(32'hb67cdf02),
	.w3(32'h369430fd),
	.w4(32'h360af212),
	.w5(32'h3536f62d),
	.w6(32'h3588c496),
	.w7(32'hb5515292),
	.w8(32'hb566f7f4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f9d05a),
	.w1(32'h37937136),
	.w2(32'h37ffa11f),
	.w3(32'h369cde9d),
	.w4(32'hb6076d04),
	.w5(32'h370444ca),
	.w6(32'h36b42b33),
	.w7(32'hb79b8e31),
	.w8(32'h37320efd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41de8d),
	.w1(32'h3a2e38d1),
	.w2(32'h391b1876),
	.w3(32'hb88277fd),
	.w4(32'hb9679055),
	.w5(32'hb8a6eab0),
	.w6(32'hb89948ed),
	.w7(32'hb871d06a),
	.w8(32'hb927372d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7939254),
	.w1(32'hb8a82baa),
	.w2(32'hb8b2fe1a),
	.w3(32'h37abd53a),
	.w4(32'hb8c43afc),
	.w5(32'hb83b291e),
	.w6(32'h381e7c43),
	.w7(32'hb8535110),
	.w8(32'hb8481517),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d84a8),
	.w1(32'hba96de84),
	.w2(32'hb9ca6c7b),
	.w3(32'hba27a174),
	.w4(32'hb93bfd7f),
	.w5(32'hb9c11c5b),
	.w6(32'h3a3f5cf4),
	.w7(32'h39efa94c),
	.w8(32'h3965355a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2623b),
	.w1(32'h3aa7ebf3),
	.w2(32'hb7374ecb),
	.w3(32'hba2ae8ad),
	.w4(32'h39dc7ac5),
	.w5(32'hba1fdd97),
	.w6(32'hba3c82d5),
	.w7(32'h3a31ed3d),
	.w8(32'hb904d0eb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3737b6fd),
	.w1(32'h37135015),
	.w2(32'hb6450dc3),
	.w3(32'hb65d3f7c),
	.w4(32'h33b551d8),
	.w5(32'hb74fe44f),
	.w6(32'hb674e41b),
	.w7(32'hb5b9ac3d),
	.w8(32'hb60fd026),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h335bd611),
	.w1(32'hb7755eb4),
	.w2(32'h3668b150),
	.w3(32'hb7b0cd3a),
	.w4(32'hb7672430),
	.w5(32'hb5d9a0bb),
	.w6(32'hb7a32546),
	.w7(32'hb7c58c4c),
	.w8(32'hb7065400),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71457ce),
	.w1(32'hb6e88113),
	.w2(32'hb7ed5d97),
	.w3(32'hb5d4568f),
	.w4(32'hb718e2db),
	.w5(32'hb7ed22e2),
	.w6(32'h36cb2f85),
	.w7(32'hb67ced23),
	.w8(32'hb782361d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38432872),
	.w1(32'hba2eedd5),
	.w2(32'hba3dad82),
	.w3(32'h37c3a93b),
	.w4(32'hba19dcd1),
	.w5(32'hba587bcc),
	.w6(32'hba4b87f7),
	.w7(32'hba44bf1b),
	.w8(32'hb9bf9b36),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fc438),
	.w1(32'hbb1d043c),
	.w2(32'hbb032524),
	.w3(32'h3a812be3),
	.w4(32'h3a908dd0),
	.w5(32'h3a9c90ab),
	.w6(32'hba4af8a0),
	.w7(32'hb9801553),
	.w8(32'h3a4605ff),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb573d73),
	.w1(32'hbb1150c4),
	.w2(32'hba0f1d3e),
	.w3(32'hbace82d3),
	.w4(32'hba69ce52),
	.w5(32'hba2ae7e9),
	.w6(32'hba239f97),
	.w7(32'hb986459c),
	.w8(32'hb7c8adab),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5582c),
	.w1(32'h38c3ad6b),
	.w2(32'h3a1701c4),
	.w3(32'hbaf83993),
	.w4(32'hb66a5338),
	.w5(32'h396909d6),
	.w6(32'h39e5951d),
	.w7(32'h3a0d2be8),
	.w8(32'h39903256),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c7dfe),
	.w1(32'h3973b83a),
	.w2(32'h3a091a93),
	.w3(32'h3a247d81),
	.w4(32'h3a952d35),
	.w5(32'h3a6b239d),
	.w6(32'hb88b746b),
	.w7(32'h39a81cbd),
	.w8(32'h3a40f52f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a6aee),
	.w1(32'h39d667e3),
	.w2(32'hb871bb13),
	.w3(32'h3a0f864e),
	.w4(32'hba3808f7),
	.w5(32'hbad8bdcf),
	.w6(32'h38d1e52c),
	.w7(32'hb9a16528),
	.w8(32'hb9e11e95),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0499b7),
	.w1(32'hba88f501),
	.w2(32'hb9879a42),
	.w3(32'hbabb7ee8),
	.w4(32'h3828f06f),
	.w5(32'h361016b7),
	.w6(32'hba8ad7ce),
	.w7(32'hb903c25c),
	.w8(32'hb9e646ad),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46e8d9),
	.w1(32'hba1ea710),
	.w2(32'hb9c011de),
	.w3(32'hba9b561c),
	.w4(32'hba7f7f33),
	.w5(32'hba7b3f27),
	.w6(32'hbaef7e2f),
	.w7(32'hb9c91701),
	.w8(32'hba1d65d5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb844f),
	.w1(32'hbae548ca),
	.w2(32'h392ffd04),
	.w3(32'hbb04e2cd),
	.w4(32'h391ab59f),
	.w5(32'h3984eb37),
	.w6(32'h3ad40dbd),
	.w7(32'h3a178746),
	.w8(32'h3a662a24),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d9b30),
	.w1(32'hb753f77f),
	.w2(32'hba24c9b2),
	.w3(32'hb7d0a641),
	.w4(32'hb9f6dd2a),
	.w5(32'hba3c2cd0),
	.w6(32'hba29eb96),
	.w7(32'hb9da5fd8),
	.w8(32'hb9bb41aa),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a9e83),
	.w1(32'hba11d92d),
	.w2(32'hb9b62c97),
	.w3(32'hba790f4f),
	.w4(32'hb9c251fb),
	.w5(32'hb91bcc50),
	.w6(32'hb9190a73),
	.w7(32'hb9aae88e),
	.w8(32'hb84a0256),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75cca7),
	.w1(32'hb964d036),
	.w2(32'h39bcd39e),
	.w3(32'hbaf7d4da),
	.w4(32'h3a90b3ef),
	.w5(32'h3a7e5aa6),
	.w6(32'h3b0349ce),
	.w7(32'h3ae3ffbd),
	.w8(32'h3aeec036),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2e8c8),
	.w1(32'hb91d2e25),
	.w2(32'hb99bff4d),
	.w3(32'h3ae81cbe),
	.w4(32'h39e1d3b7),
	.w5(32'hba19b6d3),
	.w6(32'hb9ab7926),
	.w7(32'h3a362394),
	.w8(32'h398c6cb4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2e3aa),
	.w1(32'hbb162262),
	.w2(32'hbacbe207),
	.w3(32'hba400f45),
	.w4(32'hbacc7e0b),
	.w5(32'hbaa38a6a),
	.w6(32'h3a529276),
	.w7(32'h39c8cb77),
	.w8(32'hb8b8b558),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad50a6f),
	.w1(32'hb94fa93e),
	.w2(32'hb8aff288),
	.w3(32'hbab43226),
	.w4(32'hb9ea9d57),
	.w5(32'hba1bf51d),
	.w6(32'hb9add499),
	.w7(32'hb98caa98),
	.w8(32'hb9177421),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26b825),
	.w1(32'h3a7fae44),
	.w2(32'hbad6e2df),
	.w3(32'hbb28bdad),
	.w4(32'h39daae6d),
	.w5(32'hba176bf7),
	.w6(32'hbb37071f),
	.w7(32'h39c1e8fc),
	.w8(32'h3710aa2d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ab1af),
	.w1(32'hbb0ef6de),
	.w2(32'hbb0c0a2f),
	.w3(32'hb9df27c4),
	.w4(32'hbaa2b9f3),
	.w5(32'hbae2c0ca),
	.w6(32'hb9af8b30),
	.w7(32'h39adb14a),
	.w8(32'hba0a0d12),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae12fb8),
	.w1(32'hba222a6c),
	.w2(32'hb9e46db0),
	.w3(32'hba6de1bc),
	.w4(32'hba50a9a6),
	.w5(32'hba457555),
	.w6(32'hba46c97c),
	.w7(32'hba37020a),
	.w8(32'hb9d9d878),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c46cb),
	.w1(32'h399a063c),
	.w2(32'h394aa9e7),
	.w3(32'hba6bb05d),
	.w4(32'h3a8b7bf6),
	.w5(32'h3ab6c819),
	.w6(32'h3a0233e4),
	.w7(32'h39482777),
	.w8(32'h3a3bcc8e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939a5bf),
	.w1(32'hba06a0e9),
	.w2(32'h39cabd98),
	.w3(32'h3a5c2065),
	.w4(32'hb93ef45c),
	.w5(32'h38eecebc),
	.w6(32'h3a214122),
	.w7(32'h39ea760b),
	.w8(32'h399f9140),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6e6ca),
	.w1(32'hb9504ea7),
	.w2(32'hb924042a),
	.w3(32'hb9131b74),
	.w4(32'hb9e54276),
	.w5(32'hba028886),
	.w6(32'hb99d7348),
	.w7(32'hb98f74c0),
	.w8(32'hb948343f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da97b5),
	.w1(32'hba13829a),
	.w2(32'h3987f9df),
	.w3(32'hb984c029),
	.w4(32'hba5408f4),
	.w5(32'hb8ae5a0c),
	.w6(32'hb9948a61),
	.w7(32'hb9d1e3c4),
	.w8(32'h38aea529),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8935fdd),
	.w1(32'hba12e207),
	.w2(32'hba58cf93),
	.w3(32'hb9467d42),
	.w4(32'hba250970),
	.w5(32'hba1f3ed9),
	.w6(32'hb9e28c65),
	.w7(32'hba1e7214),
	.w8(32'hb9dc72f9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd5a40),
	.w1(32'hb8bfda10),
	.w2(32'h3a9f0767),
	.w3(32'hbaa3c0a3),
	.w4(32'hba54b260),
	.w5(32'hb989d637),
	.w6(32'h3a981953),
	.w7(32'h3aed95e2),
	.w8(32'h3ac675f6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37db1dbf),
	.w1(32'h3a10683c),
	.w2(32'h39f5a7e5),
	.w3(32'hba08df98),
	.w4(32'h3a21269b),
	.w5(32'h39708c32),
	.w6(32'h39dc6bcb),
	.w7(32'hb9530c45),
	.w8(32'h3a61121d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f5c58),
	.w1(32'hbb16745c),
	.w2(32'hba800e48),
	.w3(32'hba7e386a),
	.w4(32'hbaa5f852),
	.w5(32'hba9b13f7),
	.w6(32'h3ab6b1f4),
	.w7(32'h3a0e2663),
	.w8(32'h397241fc),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e012ce),
	.w1(32'h3ab7b0ee),
	.w2(32'h3a9377d8),
	.w3(32'hbb065318),
	.w4(32'hbb0c6fd2),
	.w5(32'hbab29cf9),
	.w6(32'hba643fd5),
	.w7(32'h3a10c025),
	.w8(32'h391e9191),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6125b),
	.w1(32'h398d2cfb),
	.w2(32'hb91fc0cf),
	.w3(32'hba066258),
	.w4(32'h3a11fbad),
	.w5(32'h3a6bf522),
	.w6(32'h3a1076c8),
	.w7(32'h3a433d47),
	.w8(32'h3a51f15a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db918b),
	.w1(32'h396dc0b0),
	.w2(32'h399cd605),
	.w3(32'h3906b673),
	.w4(32'hb8891bb8),
	.w5(32'h3a2c0874),
	.w6(32'hb9aa25b1),
	.w7(32'hb94e8539),
	.w8(32'h39cfa048),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c857a),
	.w1(32'h3a05caf6),
	.w2(32'h37f5fe7f),
	.w3(32'h397d7fb1),
	.w4(32'hba3ef738),
	.w5(32'hba98d29f),
	.w6(32'h39b6de30),
	.w7(32'h399f3f9b),
	.w8(32'hb89e88a1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeeeb9c),
	.w1(32'h3aba6022),
	.w2(32'hb99ece66),
	.w3(32'hb7c26cc0),
	.w4(32'h3a881922),
	.w5(32'hb8a0b61d),
	.w6(32'h3a0b5543),
	.w7(32'hba29040e),
	.w8(32'hb921e0b0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c32291),
	.w1(32'h3a09f5ce),
	.w2(32'hba1ca855),
	.w3(32'h3a08384a),
	.w4(32'h3a1f87a5),
	.w5(32'hb9b383cf),
	.w6(32'hb8858888),
	.w7(32'hba1e36c8),
	.w8(32'hba2bea68),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c9fb9),
	.w1(32'hb9b2c512),
	.w2(32'hb7ba8f4f),
	.w3(32'hba31b828),
	.w4(32'hb97ba02a),
	.w5(32'hb97fd5f6),
	.w6(32'hb80aaf63),
	.w7(32'hb96cbb5f),
	.w8(32'hb9457478),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b820cc),
	.w1(32'hb9d0a6c4),
	.w2(32'hb97cc071),
	.w3(32'hb81a9d4f),
	.w4(32'hb9ff0aa0),
	.w5(32'hb9f7a747),
	.w6(32'hb9a91b08),
	.w7(32'hb98ce294),
	.w8(32'hb86911bf),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34f5d9),
	.w1(32'hbad805f2),
	.w2(32'h3981d08e),
	.w3(32'hbab3bdb5),
	.w4(32'h39f7e59c),
	.w5(32'h3aa27f2c),
	.w6(32'h3a4e4f15),
	.w7(32'h39d8a3fc),
	.w8(32'h3a1c1de1),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39532ded),
	.w1(32'hba956420),
	.w2(32'hbaa3c55f),
	.w3(32'h39b4755d),
	.w4(32'hba748987),
	.w5(32'hba2c90a5),
	.w6(32'hba87f2c6),
	.w7(32'hba8c6a73),
	.w8(32'h390e3e42),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3daf5f),
	.w1(32'h39dd3a98),
	.w2(32'h3922f653),
	.w3(32'h393c4b1e),
	.w4(32'h39b88788),
	.w5(32'h39e38128),
	.w6(32'hb9e40e00),
	.w7(32'h39c94887),
	.w8(32'h3997e4e6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c4bfd),
	.w1(32'hb9cf6f8d),
	.w2(32'hb9d9258a),
	.w3(32'h3a51da1e),
	.w4(32'hb9e86432),
	.w5(32'hb9a6c535),
	.w6(32'hb91e8a6e),
	.w7(32'hb946e23b),
	.w8(32'h391a208c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2494d8),
	.w1(32'hba1ea8a1),
	.w2(32'h39a9a9a4),
	.w3(32'h39570708),
	.w4(32'h3a8ad909),
	.w5(32'h3a7cb94c),
	.w6(32'hb7c6bb9f),
	.w7(32'h3a19e06a),
	.w8(32'h3a5ae7e8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d2956),
	.w1(32'h390ba537),
	.w2(32'h394b8bb5),
	.w3(32'h3973c9e9),
	.w4(32'h3973cc23),
	.w5(32'h39bdd78e),
	.w6(32'hb95c718c),
	.w7(32'hb91ac2d0),
	.w8(32'hb954241b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c1a35),
	.w1(32'hba29aeed),
	.w2(32'hba15d5d5),
	.w3(32'h39cf70f0),
	.w4(32'hba31b826),
	.w5(32'hba3ff50a),
	.w6(32'hba39fb5e),
	.w7(32'hba32b1e8),
	.w8(32'hb9910526),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994ab4d),
	.w1(32'h39516e4b),
	.w2(32'hb94b1cdc),
	.w3(32'hba62af7a),
	.w4(32'hb90b3849),
	.w5(32'hb92b1277),
	.w6(32'hb98229af),
	.w7(32'hb9847389),
	.w8(32'hb9f25aa5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabde48e),
	.w1(32'hbaf9d418),
	.w2(32'hba5cfd76),
	.w3(32'h3aad45c3),
	.w4(32'h3a5979db),
	.w5(32'h39bcd485),
	.w6(32'hba2b31b9),
	.w7(32'hba6d75a2),
	.w8(32'hb9147e49),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83ff1d),
	.w1(32'hb9c53674),
	.w2(32'hb9c3a837),
	.w3(32'hba0e6643),
	.w4(32'hb9321fd5),
	.w5(32'hb89659d9),
	.w6(32'hb96ae1e5),
	.w7(32'hb9b1aa5d),
	.w8(32'hb9a4ea95),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9579eff),
	.w1(32'hba1421ba),
	.w2(32'hba40589e),
	.w3(32'hb9b08449),
	.w4(32'hba5b9c8c),
	.w5(32'hba8af00e),
	.w6(32'hba8700e6),
	.w7(32'hba3e51d4),
	.w8(32'hba4a7ddf),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e55f7),
	.w1(32'h3aa40152),
	.w2(32'h3ace4444),
	.w3(32'hba5b7de3),
	.w4(32'h3a62f37e),
	.w5(32'h3aa4d715),
	.w6(32'h3a5432f5),
	.w7(32'h3a6446b0),
	.w8(32'h3a3e382a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7816390),
	.w1(32'h3ad77a61),
	.w2(32'h3b48ead5),
	.w3(32'h3b063724),
	.w4(32'h39efbea0),
	.w5(32'h3abdfdd5),
	.w6(32'h3a96450d),
	.w7(32'hb9be6806),
	.w8(32'hb7d884a2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fb8bb),
	.w1(32'hba7749a7),
	.w2(32'h3938f0dc),
	.w3(32'hba760bff),
	.w4(32'hb9f021a8),
	.w5(32'h38abf1b0),
	.w6(32'hb93bcf22),
	.w7(32'h39c0f22b),
	.w8(32'h3a60945f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1f92d),
	.w1(32'hbaf6d913),
	.w2(32'hbaad6183),
	.w3(32'hb9d4338d),
	.w4(32'hb9665c5e),
	.w5(32'h37b2e0b0),
	.w6(32'h39eb1a3c),
	.w7(32'hba23b9a4),
	.w8(32'hba206622),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08be12),
	.w1(32'h3a8ddab9),
	.w2(32'hb889442b),
	.w3(32'hba552804),
	.w4(32'h3acb4121),
	.w5(32'h3a1a2e7c),
	.w6(32'h3aa8130f),
	.w7(32'h39b052b2),
	.w8(32'h3a0cc7c7),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba120fe3),
	.w1(32'hba5cbf51),
	.w2(32'hb968a8cd),
	.w3(32'h3a839cfa),
	.w4(32'hb98ec609),
	.w5(32'h3818cba6),
	.w6(32'hb8f8692d),
	.w7(32'h399d8d40),
	.w8(32'h3a150c89),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2ed9f),
	.w1(32'hb9aca410),
	.w2(32'hb95d2d83),
	.w3(32'hba114633),
	.w4(32'hb9b43e17),
	.w5(32'hb9a70d13),
	.w6(32'hb9ab056c),
	.w7(32'hb9a08638),
	.w8(32'hb8f1d53a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bddec5),
	.w1(32'h39f09ab9),
	.w2(32'h3961b69b),
	.w3(32'hba0137f6),
	.w4(32'h3a8d12fa),
	.w5(32'h3a5385e4),
	.w6(32'h39c85191),
	.w7(32'h39a9539d),
	.w8(32'h3991e544),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2ca19),
	.w1(32'h3817aad4),
	.w2(32'h39c321ce),
	.w3(32'h3a55eb2b),
	.w4(32'hba183f09),
	.w5(32'hba690419),
	.w6(32'h3991774f),
	.w7(32'hb906b8e3),
	.w8(32'hba5f688d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d4844),
	.w1(32'hba2f824c),
	.w2(32'h3aacbfd3),
	.w3(32'hbb146dc8),
	.w4(32'hba335d62),
	.w5(32'h3a83df84),
	.w6(32'hb9b0be6e),
	.w7(32'h3a294456),
	.w8(32'h3a6ca621),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39996e6e),
	.w1(32'hba492be8),
	.w2(32'h391ad367),
	.w3(32'hb9ad5abf),
	.w4(32'hba1a8c9d),
	.w5(32'hb9a2d0bd),
	.w6(32'hb9760574),
	.w7(32'hb90e5f33),
	.w8(32'hb9cd454b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb705065e),
	.w1(32'h386ae18d),
	.w2(32'hb8b4597b),
	.w3(32'hb9907a09),
	.w4(32'h3934dc29),
	.w5(32'h36891c53),
	.w6(32'h39f1892d),
	.w7(32'h3994320e),
	.w8(32'h39bd5492),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19c6d7),
	.w1(32'hb9a8a3bf),
	.w2(32'hba8dad50),
	.w3(32'h388947c6),
	.w4(32'hb91ab80c),
	.w5(32'hb90664ff),
	.w6(32'hba84b1d0),
	.w7(32'hba32f41b),
	.w8(32'hb97bf614),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1300ba),
	.w1(32'h3ac5c22c),
	.w2(32'h3b412fd2),
	.w3(32'hba72dfa5),
	.w4(32'h395ce553),
	.w5(32'h3b1f99b8),
	.w6(32'h3a14366c),
	.w7(32'h3a865dd7),
	.w8(32'h3ad51fdf),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00961d),
	.w1(32'hbb846220),
	.w2(32'hbacdeb24),
	.w3(32'h39fe6ff5),
	.w4(32'hba32ab4e),
	.w5(32'hbadc3a50),
	.w6(32'hba9743ec),
	.w7(32'hba92bd7e),
	.w8(32'hbaccd6c1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ab105),
	.w1(32'h39ccbb86),
	.w2(32'h391d1449),
	.w3(32'hba9dd65c),
	.w4(32'h3a011021),
	.w5(32'h39c94bd9),
	.w6(32'hb851100d),
	.w7(32'hb93a2c9d),
	.w8(32'hb9176d77),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb642d5a),
	.w1(32'hbb02b3c1),
	.w2(32'h39baa853),
	.w3(32'h3aafe660),
	.w4(32'h3a08d613),
	.w5(32'h3a84558c),
	.w6(32'h3a4e8555),
	.w7(32'hba1a9d41),
	.w8(32'h3a5a488d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4125a2),
	.w1(32'hba6e0eb3),
	.w2(32'hb9ff8645),
	.w3(32'hbb20d21d),
	.w4(32'hbb0eb2fc),
	.w5(32'hbaa06e57),
	.w6(32'hbae15b5a),
	.w7(32'hb9d0be80),
	.w8(32'hbaac82c4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cd6d7),
	.w1(32'hbaa16b2d),
	.w2(32'hb8b1afa2),
	.w3(32'h391a71a3),
	.w4(32'hb9712f3a),
	.w5(32'h38ee75b0),
	.w6(32'hb8e511a0),
	.w7(32'hb98088d4),
	.w8(32'hb9eb31c4),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394906e6),
	.w1(32'h399da6a9),
	.w2(32'h3a999cee),
	.w3(32'h39bb71de),
	.w4(32'h37b71208),
	.w5(32'h3a8e8b16),
	.w6(32'hb87f4555),
	.w7(32'h37ef0a02),
	.w8(32'h3a19e966),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a759c8b),
	.w1(32'h3a541796),
	.w2(32'h3a2de442),
	.w3(32'h39f55f8b),
	.w4(32'h3a51fee5),
	.w5(32'h3a57a91b),
	.w6(32'h3a24d59f),
	.w7(32'h3a0c89f5),
	.w8(32'h3a09d033),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a674863),
	.w1(32'h39816865),
	.w2(32'h35f67e12),
	.w3(32'h3a81ceed),
	.w4(32'h3992b2a3),
	.w5(32'h38f45f6d),
	.w6(32'h38aa3fe7),
	.w7(32'hb91483fd),
	.w8(32'h3990e1f2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95b8d0),
	.w1(32'hbaca3feb),
	.w2(32'hbaa03add),
	.w3(32'h3a18ca0c),
	.w4(32'hb9dbe787),
	.w5(32'hba875ba6),
	.w6(32'hba4f68c4),
	.w7(32'hba919002),
	.w8(32'hb904d287),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba756b89),
	.w1(32'hb98ceb69),
	.w2(32'h37268407),
	.w3(32'hba67602f),
	.w4(32'h39dae97c),
	.w5(32'h3a3532bf),
	.w6(32'hb7c371a7),
	.w7(32'hb90496c9),
	.w8(32'hb93ca698),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a139614),
	.w1(32'h39bc8025),
	.w2(32'h38824f3a),
	.w3(32'h39518eec),
	.w4(32'h39a625ec),
	.w5(32'hb7a74b93),
	.w6(32'hb912dc56),
	.w7(32'h391ffeba),
	.w8(32'hb8b9cbd2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986b184),
	.w1(32'hb9d4d583),
	.w2(32'hb9b0c202),
	.w3(32'h39deab18),
	.w4(32'hba32d5d4),
	.w5(32'hba50965e),
	.w6(32'hba2fe073),
	.w7(32'hba1974db),
	.w8(32'hba015e5d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16d2f6),
	.w1(32'hb9e2fe39),
	.w2(32'h39ad7807),
	.w3(32'hbaa82629),
	.w4(32'h3a58473f),
	.w5(32'h39db4a6f),
	.w6(32'h39afe600),
	.w7(32'hb919db81),
	.w8(32'h39c3236a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca3935),
	.w1(32'h39a048be),
	.w2(32'h3a3b965f),
	.w3(32'h3a0f6749),
	.w4(32'hb92a4b28),
	.w5(32'h3a2bab7a),
	.w6(32'hb91f3d59),
	.w7(32'hb9f2391d),
	.w8(32'h38da97ca),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2b323),
	.w1(32'hba29e0fc),
	.w2(32'hba13c4a9),
	.w3(32'h3a09fb7a),
	.w4(32'hba134b8a),
	.w5(32'hba08759c),
	.w6(32'hba1944bc),
	.w7(32'hba4abe8f),
	.w8(32'hb9b0eee0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa00c28),
	.w1(32'hbaaad679),
	.w2(32'h3a6ef022),
	.w3(32'hba9da28d),
	.w4(32'h38a13931),
	.w5(32'h392f65b8),
	.w6(32'hba092d4c),
	.w7(32'h397a010f),
	.w8(32'h3a73376a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f575c5),
	.w1(32'hba16325d),
	.w2(32'hba0af383),
	.w3(32'hba2306cf),
	.w4(32'hba35b13b),
	.w5(32'hba1b6d63),
	.w6(32'hb99da683),
	.w7(32'hb9b6db54),
	.w8(32'hb96faa6a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ec8b4),
	.w1(32'h3a2ade5c),
	.w2(32'h3a659080),
	.w3(32'hba4413f9),
	.w4(32'h3a141ef7),
	.w5(32'h39b46427),
	.w6(32'h3a138d91),
	.w7(32'h395b7505),
	.w8(32'h394314ff),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace79a6),
	.w1(32'hb9932612),
	.w2(32'hbac4355f),
	.w3(32'hb955d320),
	.w4(32'hbad7e81e),
	.w5(32'hbb02aa18),
	.w6(32'h3aa682a7),
	.w7(32'h3a9cd051),
	.w8(32'hba031ab2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6627e),
	.w1(32'h39692952),
	.w2(32'hb85c8f48),
	.w3(32'hbab49ab6),
	.w4(32'hb9cc87f4),
	.w5(32'hba2d3068),
	.w6(32'hba53340e),
	.w7(32'hba7913bb),
	.w8(32'hba02e51e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8efe73e),
	.w1(32'h3a286ffd),
	.w2(32'h399da25e),
	.w3(32'hb9987585),
	.w4(32'h3a03a9a1),
	.w5(32'h3a1522cf),
	.w6(32'h3a2bc929),
	.w7(32'h39747581),
	.w8(32'h3988ce42),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fe0c6),
	.w1(32'h3a5b2fa1),
	.w2(32'h39555962),
	.w3(32'h39954a1b),
	.w4(32'hb912b38f),
	.w5(32'h39229659),
	.w6(32'h39becc5c),
	.w7(32'h3a9d485c),
	.w8(32'h3a21f6ce),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46afe9),
	.w1(32'hba8ea32d),
	.w2(32'hb9909f34),
	.w3(32'h3959183c),
	.w4(32'hb94761c2),
	.w5(32'hb9f18529),
	.w6(32'hb9a41274),
	.w7(32'hb93c8105),
	.w8(32'hb8a17b37),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0674ec),
	.w1(32'hb9e7c7c9),
	.w2(32'h39cc9d6b),
	.w3(32'hb9fcadbb),
	.w4(32'hb9838167),
	.w5(32'h3a1c6734),
	.w6(32'h39b7e63c),
	.w7(32'h37c02e5c),
	.w8(32'h3791e4b2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9884842),
	.w1(32'h39d53c48),
	.w2(32'h3a5018ae),
	.w3(32'h3a0f94c9),
	.w4(32'h39dd0d4a),
	.w5(32'h3a3916d4),
	.w6(32'h39baecf5),
	.w7(32'h3a2f5309),
	.w8(32'h39c91aca),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af7a80),
	.w1(32'h39a09df0),
	.w2(32'h392014c0),
	.w3(32'h39a772f7),
	.w4(32'h39f682b0),
	.w5(32'h39e68a25),
	.w6(32'h3a162d42),
	.w7(32'h39a50530),
	.w8(32'h39b5eb15),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6f699),
	.w1(32'h370d25cb),
	.w2(32'hb9984559),
	.w3(32'h3a1bed20),
	.w4(32'h39c58b9b),
	.w5(32'h3a9fffd6),
	.w6(32'h37e2f807),
	.w7(32'hb86a0a4e),
	.w8(32'h3a7df8b6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85f7a3),
	.w1(32'hb9c4869b),
	.w2(32'h3a4fbf00),
	.w3(32'h3abc69bb),
	.w4(32'h3ab82610),
	.w5(32'h3ab88023),
	.w6(32'h384a671d),
	.w7(32'h3a3291bc),
	.w8(32'h3ac135c9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5d315),
	.w1(32'h3af349de),
	.w2(32'h3a973e3e),
	.w3(32'h39fe4e8f),
	.w4(32'h3a889a74),
	.w5(32'h3a94e07c),
	.w6(32'h3a3efd09),
	.w7(32'h3a9c5ffe),
	.w8(32'h3a1bc93c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8e824),
	.w1(32'hbb687179),
	.w2(32'hbacf243e),
	.w3(32'hbaa1a591),
	.w4(32'hb9c00800),
	.w5(32'hbaf25f1f),
	.w6(32'h3b145683),
	.w7(32'h3a58bdf4),
	.w8(32'h3a948b58),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba432e90),
	.w1(32'hb9b62c3f),
	.w2(32'hb9ed98f1),
	.w3(32'h3938a732),
	.w4(32'hb9678d05),
	.w5(32'hb91c5507),
	.w6(32'hb91b2915),
	.w7(32'hb843b6f2),
	.w8(32'h390c5d1a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba162ec7),
	.w1(32'hba1757ef),
	.w2(32'h37b9302c),
	.w3(32'h39313d5c),
	.w4(32'h3934e685),
	.w5(32'h39e755ea),
	.w6(32'hb8745e47),
	.w7(32'h39dc45db),
	.w8(32'h3a4707de),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d2819),
	.w1(32'hbb159e14),
	.w2(32'hbb46bca5),
	.w3(32'h3a845d08),
	.w4(32'hba774c06),
	.w5(32'hbb02823b),
	.w6(32'h3a2f4947),
	.w7(32'hbaf3a7f5),
	.w8(32'hba0b542b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb691312),
	.w1(32'hbac63e7d),
	.w2(32'hb8fda2c2),
	.w3(32'hb7af32a5),
	.w4(32'h398206fe),
	.w5(32'h3a0791ec),
	.w6(32'h3a8af1f6),
	.w7(32'hb996b609),
	.w8(32'h3a3903a6),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0d25),
	.w1(32'hba813727),
	.w2(32'h37426a62),
	.w3(32'hba9bb9d5),
	.w4(32'h39f38a58),
	.w5(32'h39b9492d),
	.w6(32'h3aa58094),
	.w7(32'h3a8ee9b8),
	.w8(32'h39d03311),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68f655),
	.w1(32'h3ad29b00),
	.w2(32'h3a8eb82c),
	.w3(32'h3a1bc47c),
	.w4(32'h3a30dbf3),
	.w5(32'h38940988),
	.w6(32'h39cf5d3c),
	.w7(32'h3aa527a2),
	.w8(32'h3a267d71),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e1f48),
	.w1(32'h3a8cd0c2),
	.w2(32'h38c5d356),
	.w3(32'h39681d3a),
	.w4(32'h39c0ec13),
	.w5(32'hb857e972),
	.w6(32'hba43f0aa),
	.w7(32'hba0dd229),
	.w8(32'hb9d63df6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1aeb2),
	.w1(32'h38ae27dd),
	.w2(32'h38b22ad8),
	.w3(32'h39c2c052),
	.w4(32'h397db788),
	.w5(32'h396fb519),
	.w6(32'hb96a4000),
	.w7(32'hb9c04232),
	.w8(32'hb95160d8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3874417c),
	.w1(32'hba8dc9d3),
	.w2(32'hba382f17),
	.w3(32'h392f3b68),
	.w4(32'hba51edaa),
	.w5(32'hba3b00b5),
	.w6(32'hba8486a7),
	.w7(32'hba5edc17),
	.w8(32'hba290078),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf44a1),
	.w1(32'hbab38867),
	.w2(32'hbaaf2030),
	.w3(32'hb903f8a4),
	.w4(32'h38b66d46),
	.w5(32'h387ad784),
	.w6(32'h3a1b242b),
	.w7(32'hba337ddf),
	.w8(32'h3a706dc6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5f951),
	.w1(32'h399fac9e),
	.w2(32'h375a638e),
	.w3(32'h3a4cef23),
	.w4(32'h382d5f62),
	.w5(32'hb90ca21e),
	.w6(32'h3923050b),
	.w7(32'hb7db79e0),
	.w8(32'h398b212b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be9f16),
	.w1(32'hb9575a21),
	.w2(32'h3980f2f2),
	.w3(32'h3a150665),
	.w4(32'h3a33a5cc),
	.w5(32'h3aa6d35b),
	.w6(32'hb92f4dbd),
	.w7(32'hb7b47f80),
	.w8(32'h39f7a6e7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa27ec4),
	.w1(32'h39279530),
	.w2(32'h39840e11),
	.w3(32'h3a9ad73a),
	.w4(32'h3ade19a1),
	.w5(32'h3a55858d),
	.w6(32'h39b2ad76),
	.w7(32'h3abec712),
	.w8(32'h3aeff5a1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ec4ba),
	.w1(32'hbaa18689),
	.w2(32'hb9a21ef3),
	.w3(32'hb7c2e98b),
	.w4(32'hb9fb0bb4),
	.w5(32'hb68dae23),
	.w6(32'hba971e0a),
	.w7(32'hba3ec279),
	.w8(32'h3984ea8f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cd3b3),
	.w1(32'hb7b00b7f),
	.w2(32'h3a04c802),
	.w3(32'hb9da39f2),
	.w4(32'h38a12754),
	.w5(32'h391cad73),
	.w6(32'h38bfceb8),
	.w7(32'h38adeacb),
	.w8(32'h3a256ab3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb918468),
	.w1(32'hbb7d652d),
	.w2(32'hbabb0656),
	.w3(32'h388bef82),
	.w4(32'hba001e32),
	.w5(32'hb8f671f1),
	.w6(32'h39df4084),
	.w7(32'hba01677a),
	.w8(32'h3a90783c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb79da),
	.w1(32'hba8d87c9),
	.w2(32'hba1e452c),
	.w3(32'hba289701),
	.w4(32'hb9af37bc),
	.w5(32'hb9b1a9b5),
	.w6(32'hb9f8aec3),
	.w7(32'hba2c100f),
	.w8(32'h397a186a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a5fb3),
	.w1(32'hb964a421),
	.w2(32'hb98dea61),
	.w3(32'hb9d60c7c),
	.w4(32'hb987dca0),
	.w5(32'hb9d350ea),
	.w6(32'hba0119ad),
	.w7(32'hba24dfc2),
	.w8(32'hb95a10ab),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb206fb6),
	.w1(32'hbabf26dc),
	.w2(32'hba3f94f9),
	.w3(32'hba924e1d),
	.w4(32'hba69ca4b),
	.w5(32'hba101fce),
	.w6(32'h39ada542),
	.w7(32'hb9b5aab9),
	.w8(32'hb8fac80c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d4db8),
	.w1(32'h3a036542),
	.w2(32'h3a0e44b8),
	.w3(32'hb96060e7),
	.w4(32'h39cce3a2),
	.w5(32'h3a2d2ba6),
	.w6(32'hb92578f6),
	.w7(32'hb9801ae8),
	.w8(32'hb952a5d6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a41911),
	.w1(32'hb991013e),
	.w2(32'hb9520605),
	.w3(32'h3a1ac30a),
	.w4(32'hb9c76db7),
	.w5(32'hb93fa74f),
	.w6(32'hb89048a4),
	.w7(32'hb95f214f),
	.w8(32'hb943024f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976e587),
	.w1(32'hb958d382),
	.w2(32'hb98a1c80),
	.w3(32'hb9886f74),
	.w4(32'hb93b93fb),
	.w5(32'hb9a9061c),
	.w6(32'hba1bca7e),
	.w7(32'hba427a96),
	.w8(32'hb9ac76e9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91062c5),
	.w1(32'h398e6b9d),
	.w2(32'hb91f4c81),
	.w3(32'hb97d548b),
	.w4(32'h39d912ff),
	.w5(32'h3944f026),
	.w6(32'h3a132ef0),
	.w7(32'hb78b7ca0),
	.w8(32'hb98c2838),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9494a80),
	.w1(32'hba592e61),
	.w2(32'hba4741a5),
	.w3(32'hb96412d2),
	.w4(32'hba9b0048),
	.w5(32'hbab3d2ea),
	.w6(32'hba610b00),
	.w7(32'hba7de32f),
	.w8(32'hba5b45cb),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889c52),
	.w1(32'hba46bd55),
	.w2(32'h3ab22c9d),
	.w3(32'hbb6c4ef4),
	.w4(32'hba961db2),
	.w5(32'h39a71567),
	.w6(32'h3a4c1e35),
	.w7(32'h39ebcb6c),
	.w8(32'hb90f27b4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ce102),
	.w1(32'hbae729e1),
	.w2(32'hba1fc080),
	.w3(32'hbb0c7996),
	.w4(32'hba988852),
	.w5(32'hba91b16e),
	.w6(32'hb7ce3cf5),
	.w7(32'hb982b3c9),
	.w8(32'h3958dd91),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7277d5),
	.w1(32'hbab2a6e5),
	.w2(32'hb8ed0f6e),
	.w3(32'hbb1d3f7f),
	.w4(32'hba1b077b),
	.w5(32'hba0a252e),
	.w6(32'h3a88350e),
	.w7(32'hb8f40007),
	.w8(32'h39d54623),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0f4c4),
	.w1(32'hba162039),
	.w2(32'hb8c0d687),
	.w3(32'hb993ea69),
	.w4(32'hba01269a),
	.w5(32'hba17276f),
	.w6(32'hb9f3549d),
	.w7(32'hb9aa1d99),
	.w8(32'hb8cd2e1a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e45d2e),
	.w1(32'hb989f26d),
	.w2(32'hb8c083b6),
	.w3(32'hb954dbd5),
	.w4(32'hb93a84d0),
	.w5(32'hb9957c83),
	.w6(32'hba681c3c),
	.w7(32'hba57ac1d),
	.w8(32'hb949b7b2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900385a),
	.w1(32'hb9ba98e3),
	.w2(32'hb99a7b20),
	.w3(32'hb99730b1),
	.w4(32'hb9bf6da3),
	.w5(32'hb9a0344a),
	.w6(32'hba1c42ed),
	.w7(32'hba253bbe),
	.w8(32'hb9a727cf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fcf631),
	.w1(32'hb9901394),
	.w2(32'hb94f56dd),
	.w3(32'hb9694c35),
	.w4(32'hb9e84c7d),
	.w5(32'hb9d5bee4),
	.w6(32'hba118fbc),
	.w7(32'hba0fe40d),
	.w8(32'hb97646ea),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8996ca),
	.w1(32'h3a26e38d),
	.w2(32'h3ace12f8),
	.w3(32'hb80d4159),
	.w4(32'h3a52d88d),
	.w5(32'h3aa8b4fd),
	.w6(32'h38d5ec67),
	.w7(32'h3a9df78d),
	.w8(32'h3a810d68),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999f414),
	.w1(32'hb99082ad),
	.w2(32'hb9a4152a),
	.w3(32'h369db6f0),
	.w4(32'h389b692a),
	.w5(32'hb9df6f0e),
	.w6(32'hb9a17076),
	.w7(32'hba32e10e),
	.w8(32'h39a74512),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901e35b),
	.w1(32'hba046c56),
	.w2(32'h38c85ab3),
	.w3(32'hb91c0cbc),
	.w4(32'hba566d1a),
	.w5(32'hba194c2d),
	.w6(32'hb95b4259),
	.w7(32'hb81752e8),
	.w8(32'h39e80dbf),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b8393),
	.w1(32'h39ac7671),
	.w2(32'h3a8adb0e),
	.w3(32'hb9e4ce39),
	.w4(32'hb9747b98),
	.w5(32'h39c9e5cd),
	.w6(32'h3984d10b),
	.w7(32'h39e99f58),
	.w8(32'h3a11949a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397244fc),
	.w1(32'hba13c976),
	.w2(32'hb9f12113),
	.w3(32'hb98e03e1),
	.w4(32'hba0d1e0f),
	.w5(32'hba05f327),
	.w6(32'hba3e7170),
	.w7(32'hba4d0727),
	.w8(32'hb9c974e4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dfb73),
	.w1(32'hb8e6d2b7),
	.w2(32'h39a0a109),
	.w3(32'hba10ef7d),
	.w4(32'h3a6386d9),
	.w5(32'h3ab732bb),
	.w6(32'hb98595b9),
	.w7(32'hb97424c8),
	.w8(32'hb9cbf0b9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980c163),
	.w1(32'hb9696f26),
	.w2(32'h3a48ae29),
	.w3(32'h3a36b98e),
	.w4(32'hb9c72c5d),
	.w5(32'hb9253cbd),
	.w6(32'hba33573d),
	.w7(32'h39a60547),
	.w8(32'h3a39cf4f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafab7d5),
	.w1(32'hbab513bc),
	.w2(32'h3a3c7e6c),
	.w3(32'hbb2fcb02),
	.w4(32'hba989c0a),
	.w5(32'h3a11a1f3),
	.w6(32'h3a94d74c),
	.w7(32'h3ae2885d),
	.w8(32'h3a93b30a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f9fe7),
	.w1(32'h3675d114),
	.w2(32'h388ef750),
	.w3(32'hb96f18fe),
	.w4(32'h379ac21a),
	.w5(32'h38b51fa8),
	.w6(32'hb84d658a),
	.w7(32'hb6026bb2),
	.w8(32'h389b98c1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91f08c),
	.w1(32'h39978bc5),
	.w2(32'hb9f39c1f),
	.w3(32'h3a50e89a),
	.w4(32'hb7b1c99c),
	.w5(32'h38a30d2e),
	.w6(32'h39ed7e3c),
	.w7(32'h3a1a06bf),
	.w8(32'h39f307cd),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule