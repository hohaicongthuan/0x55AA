module layer_10_featuremap_67(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6b282),
	.w1(32'h3bc3609d),
	.w2(32'h3c9980d5),
	.w3(32'h3bd33c2f),
	.w4(32'hbb51c4d7),
	.w5(32'h3c8d8552),
	.w6(32'h3c4b4267),
	.w7(32'h3a9652b6),
	.w8(32'h3c11012d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d362c),
	.w1(32'h3ba64db0),
	.w2(32'hbc1bf955),
	.w3(32'h3cb90895),
	.w4(32'h3bcb64e2),
	.w5(32'hbbad4089),
	.w6(32'h3c84ac1d),
	.w7(32'h3cafdb51),
	.w8(32'hbb7fc723),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9a5a2),
	.w1(32'hbbcb69d4),
	.w2(32'hbcadf9ab),
	.w3(32'hbc07661f),
	.w4(32'hbbfaae00),
	.w5(32'hbd1a83e5),
	.w6(32'h39cbd280),
	.w7(32'hbb4d09c5),
	.w8(32'hbc8a5f1d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d85a5),
	.w1(32'hbc05d7f0),
	.w2(32'hbc3a0a01),
	.w3(32'hbce697fe),
	.w4(32'hbc11001d),
	.w5(32'hbcb7cc6a),
	.w6(32'hbcc71490),
	.w7(32'hbbbbb60f),
	.w8(32'hbc9eb5e7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e6f94),
	.w1(32'h3a9a0f9e),
	.w2(32'hbc1ada16),
	.w3(32'hbaadc446),
	.w4(32'h3a87be08),
	.w5(32'hbc5d7e58),
	.w6(32'hbc894e7c),
	.w7(32'hbbb014b7),
	.w8(32'hbc11ef66),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce3e486),
	.w1(32'hbcb285aa),
	.w2(32'hbba64b23),
	.w3(32'hbcc29485),
	.w4(32'hbce6de49),
	.w5(32'hbb94584b),
	.w6(32'hbc6e6e8f),
	.w7(32'hbcbf8cb2),
	.w8(32'hbb43cae2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad716ec),
	.w1(32'hbbe5d643),
	.w2(32'hbb4fc35d),
	.w3(32'h3b8a34c0),
	.w4(32'h3a8a4c3e),
	.w5(32'hbc299d4b),
	.w6(32'h3b91e5a2),
	.w7(32'hbb8cb5a5),
	.w8(32'hbc4696bc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ffa84),
	.w1(32'hbc73e2c5),
	.w2(32'hbc0e40e8),
	.w3(32'hbc69e18a),
	.w4(32'hbc78c4af),
	.w5(32'hbc26e4aa),
	.w6(32'hbc7b222c),
	.w7(32'hbc31cc12),
	.w8(32'h3bd971b3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8788156),
	.w1(32'h3b3444bf),
	.w2(32'h3ad923fd),
	.w3(32'hbb8b0edd),
	.w4(32'hbb85c05a),
	.w5(32'h3abb6e0e),
	.w6(32'h3b96a787),
	.w7(32'h3aafc71e),
	.w8(32'h3bb72db3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d7fc2),
	.w1(32'h3a1b880a),
	.w2(32'h3b3eed2c),
	.w3(32'h3adb7d63),
	.w4(32'hba382193),
	.w5(32'h3aded0b0),
	.w6(32'hbb376a6a),
	.w7(32'hbbaa3a36),
	.w8(32'h3b0914a9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38838dac),
	.w1(32'h3aab956e),
	.w2(32'hbc3fff81),
	.w3(32'h3b25c81f),
	.w4(32'h3b08ff68),
	.w5(32'hbcfdbe9c),
	.w6(32'h3b8110c2),
	.w7(32'h3b5b1e0f),
	.w8(32'hbcaa02bc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a15da),
	.w1(32'hbc1f7a5a),
	.w2(32'hbbb8fe06),
	.w3(32'hbd0c19d5),
	.w4(32'hbc3512bc),
	.w5(32'hbba7bcfb),
	.w6(32'hbc9c14c4),
	.w7(32'hbc18727c),
	.w8(32'hbbbf65bc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cb238),
	.w1(32'hbc24e769),
	.w2(32'hbb33ce35),
	.w3(32'hbb0f54b7),
	.w4(32'hbbcacb29),
	.w5(32'hbaab9f0a),
	.w6(32'hbbc90121),
	.w7(32'hbb986858),
	.w8(32'hba99a53f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7aa63c),
	.w1(32'hbbdebd33),
	.w2(32'hbcadb23c),
	.w3(32'hba8c146c),
	.w4(32'h3aba40f7),
	.w5(32'hbd04d541),
	.w6(32'hbb549f87),
	.w7(32'hbb352bc3),
	.w8(32'hbc2bfb32),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b681e),
	.w1(32'hbb25d9b3),
	.w2(32'hbbe05770),
	.w3(32'hbcfb1fd8),
	.w4(32'hbbb725de),
	.w5(32'hbbd465c8),
	.w6(32'hbc73936a),
	.w7(32'hbbf095cd),
	.w8(32'hbb2433f6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25acc8),
	.w1(32'hba8f5991),
	.w2(32'h3b2b50fe),
	.w3(32'hbc038e89),
	.w4(32'hba7d8a74),
	.w5(32'h3b1e6668),
	.w6(32'hbb8b4ad7),
	.w7(32'h3b35027e),
	.w8(32'h3bb373d2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb73a4),
	.w1(32'h3a01e7b0),
	.w2(32'hbacdf729),
	.w3(32'h3b92f6b5),
	.w4(32'h3b145c34),
	.w5(32'hbaf61f50),
	.w6(32'h3bbf4631),
	.w7(32'h3ba0fe15),
	.w8(32'h3c30f5bb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50a4e5),
	.w1(32'hbc5bbb63),
	.w2(32'hb950986e),
	.w3(32'hbc1b54e7),
	.w4(32'hbc01e738),
	.w5(32'hbb868812),
	.w6(32'hbbbb75a8),
	.w7(32'hbbbc6d1c),
	.w8(32'h3b6d7969),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01626a),
	.w1(32'hbc19cac8),
	.w2(32'hbbe96fa1),
	.w3(32'hbc088a9d),
	.w4(32'hbc17e816),
	.w5(32'h3acce645),
	.w6(32'hbc0070db),
	.w7(32'hbc0cdfd9),
	.w8(32'h3c1af56e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002d71),
	.w1(32'hbb7022e6),
	.w2(32'h3bd2131d),
	.w3(32'h3bad7333),
	.w4(32'h3bf1a348),
	.w5(32'h3b71662c),
	.w6(32'h3c32b3e5),
	.w7(32'h3ca82405),
	.w8(32'h3adc3737),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840804),
	.w1(32'h3b03de26),
	.w2(32'hbbb4c0b3),
	.w3(32'hbb241f99),
	.w4(32'h3accaf86),
	.w5(32'hbba1e781),
	.w6(32'hbb3331f0),
	.w7(32'h3aed4407),
	.w8(32'hbb6b6bda),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac78bdb),
	.w1(32'h3bd563d6),
	.w2(32'h3b941593),
	.w3(32'h3c7488c5),
	.w4(32'h3c9059e4),
	.w5(32'hbbc0cb7b),
	.w6(32'h3c7f04e4),
	.w7(32'h3ca5b76d),
	.w8(32'hba04aad7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfec79),
	.w1(32'hbc5fe649),
	.w2(32'hbb35d922),
	.w3(32'h3b769521),
	.w4(32'hbc2125c1),
	.w5(32'hbb832d86),
	.w6(32'hbc43478f),
	.w7(32'hbc26d0bd),
	.w8(32'hbaa6bd3f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac03637),
	.w1(32'h3b18aec8),
	.w2(32'h3a5ad66d),
	.w3(32'h3ae844c9),
	.w4(32'hb8fc55f6),
	.w5(32'h3b06dcc5),
	.w6(32'h3ad87e79),
	.w7(32'h3b09f008),
	.w8(32'h3bccc340),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd266c),
	.w1(32'h3a1f996d),
	.w2(32'hbc965c35),
	.w3(32'hbb94e5f0),
	.w4(32'h3b13211d),
	.w5(32'hbb9c72fa),
	.w6(32'hbc15b846),
	.w7(32'h3a87053e),
	.w8(32'h3b3119a1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f673e),
	.w1(32'hbafebd64),
	.w2(32'hba346a48),
	.w3(32'h3c16c9c0),
	.w4(32'h3c13e6d1),
	.w5(32'hbcdc652f),
	.w6(32'h3c89139b),
	.w7(32'h3c40a0de),
	.w8(32'hbcdbbfd5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba80489),
	.w1(32'h3c647aec),
	.w2(32'hba8e49f3),
	.w3(32'hbba3783d),
	.w4(32'h3c7c51f0),
	.w5(32'h39c897db),
	.w6(32'hbbe4896d),
	.w7(32'h3b4bbd5b),
	.w8(32'hbae61242),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73e057),
	.w1(32'hbb31568c),
	.w2(32'hbaf16ad7),
	.w3(32'h3bf4fe40),
	.w4(32'h3bbedfe5),
	.w5(32'hbc838721),
	.w6(32'h39ccfca9),
	.w7(32'h3856bdd8),
	.w8(32'hbc13056f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04c8e9),
	.w1(32'h3b5824af),
	.w2(32'hb977da18),
	.w3(32'hba5a025a),
	.w4(32'h3bbd02d3),
	.w5(32'hbc103e92),
	.w6(32'hb9f8ec3a),
	.w7(32'hbbe4204b),
	.w8(32'hbbb1eaf4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68f03c),
	.w1(32'hbb059c68),
	.w2(32'h3b9172d1),
	.w3(32'hbca28404),
	.w4(32'hba4938e0),
	.w5(32'hba18ea95),
	.w6(32'h3acaa914),
	.w7(32'h3a7b52db),
	.w8(32'hbbc46de7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2acf94),
	.w1(32'hbaf61a36),
	.w2(32'hbc40e5e6),
	.w3(32'hbb7c5c7c),
	.w4(32'hbb35dfed),
	.w5(32'hbbfc7bda),
	.w6(32'hbb55f8c4),
	.w7(32'h3a23a220),
	.w8(32'hbbda38fc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3396b1),
	.w1(32'hbbf31190),
	.w2(32'hbc1ccc5c),
	.w3(32'hbb68e213),
	.w4(32'hbbd3ed7e),
	.w5(32'hbc64e990),
	.w6(32'hbad00a8d),
	.w7(32'hbbcaff17),
	.w8(32'h3b899d9e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25612b),
	.w1(32'hbbbefb9c),
	.w2(32'h3b9039d5),
	.w3(32'h3bcd2ea5),
	.w4(32'h3c09c8fd),
	.w5(32'h3a09fa59),
	.w6(32'h3c056846),
	.w7(32'hbba9ca32),
	.w8(32'h3ba6b8aa),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83557e),
	.w1(32'h3b738e2d),
	.w2(32'h3c88c333),
	.w3(32'h3b6a554f),
	.w4(32'hbb48f7fe),
	.w5(32'h3c557b95),
	.w6(32'h3a9ff2ee),
	.w7(32'hbbe592d6),
	.w8(32'hbb8cb1d2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c465f36),
	.w1(32'hbb9947f3),
	.w2(32'h3b0871b5),
	.w3(32'h3adeedcd),
	.w4(32'hbc3eb226),
	.w5(32'h3bbd233a),
	.w6(32'h3b57e4ae),
	.w7(32'hbb4fd962),
	.w8(32'h3c3202c8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be04edb),
	.w1(32'h3bf72e5b),
	.w2(32'h3c2fba0d),
	.w3(32'h3c38bca6),
	.w4(32'h3b2889d2),
	.w5(32'h3a8bd172),
	.w6(32'h3bd64435),
	.w7(32'hbbcef1f1),
	.w8(32'hbb862f35),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b124a1d),
	.w1(32'hbca270d0),
	.w2(32'hb93c8e10),
	.w3(32'hbbf40866),
	.w4(32'hbc1053a5),
	.w5(32'h3be81297),
	.w6(32'h3b75089b),
	.w7(32'h3b1b94c9),
	.w8(32'h3c803b9d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba128b72),
	.w1(32'h3891f083),
	.w2(32'h3aa0905f),
	.w3(32'hbad62502),
	.w4(32'hbb9f1098),
	.w5(32'hbbb74f1d),
	.w6(32'hbc27a5b7),
	.w7(32'hbc599086),
	.w8(32'h3bd1b8a4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0852cc),
	.w1(32'h3c437dc4),
	.w2(32'hba581777),
	.w3(32'h3c496be4),
	.w4(32'h3b5fe71d),
	.w5(32'h3c3ceeca),
	.w6(32'h3c62f071),
	.w7(32'hbc19404c),
	.w8(32'h3b84ca81),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf07c45),
	.w1(32'hbb1f354a),
	.w2(32'h3a340225),
	.w3(32'h3bdee1e1),
	.w4(32'h3b510401),
	.w5(32'hbaa0cc4c),
	.w6(32'hbb28ba03),
	.w7(32'hbc06d871),
	.w8(32'h3c1a3228),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afa5c0),
	.w1(32'h3bb48311),
	.w2(32'h3b756c03),
	.w3(32'h3a0058dd),
	.w4(32'h3b661a0a),
	.w5(32'hbca11422),
	.w6(32'h3be067a3),
	.w7(32'h3c0aecd9),
	.w8(32'hbb9ce3af),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cd0a1),
	.w1(32'hbbb51329),
	.w2(32'h3a7da361),
	.w3(32'hbc21694d),
	.w4(32'h3bf77cae),
	.w5(32'h39805e1e),
	.w6(32'h3c81cde0),
	.w7(32'h3c6b92c8),
	.w8(32'h3b071a2e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e5899),
	.w1(32'hbc072962),
	.w2(32'hbc01127e),
	.w3(32'hbaa678bc),
	.w4(32'hbaf0352b),
	.w5(32'hb6b98f64),
	.w6(32'h3bf05e21),
	.w7(32'hbb361c60),
	.w8(32'h3b969959),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c0f3a),
	.w1(32'hba904f84),
	.w2(32'h3c417703),
	.w3(32'h3a48dd8e),
	.w4(32'hbbf983f7),
	.w5(32'h3a8902cb),
	.w6(32'hbbf4fd90),
	.w7(32'hbbc491f3),
	.w8(32'h3c81dc01),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf38edc),
	.w1(32'h3bd1bcb2),
	.w2(32'h3a80eced),
	.w3(32'h39efee5c),
	.w4(32'h3c8ca7ef),
	.w5(32'h3c67bfa2),
	.w6(32'h3c55ac12),
	.w7(32'h3bd6ef36),
	.w8(32'h3cb876d4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40c752),
	.w1(32'h3bddd645),
	.w2(32'hbbb49df6),
	.w3(32'h3c33f323),
	.w4(32'h3c133b69),
	.w5(32'h3b329673),
	.w6(32'h3c4c57f2),
	.w7(32'h38c74cc1),
	.w8(32'h3a16b21a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56bc65),
	.w1(32'h3bcec868),
	.w2(32'h3c21b674),
	.w3(32'h3be2490a),
	.w4(32'h3b8c0597),
	.w5(32'h3cb1ff35),
	.w6(32'h3a8a9ae1),
	.w7(32'hbbb3d8df),
	.w8(32'hbb94da4a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbe8c9),
	.w1(32'hbc48a041),
	.w2(32'hbbdbbae8),
	.w3(32'hbc03dd56),
	.w4(32'hbccd1214),
	.w5(32'h3ac53c84),
	.w6(32'hbcc0dae3),
	.w7(32'hbc92da29),
	.w8(32'h3b734373),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e9a43),
	.w1(32'h371848a3),
	.w2(32'hbc5a2bf7),
	.w3(32'h3b6a4c60),
	.w4(32'hb8e713ec),
	.w5(32'hbc7be4e6),
	.w6(32'h3a266c73),
	.w7(32'hbb045e2d),
	.w8(32'h3c2555ed),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64087d),
	.w1(32'h3c55e03e),
	.w2(32'hbafa7af7),
	.w3(32'h3bf4168a),
	.w4(32'h3ade161a),
	.w5(32'hbbaa1f20),
	.w6(32'h3c0326be),
	.w7(32'hbccf907c),
	.w8(32'h3ad39d02),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc008f53),
	.w1(32'hbbab27a6),
	.w2(32'h3bfa24d7),
	.w3(32'h3b333ab1),
	.w4(32'h3c2a18f1),
	.w5(32'hbbf25da3),
	.w6(32'h3ca741c1),
	.w7(32'h3c3ab6bd),
	.w8(32'hbc8cf034),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d3b61),
	.w1(32'hbc918227),
	.w2(32'hbbb0dc8b),
	.w3(32'hbc992dd3),
	.w4(32'h3c10c43b),
	.w5(32'h3b057d4f),
	.w6(32'h3bcc250b),
	.w7(32'h3cd49d0b),
	.w8(32'h3c0949f5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa30d8d),
	.w1(32'hbb624392),
	.w2(32'h3b94555c),
	.w3(32'h3c69af3c),
	.w4(32'h3a1610ad),
	.w5(32'h3c102210),
	.w6(32'h3a085e95),
	.w7(32'h3b84bcd6),
	.w8(32'hbc0041a1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfdf09),
	.w1(32'hbc34e216),
	.w2(32'h3bab896f),
	.w3(32'hbbc0cfb8),
	.w4(32'hbc840615),
	.w5(32'h3c94c99e),
	.w6(32'hbc9594fa),
	.w7(32'hbc43bd71),
	.w8(32'h3b70a53b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c587dfe),
	.w1(32'hbbada6bd),
	.w2(32'h3bef90a0),
	.w3(32'hbaad202b),
	.w4(32'hbc771915),
	.w5(32'h3c020b60),
	.w6(32'hbc7c6b99),
	.w7(32'hbbae96e3),
	.w8(32'h3acfe0da),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af00132),
	.w1(32'hbad9ffb6),
	.w2(32'hbba48068),
	.w3(32'h3ba16b27),
	.w4(32'hbb7daf86),
	.w5(32'h3be6e47b),
	.w6(32'hbb2862e5),
	.w7(32'hbc30b11a),
	.w8(32'h3bc56881),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c548b0c),
	.w1(32'h3bb69ccb),
	.w2(32'h3b7592ea),
	.w3(32'h3c26c84b),
	.w4(32'h3b41bd2e),
	.w5(32'hbc3e2f7f),
	.w6(32'h39908c7f),
	.w7(32'h3ab181f0),
	.w8(32'h3b6076d3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80d2e9),
	.w1(32'hbaabca48),
	.w2(32'hbb82b1e2),
	.w3(32'hbac93be2),
	.w4(32'h3c345819),
	.w5(32'hbc0006e9),
	.w6(32'h3c86a4af),
	.w7(32'hbbeff8d8),
	.w8(32'hbabd6487),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26128e),
	.w1(32'hbaa30687),
	.w2(32'hbc07e0e9),
	.w3(32'hbaf02bf1),
	.w4(32'hbb4919c5),
	.w5(32'hbcab1faa),
	.w6(32'h393d1af3),
	.w7(32'hbb262145),
	.w8(32'h3af4908c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e5c74),
	.w1(32'hba037db7),
	.w2(32'h3b903edc),
	.w3(32'h3ad0aaa7),
	.w4(32'h3c3ab6bd),
	.w5(32'hba75d946),
	.w6(32'h3cb09e52),
	.w7(32'hbb69677f),
	.w8(32'hbc7528d9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b517b3c),
	.w1(32'hbc2f7ebc),
	.w2(32'hbc202804),
	.w3(32'hbca46f88),
	.w4(32'hbc488fec),
	.w5(32'hbc226271),
	.w6(32'hbb8d5121),
	.w7(32'h3b82c923),
	.w8(32'hb8e5c15f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb4e2d),
	.w1(32'hbb82a850),
	.w2(32'hba934769),
	.w3(32'hb9a2d833),
	.w4(32'hbc145b9c),
	.w5(32'h3b19e44b),
	.w6(32'hbb0498be),
	.w7(32'hbc18d544),
	.w8(32'h3b6a1795),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbe954),
	.w1(32'hbb3b559f),
	.w2(32'hbc0464c3),
	.w3(32'h3c18b0d5),
	.w4(32'hba2f8486),
	.w5(32'hbca8b7e0),
	.w6(32'h3a20dcf7),
	.w7(32'hbba5e283),
	.w8(32'h3a73ccba),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1825e0),
	.w1(32'hb9d02978),
	.w2(32'h3bcefabc),
	.w3(32'h3a680c03),
	.w4(32'h3ad88db6),
	.w5(32'hbb94fdf6),
	.w6(32'h3c6663bd),
	.w7(32'hb8dc25af),
	.w8(32'h3c14b027),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a791805),
	.w1(32'h3bfc4196),
	.w2(32'h3b73cddd),
	.w3(32'hbb1af746),
	.w4(32'hbbbfa096),
	.w5(32'h3bc3bb1b),
	.w6(32'h3b988352),
	.w7(32'h3b1ee6f3),
	.w8(32'h3c00c423),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29acb9),
	.w1(32'hb9b978bb),
	.w2(32'hbb87e2a0),
	.w3(32'h3b53686f),
	.w4(32'h3b21a8e6),
	.w5(32'hbad95dfb),
	.w6(32'h3bc957da),
	.w7(32'h3b9efc22),
	.w8(32'h3bad07f6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf0201),
	.w1(32'h3ab9fea3),
	.w2(32'h3b9e0f75),
	.w3(32'hbb938651),
	.w4(32'h38e05794),
	.w5(32'hbb3f4dd2),
	.w6(32'hbc73cea6),
	.w7(32'hbb3ef577),
	.w8(32'h3b0dead7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab27f98),
	.w1(32'h3b5d0aec),
	.w2(32'h39cf2e08),
	.w3(32'hbb03ac45),
	.w4(32'h3b2a5a99),
	.w5(32'h3b8b681b),
	.w6(32'hbbbca43c),
	.w7(32'h3b50b4ec),
	.w8(32'h3a8df57d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff98c9),
	.w1(32'hbbfb3e1b),
	.w2(32'h3b01b9b6),
	.w3(32'h398a3e5d),
	.w4(32'hbc00301c),
	.w5(32'h3bca178e),
	.w6(32'hba7371fa),
	.w7(32'hba98cd2a),
	.w8(32'h3aa7cef1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c040c7f),
	.w1(32'h3c429f08),
	.w2(32'h3c2194aa),
	.w3(32'h3c2f1ecb),
	.w4(32'h3c6f0ad7),
	.w5(32'h3c7600c5),
	.w6(32'h3bea55f5),
	.w7(32'h3c322357),
	.w8(32'hbb8de947),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53e346),
	.w1(32'hbc081f53),
	.w2(32'hbaf4e665),
	.w3(32'hbc80513f),
	.w4(32'hbc866a93),
	.w5(32'h3b563825),
	.w6(32'hbccb50ed),
	.w7(32'h3af4c343),
	.w8(32'h3c0302da),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93db49),
	.w1(32'h3b936f1f),
	.w2(32'h3b98289c),
	.w3(32'h3c21c810),
	.w4(32'h3c209049),
	.w5(32'h3b9bc92d),
	.w6(32'h3c2bddb2),
	.w7(32'h3b4316dd),
	.w8(32'h3c40f10b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbce3a7),
	.w1(32'h3b69e20b),
	.w2(32'hbbc5ea81),
	.w3(32'h3b83ade3),
	.w4(32'h3ae6808a),
	.w5(32'hbb8036c6),
	.w6(32'hbb60951d),
	.w7(32'h3b018957),
	.w8(32'hbbaaee6b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d3f55),
	.w1(32'hbb97e040),
	.w2(32'hba150b8f),
	.w3(32'hbbf4326f),
	.w4(32'hbc0d642d),
	.w5(32'h3b8b3577),
	.w6(32'hbc870ba9),
	.w7(32'hbbd046f1),
	.w8(32'h3b8b92b5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a215231),
	.w1(32'h3ad0a44c),
	.w2(32'hbb256d8f),
	.w3(32'h3b70bc0b),
	.w4(32'h38dca410),
	.w5(32'h3b93aa91),
	.w6(32'hbb03390c),
	.w7(32'hbb3d003a),
	.w8(32'h3be94c5e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa75387),
	.w1(32'h3a33c9bb),
	.w2(32'hb9b70fb4),
	.w3(32'h3c179902),
	.w4(32'hbbed4e53),
	.w5(32'hbaaaa7b4),
	.w6(32'hba82dc8f),
	.w7(32'hbc18034b),
	.w8(32'h3b0db679),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbbbc4),
	.w1(32'hbc8dce10),
	.w2(32'hbb90b2f5),
	.w3(32'hbbd4c6d4),
	.w4(32'hbc2c247b),
	.w5(32'hbc2a0c64),
	.w6(32'h3b9e37b6),
	.w7(32'hbc712299),
	.w8(32'hb91cdde7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e85c7),
	.w1(32'hba9828f5),
	.w2(32'hbae5739f),
	.w3(32'h3bbaa181),
	.w4(32'h3b577ca1),
	.w5(32'h3b8d3fce),
	.w6(32'hbb03f4ab),
	.w7(32'h3c456725),
	.w8(32'h3c2e02de),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7b345),
	.w1(32'h3c17a911),
	.w2(32'h3a3a7dc2),
	.w3(32'h3ce69f27),
	.w4(32'hbb7f3a18),
	.w5(32'h3c20dd10),
	.w6(32'h3bb6ded3),
	.w7(32'hbcb62189),
	.w8(32'hbb2222c2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc487f3),
	.w1(32'hbb25c137),
	.w2(32'h3bf1b014),
	.w3(32'h3c65fd40),
	.w4(32'h3c1d4a1b),
	.w5(32'h3bf32257),
	.w6(32'h3a64bc76),
	.w7(32'hbb8b849c),
	.w8(32'hbb29ddff),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb52bc),
	.w1(32'h3b84c2f6),
	.w2(32'hbb21878c),
	.w3(32'h3b8b2f23),
	.w4(32'hbba785b7),
	.w5(32'hbb9591a8),
	.w6(32'hbb2319e6),
	.w7(32'hb9131eae),
	.w8(32'hbb7639a7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe4fda),
	.w1(32'hbbf894eb),
	.w2(32'h3b822c4d),
	.w3(32'hbbed9ed9),
	.w4(32'hbbe379c8),
	.w5(32'h3b89871d),
	.w6(32'hbc05e631),
	.w7(32'hbbb728a9),
	.w8(32'h3a326c95),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda4358),
	.w1(32'hbc07b9f1),
	.w2(32'hbb7b68ac),
	.w3(32'hbc3f0b5f),
	.w4(32'hbc26f643),
	.w5(32'h3c229ce7),
	.w6(32'hbc0146db),
	.w7(32'hbb140b43),
	.w8(32'h3af9b942),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba65491),
	.w1(32'hb9131c9e),
	.w2(32'h3a47b249),
	.w3(32'hba0705ef),
	.w4(32'hbb2bac45),
	.w5(32'h3b97cb94),
	.w6(32'h3a44797f),
	.w7(32'hbaf1e032),
	.w8(32'h3be07f57),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4252d),
	.w1(32'h3c184ba0),
	.w2(32'hbba3e387),
	.w3(32'h3bca95e1),
	.w4(32'hb8cb3b4d),
	.w5(32'h3af4a5bf),
	.w6(32'h3c60a0a6),
	.w7(32'h3b7fc232),
	.w8(32'h3c80ec6d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46eca4),
	.w1(32'hbaff7ae2),
	.w2(32'hbae0e903),
	.w3(32'h3bbe2c04),
	.w4(32'hbc499710),
	.w5(32'hb9debe06),
	.w6(32'hbb87b28f),
	.w7(32'hbc12998f),
	.w8(32'h3c193585),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb382dc1),
	.w1(32'h3bec51c8),
	.w2(32'hbb5fbf96),
	.w3(32'h3c2e039f),
	.w4(32'h3c38cffc),
	.w5(32'hbb54d0c1),
	.w6(32'h3c3d9020),
	.w7(32'h3b85cebb),
	.w8(32'hbb5b4504),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89a389),
	.w1(32'hbb55a9d5),
	.w2(32'h3ac625b4),
	.w3(32'hbad6d3c2),
	.w4(32'hbb3cf277),
	.w5(32'hbc122b49),
	.w6(32'hbb454fd8),
	.w7(32'hbbc73888),
	.w8(32'hbaaee092),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ef6b2),
	.w1(32'h3a8fead1),
	.w2(32'h3b5582d2),
	.w3(32'h3c54c19c),
	.w4(32'h3b875f25),
	.w5(32'h3cc55a0a),
	.w6(32'h3bbc6004),
	.w7(32'h3c40406c),
	.w8(32'h3b1fe74f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1364a),
	.w1(32'hb9eabebe),
	.w2(32'hbba7ae1c),
	.w3(32'h3b18ac11),
	.w4(32'hbcd0e5b1),
	.w5(32'h3c0bc117),
	.w6(32'hbd27d37f),
	.w7(32'hbcb20cb6),
	.w8(32'h3bfd2deb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c9098),
	.w1(32'hb9673db0),
	.w2(32'h3c6c9856),
	.w3(32'hbb41b276),
	.w4(32'hbc129025),
	.w5(32'hbb3860b1),
	.w6(32'hbc5d5c95),
	.w7(32'h3ac34a04),
	.w8(32'hbc2d79ed),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adeacd7),
	.w1(32'hba88a976),
	.w2(32'h3be73b63),
	.w3(32'hbc06f0fc),
	.w4(32'h3bdd54e9),
	.w5(32'h3bf391ec),
	.w6(32'h3bdd05fb),
	.w7(32'h3c32f0db),
	.w8(32'h3c2a0a96),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01a9f3),
	.w1(32'h3b97fda4),
	.w2(32'h3b0a1184),
	.w3(32'h3bab67f9),
	.w4(32'h3b7f8131),
	.w5(32'hb99d7c96),
	.w6(32'h3b779a99),
	.w7(32'h3aaae4cf),
	.w8(32'hbaeefccc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e2fb5),
	.w1(32'h3a9d916e),
	.w2(32'h3b0c0e8a),
	.w3(32'h3981d6e8),
	.w4(32'h3c177981),
	.w5(32'h3b32f844),
	.w6(32'h3b4ec5f1),
	.w7(32'h3c27b143),
	.w8(32'h3b8d9189),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb252a50),
	.w1(32'hba91e119),
	.w2(32'hbb33faa9),
	.w3(32'hbb3d115a),
	.w4(32'hba99e37b),
	.w5(32'hbc9c9ba2),
	.w6(32'hbb808cb2),
	.w7(32'h3b338e9b),
	.w8(32'hbc36c57f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc845cbf),
	.w1(32'h3ba39e96),
	.w2(32'hbc4c1543),
	.w3(32'hbc843bd8),
	.w4(32'h3b6067a6),
	.w5(32'h3c242090),
	.w6(32'h3b0ce608),
	.w7(32'h3b080609),
	.w8(32'h3b0bdd19),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cee38),
	.w1(32'hbb26fcff),
	.w2(32'hbb68cbae),
	.w3(32'h3bbaf0c8),
	.w4(32'hbc3c475b),
	.w5(32'hba5bbd08),
	.w6(32'hbc6aa2fb),
	.w7(32'hbc1ae79f),
	.w8(32'h3a6cff01),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398176b7),
	.w1(32'hbc473701),
	.w2(32'h3a5f5603),
	.w3(32'h3c25c899),
	.w4(32'hba988938),
	.w5(32'h3c98f01f),
	.w6(32'hbbadd807),
	.w7(32'hbc4a9e68),
	.w8(32'h3be20d44),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84e709),
	.w1(32'h3b6671b7),
	.w2(32'h3a0e3d36),
	.w3(32'h3cd73400),
	.w4(32'h3d29fa15),
	.w5(32'h3c4f221a),
	.w6(32'h3d00fdbf),
	.w7(32'h3af2efd0),
	.w8(32'h3b3201ed),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21c111),
	.w1(32'hbc747678),
	.w2(32'hbc1bfda4),
	.w3(32'h3b68d05b),
	.w4(32'hbc927e01),
	.w5(32'h3abae8da),
	.w6(32'hbc7610de),
	.w7(32'hbb59b134),
	.w8(32'h3b2c95c9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e604d),
	.w1(32'h3bccf058),
	.w2(32'hbbd7734a),
	.w3(32'h3b6f8245),
	.w4(32'hbb31a10c),
	.w5(32'hbaf9a8b6),
	.w6(32'hbb283ba4),
	.w7(32'hbc05e111),
	.w8(32'hbc043b29),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafef41),
	.w1(32'hbc070e93),
	.w2(32'hbc22958e),
	.w3(32'hbb8d4c78),
	.w4(32'hbb573f65),
	.w5(32'hbc4b0e33),
	.w6(32'hbb92ecda),
	.w7(32'h3bd428a5),
	.w8(32'h3b8a583e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95f993),
	.w1(32'hbb2f5b9a),
	.w2(32'hba2cb4d0),
	.w3(32'h3b875e7a),
	.w4(32'h3c3730a6),
	.w5(32'h3af6a0ac),
	.w6(32'h3c143ca6),
	.w7(32'hbbf0cd8b),
	.w8(32'h3965178b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb698051),
	.w1(32'hbc163748),
	.w2(32'hbc06d020),
	.w3(32'hbc443a7c),
	.w4(32'hbcb64804),
	.w5(32'h3bcc5b14),
	.w6(32'hbca771b1),
	.w7(32'hbc02c200),
	.w8(32'hbb0d6b3c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0388d6),
	.w1(32'hbc970e6e),
	.w2(32'hbcdeda1d),
	.w3(32'h3c1d3b01),
	.w4(32'hbbd09ade),
	.w5(32'hbc7203cc),
	.w6(32'h3b3b8301),
	.w7(32'hbb9f6897),
	.w8(32'hbb188cad),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbead075),
	.w1(32'hba7cf228),
	.w2(32'hbc579035),
	.w3(32'h3a3c366d),
	.w4(32'h3b9f3cc6),
	.w5(32'hbc330073),
	.w6(32'h3bb89421),
	.w7(32'hbba3af54),
	.w8(32'hbaee5945),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe70816),
	.w1(32'hbb731cb3),
	.w2(32'h37d8d52b),
	.w3(32'h39bd7ed8),
	.w4(32'hbae7e40f),
	.w5(32'h3b64263c),
	.w6(32'h3b5748a9),
	.w7(32'hbc095ddd),
	.w8(32'hbc53f6c2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc870d),
	.w1(32'h3c332b60),
	.w2(32'h3af814be),
	.w3(32'h3c48f31d),
	.w4(32'h3c5a3063),
	.w5(32'h3c7ef99a),
	.w6(32'hbbd8bc85),
	.w7(32'h3b5653d3),
	.w8(32'h3c56affa),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b5a83),
	.w1(32'h3b49e675),
	.w2(32'hbc60f33b),
	.w3(32'h3bf9e012),
	.w4(32'hbbfff752),
	.w5(32'h3ba798bf),
	.w6(32'hbba96bca),
	.w7(32'hbb8b6fd3),
	.w8(32'hbb8fc534),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c47c0),
	.w1(32'hbb80924e),
	.w2(32'hbacacdee),
	.w3(32'h3beb4a04),
	.w4(32'hb9a9b2c8),
	.w5(32'h3b42e393),
	.w6(32'hbc1189b9),
	.w7(32'hbc849e5c),
	.w8(32'h3aa7063d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd273b),
	.w1(32'hbb1dc0eb),
	.w2(32'hbbc0e316),
	.w3(32'hbb51bf63),
	.w4(32'hbc7299f9),
	.w5(32'h3bf9e061),
	.w6(32'hbc36ce08),
	.w7(32'hbc15e923),
	.w8(32'hbbd80ed8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f1a1b),
	.w1(32'hbc2008e1),
	.w2(32'hbc41fc4f),
	.w3(32'hbbb66314),
	.w4(32'hbc7e5f6a),
	.w5(32'hbc5a4968),
	.w6(32'hbc609e77),
	.w7(32'hbbd70f67),
	.w8(32'h3c3ba503),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3124d9),
	.w1(32'h3b92700f),
	.w2(32'hbbfbd9d5),
	.w3(32'h3c03cb3b),
	.w4(32'h3c144634),
	.w5(32'h39b8e255),
	.w6(32'h3c2914fe),
	.w7(32'hba07ee76),
	.w8(32'h3c73f713),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc11d18),
	.w1(32'hbaeeb6e0),
	.w2(32'h3ca46c80),
	.w3(32'h3c814008),
	.w4(32'h3c7900f5),
	.w5(32'hbca4c4f9),
	.w6(32'h3c0a6c50),
	.w7(32'hbbfc3613),
	.w8(32'hbc88c7a8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f759f),
	.w1(32'hbc229382),
	.w2(32'h39d2f9dc),
	.w3(32'hbcd6d97a),
	.w4(32'h3cf71be4),
	.w5(32'hbb5a3cf4),
	.w6(32'h3cc36328),
	.w7(32'h3cb35b8b),
	.w8(32'hbb47eaf2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7e8e4),
	.w1(32'h3c0077b7),
	.w2(32'h3c83d176),
	.w3(32'h3ba2662d),
	.w4(32'h3c2d1849),
	.w5(32'h3cb191c1),
	.w6(32'h3bfcee25),
	.w7(32'h3bd3dcd7),
	.w8(32'hbb00bc7f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c686b90),
	.w1(32'hbbba7297),
	.w2(32'hbb4f79ce),
	.w3(32'hbb243b9b),
	.w4(32'hbc182fd1),
	.w5(32'hbb9ab6d0),
	.w6(32'hbc6731db),
	.w7(32'h3becda25),
	.w8(32'h3a06b102),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7acb),
	.w1(32'h3a46242e),
	.w2(32'hbb4025a1),
	.w3(32'h3baae90a),
	.w4(32'h3c0231cb),
	.w5(32'hbb1869bc),
	.w6(32'h3c69ee5c),
	.w7(32'h3b9c30a5),
	.w8(32'h3c3f8222),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2babac),
	.w1(32'h3b7e1367),
	.w2(32'h3b31a8e7),
	.w3(32'h3c2672c0),
	.w4(32'h3bf97d51),
	.w5(32'hbb4fb7c6),
	.w6(32'h3a608282),
	.w7(32'hbbee35c5),
	.w8(32'h3bb13959),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b7cac),
	.w1(32'h3b377282),
	.w2(32'h3aa58f86),
	.w3(32'h3a86391a),
	.w4(32'h3ba648e7),
	.w5(32'h3c4cbbfc),
	.w6(32'hbac40737),
	.w7(32'h3b6b7ff5),
	.w8(32'h3b834fec),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a09730),
	.w1(32'h3be3a48e),
	.w2(32'hb8bd7daa),
	.w3(32'h3c452770),
	.w4(32'h3bff5493),
	.w5(32'hba7782ad),
	.w6(32'h3baf1bdb),
	.w7(32'hbc04a1bd),
	.w8(32'hba43765c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdae33),
	.w1(32'hbb7bc687),
	.w2(32'h3b577401),
	.w3(32'hba62101f),
	.w4(32'hbb5bc28a),
	.w5(32'hba4af955),
	.w6(32'hbab67107),
	.w7(32'hbb858a66),
	.w8(32'h3b4be3a8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b153f94),
	.w1(32'h3bad77b4),
	.w2(32'hbc071356),
	.w3(32'h3b04a8d2),
	.w4(32'h3bba22e7),
	.w5(32'hbce5a90a),
	.w6(32'h3b3dfa81),
	.w7(32'h3b4987f7),
	.w8(32'h3c8f989f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ebfb1),
	.w1(32'hba54e3c6),
	.w2(32'hbbff4926),
	.w3(32'h3c6a1364),
	.w4(32'h3cf2c5d7),
	.w5(32'hbba1f552),
	.w6(32'h3d68a739),
	.w7(32'hbb7cb1b2),
	.w8(32'h3ab911d0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9de98),
	.w1(32'hbb600b56),
	.w2(32'hbc8a5014),
	.w3(32'h3b27fef6),
	.w4(32'hba91a503),
	.w5(32'h3bf861db),
	.w6(32'h3b33f75d),
	.w7(32'hbbd0d985),
	.w8(32'h3c6597ae),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfbdb8),
	.w1(32'h3bf6485f),
	.w2(32'hbbf07da5),
	.w3(32'h3cb507fe),
	.w4(32'h3cc0dde7),
	.w5(32'hbc828542),
	.w6(32'h3cbb3c1a),
	.w7(32'hbc3dd8db),
	.w8(32'hbc7d0154),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd527ce),
	.w1(32'h3b394be8),
	.w2(32'h3c04cf11),
	.w3(32'hbb846c04),
	.w4(32'h3a85aa08),
	.w5(32'hbb24c886),
	.w6(32'hbbc0c45c),
	.w7(32'h3b094918),
	.w8(32'hbb692f77),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7b670),
	.w1(32'h3948898c),
	.w2(32'h3c019009),
	.w3(32'h39485f46),
	.w4(32'hbc88285c),
	.w5(32'h3a833d2a),
	.w6(32'hbb831523),
	.w7(32'hbb05a769),
	.w8(32'hbb8b5c4b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34e495),
	.w1(32'hbca455e7),
	.w2(32'h3c01028d),
	.w3(32'hbc41dc41),
	.w4(32'hbbb7fa2f),
	.w5(32'h3b8ec1a2),
	.w6(32'hbb2fd0c9),
	.w7(32'h3a1835ca),
	.w8(32'h3c799430),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27e4a9),
	.w1(32'h3c55e561),
	.w2(32'h3c281c91),
	.w3(32'h3c898308),
	.w4(32'h3ab40508),
	.w5(32'h3b31d3d3),
	.w6(32'hb74cd651),
	.w7(32'hbc62ea96),
	.w8(32'hbb4b1642),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb545ea9),
	.w1(32'hbb3e7755),
	.w2(32'hbb8e0f71),
	.w3(32'hbc147353),
	.w4(32'h3b248be4),
	.w5(32'h3c33f04c),
	.w6(32'h3be6eee4),
	.w7(32'h3c62a758),
	.w8(32'h3beec5d2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877f97),
	.w1(32'h3b0a6db5),
	.w2(32'hbb949c35),
	.w3(32'h3b8fd3fb),
	.w4(32'h3b7920fc),
	.w5(32'h3cd29450),
	.w6(32'h3c0c703c),
	.w7(32'hbaaacd8f),
	.w8(32'hba1f8a18),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccdffe),
	.w1(32'hba057b11),
	.w2(32'h3bba8187),
	.w3(32'h3c196764),
	.w4(32'hbccdc6ae),
	.w5(32'h3bc575bf),
	.w6(32'hbcf727e5),
	.w7(32'hbb8a000b),
	.w8(32'h3bf6bd64),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cd267),
	.w1(32'h3c05d1d8),
	.w2(32'h3ad4c65f),
	.w3(32'hba4dcef8),
	.w4(32'h3afda7cb),
	.w5(32'h3b049e1b),
	.w6(32'hbaf834bb),
	.w7(32'h3c466a1e),
	.w8(32'h3b582241),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf441e),
	.w1(32'hbc10191f),
	.w2(32'hbc952e5d),
	.w3(32'hbb980713),
	.w4(32'hbaf95795),
	.w5(32'hbc6857be),
	.w6(32'hbbdb763a),
	.w7(32'hbbff1962),
	.w8(32'hbbef720f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3582b),
	.w1(32'hbbbc7e04),
	.w2(32'h3b31e7cd),
	.w3(32'h3bc81273),
	.w4(32'h3bc8db8a),
	.w5(32'h3c87e9c4),
	.w6(32'h3c1a3fdf),
	.w7(32'hbc4f11bf),
	.w8(32'h3bc85ada),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db1b9b),
	.w1(32'hbbbc0abd),
	.w2(32'h3c6ff4db),
	.w3(32'h3c1b6355),
	.w4(32'hbc2b4e72),
	.w5(32'h3c971b47),
	.w6(32'hbb71bff5),
	.w7(32'hbc5e7953),
	.w8(32'h3c3b8783),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cc89c),
	.w1(32'h3ba207cf),
	.w2(32'h3c115173),
	.w3(32'h3b8dedad),
	.w4(32'h3b07ce52),
	.w5(32'h3b8037e5),
	.w6(32'h3b3cde9e),
	.w7(32'h3b66ee75),
	.w8(32'h382dbc7e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e3fb5),
	.w1(32'h38e5614a),
	.w2(32'h3b923990),
	.w3(32'hbb961462),
	.w4(32'h3b287395),
	.w5(32'h3c1e8a7f),
	.w6(32'hba2fe6a4),
	.w7(32'h3bf4a8f4),
	.w8(32'h3c5ba87e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c223e16),
	.w1(32'h3c1d3e94),
	.w2(32'hba287483),
	.w3(32'h3bc9332c),
	.w4(32'h3bf496ce),
	.w5(32'hb88ac94d),
	.w6(32'h3b6edc69),
	.w7(32'h3b835cd8),
	.w8(32'hbafb5a6b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f362b),
	.w1(32'hbae9d56f),
	.w2(32'h3c41409b),
	.w3(32'hbaaa5c10),
	.w4(32'h39a12cf8),
	.w5(32'h3be57b52),
	.w6(32'hb773dec1),
	.w7(32'hbaae8cd6),
	.w8(32'h3c5468a2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ac4a3),
	.w1(32'h3c167aee),
	.w2(32'h3b9a524f),
	.w3(32'h3c4ce043),
	.w4(32'h3c60f814),
	.w5(32'hbc2ff84f),
	.w6(32'h3c27d354),
	.w7(32'h3c5b47d9),
	.w8(32'hbc54641d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ffef9),
	.w1(32'hbc8469f8),
	.w2(32'h3ae25653),
	.w3(32'hbc9c036d),
	.w4(32'hbc1bee44),
	.w5(32'hba0f682f),
	.w6(32'hbb1f75b2),
	.w7(32'h3c8299be),
	.w8(32'hbae84ca0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47de02),
	.w1(32'h3c141fc6),
	.w2(32'h3bb6e75f),
	.w3(32'h3bafa867),
	.w4(32'h3c0c0bb1),
	.w5(32'h3a276d49),
	.w6(32'h3bf09a63),
	.w7(32'h3c28e51a),
	.w8(32'hbb33fa91),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bd67b),
	.w1(32'hba9d1369),
	.w2(32'h3b63b110),
	.w3(32'hbb52443e),
	.w4(32'h3ba1502b),
	.w5(32'h3b99b21c),
	.w6(32'h3b4972d3),
	.w7(32'h3c0d7e8b),
	.w8(32'hbbb691a4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9c138),
	.w1(32'h3b5c886a),
	.w2(32'h3c3967dd),
	.w3(32'hb9eb6546),
	.w4(32'hbb5f308e),
	.w5(32'h3c080127),
	.w6(32'hbc942c18),
	.w7(32'hbc0dcbe2),
	.w8(32'h3bea64b6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc80e39),
	.w1(32'h3c3c6440),
	.w2(32'hbc23babb),
	.w3(32'h3c1d0804),
	.w4(32'h3c01c4b0),
	.w5(32'h3b0ffc98),
	.w6(32'h3c1e0f52),
	.w7(32'h3bca8fc8),
	.w8(32'hbb855ded),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad6a67),
	.w1(32'h37b52eb5),
	.w2(32'h3be67aed),
	.w3(32'h3b65140e),
	.w4(32'hbc085a21),
	.w5(32'h3c481d45),
	.w6(32'hbc4e2d92),
	.w7(32'hbc7a40a1),
	.w8(32'h3b12620e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeca058),
	.w1(32'hbbcfdfb6),
	.w2(32'hbc1efe8a),
	.w3(32'hbb84eff4),
	.w4(32'hbc437258),
	.w5(32'h38f86458),
	.w6(32'hbc3238f9),
	.w7(32'hbbb2dbcc),
	.w8(32'h3a499c6a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba07a41),
	.w1(32'hbb1a3a06),
	.w2(32'hbb6e0dc0),
	.w3(32'h3b000044),
	.w4(32'hbc18144a),
	.w5(32'h3a232630),
	.w6(32'hbc880b8e),
	.w7(32'hbc60ea4b),
	.w8(32'h3ba95224),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f7e14),
	.w1(32'h3b902e7a),
	.w2(32'h3aead42e),
	.w3(32'h3b5af503),
	.w4(32'hbbd6b057),
	.w5(32'hbac8fec3),
	.w6(32'hbc122283),
	.w7(32'hbc4a7774),
	.w8(32'hbb1a0fcf),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad87bf7),
	.w1(32'hbbd10241),
	.w2(32'h3c43acff),
	.w3(32'hbb9b3529),
	.w4(32'hbc034205),
	.w5(32'h3bb3cc07),
	.w6(32'hbbd2f32e),
	.w7(32'hbbe28c05),
	.w8(32'h3c08d140),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00d4e8),
	.w1(32'h3bd78397),
	.w2(32'hb90f043d),
	.w3(32'h3aed897c),
	.w4(32'h3b4c26a2),
	.w5(32'h3bd776f9),
	.w6(32'h3b3d9172),
	.w7(32'h3c484fab),
	.w8(32'hbb45865f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b845ba1),
	.w1(32'h3c0ae597),
	.w2(32'hbb35ab0e),
	.w3(32'h3c16e11f),
	.w4(32'hbba2277b),
	.w5(32'hbbef87b9),
	.w6(32'hbb8c3ca5),
	.w7(32'hbc1bf23f),
	.w8(32'h3ac671fc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafc619),
	.w1(32'hbbab35d0),
	.w2(32'hba32bae3),
	.w3(32'hbb1a48ef),
	.w4(32'hba0beabc),
	.w5(32'hbadd76ea),
	.w6(32'hbb9685aa),
	.w7(32'h3b7d40a5),
	.w8(32'h3aa854bc),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaa174),
	.w1(32'hba4d2ba7),
	.w2(32'hbce9d547),
	.w3(32'hbb89e7e4),
	.w4(32'h39597960),
	.w5(32'hbd3dff3f),
	.w6(32'hbb2e6bdc),
	.w7(32'h3a72edab),
	.w8(32'hbcba455e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcccad36),
	.w1(32'hbb9e597b),
	.w2(32'hbb30c1ca),
	.w3(32'hbca64556),
	.w4(32'h3c2c0083),
	.w5(32'hba0cbe4e),
	.w6(32'hba6a2699),
	.w7(32'h3cb19ad9),
	.w8(32'h3a270be5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84acf8),
	.w1(32'h39f47217),
	.w2(32'hb9e3ffa3),
	.w3(32'hbc3630cb),
	.w4(32'hb991ef58),
	.w5(32'h3b9d7ff5),
	.w6(32'hbb37b358),
	.w7(32'hbb58496e),
	.w8(32'h3adcb873),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15ca59),
	.w1(32'hbac58021),
	.w2(32'h3c52e9e0),
	.w3(32'hb983c25e),
	.w4(32'h3ac7531a),
	.w5(32'h3cc143e3),
	.w6(32'h3b01c498),
	.w7(32'h3ae28649),
	.w8(32'h3be89be7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b744bfa),
	.w1(32'hbbc2d729),
	.w2(32'h3ba85085),
	.w3(32'h3b407a62),
	.w4(32'hbc0ed870),
	.w5(32'h3c85c8da),
	.w6(32'h3b65e11e),
	.w7(32'hbbf30c91),
	.w8(32'h3c2bad1a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49611d),
	.w1(32'h3bdc3f0c),
	.w2(32'hbbdcc747),
	.w3(32'h3be453db),
	.w4(32'hbbec4729),
	.w5(32'hbc2c07fe),
	.w6(32'h3b6adccf),
	.w7(32'hbc246b03),
	.w8(32'hbacd0d2c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919310),
	.w1(32'h3b9e19de),
	.w2(32'h3cd4c7e0),
	.w3(32'hb9ae578f),
	.w4(32'h3c1da2c5),
	.w5(32'h3cab0d81),
	.w6(32'h3b083753),
	.w7(32'h3ba10df4),
	.w8(32'hbb724f10),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfa137),
	.w1(32'hbc86d527),
	.w2(32'h3a6d5395),
	.w3(32'hbcb31a51),
	.w4(32'hbcb4ecc4),
	.w5(32'hba5306d1),
	.w6(32'hbccb8ad6),
	.w7(32'hbc9d9a82),
	.w8(32'hba78275d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1be4f),
	.w1(32'h3a221b35),
	.w2(32'hbadbe34b),
	.w3(32'h3857ac0e),
	.w4(32'hbaa59675),
	.w5(32'hbc136b86),
	.w6(32'hbb996d1a),
	.w7(32'hbbed14e3),
	.w8(32'hb9831a64),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6dc42),
	.w1(32'hbc0f90cb),
	.w2(32'hbc8619a1),
	.w3(32'hbccb1956),
	.w4(32'hbc9e3bc5),
	.w5(32'hbc6e81d3),
	.w6(32'hbb95c296),
	.w7(32'hbc8bcee1),
	.w8(32'hba787656),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6d52b),
	.w1(32'h3c260f1c),
	.w2(32'hbb99051e),
	.w3(32'h3bb3d982),
	.w4(32'h3c793101),
	.w5(32'hbc0f08ae),
	.w6(32'h3c22e0bc),
	.w7(32'h3c60be63),
	.w8(32'hbbffcb71),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb45924),
	.w1(32'hbc58207c),
	.w2(32'hb887e7a3),
	.w3(32'hbcaa451a),
	.w4(32'hbc41dd97),
	.w5(32'h3c0710d4),
	.w6(32'hbc5cae58),
	.w7(32'hbc89a2bf),
	.w8(32'hbaf9d530),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0da07f),
	.w1(32'h3bc7b7f5),
	.w2(32'h3a8c19aa),
	.w3(32'h3c187c2d),
	.w4(32'h3c482dd7),
	.w5(32'h3be00647),
	.w6(32'hba420e41),
	.w7(32'hba4bb663),
	.w8(32'h3bd6c954),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad22b54),
	.w1(32'h3b801cd2),
	.w2(32'h3c0817b3),
	.w3(32'hbb095a29),
	.w4(32'hba3a772c),
	.w5(32'hbab6325a),
	.w6(32'hbb41b141),
	.w7(32'h3b50e710),
	.w8(32'h3bf5ce0f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b771eae),
	.w1(32'h3b4a1488),
	.w2(32'h3c252902),
	.w3(32'hbc2f40a0),
	.w4(32'hbc3255b1),
	.w5(32'h3be78555),
	.w6(32'hbbafe8b3),
	.w7(32'hbb1e1fd1),
	.w8(32'h3bb8e9cb),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f9e3d),
	.w1(32'hba5a4173),
	.w2(32'hbbc4c988),
	.w3(32'h3b80879a),
	.w4(32'hb96b4cb3),
	.w5(32'hbb2227eb),
	.w6(32'h3b1d08af),
	.w7(32'hbbc30715),
	.w8(32'h3bbb9175),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ed25d),
	.w1(32'hbb97a955),
	.w2(32'hbb918f77),
	.w3(32'h3a9fb6e4),
	.w4(32'hbb26d7f5),
	.w5(32'hba6ee98f),
	.w6(32'h3b144106),
	.w7(32'h3a5432eb),
	.w8(32'hbb0f8e68),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ba597),
	.w1(32'h3b346ed2),
	.w2(32'hb9e74ae9),
	.w3(32'hba1cd547),
	.w4(32'h3c66dcd6),
	.w5(32'hbb620a3c),
	.w6(32'h3a1ce180),
	.w7(32'h3cc666d3),
	.w8(32'hbbb2744b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6ce6d),
	.w1(32'hbc0746a7),
	.w2(32'h3b95c248),
	.w3(32'hbb5bcfd5),
	.w4(32'h3ba89ab9),
	.w5(32'h3b248b25),
	.w6(32'hbaadd865),
	.w7(32'h3c19c2cd),
	.w8(32'h3912098a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace6077),
	.w1(32'h39cce2f9),
	.w2(32'h3cfb15e8),
	.w3(32'hba406db6),
	.w4(32'hbb31ef59),
	.w5(32'h3c979074),
	.w6(32'h3a7e0dae),
	.w7(32'h3a75b00b),
	.w8(32'hbb92720b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ef861),
	.w1(32'hba881c2b),
	.w2(32'h3bab3594),
	.w3(32'hbbee8327),
	.w4(32'hbc2bc1d7),
	.w5(32'h3b0b7d0b),
	.w6(32'hbd051210),
	.w7(32'hbc7c952c),
	.w8(32'h3b58b796),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf31c28),
	.w1(32'h3b9b78eb),
	.w2(32'h3bdfaeb4),
	.w3(32'h3b02d5c9),
	.w4(32'hbaa7bc79),
	.w5(32'h3c63d617),
	.w6(32'hbb0f79a6),
	.w7(32'hbb5fde26),
	.w8(32'h3bf82632),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81f507),
	.w1(32'h3ba37ba1),
	.w2(32'h3ad48014),
	.w3(32'h3c69b0cd),
	.w4(32'h3c876c01),
	.w5(32'h3bbe4e15),
	.w6(32'h3c2a87c1),
	.w7(32'h3c1cd11d),
	.w8(32'hbbdce587),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4be09),
	.w1(32'hbc4e460e),
	.w2(32'hba9751bb),
	.w3(32'hbb96bb5f),
	.w4(32'hbc2807ba),
	.w5(32'hbc3d896a),
	.w6(32'hbc5268fd),
	.w7(32'hbbb2ac7b),
	.w8(32'hbc764f3d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c9cd3),
	.w1(32'hbc6bd8f9),
	.w2(32'h3afccd66),
	.w3(32'hbd34bab4),
	.w4(32'hbd087a40),
	.w5(32'h3a46f50b),
	.w6(32'hbd11cb97),
	.w7(32'hbca60830),
	.w8(32'h3a34a5d8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ad97),
	.w1(32'hbb1a9240),
	.w2(32'h3c4412c7),
	.w3(32'h3ad655bf),
	.w4(32'h3b2ab071),
	.w5(32'h3c64edf7),
	.w6(32'h3a6041e9),
	.w7(32'h3c400781),
	.w8(32'h3c14800e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5617d),
	.w1(32'hbbcc2b8f),
	.w2(32'h3c11b4a3),
	.w3(32'hba5acbd1),
	.w4(32'hbc30971e),
	.w5(32'h3c368964),
	.w6(32'hbbaaeba2),
	.w7(32'hbbfb2261),
	.w8(32'h3c2459fb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f63c7),
	.w1(32'hba95a29a),
	.w2(32'h3c1c4922),
	.w3(32'h3c686300),
	.w4(32'h3c04925c),
	.w5(32'h3cc3ea7f),
	.w6(32'hba6f19f1),
	.w7(32'h3a7294cc),
	.w8(32'h3c1754be),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60ff90),
	.w1(32'hb9ba9ea0),
	.w2(32'h3ba88bd4),
	.w3(32'h3c1fb5dc),
	.w4(32'hbc1c9f4f),
	.w5(32'hbbfce3a7),
	.w6(32'h39488cb2),
	.w7(32'hbc3437f6),
	.w8(32'hbbd746e1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2f2b2),
	.w1(32'h39d1074f),
	.w2(32'h3be761e6),
	.w3(32'h3a8ee336),
	.w4(32'h3c154b3a),
	.w5(32'h3b78eb2b),
	.w6(32'h3b6ef17e),
	.w7(32'h3bd7bdf4),
	.w8(32'h3ba6867a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb208916),
	.w1(32'hbb657de7),
	.w2(32'hbb0e8947),
	.w3(32'hbc0e6129),
	.w4(32'hbae125a3),
	.w5(32'hbae3be39),
	.w6(32'h3b5043d6),
	.w7(32'h3b29797b),
	.w8(32'h3bbc61c4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe20eb0),
	.w1(32'h3c174e2e),
	.w2(32'h3bd0ffde),
	.w3(32'hbba540d8),
	.w4(32'h3bc20fa0),
	.w5(32'hbc43757f),
	.w6(32'hbb966fe4),
	.w7(32'h3bf8e7c6),
	.w8(32'hbc4a4294),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13ae99),
	.w1(32'hba6263e5),
	.w2(32'h3c8912cb),
	.w3(32'hbc47fb82),
	.w4(32'hbbbab5fb),
	.w5(32'h3cbc95df),
	.w6(32'hbb939bd0),
	.w7(32'hba3db1c2),
	.w8(32'h3bec27ae),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2ed93),
	.w1(32'h3c04c951),
	.w2(32'hbb9ed659),
	.w3(32'h3a2f8ce2),
	.w4(32'h3b955cac),
	.w5(32'h3c090e7a),
	.w6(32'hbc1a0932),
	.w7(32'h3c546970),
	.w8(32'h3b8ceacd),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda7015),
	.w1(32'hb93708e2),
	.w2(32'hbc20c952),
	.w3(32'h3ba9c90b),
	.w4(32'h3c1f5eee),
	.w5(32'hbc47f75a),
	.w6(32'h3c5ba543),
	.w7(32'hbb17d07b),
	.w8(32'hbc1a0060),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39ada),
	.w1(32'hbbc70bb3),
	.w2(32'hbc539e13),
	.w3(32'hbc6bf76d),
	.w4(32'h396a7143),
	.w5(32'hbcecdc25),
	.w6(32'hbbdc5736),
	.w7(32'hbc04dc6d),
	.w8(32'h3b819227),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc664a7d),
	.w1(32'h3b098527),
	.w2(32'h3bcb1661),
	.w3(32'hbc6d2efe),
	.w4(32'h3bd8153d),
	.w5(32'h3b196b92),
	.w6(32'h3c350e66),
	.w7(32'h3cb4b383),
	.w8(32'h3b2d8719),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ed5a8),
	.w1(32'hb83ef852),
	.w2(32'hbbabaf86),
	.w3(32'hbb6ac293),
	.w4(32'hbb1c2c6e),
	.w5(32'hbac4f7d6),
	.w6(32'h3b8cda65),
	.w7(32'hbb70b20f),
	.w8(32'h3b83130e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4755ce),
	.w1(32'hbb049241),
	.w2(32'hbc91e89c),
	.w3(32'hba83cde7),
	.w4(32'h3ae3a7cc),
	.w5(32'hbc0fc42c),
	.w6(32'h3bb5d040),
	.w7(32'h3b9ebfe0),
	.w8(32'h3c0f27de),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1049a9),
	.w1(32'hbb5a6b31),
	.w2(32'h3ba9caa2),
	.w3(32'h3bf76db1),
	.w4(32'h3c2475e2),
	.w5(32'hbafee276),
	.w6(32'h3c84e918),
	.w7(32'h3c62155f),
	.w8(32'h3b61d470),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb136f31),
	.w1(32'hbba35272),
	.w2(32'h3bb3732e),
	.w3(32'hbbbc9665),
	.w4(32'h3ac5b9ce),
	.w5(32'h3b8b3998),
	.w6(32'hbb6cf002),
	.w7(32'h3bbc6d6d),
	.w8(32'hbb9a6fdf),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f4605),
	.w1(32'hba8025f8),
	.w2(32'h3b274410),
	.w3(32'h3b9307d3),
	.w4(32'h3b855088),
	.w5(32'h3b912a5a),
	.w6(32'h3a4ac934),
	.w7(32'h3b93092a),
	.w8(32'h3bcd7cb6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf899),
	.w1(32'h3bb43c25),
	.w2(32'h3c5461ce),
	.w3(32'h3bd605d9),
	.w4(32'h3be1e57e),
	.w5(32'h3c832a0e),
	.w6(32'h3bf245e0),
	.w7(32'h3c340d0a),
	.w8(32'hbb4bbfb7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23f24f),
	.w1(32'hb9d71f95),
	.w2(32'hbb7688fb),
	.w3(32'h3c1ee4d4),
	.w4(32'hbb860d94),
	.w5(32'hbba1fac2),
	.w6(32'hbb2bfdaf),
	.w7(32'hbc08cb63),
	.w8(32'hba8a0d50),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af665fe),
	.w1(32'hbadb77de),
	.w2(32'h3c545b74),
	.w3(32'hbba7243a),
	.w4(32'hbb6245db),
	.w5(32'h3c370df6),
	.w6(32'hbaa7dda7),
	.w7(32'h3b5b25bd),
	.w8(32'h3be450bd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a771f19),
	.w1(32'h3b6458f7),
	.w2(32'hbb2f67a8),
	.w3(32'h3b917c1a),
	.w4(32'hbb818494),
	.w5(32'hbbcc505d),
	.w6(32'h3b2bbe22),
	.w7(32'h3a79d268),
	.w8(32'h3a0aafbb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfe9bb),
	.w1(32'hbb9409cf),
	.w2(32'h3c1acbc3),
	.w3(32'hbba273c1),
	.w4(32'hbc4194be),
	.w5(32'h3c0d3940),
	.w6(32'h3b9c4280),
	.w7(32'h3a08c965),
	.w8(32'h3bb10f88),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7f21b),
	.w1(32'h3b39c931),
	.w2(32'h3c3cac3d),
	.w3(32'h3bd01001),
	.w4(32'h39028db0),
	.w5(32'h3b6771dc),
	.w6(32'h39de2cf9),
	.w7(32'hbb7417c9),
	.w8(32'hbb31ed70),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0984a9),
	.w1(32'hbbbd11e4),
	.w2(32'hb87459d3),
	.w3(32'hbc57000c),
	.w4(32'hbc89574e),
	.w5(32'hbb56fbd8),
	.w6(32'hbcb89dab),
	.w7(32'hbcad7115),
	.w8(32'hbaa8b39e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2da66),
	.w1(32'hbbf76a2f),
	.w2(32'h3b354c90),
	.w3(32'hbb9a2a28),
	.w4(32'hbb0e612f),
	.w5(32'hbb1c6310),
	.w6(32'hba9a0590),
	.w7(32'h3a988e04),
	.w8(32'hbbd3db0d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d59826),
	.w1(32'hbc5dc6d6),
	.w2(32'h3bbb9f36),
	.w3(32'hbc271c0a),
	.w4(32'hbc814aec),
	.w5(32'h3b65c1fc),
	.w6(32'hbc66bc01),
	.w7(32'hbc70afc9),
	.w8(32'hbb1f031c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3c649),
	.w1(32'h3c16ed8c),
	.w2(32'hb89e4f2b),
	.w3(32'h3c0494bb),
	.w4(32'h3b99e88d),
	.w5(32'h3baacb1c),
	.w6(32'h3b879f4f),
	.w7(32'h3c3bdc48),
	.w8(32'hb7ca2e50),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dd39a0),
	.w1(32'hbb0e861a),
	.w2(32'h3c7c3911),
	.w3(32'h3b006c13),
	.w4(32'hba360545),
	.w5(32'h3c88fdab),
	.w6(32'h39d9f2b9),
	.w7(32'h3a9fca1c),
	.w8(32'h3acf32be),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fc8d7),
	.w1(32'h3ba24b12),
	.w2(32'hbc0095dd),
	.w3(32'h3bfafc74),
	.w4(32'hba399a3f),
	.w5(32'hbb89b458),
	.w6(32'hbbc51536),
	.w7(32'hbc4c5f84),
	.w8(32'h3a8cf31c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d68d3),
	.w1(32'hbbbb6b8b),
	.w2(32'h3ba4fc36),
	.w3(32'h3a2c9f3a),
	.w4(32'h3b8f8192),
	.w5(32'h3b992f55),
	.w6(32'h3bd610bd),
	.w7(32'h3beb3414),
	.w8(32'h3b161161),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb27998),
	.w1(32'hbc958290),
	.w2(32'hbb9a5af8),
	.w3(32'hbcef1db1),
	.w4(32'hbc62777b),
	.w5(32'hbbed3aa3),
	.w6(32'hbc9d642f),
	.w7(32'hbc015eb7),
	.w8(32'h3b69759b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a3f81),
	.w1(32'h3baff44a),
	.w2(32'h3b5d1965),
	.w3(32'h3bbcc27c),
	.w4(32'h3c521436),
	.w5(32'h3baf8ba2),
	.w6(32'h3a69da2a),
	.w7(32'h3b9ef7f9),
	.w8(32'h3c22da87),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03e51e),
	.w1(32'h3c012a09),
	.w2(32'hbb34fdbd),
	.w3(32'h3c57ac72),
	.w4(32'hbac5dba2),
	.w5(32'hbcc1f854),
	.w6(32'h3c135997),
	.w7(32'hbb3ffa66),
	.w8(32'hbc8c982d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc208c50),
	.w1(32'hbbf09f99),
	.w2(32'hbbe4ee9a),
	.w3(32'hbc858f08),
	.w4(32'hbb2f4615),
	.w5(32'hbc1a79ea),
	.w6(32'hbb108a68),
	.w7(32'hb941dfc0),
	.w8(32'hbb07c163),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc516ed4),
	.w1(32'h3aef529d),
	.w2(32'h3c245720),
	.w3(32'hbc1674f5),
	.w4(32'h3c0a76fc),
	.w5(32'h3bd62af6),
	.w6(32'hba1e9b3e),
	.w7(32'h3c20aa01),
	.w8(32'h3bdd21f2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96e64d),
	.w1(32'hb93e0d4d),
	.w2(32'h3be7ff21),
	.w3(32'h3b0ffcc8),
	.w4(32'hba5997b7),
	.w5(32'hbb20beeb),
	.w6(32'h3ac93f71),
	.w7(32'h3aa1faa1),
	.w8(32'hbc4ea433),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc538724),
	.w1(32'hbc38d300),
	.w2(32'h3c7d3f14),
	.w3(32'hbc1699d0),
	.w4(32'hbbd43008),
	.w5(32'h3c8de766),
	.w6(32'h3a48126d),
	.w7(32'hbc03124f),
	.w8(32'h3ba0d337),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29aab6),
	.w1(32'hbc4e665a),
	.w2(32'hbc3a25a2),
	.w3(32'h3b42d823),
	.w4(32'hbc98f081),
	.w5(32'h3c056233),
	.w6(32'hbaaec12e),
	.w7(32'hbcdd7c9d),
	.w8(32'h3ca7db80),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c4108),
	.w1(32'h3b6030ba),
	.w2(32'hbc2cccf2),
	.w3(32'h3c7b2d1a),
	.w4(32'h3b5a667b),
	.w5(32'hbba2f2c9),
	.w6(32'h3c168b1d),
	.w7(32'h3b443405),
	.w8(32'hb9edf785),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18d757),
	.w1(32'h3b7de259),
	.w2(32'h3c0daf5e),
	.w3(32'h3be62527),
	.w4(32'h3c9eed3d),
	.w5(32'h3bbd882a),
	.w6(32'h3c2939ad),
	.w7(32'h3c3f6544),
	.w8(32'h3b9960ae),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d8818),
	.w1(32'h3b28de24),
	.w2(32'h3bbf2bea),
	.w3(32'hbacc7da7),
	.w4(32'hbb13695c),
	.w5(32'h3befd6a9),
	.w6(32'hbb914448),
	.w7(32'hbb6ea772),
	.w8(32'h3b562062),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf400d1),
	.w1(32'hbbd08fac),
	.w2(32'hba2c4829),
	.w3(32'h3a735815),
	.w4(32'hba7c511f),
	.w5(32'h3b04c9e6),
	.w6(32'hba5cc929),
	.w7(32'h37db6abc),
	.w8(32'hbac623e6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa04bc),
	.w1(32'hba9ddf46),
	.w2(32'hbb2b3ef2),
	.w3(32'hbb7b0e2b),
	.w4(32'h3c0b02cf),
	.w5(32'hbb8de1f0),
	.w6(32'h3b4152cb),
	.w7(32'h3c049419),
	.w8(32'hbb9d8453),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a8922),
	.w1(32'hbbbca9fe),
	.w2(32'h3c250ed9),
	.w3(32'hbc650e9c),
	.w4(32'hbbb108f2),
	.w5(32'h3b492a1f),
	.w6(32'hbaf28689),
	.w7(32'h3b2d96c0),
	.w8(32'h3c45bb66),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95b5eb),
	.w1(32'h3bcca1dd),
	.w2(32'hbb940cfe),
	.w3(32'h3c05ef81),
	.w4(32'hbb249317),
	.w5(32'h3b9d039b),
	.w6(32'h3b964830),
	.w7(32'hbbc534f2),
	.w8(32'h3af95679),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baad328),
	.w1(32'h3c265303),
	.w2(32'h3ac5e61b),
	.w3(32'h3aa1d1a1),
	.w4(32'hb9099e17),
	.w5(32'h3bc86ca3),
	.w6(32'hbb4ef820),
	.w7(32'hbb9e99af),
	.w8(32'h3b0245e2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbae9a6),
	.w1(32'hbc50f6e7),
	.w2(32'hbbfdab93),
	.w3(32'hbbe66361),
	.w4(32'hbcd661f9),
	.w5(32'h3bad7193),
	.w6(32'hbcaf5d09),
	.w7(32'hbce5e74b),
	.w8(32'h3c06cce8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e3b91),
	.w1(32'h3b57a0fd),
	.w2(32'h3c58ed77),
	.w3(32'h3ccc6dbd),
	.w4(32'h3bf19de6),
	.w5(32'h3c51ebf6),
	.w6(32'h3c5b7b3e),
	.w7(32'h3b822b40),
	.w8(32'h3b3e6d6a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e5bb4),
	.w1(32'h3ab51a6d),
	.w2(32'h3c971dd6),
	.w3(32'h3ad54d2b),
	.w4(32'hbbae7bf3),
	.w5(32'h3c6400c0),
	.w6(32'h3b6617e3),
	.w7(32'hbb508d0e),
	.w8(32'h3b88d4e6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4aad99),
	.w1(32'h3a903a2f),
	.w2(32'hbc124651),
	.w3(32'h3b9cfdc9),
	.w4(32'hbbad56e1),
	.w5(32'hbc63ba9e),
	.w6(32'hbbc5bd83),
	.w7(32'hbc0d86a4),
	.w8(32'hba3f6b8f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55887a),
	.w1(32'hbbb67c2a),
	.w2(32'h3c812b1b),
	.w3(32'hbbdf9cda),
	.w4(32'h3b06d764),
	.w5(32'h3c8ae51b),
	.w6(32'h3b32242a),
	.w7(32'hbbb1dd09),
	.w8(32'h3c5c7143),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ee04c),
	.w1(32'hbb0d7e8c),
	.w2(32'hbb8d69ed),
	.w3(32'h3cad2519),
	.w4(32'hbc0e7ecc),
	.w5(32'hb8d2f416),
	.w6(32'h3b38a7ab),
	.w7(32'hbca6cabe),
	.w8(32'hbb1d3133),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54202a),
	.w1(32'hbc5e2c81),
	.w2(32'h39857c9a),
	.w3(32'hbc4e766c),
	.w4(32'hbc89c9d5),
	.w5(32'hbc31c048),
	.w6(32'hbc094828),
	.w7(32'hbc01f482),
	.w8(32'hbb116deb),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc037786),
	.w1(32'hbac49226),
	.w2(32'hbbecc818),
	.w3(32'hbb731268),
	.w4(32'h3ae7b60c),
	.w5(32'hbc7978f3),
	.w6(32'h3ab945bf),
	.w7(32'h3b92c1e8),
	.w8(32'hbc0b4925),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12b44f),
	.w1(32'hbbadee69),
	.w2(32'h3ba17592),
	.w3(32'hbc6a0cd9),
	.w4(32'hbba91bca),
	.w5(32'hb88886cb),
	.w6(32'hbc2971d0),
	.w7(32'hbad6a0e3),
	.w8(32'hbbba5cec),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53aa41),
	.w1(32'hbb0a656f),
	.w2(32'h3ae399ea),
	.w3(32'hbbc08369),
	.w4(32'hbbcbc03d),
	.w5(32'h3bfcd2e4),
	.w6(32'hbbbd15ca),
	.w7(32'hba0a5539),
	.w8(32'h3b558278),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c3435),
	.w1(32'h3c520373),
	.w2(32'h3c724c18),
	.w3(32'h3c416743),
	.w4(32'h3c3935d6),
	.w5(32'h3c726096),
	.w6(32'h3b92a970),
	.w7(32'h3bb2742d),
	.w8(32'h3c15a7ab),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c371f52),
	.w1(32'h3b5d3b38),
	.w2(32'h3b20da7d),
	.w3(32'h3b9a4cbb),
	.w4(32'hbbe5bde6),
	.w5(32'h3be4be7c),
	.w6(32'h3bdc5090),
	.w7(32'hbbf179bd),
	.w8(32'h3bc95092),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c358da9),
	.w1(32'h3b872f6c),
	.w2(32'h3c5f0801),
	.w3(32'h3c59216f),
	.w4(32'h3b6089e6),
	.w5(32'h3c278e0a),
	.w6(32'h3bafcbf4),
	.w7(32'hb9dee32c),
	.w8(32'h3b05b55f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fca1f),
	.w1(32'hbbde27d3),
	.w2(32'h3bb48ca9),
	.w3(32'hbc60c328),
	.w4(32'hbc91446e),
	.w5(32'h3c544f03),
	.w6(32'hbc4a218e),
	.w7(32'hbb91825d),
	.w8(32'h3be11f6f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d29ce),
	.w1(32'hbb83b0aa),
	.w2(32'h3cd41ce5),
	.w3(32'h3c1645bd),
	.w4(32'hbbddecec),
	.w5(32'h3be8dbdb),
	.w6(32'hbb635357),
	.w7(32'hb9059bcb),
	.w8(32'h3c334fbd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b63b3),
	.w1(32'h3b64a473),
	.w2(32'h3c4f5c03),
	.w3(32'h3b763296),
	.w4(32'hbb1c7a43),
	.w5(32'hbb75a095),
	.w6(32'hbb9ff41f),
	.w7(32'hbc44913a),
	.w8(32'hbb92e71a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c292a99),
	.w1(32'h3ac7c8b9),
	.w2(32'hbb997837),
	.w3(32'hbc3857f9),
	.w4(32'hbbe897f3),
	.w5(32'hbc2ca983),
	.w6(32'hbc291b02),
	.w7(32'hbb68cc33),
	.w8(32'hbb8ca909),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37edba),
	.w1(32'hbbee00e3),
	.w2(32'hbb5981d4),
	.w3(32'hbc375703),
	.w4(32'h3a80b2a9),
	.w5(32'h3c8db86b),
	.w6(32'h39981ca3),
	.w7(32'h3c571178),
	.w8(32'h3c0fe80f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf9c7a),
	.w1(32'hbbb26e30),
	.w2(32'hbb955439),
	.w3(32'h3b073166),
	.w4(32'hbbab594f),
	.w5(32'hbc9fd955),
	.w6(32'h390b1a84),
	.w7(32'hbc0e664a),
	.w8(32'hbbceaa92),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3db737),
	.w1(32'hbc239870),
	.w2(32'h3bb8336f),
	.w3(32'hbcb141e0),
	.w4(32'hbc341083),
	.w5(32'h3bb1da12),
	.w6(32'hbaff33a7),
	.w7(32'h3bedcb5b),
	.w8(32'hb9a1f54f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06ece0),
	.w1(32'hbc0cf216),
	.w2(32'h3bf2b59b),
	.w3(32'hbc6edc87),
	.w4(32'hbcc10592),
	.w5(32'h3c047ef0),
	.w6(32'hbc3a5b35),
	.w7(32'hbc5ca1e4),
	.w8(32'h3bd01913),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d5375),
	.w1(32'h3aa34163),
	.w2(32'hbc2d7e6c),
	.w3(32'hba0761e8),
	.w4(32'hbc07014d),
	.w5(32'hbbc4e793),
	.w6(32'hba4adb8d),
	.w7(32'hbb9059cd),
	.w8(32'hbbcd3bcf),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf71d7),
	.w1(32'hb8b92a33),
	.w2(32'h3b749869),
	.w3(32'hbb8c6cff),
	.w4(32'hbbcdfc5e),
	.w5(32'h3a95980e),
	.w6(32'hbc113305),
	.w7(32'hbc1d37be),
	.w8(32'hbb16a24d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fbcc7),
	.w1(32'h3ae29103),
	.w2(32'h3bd2b473),
	.w3(32'h39ec1e9c),
	.w4(32'hb9f1a899),
	.w5(32'h3befea02),
	.w6(32'hba1df972),
	.w7(32'hbb151270),
	.w8(32'h3ad698ce),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b765c),
	.w1(32'hbad242f0),
	.w2(32'hbc35a8dd),
	.w3(32'hbb5a10ae),
	.w4(32'hbb796470),
	.w5(32'hbc10b1cb),
	.w6(32'hbb95bfd2),
	.w7(32'hbb71d6bf),
	.w8(32'h3b833838),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca65f3f),
	.w1(32'hbc0d363f),
	.w2(32'hbc95175b),
	.w3(32'hbc92adf9),
	.w4(32'h39bf37f2),
	.w5(32'hbcc3974d),
	.w6(32'h3a13eaaf),
	.w7(32'h3c818277),
	.w8(32'hbc111e28),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57c8de),
	.w1(32'hb9819f62),
	.w2(32'h3c2c33bb),
	.w3(32'hbc3d1ff4),
	.w4(32'h3bbc8d7f),
	.w5(32'h3b8722fe),
	.w6(32'h3babc868),
	.w7(32'h3c6ffc81),
	.w8(32'h3a8245a1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc577723),
	.w1(32'hbbee4432),
	.w2(32'h3c637d6a),
	.w3(32'hbae6a632),
	.w4(32'hbbb52311),
	.w5(32'h3b08a6a6),
	.w6(32'hbbfc978d),
	.w7(32'h3b42eef8),
	.w8(32'hbb0d04a7),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e64f92),
	.w1(32'hbbced3d7),
	.w2(32'h3bea03c0),
	.w3(32'hbb73c404),
	.w4(32'hbc1f658a),
	.w5(32'h3b86164a),
	.w6(32'hba80a2d0),
	.w7(32'hbb399bef),
	.w8(32'hbb3d788c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d29977),
	.w1(32'hbb031b0b),
	.w2(32'h3c096fa5),
	.w3(32'hbbafa322),
	.w4(32'hbc3198af),
	.w5(32'hbba2ec7c),
	.w6(32'hbbf1cf99),
	.w7(32'hbb7ab489),
	.w8(32'hbb10dbcd),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule