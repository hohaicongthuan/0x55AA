module layer_10_featuremap_465(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba903952),
	.w1(32'h3a2b5fd5),
	.w2(32'hbad6c92f),
	.w3(32'h3b98c67e),
	.w4(32'h3abfba50),
	.w5(32'hbc175ce6),
	.w6(32'h3c34027a),
	.w7(32'h3abb40df),
	.w8(32'hbb455738),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ba089),
	.w1(32'hbb6951b6),
	.w2(32'hbb0ef1e4),
	.w3(32'hbaba2766),
	.w4(32'hbb171c91),
	.w5(32'h3b2595fe),
	.w6(32'hbaadec36),
	.w7(32'hba41ddb7),
	.w8(32'h396d11b0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5bccf),
	.w1(32'h3b9a1099),
	.w2(32'h3c5932f7),
	.w3(32'h3be05477),
	.w4(32'h3c119121),
	.w5(32'h3c847eb0),
	.w6(32'h3b3a8e49),
	.w7(32'h3c810536),
	.w8(32'h3c44a9c6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b92f),
	.w1(32'h3c20410c),
	.w2(32'hbae350bb),
	.w3(32'hbc64200c),
	.w4(32'h3c1b74db),
	.w5(32'h3bbb623f),
	.w6(32'hbc399af3),
	.w7(32'h3c0f2bf9),
	.w8(32'hbb9f33ad),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20255),
	.w1(32'hbab6fb1e),
	.w2(32'hba42d4c4),
	.w3(32'h39da9f56),
	.w4(32'h3b53fdaa),
	.w5(32'h389ff687),
	.w6(32'h3b975b4d),
	.w7(32'hba53d3dc),
	.w8(32'h3a5afd38),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd500a0),
	.w1(32'hbb202abf),
	.w2(32'h3a842ea4),
	.w3(32'hbab949dc),
	.w4(32'h3b0a09ed),
	.w5(32'h3b2aa066),
	.w6(32'h3b20d583),
	.w7(32'hba1c32b8),
	.w8(32'h3b40ca74),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc6fdf),
	.w1(32'hbc156795),
	.w2(32'h3aa46b0a),
	.w3(32'hbb552671),
	.w4(32'hbbf5f136),
	.w5(32'h3a8b5ccc),
	.w6(32'hbbb08d2c),
	.w7(32'hbb9162f5),
	.w8(32'h3af34569),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6f74b),
	.w1(32'hbca75497),
	.w2(32'hbae94fe5),
	.w3(32'h3b8ab71a),
	.w4(32'hbc7408bf),
	.w5(32'hbc33e16a),
	.w6(32'hbb189003),
	.w7(32'hbb47e5b2),
	.w8(32'hbc359ea2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d5e19),
	.w1(32'h3ad33e64),
	.w2(32'hbc1b168e),
	.w3(32'hbb67fa22),
	.w4(32'h3c7aed1f),
	.w5(32'h3d5bd702),
	.w6(32'hbbffc04d),
	.w7(32'h3a9d2769),
	.w8(32'hbb9578e9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c2e7a),
	.w1(32'h3bf00953),
	.w2(32'h3ad24cbc),
	.w3(32'hbc81698b),
	.w4(32'h3b08e95f),
	.w5(32'h3afd1c5b),
	.w6(32'hbc924d71),
	.w7(32'h396f243c),
	.w8(32'h3ab6afc0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08db4f),
	.w1(32'hbad12240),
	.w2(32'hbb7a9a13),
	.w3(32'h3abf42f0),
	.w4(32'hbc0240ca),
	.w5(32'hba8b4822),
	.w6(32'h3c0532ac),
	.w7(32'hbbc9596b),
	.w8(32'hbac12b31),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2b772),
	.w1(32'h3a80bc5e),
	.w2(32'hba342e88),
	.w3(32'h3b6a5b5b),
	.w4(32'hbaa0f434),
	.w5(32'h3acd6a5f),
	.w6(32'h3a6249bf),
	.w7(32'h3ab398d8),
	.w8(32'h3b44082d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a1995),
	.w1(32'h3a5d8756),
	.w2(32'hbc710518),
	.w3(32'hbaf3bc57),
	.w4(32'hbb111297),
	.w5(32'hbc036b19),
	.w6(32'h3b18de4b),
	.w7(32'hbb5739c4),
	.w8(32'hbc28a26c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea72a9),
	.w1(32'h3c2cc40c),
	.w2(32'hbb157639),
	.w3(32'h3c040f6c),
	.w4(32'h3bcc75f5),
	.w5(32'h3bccc0e6),
	.w6(32'h3bb69e56),
	.w7(32'hbc0839a2),
	.w8(32'h3c72e7b8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93b1cd),
	.w1(32'h3b09894d),
	.w2(32'h3b9d8f0c),
	.w3(32'hbbe56fd6),
	.w4(32'h3b3e2503),
	.w5(32'h3b8475ae),
	.w6(32'h3ba131ab),
	.w7(32'hb94f36fc),
	.w8(32'h3a9a91a2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43239c),
	.w1(32'hbbdd0d51),
	.w2(32'hb975dcc0),
	.w3(32'h3c483f5b),
	.w4(32'hbbc26f0c),
	.w5(32'h3a968fc3),
	.w6(32'h3b5b0a79),
	.w7(32'hbb564bf9),
	.w8(32'hbb3585fb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b906d9a),
	.w1(32'hbaedcc06),
	.w2(32'hb9d7bb3b),
	.w3(32'h3c224c6c),
	.w4(32'hbb143f32),
	.w5(32'hbb168bf7),
	.w6(32'h3ba21e1e),
	.w7(32'h3b8358ad),
	.w8(32'h3aaf003b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15bd30),
	.w1(32'hba0dbf98),
	.w2(32'hbb154284),
	.w3(32'h39c4353b),
	.w4(32'hbbb8736f),
	.w5(32'hbb7e720f),
	.w6(32'h3a862845),
	.w7(32'hb98e42a4),
	.w8(32'hbb1ff70c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0db40),
	.w1(32'hbbdcf24f),
	.w2(32'hbb899154),
	.w3(32'hb701802d),
	.w4(32'hbbb63aaa),
	.w5(32'h3c564d31),
	.w6(32'h3abda592),
	.w7(32'hbb3fc170),
	.w8(32'h3a859d67),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f2cca),
	.w1(32'h3aa97add),
	.w2(32'hbb6053bb),
	.w3(32'h3a8c1477),
	.w4(32'hba9f5027),
	.w5(32'hbbe6caad),
	.w6(32'h3b40aab7),
	.w7(32'hbb1fb597),
	.w8(32'hbb95bff8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b513b1b),
	.w1(32'hbb32a24f),
	.w2(32'h3ae102d4),
	.w3(32'hbba765bc),
	.w4(32'hbb98f931),
	.w5(32'h3c14ac44),
	.w6(32'hbb1cd969),
	.w7(32'hbbdd0c4d),
	.w8(32'h3b4dddc5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac39505),
	.w1(32'h3aa85021),
	.w2(32'hb9f90d57),
	.w3(32'h3b341b27),
	.w4(32'h3a43269d),
	.w5(32'hbb83b4d6),
	.w6(32'hba530917),
	.w7(32'hba58abde),
	.w8(32'h3a1c846b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706cb8),
	.w1(32'h3a85a682),
	.w2(32'h3a2d7bb8),
	.w3(32'hbbdd8253),
	.w4(32'h3be6342f),
	.w5(32'h3b0440bb),
	.w6(32'hbb4d9f55),
	.w7(32'h3baf1094),
	.w8(32'h3b1645fe),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2539f8),
	.w1(32'hbb79481b),
	.w2(32'hbae68d76),
	.w3(32'h3b9de97e),
	.w4(32'hbc173593),
	.w5(32'hbb0ed8b0),
	.w6(32'hbb59caa9),
	.w7(32'hbbc1ef8b),
	.w8(32'hbae51b87),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfe983),
	.w1(32'hb9e46a71),
	.w2(32'hba0003b3),
	.w3(32'h3a644e2c),
	.w4(32'hbba8c5c4),
	.w5(32'h39db2900),
	.w6(32'h3b6e1b11),
	.w7(32'hbaf7ec13),
	.w8(32'hbb18b6ef),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfb5a1),
	.w1(32'hbab8589d),
	.w2(32'h3b318f43),
	.w3(32'h3b0860f0),
	.w4(32'hbb86d2c2),
	.w5(32'h3bcbb9a2),
	.w6(32'hbaad7e95),
	.w7(32'hbbab07ef),
	.w8(32'h3bd035e1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67d315),
	.w1(32'h3bb92856),
	.w2(32'h3badecf8),
	.w3(32'h3c2c4fea),
	.w4(32'h39958a0b),
	.w5(32'h3bbf83a5),
	.w6(32'h3b3c58e9),
	.w7(32'h3b60d179),
	.w8(32'hbb360277),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25aaa2),
	.w1(32'hbba6cd34),
	.w2(32'h3955e480),
	.w3(32'hbb4d6154),
	.w4(32'hbb568f7a),
	.w5(32'h3bbecdc3),
	.w6(32'h39e07355),
	.w7(32'hbb2409db),
	.w8(32'h3b11de74),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd841b),
	.w1(32'h3c03da6f),
	.w2(32'h3adecb70),
	.w3(32'h393cac57),
	.w4(32'hb81f5054),
	.w5(32'hbad8e1b9),
	.w6(32'hbb03c28c),
	.w7(32'hba6eae99),
	.w8(32'hbacd3a4c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c57d6),
	.w1(32'hbbdce4d8),
	.w2(32'hbbb1300d),
	.w3(32'h3b36e052),
	.w4(32'hbb73c799),
	.w5(32'hbb7dffba),
	.w6(32'h3be23aa9),
	.w7(32'hbb9b1e64),
	.w8(32'hbb6af2db),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb606f59),
	.w1(32'h39c3e2f2),
	.w2(32'hbb6e9062),
	.w3(32'hbb9481a9),
	.w4(32'h39475477),
	.w5(32'hbb8789f8),
	.w6(32'hbb8957e6),
	.w7(32'hbb40d49f),
	.w8(32'h3b3db019),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d714f),
	.w1(32'h3a9255dc),
	.w2(32'h3b48794d),
	.w3(32'hba0b71ea),
	.w4(32'hbb749f8b),
	.w5(32'hbb0537ff),
	.w6(32'hbaa8fb2d),
	.w7(32'h3b0e10d3),
	.w8(32'hbb205e2a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b501fae),
	.w1(32'hbb667d43),
	.w2(32'hb926d1e7),
	.w3(32'h3c4a422c),
	.w4(32'hbc0077e4),
	.w5(32'hba9741cd),
	.w6(32'hbb3d1f8f),
	.w7(32'hbb654589),
	.w8(32'h3b3cbb3f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fd459),
	.w1(32'hbb64596e),
	.w2(32'hbb774fa8),
	.w3(32'hbbfe65ed),
	.w4(32'hbbd68c56),
	.w5(32'hbafadf59),
	.w6(32'h3aa4c145),
	.w7(32'hbb968ab9),
	.w8(32'hbac8ef84),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d45bd),
	.w1(32'h3c44b6e5),
	.w2(32'h3bca571d),
	.w3(32'h3a33c928),
	.w4(32'hbb5ed176),
	.w5(32'h3c0b944f),
	.w6(32'h3b799d14),
	.w7(32'hbc67637a),
	.w8(32'h3c7f0955),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8ed52),
	.w1(32'h3b095b5f),
	.w2(32'h3b04b1b4),
	.w3(32'h3c6a7344),
	.w4(32'h3b32311c),
	.w5(32'h3ca2a64f),
	.w6(32'h3cb3e9e9),
	.w7(32'h3b6c0f27),
	.w8(32'h3bbf928d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6468),
	.w1(32'hbcdca8bf),
	.w2(32'hbcad55bb),
	.w3(32'hbbc6aa2d),
	.w4(32'hbcfdc525),
	.w5(32'hbc9f1546),
	.w6(32'hbae8c7e2),
	.w7(32'hbcd3b1a9),
	.w8(32'hbc8da4f5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8157659),
	.w1(32'hbacbad2c),
	.w2(32'hba42ce8e),
	.w3(32'hbba436f2),
	.w4(32'h3b028314),
	.w5(32'h3ada6979),
	.w6(32'hbc0e02c4),
	.w7(32'h3919de95),
	.w8(32'hbb2fbc22),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cf817),
	.w1(32'hbbedd1fc),
	.w2(32'hbc19ff1e),
	.w3(32'hbb7d26ef),
	.w4(32'hbb271ee1),
	.w5(32'hbc7a9ece),
	.w6(32'hbc3b829c),
	.w7(32'hbadbb40e),
	.w8(32'hbc19c906),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6c70c),
	.w1(32'h3bef4968),
	.w2(32'hb96246b4),
	.w3(32'hbc35fe68),
	.w4(32'h3c33790e),
	.w5(32'h3c135763),
	.w6(32'hbc23a308),
	.w7(32'h3bf8e8a8),
	.w8(32'h3b811702),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdf4b7),
	.w1(32'h39aedab3),
	.w2(32'hbb782ebd),
	.w3(32'hb98fa157),
	.w4(32'h3cd759f4),
	.w5(32'hbca1f76f),
	.w6(32'h3a92f587),
	.w7(32'hbbd53567),
	.w8(32'hbbb89b3c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf684e),
	.w1(32'hbabaa344),
	.w2(32'h3b8ea3d3),
	.w3(32'hbbc669f3),
	.w4(32'h3b6cbafa),
	.w5(32'h3c08a3d5),
	.w6(32'hbc279ecd),
	.w7(32'h3a9aee64),
	.w8(32'h3a30dbec),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc270802),
	.w1(32'hbb5c526c),
	.w2(32'hbc057e78),
	.w3(32'hbb4e72dc),
	.w4(32'hbbe39c46),
	.w5(32'hbbf2870d),
	.w6(32'hbc404961),
	.w7(32'hbbce9cab),
	.w8(32'hbc0fcfbe),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae8c65),
	.w1(32'h3b04ca0e),
	.w2(32'h397f7d71),
	.w3(32'h393fe25b),
	.w4(32'h3b01480a),
	.w5(32'hbc2d4a6e),
	.w6(32'hb865b643),
	.w7(32'hba3eeb9a),
	.w8(32'hbb2079b9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc2a10),
	.w1(32'h3a0425fe),
	.w2(32'h3b9bdbaa),
	.w3(32'h3b91439a),
	.w4(32'h3b5c0d11),
	.w5(32'h3c1a828e),
	.w6(32'h3b04c034),
	.w7(32'h3a89c91e),
	.w8(32'h39a6fcd4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa22900),
	.w1(32'hbb996758),
	.w2(32'hbb83f538),
	.w3(32'hbb85d558),
	.w4(32'hbb5eaa91),
	.w5(32'hbad9309a),
	.w6(32'hb9350292),
	.w7(32'hbb7e6d33),
	.w8(32'hbb90e9ac),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab14c57),
	.w1(32'hbadcf1e8),
	.w2(32'hbb1b895a),
	.w3(32'h3b03917d),
	.w4(32'hbbecd52e),
	.w5(32'hbb14ec6b),
	.w6(32'hbaadfd0f),
	.w7(32'hbba9a420),
	.w8(32'h3a06d051),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83eebd),
	.w1(32'h3bd4fc8c),
	.w2(32'h3be105d7),
	.w3(32'h3b0e8605),
	.w4(32'h3bc5d5fd),
	.w5(32'h3bcd6f79),
	.w6(32'hba75f445),
	.w7(32'h3a8117e3),
	.w8(32'h3ba7ca72),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ef193),
	.w1(32'h3ab2a9f2),
	.w2(32'h3c808e31),
	.w3(32'hbc1d88bb),
	.w4(32'h3c4ce067),
	.w5(32'h3d3d9fdc),
	.w6(32'hbc039686),
	.w7(32'h3b776e39),
	.w8(32'h3cd99645),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc92de1),
	.w1(32'hbc284d4f),
	.w2(32'hbc7467eb),
	.w3(32'h3b8bf52d),
	.w4(32'hbc85543e),
	.w5(32'hbd108e1d),
	.w6(32'h3c12062e),
	.w7(32'hbc3784f7),
	.w8(32'hbc88ac1e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27ca7d),
	.w1(32'h39be04d0),
	.w2(32'hbb9c22c5),
	.w3(32'hbb85587f),
	.w4(32'h3b6dbf82),
	.w5(32'hbb7b358b),
	.w6(32'hbbcf5410),
	.w7(32'h3ba13497),
	.w8(32'hbb5f9721),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e3e94),
	.w1(32'hbb5c3ec4),
	.w2(32'h39b86009),
	.w3(32'hbba51117),
	.w4(32'hbbc4b61e),
	.w5(32'h3b8f9d7c),
	.w6(32'hbbd4de77),
	.w7(32'h3b22fcd6),
	.w8(32'h3babe249),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab6ab7),
	.w1(32'h3b960a5c),
	.w2(32'h39ae60ff),
	.w3(32'hba8c524d),
	.w4(32'h3a3b03c3),
	.w5(32'h3a0ed3f3),
	.w6(32'h3a74b7c7),
	.w7(32'hbad5e9aa),
	.w8(32'h39ea5706),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7313f6),
	.w1(32'h3be16ada),
	.w2(32'h3b8b04fa),
	.w3(32'hbbc20bad),
	.w4(32'hb9508d09),
	.w5(32'h3c7956f2),
	.w6(32'hbb3f1856),
	.w7(32'hbbea7319),
	.w8(32'h3b569d46),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89414b),
	.w1(32'hb9cd72f3),
	.w2(32'hbbd0b78b),
	.w3(32'h3b64b1b3),
	.w4(32'h3aecbdf6),
	.w5(32'hbb4bb29c),
	.w6(32'h3bac5643),
	.w7(32'h3b1df4ec),
	.w8(32'hbbdb505d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6821a2),
	.w1(32'h3b007400),
	.w2(32'hbb7cb18a),
	.w3(32'hbb88943c),
	.w4(32'h3af44ae9),
	.w5(32'h3d002c43),
	.w6(32'hbbd8dc7b),
	.w7(32'hbb8c9512),
	.w8(32'h3b5f4fcf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbf901),
	.w1(32'h3980875a),
	.w2(32'hbb3af328),
	.w3(32'h3c055303),
	.w4(32'h38c3d393),
	.w5(32'hbb8a2e91),
	.w6(32'h3b78b000),
	.w7(32'h3ae2f8d8),
	.w8(32'hba9b667f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceaadf),
	.w1(32'hbb1582a8),
	.w2(32'h394911b4),
	.w3(32'hbae5495b),
	.w4(32'hbb61d021),
	.w5(32'h3b2c18e7),
	.w6(32'h37d02494),
	.w7(32'h3b39a85d),
	.w8(32'hbb2813c2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03cf29),
	.w1(32'hbb99eae8),
	.w2(32'hbbf01c30),
	.w3(32'h3a075308),
	.w4(32'hbbd62349),
	.w5(32'hbc881a26),
	.w6(32'hbb8860cb),
	.w7(32'hbb7fe4b2),
	.w8(32'hbbffff4b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef5fb8),
	.w1(32'hbae7397b),
	.w2(32'hbb1633c1),
	.w3(32'hb9ff1ffc),
	.w4(32'hbb006b8b),
	.w5(32'h3b62f80f),
	.w6(32'hba9d2d58),
	.w7(32'hbb9416d1),
	.w8(32'hbb9af1f7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb181e),
	.w1(32'h38d3596d),
	.w2(32'h3b096a88),
	.w3(32'hba6ca22f),
	.w4(32'h3a865cb7),
	.w5(32'h3b4f3f81),
	.w6(32'hbb91d909),
	.w7(32'hbb9381f8),
	.w8(32'hbb9913fe),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b250dc5),
	.w1(32'hbb68f177),
	.w2(32'h39af8087),
	.w3(32'hbb1fe03a),
	.w4(32'hbb795fc0),
	.w5(32'hbafe622d),
	.w6(32'hbba38875),
	.w7(32'hbb91934c),
	.w8(32'hb92840b2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2eb14),
	.w1(32'hbc168918),
	.w2(32'hbbf59305),
	.w3(32'h3c2413d4),
	.w4(32'hbc439d03),
	.w5(32'hbc66d57f),
	.w6(32'h3b33b559),
	.w7(32'hbc4ca112),
	.w8(32'hbc319907),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc3d8),
	.w1(32'h3b908d19),
	.w2(32'hb9440aff),
	.w3(32'hbb5cbb33),
	.w4(32'h3b2c5d3a),
	.w5(32'hbac6d0f5),
	.w6(32'hbb266b3b),
	.w7(32'h3994e067),
	.w8(32'h398de698),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd2a62),
	.w1(32'h3be990b6),
	.w2(32'h3b6c56a0),
	.w3(32'hbaec3cfd),
	.w4(32'h3bf5dcb8),
	.w5(32'h3b8af6d2),
	.w6(32'h3b59c624),
	.w7(32'h3c0cedd1),
	.w8(32'h3bb5806e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b907cc3),
	.w1(32'h3b8dc0c0),
	.w2(32'h3b02dc1c),
	.w3(32'h3b3e32a6),
	.w4(32'h3bf9461d),
	.w5(32'h3b996a33),
	.w6(32'h3ba9fd12),
	.w7(32'h3b983e3e),
	.w8(32'h3c09b606),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaadb53),
	.w1(32'h39a50131),
	.w2(32'hbbb64945),
	.w3(32'hbaf06bac),
	.w4(32'h39037eb7),
	.w5(32'hbbb132bf),
	.w6(32'h3b22889e),
	.w7(32'hbc4be082),
	.w8(32'hbc1ccd29),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28b4b1),
	.w1(32'h3bc13512),
	.w2(32'h3bbeea81),
	.w3(32'hbc832485),
	.w4(32'hbace2c05),
	.w5(32'h3c73682a),
	.w6(32'hbc0e869d),
	.w7(32'hbad54580),
	.w8(32'h3b904041),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2baff2),
	.w1(32'hbb8808ea),
	.w2(32'hbb8e4f2e),
	.w3(32'h3a6ddb49),
	.w4(32'hbbd14579),
	.w5(32'hbb4478d4),
	.w6(32'h3b2e3fb2),
	.w7(32'hbb878972),
	.w8(32'hbbb16763),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b437618),
	.w1(32'hbc043714),
	.w2(32'hbc2fefdc),
	.w3(32'h39e87253),
	.w4(32'hbbeb0c7f),
	.w5(32'hbc2ca690),
	.w6(32'hba4ac7bb),
	.w7(32'hbba17cef),
	.w8(32'hbb442046),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55c62e),
	.w1(32'h3c869ef9),
	.w2(32'hbbccea87),
	.w3(32'hbc7473c1),
	.w4(32'h3cc7043b),
	.w5(32'h3bd0f0de),
	.w6(32'hbc7cc362),
	.w7(32'h3c4fb66f),
	.w8(32'hbc16f50c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1db51b),
	.w1(32'h3c2842f4),
	.w2(32'hbac8e162),
	.w3(32'hbc3d226b),
	.w4(32'h3ae256e8),
	.w5(32'h3bd0f801),
	.w6(32'hbc6e2792),
	.w7(32'hbc14153f),
	.w8(32'hbb9ea8fe),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2993e6),
	.w1(32'h3bcd787e),
	.w2(32'hbc1798c8),
	.w3(32'hbc2d2d07),
	.w4(32'h3c62b119),
	.w5(32'hbba2a6cd),
	.w6(32'hbb5e80fe),
	.w7(32'h3c56f952),
	.w8(32'h3c198b0d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6abdc4),
	.w1(32'hbb7cd75d),
	.w2(32'hba88215c),
	.w3(32'hbc070d46),
	.w4(32'hbb5c2ed9),
	.w5(32'h3c068090),
	.w6(32'hbc4d1399),
	.w7(32'hbbe90a3b),
	.w8(32'hbbb4cd99),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47d6f8),
	.w1(32'hbb616be2),
	.w2(32'h3bf7f932),
	.w3(32'h3ab3b693),
	.w4(32'hbbc973a9),
	.w5(32'h3b89ad9d),
	.w6(32'h3a1f2817),
	.w7(32'h3bdd98bc),
	.w8(32'h3c0743cf),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc82a50),
	.w1(32'h3c0b66b9),
	.w2(32'hba8c6a20),
	.w3(32'hbb9db6c8),
	.w4(32'h3ba937e6),
	.w5(32'h3bdfc8ca),
	.w6(32'h3bc04862),
	.w7(32'h3be89208),
	.w8(32'h3b796260),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6891),
	.w1(32'h3ae617b6),
	.w2(32'hbad5a756),
	.w3(32'hba50692b),
	.w4(32'h3a889798),
	.w5(32'hbb9cc7fa),
	.w6(32'hbb4528e4),
	.w7(32'h3b31620a),
	.w8(32'hbb274c7d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7e35f),
	.w1(32'h3b8fdd0f),
	.w2(32'hbc65fb34),
	.w3(32'h3b61b093),
	.w4(32'h3cc40cf3),
	.w5(32'hbb36ec4d),
	.w6(32'hbb2b7d4a),
	.w7(32'h3c9e328b),
	.w8(32'hbc2957d4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70076c),
	.w1(32'hbbe3aa0e),
	.w2(32'h3bd0d5eb),
	.w3(32'hbc7b6f9f),
	.w4(32'hbc8ce107),
	.w5(32'h3c529659),
	.w6(32'hbc5eb3da),
	.w7(32'hbc4cbaea),
	.w8(32'h3bb1a84f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9dc31a),
	.w1(32'h3ae73ffb),
	.w2(32'hbbf49325),
	.w3(32'h3d15eefa),
	.w4(32'h3c88cc0d),
	.w5(32'hbc8220a7),
	.w6(32'h3c39f180),
	.w7(32'h3c3c7002),
	.w8(32'h3c05200b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bcbb8),
	.w1(32'hbd2e2c0b),
	.w2(32'h3c013527),
	.w3(32'hbbbba2b9),
	.w4(32'hbd991f34),
	.w5(32'h3c5298cf),
	.w6(32'hbc2a0365),
	.w7(32'hbd61aea5),
	.w8(32'hbabdabfd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d56042d),
	.w1(32'h3b064fd7),
	.w2(32'h3a9f430b),
	.w3(32'h3db75b4b),
	.w4(32'h3c0dae1a),
	.w5(32'h3b069b45),
	.w6(32'h3d491c9a),
	.w7(32'hba4d3335),
	.w8(32'hbbb84865),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beef57a),
	.w1(32'hbb77dff8),
	.w2(32'hba5ef614),
	.w3(32'hbb05e3cf),
	.w4(32'hbb27a9cf),
	.w5(32'hbb043230),
	.w6(32'h3b61f791),
	.w7(32'h3ba9a761),
	.w8(32'h3b690a24),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05aa8d),
	.w1(32'hbbdf049a),
	.w2(32'h3c0b0913),
	.w3(32'h3b8000e2),
	.w4(32'hbbcde3b4),
	.w5(32'h3c111c54),
	.w6(32'h3aa45888),
	.w7(32'hbb7be959),
	.w8(32'hbc07411a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf18f0),
	.w1(32'h38795dac),
	.w2(32'hbc30d662),
	.w3(32'hbc237c71),
	.w4(32'h3be343b1),
	.w5(32'hbb519af1),
	.w6(32'h3a4981bc),
	.w7(32'h3b9f172e),
	.w8(32'h3ba720de),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc687442),
	.w1(32'h3c4049f7),
	.w2(32'h3b702ee9),
	.w3(32'hbc4b5741),
	.w4(32'h3cf130da),
	.w5(32'hbbacb27a),
	.w6(32'hbbb8fe0d),
	.w7(32'h3bb081c3),
	.w8(32'hbc1d18d6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90b0c1),
	.w1(32'h3c6642f1),
	.w2(32'hbbeecd86),
	.w3(32'hbc9ee0a6),
	.w4(32'h3c9bfb87),
	.w5(32'hbb110b9e),
	.w6(32'hbc04ba65),
	.w7(32'h3c92b802),
	.w8(32'h3be5bf43),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc185da0),
	.w1(32'hbb2fd376),
	.w2(32'h3abe5698),
	.w3(32'hbc8918c7),
	.w4(32'hbb0acfc0),
	.w5(32'h3be14e93),
	.w6(32'hbc461068),
	.w7(32'h3b737911),
	.w8(32'h3a25929a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6311dc),
	.w1(32'h3b073ff7),
	.w2(32'h3b5a8ff5),
	.w3(32'hb921af03),
	.w4(32'h3bdede95),
	.w5(32'h3b7de0d3),
	.w6(32'hbb99e0f5),
	.w7(32'h3b34c32a),
	.w8(32'h3a0db0a8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19a150),
	.w1(32'h3a040766),
	.w2(32'h39ee173c),
	.w3(32'hbc12760f),
	.w4(32'h3c41a773),
	.w5(32'hb99c026d),
	.w6(32'hbc6af0a5),
	.w7(32'h3c23adb4),
	.w8(32'hba2a9b69),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc125ac6),
	.w1(32'h3c034840),
	.w2(32'hbc93a330),
	.w3(32'hbc9bfd77),
	.w4(32'h3c593872),
	.w5(32'hbba1a8e5),
	.w6(32'hbbb83a11),
	.w7(32'h3c3cde07),
	.w8(32'hbc44c098),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68f1c0),
	.w1(32'hbc2c93be),
	.w2(32'h3b5ff6f7),
	.w3(32'hbd071280),
	.w4(32'h3c89f397),
	.w5(32'h3c57983d),
	.w6(32'hbc8b1d67),
	.w7(32'h39607d4d),
	.w8(32'h3b13bf0a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2cf55),
	.w1(32'h3a3f9fcd),
	.w2(32'h3b8c0796),
	.w3(32'hbc7efe38),
	.w4(32'hbbb151e8),
	.w5(32'h3b75a201),
	.w6(32'h3ba6eb5f),
	.w7(32'hbb9005a9),
	.w8(32'h3bdfc33c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67ea5c),
	.w1(32'hbc1cb4e0),
	.w2(32'h3c3555b9),
	.w3(32'h3c66beba),
	.w4(32'hbc77cd05),
	.w5(32'h3bb32232),
	.w6(32'h3bcfcf61),
	.w7(32'hbbf982c1),
	.w8(32'h3b303e13),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b823),
	.w1(32'hbc1f6ac3),
	.w2(32'hbb8e3579),
	.w3(32'h3c558026),
	.w4(32'h3bb9eaa5),
	.w5(32'h38ebe97f),
	.w6(32'h3b271a84),
	.w7(32'h3c613849),
	.w8(32'h3c1a4649),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1af506),
	.w1(32'h3c897df4),
	.w2(32'hbb20f382),
	.w3(32'hbc435f09),
	.w4(32'h3c905b3a),
	.w5(32'h3b19c5ef),
	.w6(32'hbc7f734c),
	.w7(32'h3c4fbac9),
	.w8(32'hbb8be2a8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe03fc9),
	.w1(32'h3c66f06c),
	.w2(32'h3b2b320a),
	.w3(32'hbc5565d1),
	.w4(32'h3c8a0c56),
	.w5(32'h3b5ac6bc),
	.w6(32'hbc04ca36),
	.w7(32'h3c16c3de),
	.w8(32'hbbb5357b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09cd4c),
	.w1(32'hbbc3ebdd),
	.w2(32'hbc6b2c29),
	.w3(32'hbc8accb4),
	.w4(32'h3a8b179c),
	.w5(32'hbc6b222d),
	.w6(32'hbc0da9f3),
	.w7(32'hbbc383c5),
	.w8(32'hbca15e8d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59f6f5),
	.w1(32'h3a5991bb),
	.w2(32'hba9ea668),
	.w3(32'hbc8fc574),
	.w4(32'h3c3c107e),
	.w5(32'hbbb7465a),
	.w6(32'hbc917213),
	.w7(32'h3bc48241),
	.w8(32'h3bba1b27),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ee700),
	.w1(32'hbbb65709),
	.w2(32'hbb2911a8),
	.w3(32'hbc3c82d1),
	.w4(32'h3c635f21),
	.w5(32'h3b70c26a),
	.w6(32'hbb9df525),
	.w7(32'h3bcf2206),
	.w8(32'h3bbbfa0a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed38dd),
	.w1(32'h3b876faa),
	.w2(32'h3a4626cc),
	.w3(32'hbcc2f3b0),
	.w4(32'h3b81e1a0),
	.w5(32'h3bae9f46),
	.w6(32'hbbc1934b),
	.w7(32'h3b669872),
	.w8(32'hbb497b0b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c9e6),
	.w1(32'h3bcf6bcd),
	.w2(32'h3b91e09c),
	.w3(32'hbbac114e),
	.w4(32'h3c38d3b8),
	.w5(32'hbb517f45),
	.w6(32'hbc2d8f08),
	.w7(32'h3c4cb6ff),
	.w8(32'h3b9b1a56),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc208172),
	.w1(32'h3a7284e1),
	.w2(32'h3beb8bba),
	.w3(32'hbc588afe),
	.w4(32'h3be426a9),
	.w5(32'h3c867644),
	.w6(32'hbc167eb9),
	.w7(32'hbb4d1133),
	.w8(32'hbc609466),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc111dab),
	.w1(32'h3baab438),
	.w2(32'hbbdff56b),
	.w3(32'hbc41a64c),
	.w4(32'h3c5a429d),
	.w5(32'hb9766069),
	.w6(32'hbcbce8f4),
	.w7(32'h3c25aa81),
	.w8(32'h3a58ad59),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae1f78),
	.w1(32'h3c0ce463),
	.w2(32'h3b7d0138),
	.w3(32'hbce43438),
	.w4(32'hbafdf487),
	.w5(32'h3bcabeda),
	.w6(32'hbc7202ca),
	.w7(32'h3b42024e),
	.w8(32'hb971a13c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a0f56),
	.w1(32'h3c294bdf),
	.w2(32'h3bffc683),
	.w3(32'hba69826f),
	.w4(32'h3bb4b82e),
	.w5(32'h373076e9),
	.w6(32'h3a5589e1),
	.w7(32'h390ff872),
	.w8(32'h3a38fd24),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9574e2),
	.w1(32'hba810fc2),
	.w2(32'h3b4ae071),
	.w3(32'h3b8bc0ce),
	.w4(32'h3b755119),
	.w5(32'h3c05d374),
	.w6(32'h3ae23b9e),
	.w7(32'hbb85bf68),
	.w8(32'hba932475),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20bcbc),
	.w1(32'h3c1776f7),
	.w2(32'hbcb27015),
	.w3(32'h3beb624a),
	.w4(32'h3c0f5e97),
	.w5(32'hba7e451f),
	.w6(32'h3a45380b),
	.w7(32'h3c112eb1),
	.w8(32'hbb07f291),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d53de),
	.w1(32'hb944850f),
	.w2(32'hbb5364de),
	.w3(32'hbcab5369),
	.w4(32'h3a0f0a6e),
	.w5(32'hbb8357d7),
	.w6(32'hbba8bcd6),
	.w7(32'h3bea0c3e),
	.w8(32'hbb3b775f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf9b18),
	.w1(32'h3bdb416b),
	.w2(32'h39e4d0c2),
	.w3(32'h39968f0e),
	.w4(32'h3c9f512b),
	.w5(32'hbc0e0ac7),
	.w6(32'hbac9af43),
	.w7(32'h3c9ff303),
	.w8(32'h3c07b995),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74290f),
	.w1(32'hba30ac40),
	.w2(32'hbb7ecdb0),
	.w3(32'hbc834d0e),
	.w4(32'h3ca86c8e),
	.w5(32'hbb209838),
	.w6(32'hbb97cd4c),
	.w7(32'hbbb6957c),
	.w8(32'hbc58db6e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8de1cf),
	.w1(32'h3c00e59a),
	.w2(32'h39d75a2b),
	.w3(32'hbc5b7fb7),
	.w4(32'h3cb6fc89),
	.w5(32'hbc790166),
	.w6(32'hbc018c14),
	.w7(32'h3c7088cb),
	.w8(32'hbc2424bc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ca9a1),
	.w1(32'h39acad1f),
	.w2(32'hbc03c5bc),
	.w3(32'hbc9bff85),
	.w4(32'hba135fda),
	.w5(32'hbc1754a2),
	.w6(32'hbc14f0f5),
	.w7(32'h3b8607a8),
	.w8(32'h3af87449),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc36f2),
	.w1(32'h3b86e954),
	.w2(32'hbb2a25e5),
	.w3(32'h3b956f8b),
	.w4(32'h3adfe244),
	.w5(32'h3cd0f5c5),
	.w6(32'h3c2944f8),
	.w7(32'h3b1668ab),
	.w8(32'hbc36985a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba349bd),
	.w1(32'hbb05bbc5),
	.w2(32'h399fe6d9),
	.w3(32'hbb4677f0),
	.w4(32'hbb2c5748),
	.w5(32'hbc9100c1),
	.w6(32'hbc3a437c),
	.w7(32'hbad9867f),
	.w8(32'h3b8f2812),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47cb53),
	.w1(32'h3a890024),
	.w2(32'hbc24a0b2),
	.w3(32'h3c3ad3a3),
	.w4(32'h3b65c083),
	.w5(32'hbc3d4719),
	.w6(32'h3c30cdbf),
	.w7(32'h3c029014),
	.w8(32'h3b1573c1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe50f54),
	.w1(32'h3b4c6535),
	.w2(32'hbaafb2c5),
	.w3(32'hbae103de),
	.w4(32'h3c13017f),
	.w5(32'hbba6061f),
	.w6(32'h3b78f6d9),
	.w7(32'h3ac29dfa),
	.w8(32'h3b38eb25),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dd076),
	.w1(32'hbc20e8c5),
	.w2(32'hb9d1416c),
	.w3(32'h3bdcd5de),
	.w4(32'hbb980246),
	.w5(32'h39dd6bc3),
	.w6(32'hb9ab71e3),
	.w7(32'hbb9a375c),
	.w8(32'h3b3d40f0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e6a16),
	.w1(32'h3c13ce9b),
	.w2(32'hbb637226),
	.w3(32'hbbf16f01),
	.w4(32'h3bf7f0a5),
	.w5(32'h3844ce4f),
	.w6(32'h3b9ec71e),
	.w7(32'h3c97bd75),
	.w8(32'hb91c6d8f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad18bb),
	.w1(32'h3bf2e593),
	.w2(32'h3b52e5d3),
	.w3(32'hba0f695d),
	.w4(32'h3bfa18ca),
	.w5(32'h3c206e73),
	.w6(32'hbb0b290a),
	.w7(32'h3b1ed175),
	.w8(32'hbbdf25ba),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc822193),
	.w1(32'hbc5cf3ee),
	.w2(32'h3b40eb0b),
	.w3(32'hbccfd29b),
	.w4(32'hbc229647),
	.w5(32'h3c39711e),
	.w6(32'hbc96291d),
	.w7(32'hbc88324a),
	.w8(32'h3b43619d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14ffbb),
	.w1(32'h3b7ed42f),
	.w2(32'hbb75648d),
	.w3(32'h3c1c210a),
	.w4(32'h3b0112fa),
	.w5(32'hbb56017e),
	.w6(32'h3ab1afc5),
	.w7(32'h3c7c3dcb),
	.w8(32'hbc5faee8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8f630),
	.w1(32'h3bd8a711),
	.w2(32'h3b749988),
	.w3(32'hbc8ee40c),
	.w4(32'h3c78601d),
	.w5(32'h3ae24dce),
	.w6(32'hbcd1b435),
	.w7(32'h3c283d93),
	.w8(32'h3a13c065),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ef420),
	.w1(32'hbbca4712),
	.w2(32'h3c1affc8),
	.w3(32'hbbc90c3c),
	.w4(32'hbbf741f3),
	.w5(32'h3b365154),
	.w6(32'hbae35e39),
	.w7(32'hbb377b9b),
	.w8(32'hbb5b86c9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c725349),
	.w1(32'h3c499ba1),
	.w2(32'h3a8c72c2),
	.w3(32'h3cad1143),
	.w4(32'h3c510412),
	.w5(32'hbbd2329d),
	.w6(32'h3bc4a5d9),
	.w7(32'h3c0132cb),
	.w8(32'h3b77b6d7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4da44),
	.w1(32'h3c54f47d),
	.w2(32'h3ab797ab),
	.w3(32'hbb7a28d3),
	.w4(32'h3c2746ae),
	.w5(32'h3ba232f4),
	.w6(32'hbbddfb62),
	.w7(32'hb70ad3ae),
	.w8(32'hbc200ba6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12f027),
	.w1(32'h3c0ea975),
	.w2(32'hbba34f5e),
	.w3(32'hbc851e70),
	.w4(32'h3d0fdca0),
	.w5(32'hbc06eb83),
	.w6(32'hbc25532f),
	.w7(32'h3c92088e),
	.w8(32'hbb57ea0c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e73a6),
	.w1(32'h3b46d939),
	.w2(32'h3c4a1dee),
	.w3(32'hbcf6d948),
	.w4(32'h3b107fc7),
	.w5(32'h3c0b189c),
	.w6(32'hbc5ad7ad),
	.w7(32'hba9525e1),
	.w8(32'hbc93d82e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a357a),
	.w1(32'hbc00a376),
	.w2(32'h3b3d3b97),
	.w3(32'hbc5c9c18),
	.w4(32'hbb89156d),
	.w5(32'h3b8ad51e),
	.w6(32'hbb5de699),
	.w7(32'hbba289c3),
	.w8(32'h3bc95432),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7eac8),
	.w1(32'h3b5e06ea),
	.w2(32'hbb450a51),
	.w3(32'hbb184bd5),
	.w4(32'h3c7734a7),
	.w5(32'hbb5f344e),
	.w6(32'h3b0f5c54),
	.w7(32'h3c6e2aa9),
	.w8(32'h3beec3f5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc795d96),
	.w1(32'h3b89b7a9),
	.w2(32'hbc986613),
	.w3(32'hbcdf5ce9),
	.w4(32'h3c49d19b),
	.w5(32'hbc3d798b),
	.w6(32'hbc6c8d09),
	.w7(32'h3c31a642),
	.w8(32'hbbecc7d2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44a063),
	.w1(32'h3c74e355),
	.w2(32'h3a0f62c4),
	.w3(32'hbc0c87ae),
	.w4(32'h3c3c8be2),
	.w5(32'h3c8e9b75),
	.w6(32'hbc796771),
	.w7(32'h3c8dac2f),
	.w8(32'h3c1b14b5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf29ada),
	.w1(32'hbc633809),
	.w2(32'hbbf985ee),
	.w3(32'hbbf242cd),
	.w4(32'hbc304f63),
	.w5(32'hbb83938e),
	.w6(32'hbbb323f1),
	.w7(32'hbb77cb97),
	.w8(32'hba996b0e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd60aca),
	.w1(32'hbb51fc6c),
	.w2(32'h3bb9267f),
	.w3(32'hbc586abb),
	.w4(32'hbb1380b3),
	.w5(32'hbb1bcc14),
	.w6(32'hbc1b1f8a),
	.w7(32'hbae9569a),
	.w8(32'h3ac37910),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dab5c),
	.w1(32'h3c4ba484),
	.w2(32'h3b49e350),
	.w3(32'hbb37a175),
	.w4(32'h3c4410b3),
	.w5(32'h3c5a786c),
	.w6(32'h3b07a28c),
	.w7(32'h3a2716cf),
	.w8(32'hbb19e797),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2332ff),
	.w1(32'h3b0d72d5),
	.w2(32'h3b6bdafb),
	.w3(32'h39a47de6),
	.w4(32'hbba15ac3),
	.w5(32'hbb5bbe2f),
	.w6(32'hbb6352cd),
	.w7(32'h3baf19b2),
	.w8(32'hbc13c4a6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a77e1),
	.w1(32'h3b215247),
	.w2(32'hba3aed2d),
	.w3(32'h394175c4),
	.w4(32'h3bc35572),
	.w5(32'h3c530ba0),
	.w6(32'hbc17b284),
	.w7(32'hbbcba7e7),
	.w8(32'hbc0daaa0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc095576),
	.w1(32'h3c0770b6),
	.w2(32'h3b97c0aa),
	.w3(32'hbc90efbe),
	.w4(32'h3c3aa834),
	.w5(32'h3c195d12),
	.w6(32'hbc2eb2f6),
	.w7(32'h3c426628),
	.w8(32'hb9e55cf6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcceb9),
	.w1(32'hbb82e7e8),
	.w2(32'hbb836c3f),
	.w3(32'hbc26c986),
	.w4(32'h3be7ad73),
	.w5(32'hba35e8f5),
	.w6(32'hbbcfab52),
	.w7(32'h3afd5829),
	.w8(32'h3bd2c010),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a0cf8),
	.w1(32'hbbb84c40),
	.w2(32'h3bffa80c),
	.w3(32'hbc48f304),
	.w4(32'hbc14533a),
	.w5(32'hb9544db1),
	.w6(32'hbb652c7c),
	.w7(32'hbc93c956),
	.w8(32'hbc0e319a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74765e),
	.w1(32'h3c54523b),
	.w2(32'h3aad25b1),
	.w3(32'h3cb7f7c8),
	.w4(32'h3c299b45),
	.w5(32'h3b8f961e),
	.w6(32'h3bb3f619),
	.w7(32'h3baa2bea),
	.w8(32'hbbb56d3d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843712),
	.w1(32'h3bbaf0de),
	.w2(32'hbc16da59),
	.w3(32'hbc57d00a),
	.w4(32'h3c1f9749),
	.w5(32'hbba7b282),
	.w6(32'hbc3b692e),
	.w7(32'h3c42695e),
	.w8(32'h3be8a643),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b79f),
	.w1(32'h3c56db71),
	.w2(32'hbb144cba),
	.w3(32'h3ab30f20),
	.w4(32'h3cea488f),
	.w5(32'hbb95b4a7),
	.w6(32'h38be3278),
	.w7(32'h3c89f84a),
	.w8(32'h3b971385),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6c305),
	.w1(32'hba9cb445),
	.w2(32'hbb3bb1b5),
	.w3(32'hbc2dcd7b),
	.w4(32'h3b1e7d30),
	.w5(32'hb9c930ed),
	.w6(32'hbbf01a08),
	.w7(32'hbb91c1bb),
	.w8(32'hbbeb19cc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf52e8b),
	.w1(32'h3a50bfa1),
	.w2(32'hbc0f251e),
	.w3(32'h3cb0c1cf),
	.w4(32'h3b59b4a7),
	.w5(32'hbbb72209),
	.w6(32'h3bfec362),
	.w7(32'h3b989b37),
	.w8(32'h3aa625a1),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffe26c),
	.w1(32'h3b1aa524),
	.w2(32'h3b91d4e7),
	.w3(32'hbbd06c70),
	.w4(32'hbb680b22),
	.w5(32'hb9446b9b),
	.w6(32'hbafc8b4a),
	.w7(32'hbbc77166),
	.w8(32'hbb248cb8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092d1c),
	.w1(32'h3b14985c),
	.w2(32'h39b67c4e),
	.w3(32'h3c8a287d),
	.w4(32'h3bdf41ae),
	.w5(32'h3b991e8f),
	.w6(32'h3c21bd48),
	.w7(32'hbb379863),
	.w8(32'hbb830066),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af958),
	.w1(32'hbbc543f6),
	.w2(32'hbc83895e),
	.w3(32'hbbbf052a),
	.w4(32'hbb8111cc),
	.w5(32'hbb644ab2),
	.w6(32'hbb9ef91b),
	.w7(32'hbc53e469),
	.w8(32'h3c1698a2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4fc5a),
	.w1(32'hbb824553),
	.w2(32'h3c4ed04e),
	.w3(32'hbce7df63),
	.w4(32'hbc35ba52),
	.w5(32'h3c2e4008),
	.w6(32'hbc261309),
	.w7(32'hbc2e4175),
	.w8(32'h3a1840b5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e0786),
	.w1(32'h3a88cff2),
	.w2(32'h3ae518c7),
	.w3(32'h3c0963b5),
	.w4(32'hbbc75ee5),
	.w5(32'h3c24285f),
	.w6(32'hbac036fe),
	.w7(32'hbaa28abf),
	.w8(32'h3bf830fd),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b67cc),
	.w1(32'h3c23d968),
	.w2(32'h3b9aec2a),
	.w3(32'hbc8cf59a),
	.w4(32'h3c835493),
	.w5(32'hba5e7028),
	.w6(32'hbc7f21ce),
	.w7(32'hba83b534),
	.w8(32'hbc6698a3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc886fac),
	.w1(32'h3a5b4865),
	.w2(32'hbcc34bf1),
	.w3(32'hbc9e467a),
	.w4(32'h3c8ac101),
	.w5(32'hbc5a3144),
	.w6(32'h3b1b76e3),
	.w7(32'h3c3065ea),
	.w8(32'hbca6c605),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef1443),
	.w1(32'h3c69e680),
	.w2(32'hbc8522b5),
	.w3(32'hbb209826),
	.w4(32'h3ca23f25),
	.w5(32'hbad08dbb),
	.w6(32'hbc3a8381),
	.w7(32'h3c969182),
	.w8(32'hbb3ec654),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30ebbf),
	.w1(32'hbc5685b1),
	.w2(32'h3a240710),
	.w3(32'h3a100b26),
	.w4(32'hbc8b88d2),
	.w5(32'hbba753a6),
	.w6(32'h3a53e722),
	.w7(32'hbc30b0ae),
	.w8(32'hbacc07a5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7baf7),
	.w1(32'h3c15cbe9),
	.w2(32'h3bb25d2f),
	.w3(32'hbc1c4889),
	.w4(32'h3bf21d45),
	.w5(32'h3ca5e867),
	.w6(32'hbba4091c),
	.w7(32'h39d25d80),
	.w8(32'hbcb0b45b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8feea5),
	.w1(32'h3b71ebd4),
	.w2(32'hbba0da20),
	.w3(32'hbcbb01e0),
	.w4(32'h3bae692f),
	.w5(32'hba901d38),
	.w6(32'hbc88107b),
	.w7(32'h3aaf26c8),
	.w8(32'hbb646b6f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3213d3),
	.w1(32'h3c82e05a),
	.w2(32'h3b6caa03),
	.w3(32'hbc9c1eab),
	.w4(32'h3cd214b0),
	.w5(32'hbb113330),
	.w6(32'hbc7f48b1),
	.w7(32'hbbb4ea8d),
	.w8(32'hbc8b1984),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca16fb4),
	.w1(32'hba20aa3b),
	.w2(32'h3c469720),
	.w3(32'hbc6214ba),
	.w4(32'hbbc5a27b),
	.w5(32'h3bd035ea),
	.w6(32'h3bc3fafb),
	.w7(32'hbc4e6609),
	.w8(32'hbb8e1cc8),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79265d),
	.w1(32'h3b9be3e9),
	.w2(32'h3aea3be0),
	.w3(32'h3cd8fc41),
	.w4(32'h3b37a11a),
	.w5(32'h3b881f82),
	.w6(32'h3c807ca6),
	.w7(32'hbc832c33),
	.w8(32'hbb72a798),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e6a6a),
	.w1(32'h3bff6dad),
	.w2(32'hba72cd34),
	.w3(32'hbc31e3b9),
	.w4(32'h3bd96681),
	.w5(32'h3b53c8a1),
	.w6(32'hbb9dae6f),
	.w7(32'h3be7d928),
	.w8(32'h3b2f9eb1),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11c02e),
	.w1(32'h3a906f94),
	.w2(32'hbb8da9d4),
	.w3(32'hbc55a709),
	.w4(32'h3b8bdf8f),
	.w5(32'h3be5bf37),
	.w6(32'hbc696dd3),
	.w7(32'h3c3960e2),
	.w8(32'hbb8d3a6a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5671eae),
	.w1(32'hba9cc241),
	.w2(32'h3b57058b),
	.w3(32'hbb83720d),
	.w4(32'h3b1abd06),
	.w5(32'h3afe693c),
	.w6(32'hbc1e2499),
	.w7(32'h3b1eecbf),
	.w8(32'h3ba4fc1b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51c27b),
	.w1(32'hbae01fd4),
	.w2(32'hbb9f3355),
	.w3(32'hbbb4e88b),
	.w4(32'hbbb74a2b),
	.w5(32'h3a034371),
	.w6(32'h3a9ffcbf),
	.w7(32'hbbe019f1),
	.w8(32'h3c19405b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbded95),
	.w1(32'hbba14916),
	.w2(32'hbb42ac17),
	.w3(32'h3c38f27b),
	.w4(32'hbc47e78c),
	.w5(32'h3ba5ceac),
	.w6(32'h3bb4e439),
	.w7(32'hbbee443c),
	.w8(32'h3ab8e9c8),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb02a9),
	.w1(32'hbc05b358),
	.w2(32'h3ac9d63b),
	.w3(32'h3c88bc58),
	.w4(32'hbb0897f7),
	.w5(32'h3c9aa2cd),
	.w6(32'h3bb0b326),
	.w7(32'hbb1ebbfb),
	.w8(32'h3bdbcee9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa930fe),
	.w1(32'h39be91f7),
	.w2(32'hbbf07fd3),
	.w3(32'hbc3d9947),
	.w4(32'h3abfcc69),
	.w5(32'h39d22c73),
	.w6(32'hba0ce4f4),
	.w7(32'h37dc5e9d),
	.w8(32'hbb29898b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ee3ce),
	.w1(32'hbaadba5a),
	.w2(32'hba7baa56),
	.w3(32'hbc2c8212),
	.w4(32'h3bc941db),
	.w5(32'hbc24c784),
	.w6(32'hba9e6059),
	.w7(32'hbafc0d13),
	.w8(32'hbac5cb38),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a219456),
	.w1(32'hbb3e7ced),
	.w2(32'h3af53836),
	.w3(32'hbbeab033),
	.w4(32'hbba5e20d),
	.w5(32'h3bedcafe),
	.w6(32'h3b095aa0),
	.w7(32'hbbc9631d),
	.w8(32'h3b7213d7),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d24e7),
	.w1(32'h3c69bca0),
	.w2(32'h3b81ed66),
	.w3(32'hbb827945),
	.w4(32'h3c340dd9),
	.w5(32'h3c0229fd),
	.w6(32'hbb5a2626),
	.w7(32'h3c822498),
	.w8(32'hbc14269d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37442a),
	.w1(32'h3be791c8),
	.w2(32'h3be27a26),
	.w3(32'hbb3c4c0a),
	.w4(32'h3bcec230),
	.w5(32'h3c8356eb),
	.w6(32'hbc71a2fe),
	.w7(32'h3b7d9482),
	.w8(32'h3ab8602d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb761ce1),
	.w1(32'h3b55e1a1),
	.w2(32'hbc3e70e8),
	.w3(32'hbc3d801e),
	.w4(32'h39db4c9e),
	.w5(32'h3b6967c0),
	.w6(32'hbc2fff18),
	.w7(32'h3a9c3870),
	.w8(32'hbc2a7fdc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69416e),
	.w1(32'h3ae5da48),
	.w2(32'h3adcbe64),
	.w3(32'hbbdc8e4e),
	.w4(32'hbc276682),
	.w5(32'h3a176a9f),
	.w6(32'hbc1a2342),
	.w7(32'hbb2994bc),
	.w8(32'h3c229e64),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90118e),
	.w1(32'h3b5f35b9),
	.w2(32'h3b22a9e0),
	.w3(32'h3b13d450),
	.w4(32'h3aad65ca),
	.w5(32'h3bfb8b7f),
	.w6(32'h3bd620f2),
	.w7(32'h3b373cd7),
	.w8(32'hbb808a0d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c0b21),
	.w1(32'h3beaccef),
	.w2(32'hbc0db416),
	.w3(32'hbc263231),
	.w4(32'h3c4a295a),
	.w5(32'hba847966),
	.w6(32'hbc158e09),
	.w7(32'h3b8ad411),
	.w8(32'hbb9e1db0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1f30c),
	.w1(32'hbb7acaec),
	.w2(32'hbbc7bfc3),
	.w3(32'h3aa649ed),
	.w4(32'h3aeabea6),
	.w5(32'h3be17b49),
	.w6(32'hbb566cbf),
	.w7(32'h3b259811),
	.w8(32'hbbd5c577),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841831),
	.w1(32'h3b85bc1e),
	.w2(32'hbb4cbe1e),
	.w3(32'hbb785ed1),
	.w4(32'h3c2811d5),
	.w5(32'hbc212f59),
	.w6(32'hbc4e42b5),
	.w7(32'h3c254fda),
	.w8(32'hbb5e4790),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc988147),
	.w1(32'h39afa9d7),
	.w2(32'h3c29e621),
	.w3(32'hbccd8171),
	.w4(32'hbbca00a3),
	.w5(32'h3c3bd821),
	.w6(32'hbc52e521),
	.w7(32'h3b34a016),
	.w8(32'h3c26a575),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b40e2),
	.w1(32'hbbbf1e8f),
	.w2(32'h3bbd8277),
	.w3(32'h3c990bfa),
	.w4(32'hbcb3affc),
	.w5(32'h3c287a5a),
	.w6(32'h3b1bf8b0),
	.w7(32'hbc05a4ff),
	.w8(32'h3b1a8406),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d817d),
	.w1(32'h3c166be6),
	.w2(32'hbb3d8dcb),
	.w3(32'h3d433dac),
	.w4(32'h3c82cbc1),
	.w5(32'hbc1eb85e),
	.w6(32'h3bb43d28),
	.w7(32'h3c463499),
	.w8(32'hbc58cccc),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73bec7),
	.w1(32'hbbecf1c6),
	.w2(32'hbc4136ae),
	.w3(32'hbbe66d26),
	.w4(32'h3c31fc3e),
	.w5(32'h3c17ed44),
	.w6(32'hba7a44be),
	.w7(32'h3b7e0b6b),
	.w8(32'hb992cff2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9737b),
	.w1(32'hbb45217b),
	.w2(32'h3a641758),
	.w3(32'hbd032124),
	.w4(32'hbc0c7194),
	.w5(32'h3b9538e6),
	.w6(32'hbcba497e),
	.w7(32'hbc895416),
	.w8(32'h3b98685d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48cdb0),
	.w1(32'h3b21f6ed),
	.w2(32'h3b7b2fe9),
	.w3(32'h3ca3c64a),
	.w4(32'hbc0b8a34),
	.w5(32'h3bfc0e23),
	.w6(32'h3c7013fb),
	.w7(32'hbc6904a0),
	.w8(32'hbb95ce32),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed76ae),
	.w1(32'h3ba36823),
	.w2(32'hbbb74616),
	.w3(32'h3a55b76a),
	.w4(32'h3c754cd2),
	.w5(32'h3b1e27e1),
	.w6(32'hbc3ce9a6),
	.w7(32'h3c216cd9),
	.w8(32'h3abe1674),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fe3a0),
	.w1(32'h3b6d9708),
	.w2(32'hbbab3359),
	.w3(32'hbc376d98),
	.w4(32'h3bd3f674),
	.w5(32'h3b76c725),
	.w6(32'hbb347bc1),
	.w7(32'h3c04c5f6),
	.w8(32'hba8b54b1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc272ee8),
	.w1(32'h394a66df),
	.w2(32'h3bdf954b),
	.w3(32'hbc002bb0),
	.w4(32'hbbf0736e),
	.w5(32'hbb770505),
	.w6(32'hbc6ed1b9),
	.w7(32'hbc42a801),
	.w8(32'hb87000dd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2035e6),
	.w1(32'hbc427384),
	.w2(32'hbc8ccea7),
	.w3(32'hbb408775),
	.w4(32'h3c4b3b8c),
	.w5(32'hbc046455),
	.w6(32'h3bc02abc),
	.w7(32'h3c9d18c1),
	.w8(32'hbc2aa635),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc815003),
	.w1(32'hbceb2560),
	.w2(32'hbcd33499),
	.w3(32'hbc6ebc68),
	.w4(32'hbca610f0),
	.w5(32'hbcbcb730),
	.w6(32'hbc4dee41),
	.w7(32'hbcaa05b4),
	.w8(32'hbc91c730),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc083504),
	.w1(32'h3b956f7d),
	.w2(32'hbc496f60),
	.w3(32'hbc9fa0a2),
	.w4(32'h3c487931),
	.w5(32'hbc873449),
	.w6(32'hbc2e0f23),
	.w7(32'h3b5821f2),
	.w8(32'hbaa88db2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31eea1),
	.w1(32'h3b8e25ab),
	.w2(32'hbb719749),
	.w3(32'hbcc07a84),
	.w4(32'h3c6107f5),
	.w5(32'h3bd9bc21),
	.w6(32'hbbeb3f8d),
	.w7(32'h3b7575fb),
	.w8(32'hbc0a34fb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb207ef0),
	.w1(32'h3b42ace9),
	.w2(32'h3b607319),
	.w3(32'hbc5cf0d6),
	.w4(32'h3b5ca0c6),
	.w5(32'h3a9c5aa9),
	.w6(32'hbc1104da),
	.w7(32'h3bd12216),
	.w8(32'hbb612f57),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41c8ac),
	.w1(32'h3cb73e66),
	.w2(32'hbbad1ccf),
	.w3(32'hbb831d5a),
	.w4(32'h3ca338ee),
	.w5(32'h3c03d727),
	.w6(32'hbc02c8e1),
	.w7(32'h3c92c744),
	.w8(32'hbc0897d5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca3eb2),
	.w1(32'hbc038c25),
	.w2(32'hba8929d7),
	.w3(32'hbc9f0e5b),
	.w4(32'hbc068561),
	.w5(32'hbbd5489f),
	.w6(32'hbc928194),
	.w7(32'hbc2cd693),
	.w8(32'h3aff2226),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffbd16),
	.w1(32'hbcffba04),
	.w2(32'h3b4eb7e1),
	.w3(32'h3c179d50),
	.w4(32'hbd2dc4c9),
	.w5(32'h3c404020),
	.w6(32'h3c22d014),
	.w7(32'hbd113dd5),
	.w8(32'hbaacb9c4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2171f3),
	.w1(32'hbbe04d0e),
	.w2(32'h3b22c275),
	.w3(32'h3d6105d6),
	.w4(32'hbc11ff88),
	.w5(32'h3b8d89a1),
	.w6(32'h3d0c8ba3),
	.w7(32'hbb32228f),
	.w8(32'hba715ea8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f80e5),
	.w1(32'hbb97e61b),
	.w2(32'h3a8f166c),
	.w3(32'h3c7f76e1),
	.w4(32'h3ad6a006),
	.w5(32'hbbf3f39b),
	.w6(32'h3bd9888b),
	.w7(32'h3a014cdc),
	.w8(32'hba0bb65b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd111db),
	.w1(32'h3ca152ef),
	.w2(32'hbc22f80f),
	.w3(32'hbc60aabe),
	.w4(32'h3cc93f1e),
	.w5(32'hbc6371b6),
	.w6(32'hbbc505a5),
	.w7(32'h3cc05aa0),
	.w8(32'hbbadda1a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc912bc),
	.w1(32'h3bcb0b3a),
	.w2(32'hbbc4bfb8),
	.w3(32'hbcab63ed),
	.w4(32'h3c86eaec),
	.w5(32'hbc56b380),
	.w6(32'hbc2456ce),
	.w7(32'h3bbf1813),
	.w8(32'hbc2a2d25),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcacd65e),
	.w1(32'h3778138d),
	.w2(32'h3bb8d63b),
	.w3(32'hbce55ff6),
	.w4(32'hbb9f96cc),
	.w5(32'h3bf60b7c),
	.w6(32'hbcb04069),
	.w7(32'h3b8dcb91),
	.w8(32'h3bcef5f1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1775ab),
	.w1(32'h3b3fdb61),
	.w2(32'hba916199),
	.w3(32'h3c475c80),
	.w4(32'h3a884e02),
	.w5(32'hbc4bee6b),
	.w6(32'h3ae66db7),
	.w7(32'hbbae2eb0),
	.w8(32'hbb70f02e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba817a9a),
	.w1(32'h3c3ad772),
	.w2(32'h3cca00c3),
	.w3(32'h3a400b33),
	.w4(32'h3c59deae),
	.w5(32'h3cea2d0e),
	.w6(32'h3a80b6ea),
	.w7(32'h3c9272bf),
	.w8(32'h3bea3956),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cab15),
	.w1(32'h3aa35def),
	.w2(32'h3c0a7d9a),
	.w3(32'h3c2da4b2),
	.w4(32'h38480a3b),
	.w5(32'h3c743a3a),
	.w6(32'h3ad51175),
	.w7(32'h3b4635e9),
	.w8(32'h3c2ae744),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb223f78),
	.w1(32'hb98a5661),
	.w2(32'h3b1b47cf),
	.w3(32'h3a4bad6c),
	.w4(32'hbaf6be4e),
	.w5(32'h3b2f2da2),
	.w6(32'h3bac655c),
	.w7(32'hba229e92),
	.w8(32'hb9d1c9c6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb646ec5),
	.w1(32'h3b9b640a),
	.w2(32'hba14fcfa),
	.w3(32'hbbf9ea03),
	.w4(32'h3aff014c),
	.w5(32'h3c38d37f),
	.w6(32'hbb8313bd),
	.w7(32'h3a59f106),
	.w8(32'hbaa80b06),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2fe23),
	.w1(32'hbc7728d0),
	.w2(32'hbc1f4d6b),
	.w3(32'hba957c85),
	.w4(32'hbc440eac),
	.w5(32'hbb8cf6bc),
	.w6(32'h3b166929),
	.w7(32'h38eeb637),
	.w8(32'hba0cc35a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cf254),
	.w1(32'h3a942697),
	.w2(32'h3bd413df),
	.w3(32'hbadac7ea),
	.w4(32'h3bbc957f),
	.w5(32'h3bf92e61),
	.w6(32'hbb1b7c10),
	.w7(32'h3ba54698),
	.w8(32'h3c38fe08),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae62e),
	.w1(32'hbc80517e),
	.w2(32'hbb929faa),
	.w3(32'hbbda908c),
	.w4(32'hbc88e35b),
	.w5(32'hbbf79a4a),
	.w6(32'hbb5d3dd0),
	.w7(32'hbbca73ef),
	.w8(32'hbc45ab6c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb73433),
	.w1(32'hbbe8e7c9),
	.w2(32'hbaa48743),
	.w3(32'hbc9ae99c),
	.w4(32'hbc39020b),
	.w5(32'hbbc56af7),
	.w6(32'hbc700c21),
	.w7(32'hbb4fd675),
	.w8(32'hbb2d252c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa45f49),
	.w1(32'h3a88c411),
	.w2(32'hbbeb6b34),
	.w3(32'hbbbb16a5),
	.w4(32'h3b34de94),
	.w5(32'h3c0f2991),
	.w6(32'hbb95b0c1),
	.w7(32'hbbd1888b),
	.w8(32'hba8374d2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb4e77),
	.w1(32'h3b63d65b),
	.w2(32'h3b77fffa),
	.w3(32'hbb11f8a4),
	.w4(32'hb9ca7cc3),
	.w5(32'h3aaf1741),
	.w6(32'h3bb2d9d2),
	.w7(32'h3b7e6445),
	.w8(32'h3b8f89c6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838bd5),
	.w1(32'h3b3f260e),
	.w2(32'hbbcc435a),
	.w3(32'h3a9b62a2),
	.w4(32'h3b8d2852),
	.w5(32'hbbee8071),
	.w6(32'h3b33fd4b),
	.w7(32'h3bbae24a),
	.w8(32'hbb9458f8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3fcd4),
	.w1(32'hb8c5f6ba),
	.w2(32'h37fac1ea),
	.w3(32'h3bb0f8e2),
	.w4(32'hba77c3a5),
	.w5(32'hbbffd5c7),
	.w6(32'h3af3db2b),
	.w7(32'hbb4ad38a),
	.w8(32'hbaf3a96b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34c1fc),
	.w1(32'h3b6af079),
	.w2(32'h3be95a45),
	.w3(32'h3afc2a56),
	.w4(32'hbad086aa),
	.w5(32'hba05b894),
	.w6(32'h3b1c5b90),
	.w7(32'hbadf3da8),
	.w8(32'hbb0d5420),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd638aa),
	.w1(32'h3bae2173),
	.w2(32'hbbebb849),
	.w3(32'hbc10c76f),
	.w4(32'h3c3bd7a9),
	.w5(32'hbc4db638),
	.w6(32'hbb5951a5),
	.w7(32'h3c5b4770),
	.w8(32'hbc2aa8d2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c392f62),
	.w1(32'hbc158f19),
	.w2(32'h3b8f2f7c),
	.w3(32'hba9b2196),
	.w4(32'hbbb8a6de),
	.w5(32'h3bd938c7),
	.w6(32'h3a85c88f),
	.w7(32'hbc17a2d2),
	.w8(32'h3a63402b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7ee08),
	.w1(32'h3cd3eea4),
	.w2(32'h3c941d2f),
	.w3(32'h3b7d8c8b),
	.w4(32'h3c8df9ee),
	.w5(32'h3c454817),
	.w6(32'h3aa7f556),
	.w7(32'h3c38ba93),
	.w8(32'h3bb40e55),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a398c),
	.w1(32'h3c9ef346),
	.w2(32'h3c4e9c24),
	.w3(32'h3c0a7e4a),
	.w4(32'h3c4d7002),
	.w5(32'h3c80575c),
	.w6(32'h3c9b6515),
	.w7(32'h399f6001),
	.w8(32'h3cac77ce),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79b9a7),
	.w1(32'hbb16779a),
	.w2(32'h3b9c1159),
	.w3(32'h3c503ad3),
	.w4(32'h3c0952d1),
	.w5(32'hbbaac20c),
	.w6(32'h3cd19944),
	.w7(32'hba53c037),
	.w8(32'hb814fdcd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac957d),
	.w1(32'h3be0dfea),
	.w2(32'h3b5018d6),
	.w3(32'hbb35f6c4),
	.w4(32'h3b7164e0),
	.w5(32'h3be96cd6),
	.w6(32'hbb4d3608),
	.w7(32'h399d8909),
	.w8(32'h3be26d84),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab775c4),
	.w1(32'h3a08f3bd),
	.w2(32'h388f21a7),
	.w3(32'hbbc1e998),
	.w4(32'h3c03941a),
	.w5(32'h3b87f7e1),
	.w6(32'h3a025508),
	.w7(32'h39f9d5da),
	.w8(32'h3b6578d9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53b838),
	.w1(32'h3bb0f822),
	.w2(32'h3b25983d),
	.w3(32'h3a862e14),
	.w4(32'hbb1f1887),
	.w5(32'hbc225b2a),
	.w6(32'h3b873c82),
	.w7(32'h3a109898),
	.w8(32'h3b44cee2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5086b5),
	.w1(32'h3a714cff),
	.w2(32'h3b279d06),
	.w3(32'hbb76bb21),
	.w4(32'hbb236c73),
	.w5(32'h3ba4192b),
	.w6(32'hbae5550c),
	.w7(32'h3b70358b),
	.w8(32'h385c02bc),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18164e),
	.w1(32'hb8483e35),
	.w2(32'h3b186453),
	.w3(32'h3b7cb2bf),
	.w4(32'hbb26f7cc),
	.w5(32'hbb9f5877),
	.w6(32'hbac50828),
	.w7(32'h3b114f89),
	.w8(32'h3b76833c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e2166),
	.w1(32'h3bb01ea1),
	.w2(32'h3af14247),
	.w3(32'hbbd550db),
	.w4(32'h3bde8b3f),
	.w5(32'h3abbeb5f),
	.w6(32'h3ac8aa43),
	.w7(32'hbbf21a94),
	.w8(32'h3ba34c8a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14a51c),
	.w1(32'hbc9cd51b),
	.w2(32'hbadfed39),
	.w3(32'hbbc096fd),
	.w4(32'hbc500de8),
	.w5(32'h3caedc72),
	.w6(32'h3b2b44d4),
	.w7(32'hbbb87ce8),
	.w8(32'h38513c89),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bcbc7),
	.w1(32'h3bb6bc90),
	.w2(32'hbc13e30e),
	.w3(32'hbcb3a620),
	.w4(32'h3c0b077b),
	.w5(32'hbc5f48ff),
	.w6(32'hbc4f4cf8),
	.w7(32'h3baa5742),
	.w8(32'h3bc3f73a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e605),
	.w1(32'h3c17a123),
	.w2(32'h3ba736c2),
	.w3(32'h3c96de87),
	.w4(32'h3b90acef),
	.w5(32'h3c0dcda3),
	.w6(32'h3c7b6fc0),
	.w7(32'h3a13a5fc),
	.w8(32'h3b517233),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d09b1),
	.w1(32'hbb442421),
	.w2(32'h3a58b343),
	.w3(32'hbaf3ae5f),
	.w4(32'hbb6a226c),
	.w5(32'hba95ebe2),
	.w6(32'h3a998231),
	.w7(32'hbad760d5),
	.w8(32'h3b5258b3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a654d),
	.w1(32'hbaa413b0),
	.w2(32'h3ac6d085),
	.w3(32'h3c4ea00c),
	.w4(32'h39b363be),
	.w5(32'hbb2de3ba),
	.w6(32'h3af2b997),
	.w7(32'h3b46fc7b),
	.w8(32'h3b19857e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39cbb1),
	.w1(32'h3be4c4d3),
	.w2(32'h3b04616a),
	.w3(32'hbb5d499e),
	.w4(32'h3c175c53),
	.w5(32'hbb024941),
	.w6(32'hba7d2afc),
	.w7(32'h3b5f658b),
	.w8(32'h3beda953),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5baf1),
	.w1(32'h3bc1d515),
	.w2(32'h3a8dc743),
	.w3(32'hbba6275c),
	.w4(32'h3c58d7ab),
	.w5(32'hbc99d45c),
	.w6(32'h3c42e88e),
	.w7(32'h3c6e33e1),
	.w8(32'hbbd2c7ed),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97eb40),
	.w1(32'hbc6d7246),
	.w2(32'hbab750d1),
	.w3(32'h3c75d8f9),
	.w4(32'hbc3f0e99),
	.w5(32'h3c04601c),
	.w6(32'h3c362c83),
	.w7(32'hbc295515),
	.w8(32'hbb790071),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a78db),
	.w1(32'hbc2d5d11),
	.w2(32'hbb68889c),
	.w3(32'hbc06f8a2),
	.w4(32'hbb41a2e4),
	.w5(32'hbbddc97e),
	.w6(32'hbc7102aa),
	.w7(32'hb8113bed),
	.w8(32'hbb3cb7d1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0a8c6),
	.w1(32'hbc3a6da6),
	.w2(32'hbb7214cf),
	.w3(32'hbc4e7eaf),
	.w4(32'hbc78730a),
	.w5(32'hbb1eb983),
	.w6(32'hbb7facda),
	.w7(32'hbc6a8ada),
	.w8(32'hba3e31fb),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb435e5f),
	.w1(32'hbb4a5b5e),
	.w2(32'hbb9070bb),
	.w3(32'hbb534939),
	.w4(32'hba85b70a),
	.w5(32'hbbce3943),
	.w6(32'hbc2dd331),
	.w7(32'hbb98dbc6),
	.w8(32'h3a4eb4be),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb710a94),
	.w1(32'hbb4dd2c3),
	.w2(32'h3981b931),
	.w3(32'h3b44191c),
	.w4(32'hbb9e00b7),
	.w5(32'hbb4389db),
	.w6(32'h3abd1db1),
	.w7(32'hbbeb32a8),
	.w8(32'hbb801b70),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf74fb),
	.w1(32'h39d12684),
	.w2(32'hbb24d7ab),
	.w3(32'h3aa50943),
	.w4(32'hbb8ffbd2),
	.w5(32'hbb847a7a),
	.w6(32'hbc0de717),
	.w7(32'hbb8c67ba),
	.w8(32'hbbded746),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87efea),
	.w1(32'h3a074a14),
	.w2(32'hb9a9c788),
	.w3(32'h3c13f49c),
	.w4(32'hbacf331d),
	.w5(32'h3c21b791),
	.w6(32'h3aeb57c1),
	.w7(32'h3ba569b2),
	.w8(32'h3baab2ce),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb304b6),
	.w1(32'hbc3d7da9),
	.w2(32'hbb6ab5d0),
	.w3(32'h3c806bd1),
	.w4(32'hbc82a0cb),
	.w5(32'h3b4d0c8c),
	.w6(32'h3b2e9956),
	.w7(32'hbc6d39c1),
	.w8(32'hbaf8ce61),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc211cad),
	.w1(32'hbae9aa93),
	.w2(32'hbadf3d52),
	.w3(32'hbcb9a89d),
	.w4(32'hbb388802),
	.w5(32'h3b8c0728),
	.w6(32'hbc07563f),
	.w7(32'h3a52fec0),
	.w8(32'hbaf26bd4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb707d03),
	.w1(32'hbc1bf69f),
	.w2(32'hbba9a5c2),
	.w3(32'hbb1bfe40),
	.w4(32'hba9197e8),
	.w5(32'hbc01978f),
	.w6(32'hbc0ff7dd),
	.w7(32'hbba26912),
	.w8(32'hbbd74e16),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dedbfd),
	.w1(32'h3c387923),
	.w2(32'h3a77f3ed),
	.w3(32'h3b6e3381),
	.w4(32'h3c921c0b),
	.w5(32'h3c119fd7),
	.w6(32'hbae1a171),
	.w7(32'h3c29fa90),
	.w8(32'h39455d85),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7306b3),
	.w1(32'h3be19042),
	.w2(32'h3c48ae4a),
	.w3(32'h39405761),
	.w4(32'h3bf995ce),
	.w5(32'h3a7875c2),
	.w6(32'hbb05a5a1),
	.w7(32'h3b90c5d2),
	.w8(32'h3a66b056),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3ab7d),
	.w1(32'h3c1702fb),
	.w2(32'h3beb758e),
	.w3(32'h3af830f9),
	.w4(32'h3a6ab168),
	.w5(32'h3b4cf1f9),
	.w6(32'h3a86eba9),
	.w7(32'hbb20e3d0),
	.w8(32'hbb156d29),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de1665),
	.w1(32'hba446161),
	.w2(32'hbbabf81d),
	.w3(32'hbbaba363),
	.w4(32'h3a5dd4b7),
	.w5(32'hbbba5f85),
	.w6(32'hbb06610b),
	.w7(32'h3b44fa5a),
	.w8(32'h3b8b6bf1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cba65),
	.w1(32'h3ba0d8f1),
	.w2(32'hbb6b455a),
	.w3(32'h3c05f4ca),
	.w4(32'h3c504fce),
	.w5(32'h3b6d39af),
	.w6(32'h3be1f269),
	.w7(32'h3a2d53f6),
	.w8(32'h3acb372f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921c22c),
	.w1(32'h3ae1eb12),
	.w2(32'hba0453b9),
	.w3(32'hbb6538d6),
	.w4(32'hbab92150),
	.w5(32'hba5b811b),
	.w6(32'hbb0ec06d),
	.w7(32'hbbcbeb07),
	.w8(32'h3b9322ce),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad06310),
	.w1(32'h3b98b6e6),
	.w2(32'h3b26ba9d),
	.w3(32'h3b1c060b),
	.w4(32'hb9f0e2e6),
	.w5(32'h3a9f96cb),
	.w6(32'h3bb0f238),
	.w7(32'hbb790546),
	.w8(32'h39bed897),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9efb1),
	.w1(32'hbc10fd4f),
	.w2(32'h3bafa042),
	.w3(32'h371a5a79),
	.w4(32'hba4c012b),
	.w5(32'h3d0583b8),
	.w6(32'h3b511956),
	.w7(32'hb9299dfa),
	.w8(32'h3b6a6801),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5207f),
	.w1(32'h3b8496c4),
	.w2(32'hb981a8dc),
	.w3(32'hbb27c5fb),
	.w4(32'h3ab0131f),
	.w5(32'hbb7d03c1),
	.w6(32'hbbbe29e7),
	.w7(32'h3b345439),
	.w8(32'h3b7f40c5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16ae94),
	.w1(32'hbbcc9e91),
	.w2(32'hbc214773),
	.w3(32'hbbe979ca),
	.w4(32'hb748bcbe),
	.w5(32'hba897967),
	.w6(32'hba3e30bd),
	.w7(32'h3aa558c5),
	.w8(32'h3bae65c7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af29a3b),
	.w1(32'h3c4cb733),
	.w2(32'h3bada774),
	.w3(32'h3c190be9),
	.w4(32'h3c5c9d2d),
	.w5(32'hbbe54fdf),
	.w6(32'h39d8cac9),
	.w7(32'h3b823826),
	.w8(32'h3b5dc040),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dfe24),
	.w1(32'hb7e0a483),
	.w2(32'hbada87fa),
	.w3(32'h3c606568),
	.w4(32'h3be2fa2e),
	.w5(32'hbbecd3a9),
	.w6(32'h3c3fdbe8),
	.w7(32'h3b8181b7),
	.w8(32'hbbdae33a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b241d53),
	.w1(32'h3c43fe1e),
	.w2(32'h3c6b9d2a),
	.w3(32'h3bd4046d),
	.w4(32'h3c9f8bfe),
	.w5(32'h3cca02d4),
	.w6(32'hba4551de),
	.w7(32'h3cb2e8a4),
	.w8(32'h3c510981),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d81c),
	.w1(32'h3a2d189a),
	.w2(32'hbade8492),
	.w3(32'h3cb46414),
	.w4(32'h3a19a5b9),
	.w5(32'hba1ac0d0),
	.w6(32'h3c1970e2),
	.w7(32'h3bd859e8),
	.w8(32'h39e66c28),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb384f80),
	.w1(32'hbbd9e6a3),
	.w2(32'hba4c13e0),
	.w3(32'hbc13f80a),
	.w4(32'h3c071eb0),
	.w5(32'h3b03dce8),
	.w6(32'hbc4c06ef),
	.w7(32'hbb9d2356),
	.w8(32'h3b801e96),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b999725),
	.w1(32'hbbd6f09e),
	.w2(32'hba436a07),
	.w3(32'h3bef726e),
	.w4(32'hbaea78ac),
	.w5(32'h396f3eed),
	.w6(32'h3c1d49f3),
	.w7(32'hbb9332df),
	.w8(32'hbba123c3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule