module layer_10_featuremap_482(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba995004),
	.w1(32'h3ab9a405),
	.w2(32'h3af20015),
	.w3(32'hb92f1a3b),
	.w4(32'h3b06a39e),
	.w5(32'h3b05751c),
	.w6(32'hb8f82fef),
	.w7(32'h3a945a7d),
	.w8(32'h3aa5e744),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b183f39),
	.w1(32'hba6d0327),
	.w2(32'h36068997),
	.w3(32'h3b1f2b31),
	.w4(32'hba5cf483),
	.w5(32'hba7632a4),
	.w6(32'h3a8d94db),
	.w7(32'hba1870be),
	.w8(32'hba518d3a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6d658),
	.w1(32'hbad18318),
	.w2(32'hbafe4835),
	.w3(32'hba318737),
	.w4(32'hbae20250),
	.w5(32'hbb2d50e5),
	.w6(32'hb901583a),
	.w7(32'hba994def),
	.w8(32'hb8845f15),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb009ab7),
	.w1(32'hb9b2d70c),
	.w2(32'hba39380f),
	.w3(32'hba845893),
	.w4(32'hb919dece),
	.w5(32'h3a978ea6),
	.w6(32'h39d60da0),
	.w7(32'h399c85f5),
	.w8(32'h388249f5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9480947),
	.w1(32'h3a541820),
	.w2(32'h3a47ea7d),
	.w3(32'h38fe21aa),
	.w4(32'h3a183bd7),
	.w5(32'hb9017252),
	.w6(32'h393a90cb),
	.w7(32'h397cd7fa),
	.w8(32'h354a2d6a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bc8c8),
	.w1(32'hba76b5dc),
	.w2(32'h39aa8f8f),
	.w3(32'hb8b8bea6),
	.w4(32'hb92f9e9d),
	.w5(32'hbb0e3a09),
	.w6(32'h39c3c4d9),
	.w7(32'hba8553c1),
	.w8(32'hba31a360),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50226a),
	.w1(32'h3a6ed60d),
	.w2(32'hb9af0eb7),
	.w3(32'hba9bc351),
	.w4(32'hb90dde1c),
	.w5(32'h3b4a036c),
	.w6(32'hba9fa212),
	.w7(32'h392c4fbd),
	.w8(32'h3a937ab2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a417185),
	.w1(32'hb9f5c4cd),
	.w2(32'hbafbdf8b),
	.w3(32'h3accea3d),
	.w4(32'hbab5bdf8),
	.w5(32'hbb2b5469),
	.w6(32'h388fd7f2),
	.w7(32'h3ace45e3),
	.w8(32'h3aba69f6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7376dd),
	.w1(32'hbaa75648),
	.w2(32'hb9d29a52),
	.w3(32'hba5975da),
	.w4(32'hbac06de0),
	.w5(32'h3a4161d1),
	.w6(32'h3aba8c2c),
	.w7(32'h38c08ca2),
	.w8(32'h3a894e05),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963c2e1),
	.w1(32'h3b1f2754),
	.w2(32'h3afef733),
	.w3(32'hba6f0453),
	.w4(32'h3a826b76),
	.w5(32'h3b215ec9),
	.w6(32'hbad2fc7e),
	.w7(32'hb90a21ad),
	.w8(32'h3a3c7bb3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08d30d),
	.w1(32'hba820fcb),
	.w2(32'hba5678e7),
	.w3(32'hb9a4a45e),
	.w4(32'h39d46325),
	.w5(32'h398d9c0a),
	.w6(32'hb8af4893),
	.w7(32'hb99e865e),
	.w8(32'hba34c2e0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381366f2),
	.w1(32'h39b8afdf),
	.w2(32'hb90ce532),
	.w3(32'h39a09e7a),
	.w4(32'h3a3d884f),
	.w5(32'hb9f2fb85),
	.w6(32'h39a02fde),
	.w7(32'h39f3e7e0),
	.w8(32'h3a783187),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa193a0),
	.w1(32'h39700ac3),
	.w2(32'h3a8f66c1),
	.w3(32'hba4d467e),
	.w4(32'hba78d15b),
	.w5(32'h3a9409ba),
	.w6(32'hba4f8867),
	.w7(32'hbb0ecb36),
	.w8(32'hba1b0e98),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba081d02),
	.w1(32'hb9d0a4d8),
	.w2(32'hba008a8f),
	.w3(32'hb9c065e9),
	.w4(32'hba8e082e),
	.w5(32'hbace397d),
	.w6(32'h3a9be14e),
	.w7(32'hba8621f6),
	.w8(32'hba9c8b64),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66f409),
	.w1(32'hb9db849a),
	.w2(32'hba698dce),
	.w3(32'hb9e73200),
	.w4(32'hb9f2c7ca),
	.w5(32'hba84d384),
	.w6(32'hba03afa8),
	.w7(32'hba3338f7),
	.w8(32'hb7dade79),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba226894),
	.w1(32'hb9ecbf89),
	.w2(32'hb8a4085d),
	.w3(32'hbb11f50b),
	.w4(32'hba73294b),
	.w5(32'h38b609fc),
	.w6(32'hbaf3b9c8),
	.w7(32'hba811420),
	.w8(32'h3a8fa9c3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79f54a),
	.w1(32'h39dfa309),
	.w2(32'hb9490b5d),
	.w3(32'hba8bf2a3),
	.w4(32'h39b4bddf),
	.w5(32'h3a747f1b),
	.w6(32'h39e1afb4),
	.w7(32'hb944b071),
	.w8(32'h3ae2b3c1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa140d1),
	.w1(32'h3a512fd0),
	.w2(32'h3ae35bb9),
	.w3(32'hba6f7553),
	.w4(32'h3aaf41d6),
	.w5(32'h3ab47269),
	.w6(32'h3a778531),
	.w7(32'h3a70a617),
	.w8(32'h3a3d6f5f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a419618),
	.w1(32'hb8f98988),
	.w2(32'hbad71e78),
	.w3(32'h3990010a),
	.w4(32'hbaa104ed),
	.w5(32'hba986511),
	.w6(32'h3a2620d5),
	.w7(32'hba22fac6),
	.w8(32'hb91f3150),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba921ff3),
	.w1(32'h38bd58e8),
	.w2(32'hb951b8af),
	.w3(32'hba707f2c),
	.w4(32'hba68e2ac),
	.w5(32'hb98c7ee1),
	.w6(32'hba10a945),
	.w7(32'h3a22a518),
	.w8(32'h3a3a03df),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e19bee),
	.w1(32'hbabe0f4b),
	.w2(32'hbab24763),
	.w3(32'hbae5b803),
	.w4(32'hb98a45dd),
	.w5(32'hbacb0990),
	.w6(32'hbacdb094),
	.w7(32'hb9cab28c),
	.w8(32'hba51f1f2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81e4c1),
	.w1(32'hbb4758c2),
	.w2(32'hb9a67b86),
	.w3(32'hba9e3610),
	.w4(32'hbb2c3d9c),
	.w5(32'hbabef1a3),
	.w6(32'hba2fd983),
	.w7(32'hbadaf47d),
	.w8(32'hbb0d3dc5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39426431),
	.w1(32'hba2168ee),
	.w2(32'h38e6e63b),
	.w3(32'hba3584e4),
	.w4(32'hbadadb84),
	.w5(32'hba95ebe3),
	.w6(32'hba012065),
	.w7(32'hb9e3246e),
	.w8(32'h3a693970),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa09ba),
	.w1(32'hbaabdefe),
	.w2(32'hba67f8aa),
	.w3(32'hbaafcb06),
	.w4(32'hbb268771),
	.w5(32'hbac460c6),
	.w6(32'h39fe931b),
	.w7(32'hbad2ab89),
	.w8(32'hba8d4828),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fda5b),
	.w1(32'hbb00134d),
	.w2(32'h3a3cd22a),
	.w3(32'hba8636e2),
	.w4(32'hbae35a5e),
	.w5(32'hba6dfc51),
	.w6(32'hba08bf9d),
	.w7(32'hbabf5593),
	.w8(32'hba90a6f1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4860cf),
	.w1(32'h3b5774c0),
	.w2(32'h3b194e7c),
	.w3(32'hbaf5bc09),
	.w4(32'h3b4de78d),
	.w5(32'hb9d79751),
	.w6(32'hbb048bf3),
	.w7(32'h3accf463),
	.w8(32'hb8277d19),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82317b),
	.w1(32'h3acb41d7),
	.w2(32'h3ada12aa),
	.w3(32'hba52356b),
	.w4(32'h3aad28a8),
	.w5(32'h3b34a8f4),
	.w6(32'hb86a5b4a),
	.w7(32'h3a795875),
	.w8(32'h3aa905bd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac40f6e),
	.w1(32'h3a579799),
	.w2(32'hba0003c2),
	.w3(32'h3aac8ba9),
	.w4(32'h3a940fd5),
	.w5(32'h3aeaab54),
	.w6(32'h3b098889),
	.w7(32'h38396b7f),
	.w8(32'hb9be0b48),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ca06c),
	.w1(32'h3b143e1b),
	.w2(32'h3aa36beb),
	.w3(32'h3a12579d),
	.w4(32'h3ad44854),
	.w5(32'h392f6a6a),
	.w6(32'hb985d6a9),
	.w7(32'h3a81deee),
	.w8(32'h39d0f648),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91d73e),
	.w1(32'hba5cd1d5),
	.w2(32'h378aa7bb),
	.w3(32'hbaeb7110),
	.w4(32'hb98715b3),
	.w5(32'hba2cb9d1),
	.w6(32'h3978c1e8),
	.w7(32'hba2126a0),
	.w8(32'hb979c237),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba061743),
	.w1(32'h3a85c0d2),
	.w2(32'h392c7fcb),
	.w3(32'hb99bbb9d),
	.w4(32'h3913ceaf),
	.w5(32'h3a193694),
	.w6(32'h3838a454),
	.w7(32'hba8520b6),
	.w8(32'h3893065a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0471a6),
	.w1(32'hba6dfe05),
	.w2(32'hb90e04b5),
	.w3(32'hb9101287),
	.w4(32'hba824945),
	.w5(32'hb9f93384),
	.w6(32'h3870d88b),
	.w7(32'hba82dafe),
	.w8(32'hb92fbcd0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12edc3),
	.w1(32'h39b72f88),
	.w2(32'h3abcd587),
	.w3(32'hbac14291),
	.w4(32'hbacb55cc),
	.w5(32'hb9aa32c9),
	.w6(32'hb9e9a44d),
	.w7(32'h3964493a),
	.w8(32'h3a07be3d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a865926),
	.w1(32'h39b89f1a),
	.w2(32'hb9371e78),
	.w3(32'hbab7b542),
	.w4(32'hba1a6864),
	.w5(32'h3ab417ff),
	.w6(32'hbadbfd31),
	.w7(32'h39bead6d),
	.w8(32'h3a3cb5cf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c70ac),
	.w1(32'hb975d0f7),
	.w2(32'hb98091e8),
	.w3(32'h3a3db546),
	.w4(32'h37980700),
	.w5(32'hb9e955e8),
	.w6(32'h3a2a0fcf),
	.w7(32'h3910a2ab),
	.w8(32'hba27f283),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f274e6),
	.w1(32'h3a2a6c9b),
	.w2(32'h3a1cc8e7),
	.w3(32'h3a5bfa68),
	.w4(32'h3a42ad91),
	.w5(32'h39f75381),
	.w6(32'h391afbd4),
	.w7(32'h3a972529),
	.w8(32'h3a6d4ea8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25b08b),
	.w1(32'hbadfac8e),
	.w2(32'hbb111bb0),
	.w3(32'hb923b803),
	.w4(32'hbaff7bd4),
	.w5(32'hbaad7293),
	.w6(32'hb82f19b1),
	.w7(32'hbb2a18ec),
	.w8(32'hbae13e5e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba103b80),
	.w1(32'h3a98cb26),
	.w2(32'h3b2ff3fa),
	.w3(32'hb9d2cbfc),
	.w4(32'hb9f73d80),
	.w5(32'h3ae2a4cf),
	.w6(32'hba10657d),
	.w7(32'hba65200c),
	.w8(32'h3aa350c1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bb50d),
	.w1(32'hb988327d),
	.w2(32'h39b68634),
	.w3(32'h3a749be1),
	.w4(32'hb98f7834),
	.w5(32'h3a17fc5c),
	.w6(32'h3b1a8f98),
	.w7(32'h39153cd0),
	.w8(32'h3aa5669c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1534b0),
	.w1(32'h3ab5dac0),
	.w2(32'h3a0df214),
	.w3(32'h3af40265),
	.w4(32'h3a9f7a78),
	.w5(32'h3ab4a9e1),
	.w6(32'h3a7b4075),
	.w7(32'h3aa48eab),
	.w8(32'h3a845e7b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4715a0),
	.w1(32'hb94289d9),
	.w2(32'h3a1062b1),
	.w3(32'h39969f65),
	.w4(32'hba439ca8),
	.w5(32'hbb128887),
	.w6(32'h38973ae0),
	.w7(32'h3a21df12),
	.w8(32'hbb120284),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38081d1a),
	.w1(32'hbaceeffb),
	.w2(32'hbaf15961),
	.w3(32'hbaca2e3a),
	.w4(32'hbacabce6),
	.w5(32'hba205cf7),
	.w6(32'hba5663c4),
	.w7(32'hba7a8545),
	.w8(32'hba426c3e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f11d1),
	.w1(32'h38890c7d),
	.w2(32'h39bb5646),
	.w3(32'h3a522213),
	.w4(32'hba393f6d),
	.w5(32'h3a125b58),
	.w6(32'hb9a11feb),
	.w7(32'hba2f8a11),
	.w8(32'hba300ac6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1f3d2),
	.w1(32'h3a3f9618),
	.w2(32'h3b01d512),
	.w3(32'hbae40900),
	.w4(32'h3a72ff11),
	.w5(32'h3a68e8ce),
	.w6(32'hba528a57),
	.w7(32'h3aeb4fc2),
	.w8(32'h3b543b44),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b096c6a),
	.w1(32'h3a665a7b),
	.w2(32'h3a94cc45),
	.w3(32'h3ae205ae),
	.w4(32'h39f3e77c),
	.w5(32'h3b2a2c99),
	.w6(32'h3acab716),
	.w7(32'h3ab53169),
	.w8(32'h3aae204b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa7e37),
	.w1(32'hba3264b6),
	.w2(32'hb9d8ed12),
	.w3(32'hbab4ed60),
	.w4(32'hba68913c),
	.w5(32'hba6bce89),
	.w6(32'hbb06d9a9),
	.w7(32'hbaaf6fa9),
	.w8(32'hb9fc79ff),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba452e2b),
	.w1(32'h3ae324ae),
	.w2(32'h3a7a96d9),
	.w3(32'hbaea2c6c),
	.w4(32'hb8d16df9),
	.w5(32'h3ac7a50a),
	.w6(32'hba96d792),
	.w7(32'hba85a117),
	.w8(32'hb902a281),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a9972),
	.w1(32'hb96f96dc),
	.w2(32'h38c8e25b),
	.w3(32'hba888bad),
	.w4(32'hb9ac0273),
	.w5(32'h3a8cca66),
	.w6(32'hba47f135),
	.w7(32'h398b4969),
	.w8(32'h3a51758c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bdb8e),
	.w1(32'hbaa19ec8),
	.w2(32'hba8a6542),
	.w3(32'h3a3a1262),
	.w4(32'hbb1958b2),
	.w5(32'hbaee9e1c),
	.w6(32'hb9123f7c),
	.w7(32'hba7c9baf),
	.w8(32'hb9923cc6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f424b2),
	.w1(32'hb96d8001),
	.w2(32'h3a258157),
	.w3(32'hba1f712d),
	.w4(32'hba146a9e),
	.w5(32'hba89af5d),
	.w6(32'h3a54bcff),
	.w7(32'hb98e8f8a),
	.w8(32'hba8ee673),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a451e5f),
	.w1(32'h3ad8c2b6),
	.w2(32'h3a4ec63b),
	.w3(32'hb94337d3),
	.w4(32'h3932cb1b),
	.w5(32'hba8d846e),
	.w6(32'h392fca7e),
	.w7(32'h3a162ceb),
	.w8(32'hba402c28),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58e20f),
	.w1(32'hbb3e561c),
	.w2(32'hb90c4de3),
	.w3(32'hb9c5c338),
	.w4(32'hbb76695a),
	.w5(32'hba2df5c8),
	.w6(32'hb9cbfddf),
	.w7(32'hbb5ab98f),
	.w8(32'hbacef509),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd8c9b),
	.w1(32'h38e081c6),
	.w2(32'h3a4c9b7f),
	.w3(32'hb9a43be7),
	.w4(32'hba356780),
	.w5(32'h38ba15db),
	.w6(32'hbadfa8ff),
	.w7(32'h39f2c5fc),
	.w8(32'h38b433f7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f01007),
	.w1(32'h392cae98),
	.w2(32'h3a82c6f9),
	.w3(32'hba219170),
	.w4(32'hb91122df),
	.w5(32'hb83cb273),
	.w6(32'hb9f9238f),
	.w7(32'h3a869082),
	.w8(32'hb80d931d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59e233),
	.w1(32'h3a9f8d00),
	.w2(32'h38b4f2f5),
	.w3(32'h39b02164),
	.w4(32'h3aa0af39),
	.w5(32'h3a908f3c),
	.w6(32'h3a238e0d),
	.w7(32'h3a8c5316),
	.w8(32'h3a870f0a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08176c),
	.w1(32'h36f34c9b),
	.w2(32'h39a68407),
	.w3(32'hbacf3755),
	.w4(32'hb9cb54bf),
	.w5(32'hbab6e40e),
	.w6(32'hba1c1b83),
	.w7(32'hbab6e7bf),
	.w8(32'hbabd6b98),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0efb95),
	.w1(32'h3a070256),
	.w2(32'hb9ddae13),
	.w3(32'hb960d401),
	.w4(32'hb9e36038),
	.w5(32'hba7e4182),
	.w6(32'hb8597abf),
	.w7(32'hba337106),
	.w8(32'hba11d54a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1297f0),
	.w1(32'hb9b0f4f8),
	.w2(32'hba984c8a),
	.w3(32'h3a25f253),
	.w4(32'hbab9c2b0),
	.w5(32'hbb26be91),
	.w6(32'h39a1dd4b),
	.w7(32'hbab132f6),
	.w8(32'hbb096202),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e7d4af),
	.w1(32'hb96ce09a),
	.w2(32'hbaccad27),
	.w3(32'hbaa3c91f),
	.w4(32'hb9f48df8),
	.w5(32'hba9f889c),
	.w6(32'hbae98d9d),
	.w7(32'hb8364964),
	.w8(32'h392cfe60),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9907572),
	.w1(32'h39945f9f),
	.w2(32'hbad37459),
	.w3(32'h3a026f4a),
	.w4(32'hb970ae22),
	.w5(32'hbafef176),
	.w6(32'h3a38727c),
	.w7(32'hbaa38815),
	.w8(32'hbb6767f9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba191efe),
	.w1(32'h3b07bc5d),
	.w2(32'h3a8ee61d),
	.w3(32'hbb589af2),
	.w4(32'h3ae43a48),
	.w5(32'h3abaf082),
	.w6(32'hbb80cbac),
	.w7(32'h3ae169f9),
	.w8(32'h3ad6c5f8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace2068),
	.w1(32'h3a23fab2),
	.w2(32'hba0fcbef),
	.w3(32'h3a5cd687),
	.w4(32'h39933cae),
	.w5(32'hba434432),
	.w6(32'h3ab2665e),
	.w7(32'h3a64e98b),
	.w8(32'hb9c420ab),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be94ea),
	.w1(32'hba818615),
	.w2(32'hb98be197),
	.w3(32'hb9c1b2a1),
	.w4(32'hb9da2877),
	.w5(32'h3a376467),
	.w6(32'hba0647a4),
	.w7(32'hba44aeb3),
	.w8(32'hba927b64),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e6308),
	.w1(32'h3af3f161),
	.w2(32'h3a951a02),
	.w3(32'hbac6282d),
	.w4(32'h3a882be4),
	.w5(32'h38eb51a2),
	.w6(32'hbac39155),
	.w7(32'h3a5da4a0),
	.w8(32'h3a311a4f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b9722),
	.w1(32'h3af6a0a9),
	.w2(32'h3b2e3c07),
	.w3(32'hb98031f8),
	.w4(32'h3a9de71d),
	.w5(32'h3b0e4aa0),
	.w6(32'h3a245f9d),
	.w7(32'h3ae96a51),
	.w8(32'h3b2103c6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b482121),
	.w1(32'h3a494330),
	.w2(32'hb99f8923),
	.w3(32'h3b383cbb),
	.w4(32'h3a4ee0d2),
	.w5(32'h392378b3),
	.w6(32'h3b5786c1),
	.w7(32'h3a3c030b),
	.w8(32'h3a65fbe2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff2c3d),
	.w1(32'hbaebd9dd),
	.w2(32'hb8a11cc7),
	.w3(32'h3b217d2b),
	.w4(32'hbab8cd6f),
	.w5(32'h377c0ec6),
	.w6(32'h3b06d6d1),
	.w7(32'hba291c9b),
	.w8(32'hb7e67dc2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a177f),
	.w1(32'hba378e61),
	.w2(32'hb8904d1f),
	.w3(32'h3a8d7669),
	.w4(32'hbac59f51),
	.w5(32'hba563a8e),
	.w6(32'h3912e9eb),
	.w7(32'hbab5c89c),
	.w8(32'hb9fca9f4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0b2da),
	.w1(32'h3a30f096),
	.w2(32'h3ab56a13),
	.w3(32'hba9df675),
	.w4(32'h3a8241aa),
	.w5(32'h3b1ab0dd),
	.w6(32'hba38d47d),
	.w7(32'h3ad4c144),
	.w8(32'h3b1ab191),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa94171),
	.w1(32'hbb62a309),
	.w2(32'hba482843),
	.w3(32'h3aaaa5a8),
	.w4(32'hbb254b55),
	.w5(32'hba87c391),
	.w6(32'h3a8a249b),
	.w7(32'hbae1d2e3),
	.w8(32'hbaeddd8f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04e17c),
	.w1(32'hb9dca6ae),
	.w2(32'h3af6ddd7),
	.w3(32'hba95a9b1),
	.w4(32'h393aaf98),
	.w5(32'h3b66000b),
	.w6(32'h37ee3d41),
	.w7(32'h3a16c99e),
	.w8(32'h3b00452a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfd93b),
	.w1(32'h3b85ef33),
	.w2(32'h3b9643c2),
	.w3(32'h3b847092),
	.w4(32'h3723e972),
	.w5(32'h3b4aa7f9),
	.w6(32'hbace4be7),
	.w7(32'hb91988ce),
	.w8(32'h3c02c78c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad87aec),
	.w1(32'h3a5ba16b),
	.w2(32'hbb1fb902),
	.w3(32'h3b1aa3f5),
	.w4(32'h3a3cb6ff),
	.w5(32'h3b61a095),
	.w6(32'h3b27f038),
	.w7(32'h3a84c0dd),
	.w8(32'h3a3e9406),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14f543),
	.w1(32'h3b09212c),
	.w2(32'h3b46031b),
	.w3(32'hbb3a2958),
	.w4(32'h39891a2f),
	.w5(32'hbb002890),
	.w6(32'h3a801d4c),
	.w7(32'h3b6de27f),
	.w8(32'h3aab2c47),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf24f44),
	.w1(32'h3b4b7383),
	.w2(32'h3baa9148),
	.w3(32'h3c26d3c8),
	.w4(32'h3baae4f7),
	.w5(32'h3bb61463),
	.w6(32'h3bedfa5d),
	.w7(32'h3b5ccc29),
	.w8(32'h3c024c05),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94c21c),
	.w1(32'hbc32c14c),
	.w2(32'hbc1d7386),
	.w3(32'h3bfc97d7),
	.w4(32'hbc4bcae0),
	.w5(32'hbc278f1e),
	.w6(32'h3c0f914c),
	.w7(32'hbb443f01),
	.w8(32'hb8f905cb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc5574),
	.w1(32'hba40b4fe),
	.w2(32'hbb63b2db),
	.w3(32'h3b823c6c),
	.w4(32'hbaeb7851),
	.w5(32'hbb1af3f8),
	.w6(32'hbbe0298e),
	.w7(32'hbbe8abea),
	.w8(32'hbbbf5bfe),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56da3a),
	.w1(32'h3b2e7b52),
	.w2(32'h3c7b128d),
	.w3(32'hbb81454c),
	.w4(32'h3ada76d5),
	.w5(32'h3ca17577),
	.w6(32'hbb94e28c),
	.w7(32'hbb867b65),
	.w8(32'h3b085b4f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae43bfb),
	.w1(32'h3ba707e5),
	.w2(32'h3ca9c7e6),
	.w3(32'h3c6d2622),
	.w4(32'h3c5bc3ee),
	.w5(32'h3d009cef),
	.w6(32'h3c277743),
	.w7(32'h3c29233f),
	.w8(32'h3cbcc786),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12e1f9),
	.w1(32'hba3e57d2),
	.w2(32'hbb4d93a7),
	.w3(32'h3c874279),
	.w4(32'hbb04fc89),
	.w5(32'hbb4c11e9),
	.w6(32'h3c62289d),
	.w7(32'h3abe5110),
	.w8(32'hbb1300ee),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd12ba),
	.w1(32'h3c118940),
	.w2(32'h3a962079),
	.w3(32'hbad015e1),
	.w4(32'h3bf1047e),
	.w5(32'hbbbf09a7),
	.w6(32'hb9976466),
	.w7(32'h3bc5e710),
	.w8(32'hbb8140fe),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54ab5c),
	.w1(32'hbb6ce6d5),
	.w2(32'hbbe57ece),
	.w3(32'h3b32d358),
	.w4(32'hbb9e5c2d),
	.w5(32'hbc0f318d),
	.w6(32'h3b8eb789),
	.w7(32'hbba845dd),
	.w8(32'hbc0852b4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1086f),
	.w1(32'h3b1f08f8),
	.w2(32'hbbabb82b),
	.w3(32'hbbe9f9c0),
	.w4(32'hbb7e4703),
	.w5(32'hbc36242e),
	.w6(32'hbc0e64f1),
	.w7(32'hbbcd2108),
	.w8(32'hbbbbf8c2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa18a64),
	.w1(32'h3b625859),
	.w2(32'h3b73ca10),
	.w3(32'h3b7b9730),
	.w4(32'hb9a19528),
	.w5(32'h3b601816),
	.w6(32'h3bfae257),
	.w7(32'h3aa68724),
	.w8(32'h3a836171),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90db5ca),
	.w1(32'hbb446c9d),
	.w2(32'h3b15dc27),
	.w3(32'hba970849),
	.w4(32'hbb849e94),
	.w5(32'h3b065383),
	.w6(32'hbbb14c02),
	.w7(32'hbb37db3a),
	.w8(32'h3b81cc45),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc51769),
	.w1(32'h378dbd17),
	.w2(32'hb9d87872),
	.w3(32'h3b15253b),
	.w4(32'hbb3da565),
	.w5(32'hbb81f584),
	.w6(32'hb9bc871b),
	.w7(32'h3b6e529f),
	.w8(32'hbac19ffe),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b592e5c),
	.w1(32'hbb840b13),
	.w2(32'h3c42385b),
	.w3(32'hba9cbdda),
	.w4(32'h3ba1de5e),
	.w5(32'h3cd4931b),
	.w6(32'hbb7f9b8e),
	.w7(32'h3bddde95),
	.w8(32'h3c7ccbe9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf41bcf),
	.w1(32'hbaf20938),
	.w2(32'h3b48dc36),
	.w3(32'h3c590fd1),
	.w4(32'h3ba623f2),
	.w5(32'h3c1c52e7),
	.w6(32'h3bd44bc5),
	.w7(32'h3b6df3e6),
	.w8(32'h3bcab1a0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82a708),
	.w1(32'h3a9963f7),
	.w2(32'h3acd3900),
	.w3(32'hbabb73f2),
	.w4(32'h3a61d352),
	.w5(32'h3a8cb8d6),
	.w6(32'hb886ba43),
	.w7(32'hbb990026),
	.w8(32'hba73ec59),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93babb),
	.w1(32'hbc58ace9),
	.w2(32'hbc2e9b37),
	.w3(32'hbaed2b22),
	.w4(32'hbc308010),
	.w5(32'hbb3a4ec5),
	.w6(32'h3a543a96),
	.w7(32'hbbc50048),
	.w8(32'hbbe281e2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8957a),
	.w1(32'h3b081b17),
	.w2(32'h3b0fb878),
	.w3(32'hbb01ff8d),
	.w4(32'h3a8298ac),
	.w5(32'h3ad42452),
	.w6(32'hbba0a3e4),
	.w7(32'hba88c3d4),
	.w8(32'h399893cf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7138fd),
	.w1(32'hb8cab30a),
	.w2(32'hb7cf7146),
	.w3(32'h380e2bbb),
	.w4(32'hba6f1945),
	.w5(32'hbb0a7281),
	.w6(32'hbb2bdb26),
	.w7(32'hb9eba0ef),
	.w8(32'hba3ff7b0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6743f),
	.w1(32'h3ba2904b),
	.w2(32'h3bb9ad33),
	.w3(32'hbb7716b7),
	.w4(32'h3b3627e7),
	.w5(32'h3ad7ee11),
	.w6(32'hbb8b972f),
	.w7(32'h3a344472),
	.w8(32'h3b73f9db),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc41be2),
	.w1(32'hbb99d14f),
	.w2(32'hbc0ea05a),
	.w3(32'h3b942fb7),
	.w4(32'h3a3f1182),
	.w5(32'hbbfef845),
	.w6(32'h3bf00162),
	.w7(32'h3b1a2446),
	.w8(32'hbb2c4cad),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b1433),
	.w1(32'h3aa493bb),
	.w2(32'hb93a1762),
	.w3(32'hbc0b8d8f),
	.w4(32'hbb27599b),
	.w5(32'hbb5d1bda),
	.w6(32'hbbc8675f),
	.w7(32'h3963f3f8),
	.w8(32'h38d69c11),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40aacc),
	.w1(32'h3c026621),
	.w2(32'hbaf3e09b),
	.w3(32'hbb307d1a),
	.w4(32'h3c278bb0),
	.w5(32'hbbb86e5d),
	.w6(32'hbad76c55),
	.w7(32'hbab1c58f),
	.w8(32'hbc4778ee),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba48b62),
	.w1(32'hb9d91121),
	.w2(32'h3ae85920),
	.w3(32'hbc20b1be),
	.w4(32'hbb368251),
	.w5(32'h3aa328c6),
	.w6(32'hbb8a31a7),
	.w7(32'h38b908f7),
	.w8(32'h3aa76a82),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391deb9e),
	.w1(32'h3b4e9598),
	.w2(32'hb99b58d4),
	.w3(32'hbac94781),
	.w4(32'h3c04f16c),
	.w5(32'h3a85f50c),
	.w6(32'hbb1886c3),
	.w7(32'h3c573bea),
	.w8(32'h3b47c76c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6079ee),
	.w1(32'hbc057628),
	.w2(32'hbaf02bbc),
	.w3(32'hbb95b23b),
	.w4(32'hb9f5990d),
	.w5(32'h3bc3e165),
	.w6(32'hb8009a2e),
	.w7(32'h3b6eea2e),
	.w8(32'h3b9d02a4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03feb6),
	.w1(32'hbb448199),
	.w2(32'hbb9990f2),
	.w3(32'h3b9847e5),
	.w4(32'h3b6fc073),
	.w5(32'h3b4d0bb7),
	.w6(32'h3b9ae893),
	.w7(32'h3b481c4f),
	.w8(32'h3a98b1ce),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ed66),
	.w1(32'hbb568604),
	.w2(32'hba82c1bc),
	.w3(32'hbb0857a8),
	.w4(32'hbb7008bd),
	.w5(32'hbb1e7a46),
	.w6(32'hbb4f26b6),
	.w7(32'h3b69b09b),
	.w8(32'h3b1cf25d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58e495),
	.w1(32'h3b99ccdc),
	.w2(32'h3930910d),
	.w3(32'h3acb4857),
	.w4(32'h3b8b1c7f),
	.w5(32'h3ba68c63),
	.w6(32'hbb6fd670),
	.w7(32'h3b84435a),
	.w8(32'h3bb335cf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d6d9),
	.w1(32'hbb941644),
	.w2(32'h3c814d78),
	.w3(32'h3ae02b86),
	.w4(32'hbb9d5c85),
	.w5(32'h3bcdef6e),
	.w6(32'h3b3709d7),
	.w7(32'hbc8c14c9),
	.w8(32'hba8035ca),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc011aeb),
	.w1(32'hbc0cf32d),
	.w2(32'h3c19cd01),
	.w3(32'hbc59823c),
	.w4(32'hbaf035cc),
	.w5(32'h3d10d2dc),
	.w6(32'hba523837),
	.w7(32'hbc0e4a18),
	.w8(32'h3b0b0bc6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a61c6),
	.w1(32'h3b1b4d71),
	.w2(32'h3a96a049),
	.w3(32'h3c104a13),
	.w4(32'hb7f338fd),
	.w5(32'h3b73f7ec),
	.w6(32'hba547e82),
	.w7(32'h3b0d408d),
	.w8(32'h3bfebc9e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f4f54),
	.w1(32'h3b8d64c4),
	.w2(32'hbafcdc35),
	.w3(32'h3a9816e5),
	.w4(32'h3bb0dce5),
	.w5(32'hba083cc0),
	.w6(32'h3b070855),
	.w7(32'h3c070d63),
	.w8(32'h3aef4a78),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d87bc),
	.w1(32'h3b198373),
	.w2(32'hba4a74a4),
	.w3(32'hbbb016e9),
	.w4(32'h3b46ff88),
	.w5(32'h3b072508),
	.w6(32'hbaa293cb),
	.w7(32'h38ecb976),
	.w8(32'hb9e79162),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac14cd),
	.w1(32'hb8469208),
	.w2(32'h3b4967f7),
	.w3(32'h3bda2ea9),
	.w4(32'hbb8a56d6),
	.w5(32'h3a3868b9),
	.w6(32'hbb4c0245),
	.w7(32'hbb87f0c2),
	.w8(32'h39fdce08),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3420b),
	.w1(32'hb8a93150),
	.w2(32'hba23a5e9),
	.w3(32'hbab3debb),
	.w4(32'hbb4b96be),
	.w5(32'hbba3170d),
	.w6(32'hb9dc4eb1),
	.w7(32'hba9b58f1),
	.w8(32'h3b857748),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc99d6),
	.w1(32'hbb82bbd1),
	.w2(32'hbbaf888e),
	.w3(32'hbb073283),
	.w4(32'hbb10eb1a),
	.w5(32'hbb4c8d16),
	.w6(32'hbaf87a31),
	.w7(32'h3b67bf53),
	.w8(32'h3bd93fe0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf0437),
	.w1(32'hbb8142ee),
	.w2(32'hbb531b36),
	.w3(32'h3b640efd),
	.w4(32'hbafad72e),
	.w5(32'hbb47ee4d),
	.w6(32'hbbc96b24),
	.w7(32'h3b1b1074),
	.w8(32'hb884efef),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17f46f),
	.w1(32'h3b6e662f),
	.w2(32'hbb1d889f),
	.w3(32'hbbd528ed),
	.w4(32'h3b1a477f),
	.w5(32'hba07b6b0),
	.w6(32'hbb03361f),
	.w7(32'h3b0c8cdc),
	.w8(32'hba45845d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc97025),
	.w1(32'h3ab74c38),
	.w2(32'hbc31248d),
	.w3(32'hbbd9169a),
	.w4(32'hbb8c2677),
	.w5(32'hbca161e8),
	.w6(32'hbbd364c2),
	.w7(32'hbabefdae),
	.w8(32'hbc800558),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb3d09),
	.w1(32'hbca5c59b),
	.w2(32'hbc898b3e),
	.w3(32'hbc5f235a),
	.w4(32'hbcc27d01),
	.w5(32'hbcb7b1d3),
	.w6(32'hbb96fe18),
	.w7(32'hbc7a3fb1),
	.w8(32'hbc1d72de),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb04d39),
	.w1(32'hbbd43aa2),
	.w2(32'h3a97d57f),
	.w3(32'h3d4c1197),
	.w4(32'hbba2f8e7),
	.w5(32'h3bf790b0),
	.w6(32'h3c8d53e9),
	.w7(32'hbb26743c),
	.w8(32'h3bc4d87d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2181ef),
	.w1(32'h3815eaa9),
	.w2(32'hbb90a19a),
	.w3(32'h3c4284c5),
	.w4(32'hbb2485ee),
	.w5(32'hbb7fb1da),
	.w6(32'h3c12f4c8),
	.w7(32'hbb16c06f),
	.w8(32'hbba2a589),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4be3b5),
	.w1(32'hbb99e658),
	.w2(32'hbcab97ea),
	.w3(32'h3b0f6482),
	.w4(32'hbb31aef7),
	.w5(32'hbcca9ce5),
	.w6(32'h3b1a6982),
	.w7(32'h3930f053),
	.w8(32'hbc85925a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc077b35),
	.w1(32'h3a15b011),
	.w2(32'hba0d001c),
	.w3(32'hbc80d051),
	.w4(32'h3c64671e),
	.w5(32'h3c67806d),
	.w6(32'hbc980a09),
	.w7(32'h3c7b044d),
	.w8(32'h3c570677),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef8491),
	.w1(32'hbb0a48ed),
	.w2(32'h3ba58014),
	.w3(32'h3c0c0204),
	.w4(32'hbab86b73),
	.w5(32'h3ac7bdc6),
	.w6(32'h3c0dac44),
	.w7(32'hba9b2a82),
	.w8(32'h3b83cc7a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb308a25),
	.w1(32'h3a32f348),
	.w2(32'hbba4e5d4),
	.w3(32'hbb870678),
	.w4(32'hbb7e6f9f),
	.w5(32'hbc19b296),
	.w6(32'h3a1ab275),
	.w7(32'hbc0a1bfa),
	.w8(32'hbc25c50d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba60098),
	.w1(32'h3b225fb6),
	.w2(32'hbb55b2e3),
	.w3(32'hbc17b24c),
	.w4(32'h3b03dfef),
	.w5(32'hbb979e6a),
	.w6(32'hbbffcf0f),
	.w7(32'hba2866f6),
	.w8(32'hbb502ff7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7946bf),
	.w1(32'hbb1bb791),
	.w2(32'h3ab983b7),
	.w3(32'h3bc6ecc5),
	.w4(32'h394e5fa1),
	.w5(32'hbae66454),
	.w6(32'h3ae82d36),
	.w7(32'hbad3054d),
	.w8(32'h3b047916),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b233937),
	.w1(32'hbab37c29),
	.w2(32'hbbc7cd5f),
	.w3(32'h3b0dd4d6),
	.w4(32'hbbeedfd6),
	.w5(32'hbc21d895),
	.w6(32'h3a99a0fb),
	.w7(32'hbc47ea9f),
	.w8(32'hbc16d5dd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdba7e),
	.w1(32'h3b8885ca),
	.w2(32'hbb9c883c),
	.w3(32'hbbfb5211),
	.w4(32'hba784a50),
	.w5(32'hbc220027),
	.w6(32'hbb8895e7),
	.w7(32'h3b210e8e),
	.w8(32'hbba6a147),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989865),
	.w1(32'hbb79bd03),
	.w2(32'h3ab00d29),
	.w3(32'hbc4082a8),
	.w4(32'hbba071fe),
	.w5(32'h3abfeabd),
	.w6(32'hbb4c8d30),
	.w7(32'hbac449bd),
	.w8(32'h3bf1ac60),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b040518),
	.w1(32'hbc50dc7e),
	.w2(32'hb9eeb9e8),
	.w3(32'h3c0efc72),
	.w4(32'hbb8ff5fa),
	.w5(32'h3c5883e5),
	.w6(32'h3b4510e5),
	.w7(32'h3a01ee72),
	.w8(32'h3c97b8f4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83ad02),
	.w1(32'h3b0db579),
	.w2(32'h3c351d01),
	.w3(32'h3ceb2228),
	.w4(32'h3ab66e01),
	.w5(32'h3be4789f),
	.w6(32'h3c367fb1),
	.w7(32'hbb59c998),
	.w8(32'h3b1f33a2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b813a),
	.w1(32'h3b6b1718),
	.w2(32'h392f7363),
	.w3(32'h3bdb2cc8),
	.w4(32'h3a763c4f),
	.w5(32'hb97f7855),
	.w6(32'h3bcf5189),
	.w7(32'hbb89be79),
	.w8(32'h3abf0773),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9005a6c),
	.w1(32'hbbab5812),
	.w2(32'hbb51710b),
	.w3(32'hba86b310),
	.w4(32'hbb0a18ac),
	.w5(32'hbab338e8),
	.w6(32'h3bced38a),
	.w7(32'h3a520748),
	.w8(32'hbb51f5e5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f43238),
	.w1(32'hbc0c6b05),
	.w2(32'hbbdc382e),
	.w3(32'h3a042f8b),
	.w4(32'hbc56bedd),
	.w5(32'hbae73cc4),
	.w6(32'h3a4880a7),
	.w7(32'hbc64b972),
	.w8(32'hbbc3a4dd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8317c5),
	.w1(32'hbc4718b3),
	.w2(32'hb9262381),
	.w3(32'h3a8a1052),
	.w4(32'hbc01cb38),
	.w5(32'h3c00850e),
	.w6(32'hba17f2e0),
	.w7(32'hbb87b5e9),
	.w8(32'h3bfded37),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6a9ee),
	.w1(32'h3a1a5a43),
	.w2(32'hbb0f6ac8),
	.w3(32'hbb70c8ee),
	.w4(32'h3b9207ab),
	.w5(32'h3c428eee),
	.w6(32'hbc4ef263),
	.w7(32'h3b778831),
	.w8(32'h3c47be7f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bd56e),
	.w1(32'h3bb6f6b7),
	.w2(32'hbb938cda),
	.w3(32'h3cc11eb8),
	.w4(32'h3c0e05ac),
	.w5(32'h3af01a86),
	.w6(32'h3c9651d5),
	.w7(32'h3c482dc2),
	.w8(32'h3b9547e7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd30ed4),
	.w1(32'h3b857ee3),
	.w2(32'hbb319039),
	.w3(32'hbbdca1fd),
	.w4(32'h3b51bd93),
	.w5(32'hbac4a3b8),
	.w6(32'hbaa1a6db),
	.w7(32'h3b08c946),
	.w8(32'h3a982c64),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933018d),
	.w1(32'h3b0e876e),
	.w2(32'h3c0cd8fb),
	.w3(32'hbb6bc806),
	.w4(32'h3b73d66c),
	.w5(32'h3b9e1ad5),
	.w6(32'hbaf45244),
	.w7(32'hba32ff0f),
	.w8(32'hbb43d80c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d61d4),
	.w1(32'hbbc5c196),
	.w2(32'hbbf442ca),
	.w3(32'hbb13be51),
	.w4(32'hbabbe5f2),
	.w5(32'hbbe733ec),
	.w6(32'h3ac0b02c),
	.w7(32'h374bc824),
	.w8(32'hba9227e5),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ec37),
	.w1(32'hbbdca0dd),
	.w2(32'h3bc838a4),
	.w3(32'h3a5e9f87),
	.w4(32'hba2f50d4),
	.w5(32'h3cc89d02),
	.w6(32'hba519825),
	.w7(32'hba5d8216),
	.w8(32'h3c33bd7e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c412e4c),
	.w1(32'h3b611c09),
	.w2(32'h3b986084),
	.w3(32'h3cf0cb8e),
	.w4(32'h3c189938),
	.w5(32'h3c231f4d),
	.w6(32'h3c213575),
	.w7(32'h3bebedd0),
	.w8(32'h3bbe3895),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9743ee),
	.w1(32'hba02ee3d),
	.w2(32'h3b593a0f),
	.w3(32'h3b2cf85f),
	.w4(32'hbc035b55),
	.w5(32'hbc1091be),
	.w6(32'hbbbe3b6b),
	.w7(32'hbc03d5f2),
	.w8(32'hbbf2094d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d3594),
	.w1(32'h3a637c54),
	.w2(32'h3a01b51f),
	.w3(32'hbbfee4f3),
	.w4(32'hbb482723),
	.w5(32'hbba10cbb),
	.w6(32'hbc3ec8d0),
	.w7(32'hbb942f1e),
	.w8(32'hbbeb9b99),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2561ee),
	.w1(32'hbb6d42eb),
	.w2(32'hba7884d3),
	.w3(32'h3aed2399),
	.w4(32'h3b76b8c5),
	.w5(32'h3c5eda1c),
	.w6(32'hbafa2733),
	.w7(32'hbb8a6fcf),
	.w8(32'h3af80b6c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989df43),
	.w1(32'hbafea1fe),
	.w2(32'h3bfb3e8e),
	.w3(32'h3c870437),
	.w4(32'hbb18584a),
	.w5(32'h3c3b0dd3),
	.w6(32'h3bd1c062),
	.w7(32'hbbea5b3f),
	.w8(32'hba2da011),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1312fa),
	.w1(32'hbb751e6e),
	.w2(32'hbb4adedc),
	.w3(32'hba06bced),
	.w4(32'hbbac5b4c),
	.w5(32'hbc1419ff),
	.w6(32'h3b642fd8),
	.w7(32'hbbdc8c64),
	.w8(32'hbc060009),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2384aa),
	.w1(32'hbb841799),
	.w2(32'hbb478000),
	.w3(32'hbbc89b76),
	.w4(32'hbb7996a0),
	.w5(32'hbbd4d19d),
	.w6(32'hbc36d947),
	.w7(32'hbbe2b624),
	.w8(32'hbc1c546f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f69f0d),
	.w1(32'hbaf87655),
	.w2(32'hba8182ed),
	.w3(32'h3b2d08c9),
	.w4(32'h3a55a18d),
	.w5(32'hbb68b55d),
	.w6(32'hbb0f9140),
	.w7(32'h3b70ba20),
	.w8(32'hba7978af),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d38946),
	.w1(32'hbb84591a),
	.w2(32'h3ae4e38c),
	.w3(32'h3b00e61a),
	.w4(32'hbae6360a),
	.w5(32'h3b96be9f),
	.w6(32'hbb173305),
	.w7(32'hbb6c8e88),
	.w8(32'hbb845d77),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe6488),
	.w1(32'h39a39e66),
	.w2(32'hbb36e44c),
	.w3(32'h3a5589f9),
	.w4(32'hbb76abf8),
	.w5(32'hbbfa1ffb),
	.w6(32'hbb5b5ec3),
	.w7(32'hbb134202),
	.w8(32'hbb50e97b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b181744),
	.w1(32'h3ac18d5d),
	.w2(32'h3bc5417f),
	.w3(32'h3b882888),
	.w4(32'h3b0c3f17),
	.w5(32'h3bc226d2),
	.w6(32'hba879a56),
	.w7(32'hbb6bd5b4),
	.w8(32'h3bd934da),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39e231),
	.w1(32'h3bcff729),
	.w2(32'h3b7e87ba),
	.w3(32'h3b2461d6),
	.w4(32'h3bf0c32c),
	.w5(32'h3b3078db),
	.w6(32'hba9ac9d9),
	.w7(32'h3b25cf61),
	.w8(32'hba1fb626),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8603d),
	.w1(32'h38d51b24),
	.w2(32'h3b15c588),
	.w3(32'h3bb650c2),
	.w4(32'h3a37907e),
	.w5(32'h3a824a68),
	.w6(32'h384f26d5),
	.w7(32'hb9af4f10),
	.w8(32'h3b95b8b5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad183be),
	.w1(32'hbb60e262),
	.w2(32'hb7e7b589),
	.w3(32'h3abc6de0),
	.w4(32'hbb87c931),
	.w5(32'h3b3319b7),
	.w6(32'h39328f6a),
	.w7(32'hba7948bf),
	.w8(32'h3a89d672),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3159b4),
	.w1(32'hbb0e3a35),
	.w2(32'hbb9a7192),
	.w3(32'hbbd48a13),
	.w4(32'hbb336e0f),
	.w5(32'hbac0589d),
	.w6(32'hbb30a04c),
	.w7(32'hbbf4cf9d),
	.w8(32'hbbe40d8b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8f64d),
	.w1(32'h3a7d9847),
	.w2(32'hba4847ff),
	.w3(32'h3b84a858),
	.w4(32'h3b9450db),
	.w5(32'h3b498fa4),
	.w6(32'hbad8202a),
	.w7(32'h3b236ffc),
	.w8(32'hba69aa21),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addddd7),
	.w1(32'hbaf9bcf1),
	.w2(32'hbaf608f5),
	.w3(32'h3b86c948),
	.w4(32'hbab215f9),
	.w5(32'hbb54a4dc),
	.w6(32'h3aab139f),
	.w7(32'hbb304c31),
	.w8(32'hbbb7a921),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e94536),
	.w1(32'h3bd3c4a5),
	.w2(32'h3b63e9c0),
	.w3(32'hbb741f2d),
	.w4(32'h3c3c5749),
	.w5(32'hba2aef4d),
	.w6(32'hbbb479a4),
	.w7(32'h3c2bb834),
	.w8(32'hbb13d242),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9861ad),
	.w1(32'h3a9e0fc7),
	.w2(32'h3ae83cb3),
	.w3(32'hbb34775f),
	.w4(32'hbb50ef78),
	.w5(32'h3b394e69),
	.w6(32'hbae3af0b),
	.w7(32'hbbea769e),
	.w8(32'hb9c8f6f0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba252b77),
	.w1(32'h3b8d72b5),
	.w2(32'h3a2d8b20),
	.w3(32'h394a9c5d),
	.w4(32'h3b90e453),
	.w5(32'h3a811d41),
	.w6(32'hb9edd4ba),
	.w7(32'h3ab10e11),
	.w8(32'h3bb470ba),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f81c8),
	.w1(32'h3bb72f66),
	.w2(32'h3b72c79d),
	.w3(32'hba8ea08f),
	.w4(32'h3c0a416f),
	.w5(32'h3b8c0fb8),
	.w6(32'h3b501c69),
	.w7(32'h3b5cb9aa),
	.w8(32'h3b020d05),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6f047),
	.w1(32'hba933f5f),
	.w2(32'hbb2c345d),
	.w3(32'h3a1a0e7e),
	.w4(32'h3b0106ab),
	.w5(32'h3b0bf0e1),
	.w6(32'hbb0cc108),
	.w7(32'hbb873fc0),
	.w8(32'hbb01ce3d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb640a19),
	.w1(32'hbb9ea19c),
	.w2(32'hbc830d0b),
	.w3(32'h3aeef396),
	.w4(32'hbbcc9be3),
	.w5(32'hbc970d78),
	.w6(32'hbb71e519),
	.w7(32'hbbb40b6e),
	.w8(32'hbc8b55c9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea035e),
	.w1(32'hbafe6293),
	.w2(32'h3c1f35e5),
	.w3(32'hbc3e36a6),
	.w4(32'hbb5ec64e),
	.w5(32'h3ae20bfd),
	.w6(32'hbc8714d0),
	.w7(32'h3b10fa0d),
	.w8(32'hbbda34cb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba208f88),
	.w1(32'hba13c270),
	.w2(32'hbb935e90),
	.w3(32'hbba9e829),
	.w4(32'hbaadcb35),
	.w5(32'hbbd8e42d),
	.w6(32'hbbbed400),
	.w7(32'h39f11e35),
	.w8(32'hbb9dfe84),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06aa46),
	.w1(32'hb9cfcf91),
	.w2(32'h3b1969d7),
	.w3(32'hbbf74e04),
	.w4(32'hbaa443c1),
	.w5(32'hb96945fa),
	.w6(32'h3b70b530),
	.w7(32'hbbc7ac47),
	.w8(32'hbba059e2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22eee2),
	.w1(32'hbbd290cb),
	.w2(32'h3c12aae1),
	.w3(32'h3a8c24d0),
	.w4(32'h3b55de4b),
	.w5(32'h3ca65e7b),
	.w6(32'h3b887b4f),
	.w7(32'h3af79d0a),
	.w8(32'h3c4629fc),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c383372),
	.w1(32'hbc52a805),
	.w2(32'hbc0d229b),
	.w3(32'h3ccd011c),
	.w4(32'hbc62a0e5),
	.w5(32'hbc0118fb),
	.w6(32'h3c66d3b3),
	.w7(32'hbc1348cb),
	.w8(32'hbb21d794),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac47b64),
	.w1(32'hbb1425a5),
	.w2(32'h3b0d2530),
	.w3(32'h3b527ca3),
	.w4(32'hbb905870),
	.w5(32'h3c217687),
	.w6(32'h3a973c60),
	.w7(32'hbac2b925),
	.w8(32'h3bbefe99),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb00d5c),
	.w1(32'h3b867477),
	.w2(32'hbbeff432),
	.w3(32'hbaa1543b),
	.w4(32'h3ad3ce68),
	.w5(32'hbc2c911d),
	.w6(32'hbbf4b6ef),
	.w7(32'h3a44207f),
	.w8(32'hbc2f4990),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe6253),
	.w1(32'h3beadf8c),
	.w2(32'h3bddc956),
	.w3(32'hbc3e4f79),
	.w4(32'h3c0f2c62),
	.w5(32'h3c4a397e),
	.w6(32'hbc44a66f),
	.w7(32'h3c2d6ead),
	.w8(32'h3c4f67d6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba189213),
	.w1(32'h3b5b73dc),
	.w2(32'hbac8917c),
	.w3(32'h3b807f13),
	.w4(32'h3c77f71c),
	.w5(32'h3ac2bc7c),
	.w6(32'h3baddae1),
	.w7(32'hb8d128aa),
	.w8(32'hbbd69cd4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fe8a5),
	.w1(32'hbc378d12),
	.w2(32'hbbcf80a6),
	.w3(32'hbc9328b5),
	.w4(32'hbc31f6cc),
	.w5(32'hbbff5b0f),
	.w6(32'hbba94908),
	.w7(32'hbc64d16a),
	.w8(32'hbc1d1d1f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc445efa),
	.w1(32'hbb4ea553),
	.w2(32'h3b706716),
	.w3(32'hbc527c59),
	.w4(32'hba6ba8d3),
	.w5(32'h3c621516),
	.w6(32'hbc3008f6),
	.w7(32'hbb17c374),
	.w8(32'h3c26a288),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d6724),
	.w1(32'h3b3bb399),
	.w2(32'hbc0b7f5b),
	.w3(32'h3c9a1bbf),
	.w4(32'h3bdcaa41),
	.w5(32'hbc2eaf0c),
	.w6(32'h3c4aecaa),
	.w7(32'h3bbe3777),
	.w8(32'hbc2d6e48),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ef162),
	.w1(32'h3b5e7e38),
	.w2(32'h38cd4eea),
	.w3(32'hbb9ed163),
	.w4(32'hbacb0482),
	.w5(32'h3a8a4525),
	.w6(32'hbb96dc79),
	.w7(32'h3abe728d),
	.w8(32'h3a86f1d8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1d40a),
	.w1(32'hbb0c04fa),
	.w2(32'h3b8c6ad4),
	.w3(32'h3b838537),
	.w4(32'hbb91acc1),
	.w5(32'h3b55fd49),
	.w6(32'h3b32edd2),
	.w7(32'hbb8b7780),
	.w8(32'hbab501dd),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41586c),
	.w1(32'h3b2a0306),
	.w2(32'h3b0c2662),
	.w3(32'h3a74da3a),
	.w4(32'hbac1cd63),
	.w5(32'hbb7142e2),
	.w6(32'h3aa49ccc),
	.w7(32'hbb8ed288),
	.w8(32'h3aa2d305),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d4ecc),
	.w1(32'h3b894f44),
	.w2(32'h3b156850),
	.w3(32'h3bac58ba),
	.w4(32'h3b8b701d),
	.w5(32'hba2599f0),
	.w6(32'h3a64305b),
	.w7(32'h3b7e3086),
	.w8(32'hbb2f3404),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb0434),
	.w1(32'h3b9e2c84),
	.w2(32'h3c76fec2),
	.w3(32'hbbc970e2),
	.w4(32'h3c3d57a5),
	.w5(32'h3c8b74f7),
	.w6(32'hbba8e944),
	.w7(32'h3c2f5fdc),
	.w8(32'h3c86d277),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bc678),
	.w1(32'hbba183dc),
	.w2(32'hbcb1afa2),
	.w3(32'h3caa611e),
	.w4(32'hbbf1f9d7),
	.w5(32'hbd0ef35c),
	.w6(32'h3c9cf8ea),
	.w7(32'hbc46365b),
	.w8(32'hbcd2ad77),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4605c8),
	.w1(32'h3bb9c4bf),
	.w2(32'hbae0b22c),
	.w3(32'hbcab4f5c),
	.w4(32'h3bacad63),
	.w5(32'h3bc0d192),
	.w6(32'hbc85cfe5),
	.w7(32'h3be1d74d),
	.w8(32'h3b9715d5),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4d4a0),
	.w1(32'h3bb501f0),
	.w2(32'h3bcb0f26),
	.w3(32'hbb48646b),
	.w4(32'h3ba4a62d),
	.w5(32'h3b5721c4),
	.w6(32'hba87e84f),
	.w7(32'h3bbaa92f),
	.w8(32'h3bef0cc2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52dc2c),
	.w1(32'h3b9480c2),
	.w2(32'h3a9e610d),
	.w3(32'h3ba42d79),
	.w4(32'hbb65b9a5),
	.w5(32'hbb8a3c2e),
	.w6(32'h3b9c4edb),
	.w7(32'hbaea1c68),
	.w8(32'hbbb15707),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a1a1),
	.w1(32'hbaa0a17b),
	.w2(32'h3c4166b4),
	.w3(32'hbc0bcc7b),
	.w4(32'hba83c997),
	.w5(32'h3ca0fa39),
	.w6(32'hbb0a6d08),
	.w7(32'h3b7d78a8),
	.w8(32'h3c23e3d2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c315139),
	.w1(32'h3bf1e2d5),
	.w2(32'h3afc352e),
	.w3(32'h3c87ec48),
	.w4(32'h3c181127),
	.w5(32'h3c8f1189),
	.w6(32'h3c6f4a82),
	.w7(32'h3c13fea1),
	.w8(32'h3c1f1fb8),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a25b8),
	.w1(32'hbba03a15),
	.w2(32'h3ca6e307),
	.w3(32'hbc063b16),
	.w4(32'hbbb542ff),
	.w5(32'h3d27d28f),
	.w6(32'hbc0321e3),
	.w7(32'hbc196f70),
	.w8(32'h3c21a0de),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bd2ce),
	.w1(32'h3a9c1015),
	.w2(32'hbb6f54b4),
	.w3(32'h3cbe4ebb),
	.w4(32'h3bd28a3b),
	.w5(32'h3a8f38cc),
	.w6(32'h3c14166a),
	.w7(32'h3bae0f9d),
	.w8(32'hbaa09927),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb643194),
	.w1(32'h3a4bdb07),
	.w2(32'h3b429209),
	.w3(32'hbae5073c),
	.w4(32'h3bb61c96),
	.w5(32'h3b4614e9),
	.w6(32'h390963c0),
	.w7(32'h3b126885),
	.w8(32'h3a182b0b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0bcc8),
	.w1(32'hbc06d69c),
	.w2(32'hbc6f1f60),
	.w3(32'hbb41a03e),
	.w4(32'hbba95d78),
	.w5(32'hbc615439),
	.w6(32'hbb29a14f),
	.w7(32'hbbe2d496),
	.w8(32'hbc7819b5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc649728),
	.w1(32'h3a0db1bb),
	.w2(32'h3a3d4cac),
	.w3(32'hbc87b028),
	.w4(32'hb89d1973),
	.w5(32'h3b8ce9c3),
	.w6(32'hbc951237),
	.w7(32'hbb973ed3),
	.w8(32'hbb63401e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956b406),
	.w1(32'h3adcf566),
	.w2(32'h3bf9a64b),
	.w3(32'h3ac0b889),
	.w4(32'h3befbd42),
	.w5(32'h3c004135),
	.w6(32'hbab46530),
	.w7(32'h3b9763ec),
	.w8(32'h3b532ff4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b672640),
	.w1(32'hbb4c79ce),
	.w2(32'hbc134d80),
	.w3(32'hba3c4724),
	.w4(32'hbbaa3297),
	.w5(32'hbc44031e),
	.w6(32'hbb007dde),
	.w7(32'hbadcad20),
	.w8(32'hbbdc336d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5afc252),
	.w1(32'hbb476ea6),
	.w2(32'h3bbfb57e),
	.w3(32'hbbfa30fb),
	.w4(32'hbad0324e),
	.w5(32'h3c45dfb0),
	.w6(32'hbbee7f7c),
	.w7(32'hbc3ca9b0),
	.w8(32'hba678b19),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a220458),
	.w1(32'h3b94e643),
	.w2(32'hba9952f8),
	.w3(32'h3ba09302),
	.w4(32'h3b3ae933),
	.w5(32'hb9101002),
	.w6(32'hbb0f6757),
	.w7(32'hb6bc7662),
	.w8(32'hbb5059ab),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cf93f),
	.w1(32'h3ba56bea),
	.w2(32'h3b2dc65c),
	.w3(32'hbb3129ca),
	.w4(32'h3c3a0d05),
	.w5(32'h3c134fc1),
	.w6(32'hbaa204bf),
	.w7(32'h3c395f18),
	.w8(32'h3bdb420a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6b1e6),
	.w1(32'h3bf3eed9),
	.w2(32'hb8fcaab5),
	.w3(32'h3c0a2b47),
	.w4(32'h3b12012b),
	.w5(32'hbbe64c5a),
	.w6(32'h3bbb4035),
	.w7(32'h3a50e2fd),
	.w8(32'hbba14c45),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe85475),
	.w1(32'hbc07503c),
	.w2(32'h3b552bbb),
	.w3(32'hbc1db514),
	.w4(32'hbc497977),
	.w5(32'h3bcc2fea),
	.w6(32'hbb9320db),
	.w7(32'hbc190611),
	.w8(32'h3adc6e84),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7146a),
	.w1(32'hbb83e606),
	.w2(32'h3bc1551a),
	.w3(32'hbbd91727),
	.w4(32'hbbcd7217),
	.w5(32'h3b641514),
	.w6(32'hbbf94870),
	.w7(32'hb9d68e8c),
	.w8(32'h3b60e2bf),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf9d3e),
	.w1(32'hbb932ccd),
	.w2(32'hbc023f83),
	.w3(32'h3c1e3b81),
	.w4(32'hbbbbeb5f),
	.w5(32'hbb744b77),
	.w6(32'h3bdfe560),
	.w7(32'hbadc9d2a),
	.w8(32'hbb80d2bd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7972c05),
	.w1(32'hbb9b5c1c),
	.w2(32'h3c4a98c1),
	.w3(32'h3943f9b9),
	.w4(32'hbbc0ff22),
	.w5(32'h3aa67498),
	.w6(32'h39ada838),
	.w7(32'h3b27e30a),
	.w8(32'h3a9d8465),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c202429),
	.w1(32'h3a9734e6),
	.w2(32'hbb229068),
	.w3(32'h3c13e794),
	.w4(32'h3bb1cc6f),
	.w5(32'hba104a50),
	.w6(32'h3b5897cd),
	.w7(32'h3b17d2a1),
	.w8(32'hbb8e348b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde9e1b),
	.w1(32'h3b99e2bc),
	.w2(32'h3ae162cb),
	.w3(32'h39a6345c),
	.w4(32'h39d620ef),
	.w5(32'h3ac4354f),
	.w6(32'hbb5d54a6),
	.w7(32'h3c238ea7),
	.w8(32'h3bc59077),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ca9ad),
	.w1(32'hbad09f50),
	.w2(32'h3b83285e),
	.w3(32'hbc878715),
	.w4(32'h39d9396d),
	.w5(32'h3c3002e7),
	.w6(32'h3aa7a133),
	.w7(32'h39db82e5),
	.w8(32'h3c52b21f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152c0a),
	.w1(32'hbbab1345),
	.w2(32'h3a3f3408),
	.w3(32'h3aeab10c),
	.w4(32'h3bbd7da0),
	.w5(32'h3ae92b07),
	.w6(32'h3b3f1aea),
	.w7(32'h3a87ec9c),
	.w8(32'h3b709675),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86f4b6),
	.w1(32'h3b09a016),
	.w2(32'hb8971708),
	.w3(32'hbb268734),
	.w4(32'h3b256dfc),
	.w5(32'h3cdb447a),
	.w6(32'hbacf303e),
	.w7(32'hbbcb2237),
	.w8(32'h3b828be0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd261ce),
	.w1(32'hb74f5846),
	.w2(32'h3ae092f8),
	.w3(32'h3b951191),
	.w4(32'hba6c67ec),
	.w5(32'h3bec676d),
	.w6(32'hba8e246d),
	.w7(32'h3b89faea),
	.w8(32'h3b8de8ce),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b990386),
	.w1(32'h3c89bc86),
	.w2(32'h3c4be0f6),
	.w3(32'h3a84c5ee),
	.w4(32'h3c1e9d67),
	.w5(32'h3a762c52),
	.w6(32'h3a91fc94),
	.w7(32'h3bf3c3db),
	.w8(32'h3c512025),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc40714),
	.w1(32'h3a017087),
	.w2(32'hbb04c37b),
	.w3(32'h3a29b454),
	.w4(32'h3a2eefe8),
	.w5(32'hbade1aa2),
	.w6(32'h3c359cf0),
	.w7(32'h3c0a6de5),
	.w8(32'h3c34cdb9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c775e07),
	.w1(32'hba859f5d),
	.w2(32'hb68b1733),
	.w3(32'h385b3c35),
	.w4(32'hbae8fd05),
	.w5(32'h3ba855c4),
	.w6(32'h39e0204e),
	.w7(32'h3a4973a7),
	.w8(32'h3a1dc526),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b128b83),
	.w1(32'h3ca67ffa),
	.w2(32'h3cb11d47),
	.w3(32'h3bd6ac5c),
	.w4(32'h3c84d5ff),
	.w5(32'h3d23d330),
	.w6(32'h3b80f326),
	.w7(32'hbbb37cbf),
	.w8(32'h3c9fd7a7),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c2cde),
	.w1(32'h399d499d),
	.w2(32'hbbb9c4da),
	.w3(32'h3b125712),
	.w4(32'hbc0dd6e4),
	.w5(32'hbcd3d017),
	.w6(32'h3c6b953f),
	.w7(32'h3c46eb6b),
	.w8(32'hbbb0cdf8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c3379),
	.w1(32'hb979831c),
	.w2(32'h39da3968),
	.w3(32'hbbbd5f1a),
	.w4(32'hba6bd6e2),
	.w5(32'h3a0964dd),
	.w6(32'hbb2c4f36),
	.w7(32'hb9d5e750),
	.w8(32'hbb8f346a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d0c6e),
	.w1(32'h3ba9a1b2),
	.w2(32'hba8c51b3),
	.w3(32'hbb365a2c),
	.w4(32'h3bd30f56),
	.w5(32'h3a968051),
	.w6(32'hbaebc13b),
	.w7(32'h3b414491),
	.w8(32'hb8811587),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9da18),
	.w1(32'hbac4b11d),
	.w2(32'h3b88b9cc),
	.w3(32'h3bc1ad87),
	.w4(32'hbac0e6b5),
	.w5(32'h3b6a3e56),
	.w6(32'h3ae4f775),
	.w7(32'h3c3ec8ac),
	.w8(32'h3ac5d90a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f4653),
	.w1(32'hba35e55d),
	.w2(32'hba909aab),
	.w3(32'h3badeda4),
	.w4(32'h3b14af59),
	.w5(32'h3b83582b),
	.w6(32'h3afe735d),
	.w7(32'h3bc5f329),
	.w8(32'h3bfedd33),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0bc89),
	.w1(32'hbc6e0dc7),
	.w2(32'hbc044104),
	.w3(32'hbb682217),
	.w4(32'hbc387086),
	.w5(32'h3a3abb77),
	.w6(32'h3a6ec7b5),
	.w7(32'hbc11c0dc),
	.w8(32'hbc2f668f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a37c),
	.w1(32'h3bb4bb1c),
	.w2(32'h3a7531f3),
	.w3(32'hbc687eb1),
	.w4(32'h3b1d833d),
	.w5(32'h3cff86ec),
	.w6(32'hbc08c303),
	.w7(32'hbc4f6561),
	.w8(32'h3b9b2d33),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2713b4),
	.w1(32'h3b25eba9),
	.w2(32'hbc43d146),
	.w3(32'h3b440a4a),
	.w4(32'hba651423),
	.w5(32'h3c411bbe),
	.w6(32'h3c5c93a4),
	.w7(32'hbb99b26b),
	.w8(32'hbc22ec20),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bcbaa),
	.w1(32'hbad6efab),
	.w2(32'hbb4eb1fa),
	.w3(32'hbb65d8ee),
	.w4(32'hbb16637e),
	.w5(32'hbae3180f),
	.w6(32'h3bc6c39a),
	.w7(32'h3c053ed8),
	.w8(32'h3c7664ba),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b592910),
	.w1(32'hbaf24e1d),
	.w2(32'hbbd04ee8),
	.w3(32'h3b4cc7f9),
	.w4(32'hbb1a0f79),
	.w5(32'h3c1b7ae4),
	.w6(32'h3b9e4dcd),
	.w7(32'hbc05aee6),
	.w8(32'h3b57c09c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc506b34),
	.w1(32'hbc11cd5e),
	.w2(32'hbc6ff332),
	.w3(32'hbb7773aa),
	.w4(32'hbc0cd12d),
	.w5(32'hbb70db65),
	.w6(32'h3ab818cb),
	.w7(32'hbc134313),
	.w8(32'hbb5a904f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf13484),
	.w1(32'h3bb22a9d),
	.w2(32'h3be4188c),
	.w3(32'h3bd67320),
	.w4(32'h3cd8218d),
	.w5(32'h3ce57171),
	.w6(32'h39aae40e),
	.w7(32'h3b280a21),
	.w8(32'hbb6a3097),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a4729),
	.w1(32'hbb2fd9e8),
	.w2(32'hbbe76753),
	.w3(32'h3c618de9),
	.w4(32'hbbc7400e),
	.w5(32'h3c199b21),
	.w6(32'hba954b7f),
	.w7(32'hbb342ca2),
	.w8(32'hbb5aef2a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3bab2),
	.w1(32'hbad2da86),
	.w2(32'hbbf034a6),
	.w3(32'h3b121c85),
	.w4(32'hba91b5fa),
	.w5(32'hbb8b8692),
	.w6(32'h3ab60ab8),
	.w7(32'h3b487276),
	.w8(32'hbb9b8cf1),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba157573),
	.w1(32'h3c4bb50c),
	.w2(32'h3b969f84),
	.w3(32'hba2ff42c),
	.w4(32'h3d0703b2),
	.w5(32'h3cfe3514),
	.w6(32'hba140e4b),
	.w7(32'h3c8957c6),
	.w8(32'h3d0353d4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b858fbc),
	.w1(32'h3ba0a591),
	.w2(32'h3be42506),
	.w3(32'h3ca493f3),
	.w4(32'hbc7963a2),
	.w5(32'hbbc26045),
	.w6(32'h3c9e274a),
	.w7(32'hbbe0997d),
	.w8(32'h3b794405),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc507f60),
	.w1(32'hbbcc3057),
	.w2(32'hbbe67b89),
	.w3(32'hbc6fae34),
	.w4(32'hbb07be6f),
	.w5(32'hbc35b43f),
	.w6(32'h3b16827b),
	.w7(32'hbb9a7c50),
	.w8(32'hbbb6dbd6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edbf08),
	.w1(32'hbb5c3458),
	.w2(32'hbab3e1ba),
	.w3(32'hbafc9cd7),
	.w4(32'hbb0cbefe),
	.w5(32'hbb62fd86),
	.w6(32'hbb81ddce),
	.w7(32'hb9d8220c),
	.w8(32'hbc10bf06),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ea226),
	.w1(32'hbae88ac9),
	.w2(32'hbc2b9a66),
	.w3(32'h3aef2738),
	.w4(32'h3b87291f),
	.w5(32'h3b0b9940),
	.w6(32'hbb944df9),
	.w7(32'hbbce0b72),
	.w8(32'hbbd28220),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb9747),
	.w1(32'h3bb033df),
	.w2(32'h3bbafa73),
	.w3(32'h3b140285),
	.w4(32'hbc31967a),
	.w5(32'h396eb708),
	.w6(32'hbba99e5e),
	.w7(32'h3beef9ac),
	.w8(32'hbb7049fa),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00ce5),
	.w1(32'h3b5ae285),
	.w2(32'hbbd4c19e),
	.w3(32'hbac70417),
	.w4(32'h3c14b423),
	.w5(32'h3bbc7014),
	.w6(32'hba624ea3),
	.w7(32'h3c09baf5),
	.w8(32'h3c2ab3dd),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf8162),
	.w1(32'h3af766db),
	.w2(32'h3b7d4ee8),
	.w3(32'h3be97cf1),
	.w4(32'hbb073fa6),
	.w5(32'h3c330658),
	.w6(32'h3c0d5000),
	.w7(32'hba8a48dd),
	.w8(32'h3731287a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb970efa9),
	.w1(32'h3c3d2125),
	.w2(32'h3b276524),
	.w3(32'hbb5babe7),
	.w4(32'h3b6802e5),
	.w5(32'hbb9760eb),
	.w6(32'hbb6175dc),
	.w7(32'h3b96cb1c),
	.w8(32'hbb84e0c5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf86fb),
	.w1(32'hba0040d0),
	.w2(32'h3b29739d),
	.w3(32'hbb899f0c),
	.w4(32'hbae7423b),
	.w5(32'h3b41cfe1),
	.w6(32'hbb0a9576),
	.w7(32'h3bb3c6de),
	.w8(32'hba1843b9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f05b5),
	.w1(32'hbb13e45a),
	.w2(32'hbbefc326),
	.w3(32'hbbc79b63),
	.w4(32'h3a87a113),
	.w5(32'hbbe58291),
	.w6(32'h3962e3a2),
	.w7(32'h3b8df28f),
	.w8(32'hbac0d584),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2937f5),
	.w1(32'hbb8968ec),
	.w2(32'hbb5efdcb),
	.w3(32'hbbe513ef),
	.w4(32'h3bc38a8c),
	.w5(32'h3b11f7a5),
	.w6(32'hbba77892),
	.w7(32'h3bbc691d),
	.w8(32'hbad32292),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393144bb),
	.w1(32'h3b1e336a),
	.w2(32'h3bd5f8ab),
	.w3(32'h3b25bd81),
	.w4(32'hb93cfabe),
	.w5(32'h3b093009),
	.w6(32'h3a4d4721),
	.w7(32'hbb39a569),
	.w8(32'hbafdcd8b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca7e3d),
	.w1(32'hbae89f28),
	.w2(32'h3b83443d),
	.w3(32'h3990cbae),
	.w4(32'hbc204c09),
	.w5(32'hbc05b6e2),
	.w6(32'hb9242589),
	.w7(32'hba6395a4),
	.w8(32'hbb92aa96),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7017cf),
	.w1(32'hbba8df66),
	.w2(32'hb9d47b9e),
	.w3(32'h3c1aeeb5),
	.w4(32'hbbea8aa8),
	.w5(32'hbaf783cf),
	.w6(32'h3b3c26dc),
	.w7(32'hbb3f5584),
	.w8(32'hbc05af53),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab44e78),
	.w1(32'h3b49fbbf),
	.w2(32'h3b8d6e84),
	.w3(32'hbb8e0b92),
	.w4(32'h3bc0020e),
	.w5(32'h3c229784),
	.w6(32'hba4d633a),
	.w7(32'hbb8ab462),
	.w8(32'hba303a77),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e7c4),
	.w1(32'h3b535921),
	.w2(32'h3c7841c0),
	.w3(32'h3b46eac2),
	.w4(32'hba4df5c3),
	.w5(32'hbbb507d3),
	.w6(32'hb9eb3931),
	.w7(32'h3ab2b220),
	.w8(32'h3b50b9a0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba30637),
	.w1(32'hbbbd1559),
	.w2(32'hba4efab4),
	.w3(32'hba8f5d86),
	.w4(32'h3affbe82),
	.w5(32'hb9c09c4f),
	.w6(32'h39fd33a6),
	.w7(32'h3b6a0bb2),
	.w8(32'h3bfedbbd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdf585),
	.w1(32'hbb984a75),
	.w2(32'hb9f67bf7),
	.w3(32'h3a7643b6),
	.w4(32'hb9fabca2),
	.w5(32'hba67fdb7),
	.w6(32'hbbd73e1a),
	.w7(32'h39eaaabf),
	.w8(32'h3a74cf4c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14d1ba),
	.w1(32'h3b3b5306),
	.w2(32'h3c6cb3f7),
	.w3(32'h3b7cc87e),
	.w4(32'h3aac6210),
	.w5(32'h3b5ecadc),
	.w6(32'h3b900d80),
	.w7(32'h3ac49abd),
	.w8(32'hbbd72e6a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b296eab),
	.w1(32'hb9a70f92),
	.w2(32'hbb12527d),
	.w3(32'h3b8a223a),
	.w4(32'h3c6d7582),
	.w5(32'h3b8f6387),
	.w6(32'h3abdead5),
	.w7(32'h3c1a20c9),
	.w8(32'hbb1b92cb),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2d199),
	.w1(32'h3a80d1ec),
	.w2(32'hbb4a200d),
	.w3(32'hbc180e4f),
	.w4(32'h38c65aa8),
	.w5(32'hbacb29fd),
	.w6(32'hb9360e17),
	.w7(32'h3b1b170c),
	.w8(32'hbb31c39b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27b347),
	.w1(32'h3bfcc02c),
	.w2(32'h3ad83abe),
	.w3(32'h3be80383),
	.w4(32'h3bb742eb),
	.w5(32'h3c8a5c55),
	.w6(32'h3aab5543),
	.w7(32'h3b70ee0f),
	.w8(32'h3c06ade2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17b38f),
	.w1(32'h3c246954),
	.w2(32'h3b4ed47a),
	.w3(32'h3b963ea7),
	.w4(32'h3c8a5bb3),
	.w5(32'h3bc07100),
	.w6(32'h3c3501d4),
	.w7(32'h3c651747),
	.w8(32'h3b9a3824),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a94e0),
	.w1(32'hb99790ea),
	.w2(32'hbb6c8ec4),
	.w3(32'h3aae60b3),
	.w4(32'hbb9bd03a),
	.w5(32'h3bb5650e),
	.w6(32'h3bbe722b),
	.w7(32'hbbe80215),
	.w8(32'h3b2b9308),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c85c0),
	.w1(32'h3c072b49),
	.w2(32'h3c08cfa7),
	.w3(32'hbb6f36ab),
	.w4(32'hbb21bdab),
	.w5(32'h3bb63ccf),
	.w6(32'hba4a40c3),
	.w7(32'h3b247ff2),
	.w8(32'h3b84d020),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8da893),
	.w1(32'h39507515),
	.w2(32'hba912306),
	.w3(32'h3b05cc99),
	.w4(32'hbb4d0e1a),
	.w5(32'hbbfdebe3),
	.w6(32'h3bd129d0),
	.w7(32'hbb855798),
	.w8(32'hbaf71c9b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb22fe9),
	.w1(32'hbb39e01a),
	.w2(32'hbbcea990),
	.w3(32'hbae5e861),
	.w4(32'hbb594cca),
	.w5(32'hbc1004b1),
	.w6(32'hba3f0f7e),
	.w7(32'hbbbac838),
	.w8(32'hbc869605),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2719cd),
	.w1(32'h39aa6c4f),
	.w2(32'hbb883fd3),
	.w3(32'hbb037190),
	.w4(32'h3b6fd896),
	.w5(32'hbbc47cf0),
	.w6(32'hbb7761be),
	.w7(32'h3b45d424),
	.w8(32'hbb7cc9a0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc817a3),
	.w1(32'hbc067918),
	.w2(32'h3b774ca8),
	.w3(32'h3c00be94),
	.w4(32'hbb7dbbba),
	.w5(32'h3bcc4dd2),
	.w6(32'hba419f80),
	.w7(32'h3b9db5a4),
	.w8(32'h3b09d2c5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04d83c),
	.w1(32'hbb8d4ef6),
	.w2(32'hbb345ea4),
	.w3(32'h3c202c25),
	.w4(32'hbabdd74a),
	.w5(32'h3a8c5879),
	.w6(32'hba8a873f),
	.w7(32'h3c0a3b7d),
	.w8(32'h3b7b93e6),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9faf04),
	.w1(32'hbb854c76),
	.w2(32'hbbc5b3a0),
	.w3(32'hbbcbb5e9),
	.w4(32'h3c0dc247),
	.w5(32'h3c03167c),
	.w6(32'h3a8990fd),
	.w7(32'hbb4396f0),
	.w8(32'hbb5c06e2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc031adb),
	.w1(32'hbb92e7fe),
	.w2(32'hbb8ae7ff),
	.w3(32'h3a662b46),
	.w4(32'h3af466db),
	.w5(32'h3bff4a82),
	.w6(32'hbac11933),
	.w7(32'hbc738215),
	.w8(32'h3c0c4ae0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a494f6d),
	.w1(32'hbbbac849),
	.w2(32'hbbbf3897),
	.w3(32'hbb8c7935),
	.w4(32'hbacbfa06),
	.w5(32'h3b1fce80),
	.w6(32'hbc575405),
	.w7(32'h3acb6f6d),
	.w8(32'hbb17c8ea),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule