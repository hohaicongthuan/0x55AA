module layer_10_featuremap_90(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49176a),
	.w1(32'h3b1a8ff5),
	.w2(32'hbaf4a7be),
	.w3(32'hbab018be),
	.w4(32'h38b77e46),
	.w5(32'h3b839fb9),
	.w6(32'hbb92dd28),
	.w7(32'hbb3bc7a1),
	.w8(32'h3b6090e3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb4aca),
	.w1(32'hbadf20b6),
	.w2(32'h3997cf88),
	.w3(32'h3be8220c),
	.w4(32'hb8fea87c),
	.w5(32'hbb1503d4),
	.w6(32'h38d6936e),
	.w7(32'hba813262),
	.w8(32'h3a233641),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52cd3e),
	.w1(32'h3b28ee48),
	.w2(32'h3b871658),
	.w3(32'h3ac9e3a5),
	.w4(32'h3bc39365),
	.w5(32'hbb429ca5),
	.w6(32'hbc29d049),
	.w7(32'hb9267d2b),
	.w8(32'h3a82c823),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a695a6e),
	.w1(32'h3ba5046f),
	.w2(32'h3b5aee27),
	.w3(32'hbb4a34b1),
	.w4(32'hbb92f260),
	.w5(32'h3b50e8f7),
	.w6(32'h3ad893ca),
	.w7(32'h3b573349),
	.w8(32'h3a29f8ff),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c6973),
	.w1(32'h3bcd9c57),
	.w2(32'h3b4cb383),
	.w3(32'hbaf3698b),
	.w4(32'hbb4fa0b4),
	.w5(32'h39b0d9bd),
	.w6(32'hbadab070),
	.w7(32'hbb3697de),
	.w8(32'hbca101cd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0d371),
	.w1(32'h39afd925),
	.w2(32'h39fc31f7),
	.w3(32'h3b528777),
	.w4(32'h3add085b),
	.w5(32'h3ab83dfd),
	.w6(32'hbbc47d12),
	.w7(32'hba236e5d),
	.w8(32'hba1429a9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ffe62),
	.w1(32'h3b7c62d7),
	.w2(32'h39cd196d),
	.w3(32'hbac59d2a),
	.w4(32'h3c014e8a),
	.w5(32'h3cc7db6c),
	.w6(32'hbbf4cfce),
	.w7(32'hbad491ec),
	.w8(32'h3bf5f229),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6a07c),
	.w1(32'h3b919cbb),
	.w2(32'h3ab51e2a),
	.w3(32'h3af0c9d7),
	.w4(32'h3b0ec1e9),
	.w5(32'hb9e22a88),
	.w6(32'h3b288f19),
	.w7(32'h3add6282),
	.w8(32'h39f4ce7b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944b9a),
	.w1(32'h3c8e27d6),
	.w2(32'h3ba05ad7),
	.w3(32'h3b0b98ee),
	.w4(32'h3b3f1b94),
	.w5(32'hbb2cd611),
	.w6(32'hbb4241b4),
	.w7(32'hb7c6c848),
	.w8(32'h39815654),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c464f79),
	.w1(32'h3bb74325),
	.w2(32'h3b417137),
	.w3(32'h3b41b882),
	.w4(32'h3b3de795),
	.w5(32'hbb3710b3),
	.w6(32'h3bcec3b1),
	.w7(32'h3a60328a),
	.w8(32'hba4473a0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3879501b),
	.w1(32'hbb8a6e73),
	.w2(32'h3b06b529),
	.w3(32'h3a051221),
	.w4(32'hbb31d48a),
	.w5(32'hbc4b669a),
	.w6(32'hbadf027e),
	.w7(32'h39f32495),
	.w8(32'hba474134),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43606c),
	.w1(32'h3ae1c036),
	.w2(32'h3c5f75cc),
	.w3(32'hbbb38354),
	.w4(32'h3c102767),
	.w5(32'h3bae3f34),
	.w6(32'hbbe6677d),
	.w7(32'hbaaf586d),
	.w8(32'h3bacaaba),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86f255),
	.w1(32'h3be74896),
	.w2(32'h3a71254b),
	.w3(32'h3bcf00c5),
	.w4(32'h3c3bafe9),
	.w5(32'hba158650),
	.w6(32'h3c55c17e),
	.w7(32'h3c4f0036),
	.w8(32'hbb3523bf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce06433),
	.w1(32'hba5b0458),
	.w2(32'hbb200682),
	.w3(32'h3af50a00),
	.w4(32'hbc48f803),
	.w5(32'h3a91e3da),
	.w6(32'h3afae577),
	.w7(32'h3bd1085e),
	.w8(32'hba864b89),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54027c),
	.w1(32'h3c0d3937),
	.w2(32'hba9ee1a3),
	.w3(32'h3b8f7400),
	.w4(32'h3b80cdf7),
	.w5(32'hbc16e253),
	.w6(32'hba27eeef),
	.w7(32'h3b70aeb4),
	.w8(32'hbaf0b386),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83e5fd),
	.w1(32'h3b868865),
	.w2(32'h3b933689),
	.w3(32'h3cbd57cf),
	.w4(32'h3bee8fde),
	.w5(32'hbba694f1),
	.w6(32'h3c4b3c50),
	.w7(32'h3b3dcf82),
	.w8(32'h3c5fc40f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de2c1d),
	.w1(32'h3cb08a3d),
	.w2(32'hba1b1c28),
	.w3(32'hbb8cb5b4),
	.w4(32'hb9a8c038),
	.w5(32'hbc7298c3),
	.w6(32'h3b799839),
	.w7(32'hbab578ed),
	.w8(32'h3a24fdb8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b539734),
	.w1(32'hbb1d8d0b),
	.w2(32'hbc142cdb),
	.w3(32'h3b28310f),
	.w4(32'h3c1f2196),
	.w5(32'h3ba2e885),
	.w6(32'h3bad48cd),
	.w7(32'hbc00eb38),
	.w8(32'h3ae1484e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c434e),
	.w1(32'h3b58baf8),
	.w2(32'h3aea0b58),
	.w3(32'h3b946fb3),
	.w4(32'h3a41306d),
	.w5(32'hba41a096),
	.w6(32'h3b8523b2),
	.w7(32'h3ba1d5da),
	.w8(32'hba5bde11),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a286),
	.w1(32'h3af379c1),
	.w2(32'hbb86a473),
	.w3(32'hbba0fb1b),
	.w4(32'h3c1d9f82),
	.w5(32'h3b1ade81),
	.w6(32'h378f0f28),
	.w7(32'hbb0ebd16),
	.w8(32'hbb89fc14),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa94a64),
	.w1(32'hbb317c51),
	.w2(32'h3be55492),
	.w3(32'hbb27b1af),
	.w4(32'h396c41fb),
	.w5(32'hbad59f88),
	.w6(32'hb87443d8),
	.w7(32'hbaa7ae56),
	.w8(32'h3a1ad070),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad3c62),
	.w1(32'h398da9db),
	.w2(32'h3ac92292),
	.w3(32'h39d3c6db),
	.w4(32'hbaa1b308),
	.w5(32'hba491c58),
	.w6(32'h39247ff7),
	.w7(32'h3943a227),
	.w8(32'h39341560),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73146b),
	.w1(32'h3b75cddc),
	.w2(32'hbc88ba76),
	.w3(32'h3c5a5da9),
	.w4(32'h3bde4a5d),
	.w5(32'hbc617be6),
	.w6(32'h3c01a266),
	.w7(32'h3c027dd9),
	.w8(32'h3bb06e49),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17684b),
	.w1(32'h3bddac6a),
	.w2(32'hbbc0d7ce),
	.w3(32'h3c081db2),
	.w4(32'h3b6625c2),
	.w5(32'hbb318de0),
	.w6(32'h3c28a5af),
	.w7(32'h3bc97d5d),
	.w8(32'hbaebae95),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae954b),
	.w1(32'h3b43af85),
	.w2(32'hbb15a0e7),
	.w3(32'h3c18b08c),
	.w4(32'h3c05ee2e),
	.w5(32'hbb848aed),
	.w6(32'h3c4baf02),
	.w7(32'h3c6916dc),
	.w8(32'hb9b1b318),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace8b70),
	.w1(32'hbaf604b6),
	.w2(32'h3bb42bb2),
	.w3(32'hbb4de69d),
	.w4(32'hbc92731d),
	.w5(32'h3b5e6e58),
	.w6(32'hbb6ff14b),
	.w7(32'h39ab2bc2),
	.w8(32'h3a87861e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83bc14),
	.w1(32'h39cef978),
	.w2(32'h38c92b5d),
	.w3(32'h3b5aa07a),
	.w4(32'h39465195),
	.w5(32'h394a302d),
	.w6(32'hba78aa47),
	.w7(32'h3822c3de),
	.w8(32'h397d7eb3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ebc16),
	.w1(32'hbb7901ed),
	.w2(32'h3b0d952a),
	.w3(32'h3a85898d),
	.w4(32'h3b2d5205),
	.w5(32'h3ce5e90d),
	.w6(32'hbae90e80),
	.w7(32'hbb3f63d2),
	.w8(32'h3abba392),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb451822),
	.w1(32'hba9c90ba),
	.w2(32'hbcbea02d),
	.w3(32'hbb552a56),
	.w4(32'hbab2cdb2),
	.w5(32'h3aee6bfa),
	.w6(32'hbb9899ff),
	.w7(32'hbaea270c),
	.w8(32'h3a4a5374),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a349acf),
	.w1(32'h3a53b3a3),
	.w2(32'hbb6809a4),
	.w3(32'h3bdb0bc0),
	.w4(32'hbcaf3444),
	.w5(32'hbb38d747),
	.w6(32'h3c0e94ad),
	.w7(32'h3b4325e2),
	.w8(32'hbba2559b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf91964),
	.w1(32'h3b19bf6e),
	.w2(32'hba204feb),
	.w3(32'h3aa23a4f),
	.w4(32'h3abac669),
	.w5(32'hb9c68722),
	.w6(32'h393cad95),
	.w7(32'h3acec1b6),
	.w8(32'h3ad21acf),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964adba),
	.w1(32'h3ab347be),
	.w2(32'hba6e4f56),
	.w3(32'hba2da9a1),
	.w4(32'h3a6f550a),
	.w5(32'hbab63c0f),
	.w6(32'h39ee3409),
	.w7(32'h3a011945),
	.w8(32'h3ada50b1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a8c21),
	.w1(32'h3b6fde7b),
	.w2(32'hbb371e29),
	.w3(32'h3b756bb9),
	.w4(32'h3b8b7b22),
	.w5(32'hbb91de69),
	.w6(32'h3b926a73),
	.w7(32'h3acdab74),
	.w8(32'hbae9736c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97b08e),
	.w1(32'hbbbaa4a1),
	.w2(32'hbbcf7d52),
	.w3(32'h3aee4ddd),
	.w4(32'h3a927c2a),
	.w5(32'hba8f86aa),
	.w6(32'h3aef0f28),
	.w7(32'h3b0222b0),
	.w8(32'hb9f201af),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a7d56),
	.w1(32'h39ff929b),
	.w2(32'hb7b42968),
	.w3(32'hb9980d8c),
	.w4(32'h3a9cc003),
	.w5(32'h3acf0b35),
	.w6(32'h3932a2e3),
	.w7(32'h3b33008a),
	.w8(32'h3b5690cc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab48ecd),
	.w1(32'h3c28413f),
	.w2(32'hbb262d3b),
	.w3(32'h3abb8aa0),
	.w4(32'h3b895b4c),
	.w5(32'h3b73d3bd),
	.w6(32'h3bd913bd),
	.w7(32'h38c526bd),
	.w8(32'hbaee3499),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53c752),
	.w1(32'hbaaa61f0),
	.w2(32'hbb6b7df7),
	.w3(32'h3ba7c8c9),
	.w4(32'hbbb3cf23),
	.w5(32'h3bb85838),
	.w6(32'h3c21622e),
	.w7(32'h3b8952bf),
	.w8(32'hbb90a672),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f72a8),
	.w1(32'hbc0ee7ab),
	.w2(32'hbb53722d),
	.w3(32'hbb0d64f7),
	.w4(32'hbc313a8c),
	.w5(32'hbbf98963),
	.w6(32'h3a2bf8ec),
	.w7(32'hbb780ae8),
	.w8(32'hba6fb612),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe99d3f),
	.w1(32'hbaf8f836),
	.w2(32'h3a9cd2cc),
	.w3(32'hba22d0db),
	.w4(32'hbba706c3),
	.w5(32'hbbc2a49b),
	.w6(32'hba1e0e7a),
	.w7(32'hbab38056),
	.w8(32'h3bd21e5d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebf0c5),
	.w1(32'hbaa817d6),
	.w2(32'hb96f9098),
	.w3(32'hba19ef4f),
	.w4(32'hbcafe73a),
	.w5(32'hb978e615),
	.w6(32'hbcff6c04),
	.w7(32'h3a0cc145),
	.w8(32'hb8b11416),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8837253),
	.w1(32'h39153ee9),
	.w2(32'h3a6f24f1),
	.w3(32'hbb822d5f),
	.w4(32'h39fcc5bd),
	.w5(32'hbaa0cce0),
	.w6(32'hb996ea02),
	.w7(32'h3a32c535),
	.w8(32'hb9ff861e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f83c6),
	.w1(32'hb9913266),
	.w2(32'h3987d312),
	.w3(32'hba0919b3),
	.w4(32'h3cc74010),
	.w5(32'hbb59960c),
	.w6(32'hba86e17f),
	.w7(32'h3b08743a),
	.w8(32'h3b781afa),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5ba04),
	.w1(32'hba8bac22),
	.w2(32'h3a8ae7e6),
	.w3(32'hbb1dead3),
	.w4(32'hba955e52),
	.w5(32'h3a5a4190),
	.w6(32'hbb4e1ddf),
	.w7(32'hbb371f5d),
	.w8(32'h39f35348),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba639e2),
	.w1(32'h3b14b0b0),
	.w2(32'hba6a8cfa),
	.w3(32'h3bb076c9),
	.w4(32'h3b14bfd6),
	.w5(32'hb960cedc),
	.w6(32'h3bf7800a),
	.w7(32'h3b77c7a3),
	.w8(32'hbb21894d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88fadd),
	.w1(32'h3cac3eb8),
	.w2(32'hbb84969b),
	.w3(32'h3bd9db1b),
	.w4(32'h3b9bd23e),
	.w5(32'h3c9f731d),
	.w6(32'h3c292340),
	.w7(32'h3bbdff13),
	.w8(32'hbab35a04),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b21b),
	.w1(32'h3bde6028),
	.w2(32'hbb702d5d),
	.w3(32'h3c2e10a5),
	.w4(32'h3b995ac1),
	.w5(32'hbd0659eb),
	.w6(32'h3b690ffb),
	.w7(32'h3c100f98),
	.w8(32'hbb3c3bcd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb338130),
	.w1(32'h37bafea2),
	.w2(32'hbb07f4e3),
	.w3(32'hbc385336),
	.w4(32'h3b8150e5),
	.w5(32'hbc853c32),
	.w6(32'h3b327a2b),
	.w7(32'h3b4eb60f),
	.w8(32'hbaf5f870),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6d4d3),
	.w1(32'h3c19279c),
	.w2(32'h3be64d33),
	.w3(32'h3a75e98e),
	.w4(32'hbc3252b0),
	.w5(32'h3c051ad6),
	.w6(32'h3c2cda16),
	.w7(32'h3c19f907),
	.w8(32'h3c08afc3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba929e1d),
	.w1(32'h39f24a09),
	.w2(32'hbb57b792),
	.w3(32'h3b56fa6f),
	.w4(32'h3aeab3b3),
	.w5(32'h3a1a6750),
	.w6(32'h3ab3c8b5),
	.w7(32'h39c609dc),
	.w8(32'h3b0db495),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a3ed4),
	.w1(32'h3b6c62c2),
	.w2(32'hb99260a5),
	.w3(32'h3b73d028),
	.w4(32'h3bf9cdc4),
	.w5(32'h3b52b86c),
	.w6(32'h3a8cfc09),
	.w7(32'h37c1ba6d),
	.w8(32'h399dd4fd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920c169),
	.w1(32'h3a8fc048),
	.w2(32'hb8a6f825),
	.w3(32'h3a14d712),
	.w4(32'h38e6658f),
	.w5(32'h39efe5ed),
	.w6(32'h392f4d82),
	.w7(32'h3b00f6cf),
	.w8(32'hba389c45),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e2ede),
	.w1(32'h3bd86608),
	.w2(32'h39a19872),
	.w3(32'h3b1b63a5),
	.w4(32'h3b9d8784),
	.w5(32'hba342d2c),
	.w6(32'hbb8c2656),
	.w7(32'h3bf07e73),
	.w8(32'h3a99ac8a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a222c79),
	.w1(32'h39437d6c),
	.w2(32'hbac8dea4),
	.w3(32'h3a816a79),
	.w4(32'h3a2bdfcb),
	.w5(32'hbb07d9e4),
	.w6(32'h3abe64c8),
	.w7(32'h3a962ed0),
	.w8(32'h3b50ec0a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24a57d),
	.w1(32'h3c17fe4a),
	.w2(32'h3b8ddbeb),
	.w3(32'h3bd7b480),
	.w4(32'h3c003c6c),
	.w5(32'h3b8cf7f3),
	.w6(32'h3c184729),
	.w7(32'h3b4a9551),
	.w8(32'h3b60fb23),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac11a15),
	.w1(32'h3a84de9c),
	.w2(32'h3b216f67),
	.w3(32'h3858e6dd),
	.w4(32'hbaa77f28),
	.w5(32'h3b2d8e3d),
	.w6(32'h3b0ca64a),
	.w7(32'hbaf6dc25),
	.w8(32'hb7a7f6cc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a805dff),
	.w1(32'h3a8c7d1f),
	.w2(32'h3afa6ea9),
	.w3(32'hbaecf1b5),
	.w4(32'h3b483c71),
	.w5(32'h3a1e3276),
	.w6(32'h3aec759d),
	.w7(32'h3b87bd6c),
	.w8(32'hbbfd8174),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4ee42),
	.w1(32'hbac1f16c),
	.w2(32'h3aa0631a),
	.w3(32'h3b07bd13),
	.w4(32'h3b034f7b),
	.w5(32'h3b46e416),
	.w6(32'h3c8b5849),
	.w7(32'hbb299f0c),
	.w8(32'hba2fc82a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9852447),
	.w1(32'h3ad2fd13),
	.w2(32'h39ac758d),
	.w3(32'hbbe24ca9),
	.w4(32'hbb09c889),
	.w5(32'hbaa134dc),
	.w6(32'h3b146d73),
	.w7(32'hbac09184),
	.w8(32'h391f365d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5d8a8),
	.w1(32'h398fc79e),
	.w2(32'h3b931d6d),
	.w3(32'hbaed5a58),
	.w4(32'h3b746cb3),
	.w5(32'h3a9aaf04),
	.w6(32'hb9c3925f),
	.w7(32'h39889b6e),
	.w8(32'h3b42bc79),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b70c),
	.w1(32'h3a9b6d1a),
	.w2(32'hbb233a5b),
	.w3(32'hbbc279d4),
	.w4(32'hbb020d53),
	.w5(32'h3b86e7b7),
	.w6(32'hba09a2e8),
	.w7(32'h3a163631),
	.w8(32'hba079ae4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb316a0b),
	.w1(32'h3bb9b283),
	.w2(32'h3a95705f),
	.w3(32'h3b3b1753),
	.w4(32'h3af330cc),
	.w5(32'h3a84e209),
	.w6(32'h3bee029b),
	.w7(32'h3a797827),
	.w8(32'h3a263128),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cc85d),
	.w1(32'hbb073503),
	.w2(32'h3b091653),
	.w3(32'h3b2edf2e),
	.w4(32'hb91552ef),
	.w5(32'h3c904680),
	.w6(32'h3b4a0b66),
	.w7(32'h3b8e6cbc),
	.w8(32'h3a7d9c94),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30116e),
	.w1(32'h39a03713),
	.w2(32'hbb9c1a01),
	.w3(32'hbb83b5aa),
	.w4(32'hba94d9a0),
	.w5(32'h3a9b1833),
	.w6(32'hbab509fe),
	.w7(32'hba69e693),
	.w8(32'h3b1f0c6c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0531a),
	.w1(32'hbc1d1149),
	.w2(32'h3c5f86fc),
	.w3(32'h3b91d1d3),
	.w4(32'hbb84fb4a),
	.w5(32'h3b82e55e),
	.w6(32'hbaaf1d26),
	.w7(32'h3b79acd7),
	.w8(32'hbbd4d19f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cc296),
	.w1(32'h3af1c901),
	.w2(32'h3a78df33),
	.w3(32'hba453537),
	.w4(32'hbaa9db19),
	.w5(32'hb99f8cea),
	.w6(32'h39fac1ee),
	.w7(32'h3a6b62c5),
	.w8(32'hbaad6e1d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eb5f1),
	.w1(32'h38d45bf7),
	.w2(32'hb9b3829d),
	.w3(32'h3b2e785b),
	.w4(32'hb9457dd1),
	.w5(32'h3722ecd2),
	.w6(32'h3c12a300),
	.w7(32'h3c5f39ee),
	.w8(32'h3b3d252d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14ae0d),
	.w1(32'h3b26f6ce),
	.w2(32'h3b66df41),
	.w3(32'h3c3b14f4),
	.w4(32'h3a7331e2),
	.w5(32'h3bfb6eee),
	.w6(32'h3ade47b3),
	.w7(32'hbba7f491),
	.w8(32'hb94e2d66),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2bbe5),
	.w1(32'h3bb8138c),
	.w2(32'hbc8577ea),
	.w3(32'h3c566d73),
	.w4(32'h3c1a250f),
	.w5(32'hbbfbba38),
	.w6(32'h3c40db45),
	.w7(32'h3bede80d),
	.w8(32'hbc0f9d10),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b71a4),
	.w1(32'h3bd58718),
	.w2(32'h3914b762),
	.w3(32'h3b3bac3d),
	.w4(32'h3b83f603),
	.w5(32'hbb0a6212),
	.w6(32'h3bdd4048),
	.w7(32'h3c3d7fbb),
	.w8(32'h3b5e7de5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9c4b2),
	.w1(32'h3c0c8748),
	.w2(32'hbb8550eb),
	.w3(32'h3bbcba33),
	.w4(32'h3c148016),
	.w5(32'hbbb51dee),
	.w6(32'h3c61a6df),
	.w7(32'h3c91617c),
	.w8(32'h3c262998),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4e8ee),
	.w1(32'hbbe0e9dc),
	.w2(32'h3b7f445e),
	.w3(32'hbb3b2f5f),
	.w4(32'h3ac7de7c),
	.w5(32'hbb078431),
	.w6(32'hbb7d2295),
	.w7(32'h3a0d6eb4),
	.w8(32'hbb5510d5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a35a5),
	.w1(32'h3b2c344e),
	.w2(32'hba1a52c5),
	.w3(32'h3a8883e6),
	.w4(32'h3b130a80),
	.w5(32'hbab215b3),
	.w6(32'h3a29c156),
	.w7(32'hbb16c2a3),
	.w8(32'hbb8b2be5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199dfe),
	.w1(32'h3a3ed63d),
	.w2(32'h3aac102e),
	.w3(32'hbb006cc3),
	.w4(32'h3913a928),
	.w5(32'h3ba7a73f),
	.w6(32'hbb0220e6),
	.w7(32'hbac8ce92),
	.w8(32'h3b47c964),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a460515),
	.w1(32'h3a998d54),
	.w2(32'hbbfa1d41),
	.w3(32'h3ab77e84),
	.w4(32'h3bbb9ea1),
	.w5(32'hb844b399),
	.w6(32'h3c501083),
	.w7(32'h3a9817af),
	.w8(32'hbb2ba4fa),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa486d0),
	.w1(32'h3b4efa27),
	.w2(32'h38d1f2c8),
	.w3(32'hbb161395),
	.w4(32'h3c567714),
	.w5(32'h3b4ea988),
	.w6(32'h3bc12f6d),
	.w7(32'hbb9a2bc1),
	.w8(32'h3b1d426e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2a889),
	.w1(32'hba078158),
	.w2(32'h36e8b6e4),
	.w3(32'h3b4c65b8),
	.w4(32'h3ba1663c),
	.w5(32'h3ba44530),
	.w6(32'h3b7214d5),
	.w7(32'h3ba3fd7b),
	.w8(32'hbb47b9f2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb68e04),
	.w1(32'h3a36eb9e),
	.w2(32'hba8ad95e),
	.w3(32'hbb3af76b),
	.w4(32'h3bc022ac),
	.w5(32'h3b2f39b2),
	.w6(32'h3bd7bc8f),
	.w7(32'h3bdcc23f),
	.w8(32'hba53104e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa894bb),
	.w1(32'h3bb59d48),
	.w2(32'h39aacb08),
	.w3(32'h3c08fe67),
	.w4(32'h3bdf7ee6),
	.w5(32'hbb2611af),
	.w6(32'h3bf82513),
	.w7(32'hbb25c5cf),
	.w8(32'h3c112a43),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e659b),
	.w1(32'h3b3b551a),
	.w2(32'hba67d4cb),
	.w3(32'h3b68dc16),
	.w4(32'h3adbde90),
	.w5(32'hbb5b7832),
	.w6(32'h3b69c393),
	.w7(32'h3a5d99a9),
	.w8(32'hbb4539c4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf69769),
	.w1(32'h3abd6d52),
	.w2(32'hbc987282),
	.w3(32'h3b594ecc),
	.w4(32'h3ba3f632),
	.w5(32'h3b7a76c9),
	.w6(32'h3b4f4456),
	.w7(32'hbae14b9c),
	.w8(32'h38705aab),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa5b2f),
	.w1(32'h3b3ff136),
	.w2(32'h3a0dd884),
	.w3(32'h3aefcf8f),
	.w4(32'h3b33991f),
	.w5(32'hba8e064a),
	.w6(32'h3aaa696b),
	.w7(32'h3bad85b4),
	.w8(32'h3b71defb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bce70),
	.w1(32'h3be9afe1),
	.w2(32'hb88bf0af),
	.w3(32'h3b586124),
	.w4(32'h3bf12d25),
	.w5(32'h3bad9598),
	.w6(32'h3b8b2e9a),
	.w7(32'h3bfcbf31),
	.w8(32'h3bafd573),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a9f4b),
	.w1(32'hbbb5edd7),
	.w2(32'h3adb6c29),
	.w3(32'hbb8517d4),
	.w4(32'hba8d2647),
	.w5(32'h3a11cc77),
	.w6(32'h3bb37437),
	.w7(32'hbbe707bb),
	.w8(32'h3b491d61),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42778c),
	.w1(32'h38b5f9ad),
	.w2(32'h39725cc0),
	.w3(32'hbaeb2b95),
	.w4(32'h3ad44a19),
	.w5(32'h3c079664),
	.w6(32'h3b16f9d7),
	.w7(32'h3b22c58f),
	.w8(32'hbc180642),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba477ff0),
	.w1(32'h3bb7d2c8),
	.w2(32'hbc018274),
	.w3(32'h3b5ca937),
	.w4(32'h3c9b05a7),
	.w5(32'hbb4e4945),
	.w6(32'hba6bf727),
	.w7(32'hb8b07da9),
	.w8(32'h3ab4c4b6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b57cc6),
	.w1(32'h39baf12c),
	.w2(32'hbbdf50bd),
	.w3(32'hbb3c8a2c),
	.w4(32'hbaf86375),
	.w5(32'hbb9d50e6),
	.w6(32'hbb39943b),
	.w7(32'h3c990bac),
	.w8(32'h399c8390),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92c78f),
	.w1(32'h3d121a06),
	.w2(32'h3ba77f40),
	.w3(32'hba935afe),
	.w4(32'hbb4194d3),
	.w5(32'hbc220638),
	.w6(32'hba11e64a),
	.w7(32'h39670da2),
	.w8(32'h3b05ead0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891144),
	.w1(32'hbc05097d),
	.w2(32'hbb30cdf8),
	.w3(32'hbb2c78be),
	.w4(32'h3909764c),
	.w5(32'h3c1ce924),
	.w6(32'hbb3732f2),
	.w7(32'hb98886d5),
	.w8(32'h3b8ef4df),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccd922),
	.w1(32'h3b8d42c7),
	.w2(32'hbbc6ae4c),
	.w3(32'h3c209e85),
	.w4(32'h3c78298e),
	.w5(32'h3b72dedf),
	.w6(32'h3ac05e11),
	.w7(32'hb8ce97ba),
	.w8(32'hba85d453),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9963f),
	.w1(32'hb9ad5c7e),
	.w2(32'h3aa8c59f),
	.w3(32'hba6570a3),
	.w4(32'hbbc52743),
	.w5(32'h3b647916),
	.w6(32'h3bb92931),
	.w7(32'h3a954951),
	.w8(32'h3b8802d2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02bde3),
	.w1(32'hbbb8993d),
	.w2(32'hb9bae3f0),
	.w3(32'hba885762),
	.w4(32'hb9075035),
	.w5(32'hb9763bfa),
	.w6(32'hbc0cc1e8),
	.w7(32'h399c8a3b),
	.w8(32'h3a040c8b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7029be),
	.w1(32'h3b1fa251),
	.w2(32'hbb4db028),
	.w3(32'h378fbf2e),
	.w4(32'hbc0cbf33),
	.w5(32'hbc19c34f),
	.w6(32'hbb813f74),
	.w7(32'hba95422f),
	.w8(32'hbb3d1404),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e6efd),
	.w1(32'h3ad58139),
	.w2(32'hbbda8fc2),
	.w3(32'h3bbabd4d),
	.w4(32'h3b2fea06),
	.w5(32'h3a2dd561),
	.w6(32'h3ba7e1c7),
	.w7(32'h3a88a2f0),
	.w8(32'hbbe7995a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ce7a5),
	.w1(32'h3b87eaea),
	.w2(32'hbbc4c9e8),
	.w3(32'h3b08ed4d),
	.w4(32'h3abaddb7),
	.w5(32'hbb9398da),
	.w6(32'h3c2c2bfd),
	.w7(32'hbb1ef7a0),
	.w8(32'hbb1bfb8a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc41ba3),
	.w1(32'h3b4b3cba),
	.w2(32'hba95c10c),
	.w3(32'h3a13f789),
	.w4(32'h3b2b1e9f),
	.w5(32'hba81b411),
	.w6(32'h3b84e6dc),
	.w7(32'hba11e756),
	.w8(32'h3b80797c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966dfc0),
	.w1(32'hbbb69cbe),
	.w2(32'hbb40f2de),
	.w3(32'h3a8314bf),
	.w4(32'h3be1ed45),
	.w5(32'hbb7d7d66),
	.w6(32'hbb34046e),
	.w7(32'h3b400dc5),
	.w8(32'hbb0651f5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d9f68),
	.w1(32'h3c2e6fb4),
	.w2(32'h3aa43dcc),
	.w3(32'h3b18dc20),
	.w4(32'h3a332395),
	.w5(32'h3b6bc8b3),
	.w6(32'h3ba95fbd),
	.w7(32'h3badb3b4),
	.w8(32'h3a051166),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ebd6f),
	.w1(32'h3c3f49a5),
	.w2(32'hba2f7e5f),
	.w3(32'h3bb42840),
	.w4(32'h3bb61012),
	.w5(32'hbb19c379),
	.w6(32'h3c17f673),
	.w7(32'hbaca819c),
	.w8(32'h3b8e9dd5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaecb90),
	.w1(32'hbb1b2acd),
	.w2(32'hba8694cc),
	.w3(32'hbbf8a15e),
	.w4(32'h3c23b2bc),
	.w5(32'h3cac8dbc),
	.w6(32'h3b003554),
	.w7(32'hbaa72291),
	.w8(32'hbb8841ba),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c876ed0),
	.w1(32'h3ca661e8),
	.w2(32'h3b446a03),
	.w3(32'h3c1c531a),
	.w4(32'h3bbe3dc8),
	.w5(32'h3b6a0701),
	.w6(32'h3c785ef8),
	.w7(32'h3c21ce60),
	.w8(32'h3b9d4e38),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba24ee5),
	.w1(32'hbc57d07c),
	.w2(32'h3a37e784),
	.w3(32'hbb309528),
	.w4(32'hbc8a48ad),
	.w5(32'hbc12ee67),
	.w6(32'hbbf0f784),
	.w7(32'hbc33e15c),
	.w8(32'hb98ebecb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a6a51),
	.w1(32'h3b5b49bc),
	.w2(32'hbba5726d),
	.w3(32'h3c2a58f0),
	.w4(32'h3b0db770),
	.w5(32'hbbcac458),
	.w6(32'h3c888bdf),
	.w7(32'h3c0db599),
	.w8(32'hbbc1a9fe),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0090a5),
	.w1(32'h3a7837ec),
	.w2(32'hbaeac12a),
	.w3(32'h3bf7eb0d),
	.w4(32'h3b1dfd3a),
	.w5(32'h3b169f67),
	.w6(32'h3ae0e4cd),
	.w7(32'h3ba93bc1),
	.w8(32'h3af8ce34),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc42aaa),
	.w1(32'hbaf979c4),
	.w2(32'h3beb1bf4),
	.w3(32'h3a4dc910),
	.w4(32'h3b56d1e0),
	.w5(32'hbb1ed42a),
	.w6(32'hbbdd45a8),
	.w7(32'hba46704c),
	.w8(32'h3ba136b5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5511b0),
	.w1(32'h3c4dbc87),
	.w2(32'h3bede055),
	.w3(32'h3cde84d6),
	.w4(32'h3c351d0f),
	.w5(32'hbbac8063),
	.w6(32'h3c0eb6b9),
	.w7(32'h3c1ef5f6),
	.w8(32'hbab3cf4e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d3dbd),
	.w1(32'h3c2960ea),
	.w2(32'h3b535425),
	.w3(32'hbb64a2bb),
	.w4(32'h3b72fdf4),
	.w5(32'h3b4d1eaf),
	.w6(32'hbbf41d56),
	.w7(32'hbb1dda29),
	.w8(32'h3c2f1d12),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19f8e9),
	.w1(32'h3b857ba2),
	.w2(32'h3b897b9b),
	.w3(32'h3b46afdd),
	.w4(32'hb91d38e8),
	.w5(32'h39790c49),
	.w6(32'h39313553),
	.w7(32'hba97644d),
	.w8(32'hb79758ae),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fee92),
	.w1(32'h3b139ae7),
	.w2(32'h39ab0d71),
	.w3(32'h3afd544d),
	.w4(32'hb9ce7577),
	.w5(32'h39476215),
	.w6(32'h3ab97104),
	.w7(32'h3a87efbd),
	.w8(32'h3b49ab8e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d15cbd5),
	.w1(32'h3b4424d2),
	.w2(32'h3b3a1056),
	.w3(32'h3a492ed9),
	.w4(32'hbae08955),
	.w5(32'hbb40cc66),
	.w6(32'h3b43b26c),
	.w7(32'h3b08b961),
	.w8(32'h3c262f1b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec99b2),
	.w1(32'h3a9cfec4),
	.w2(32'hbb9fa45a),
	.w3(32'h3bf2077e),
	.w4(32'h3bbd980f),
	.w5(32'hba73b1de),
	.w6(32'h3c2c9bd8),
	.w7(32'h3ba689b4),
	.w8(32'hbbbbafab),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8329b1),
	.w1(32'h3bb304fa),
	.w2(32'hbb9e9749),
	.w3(32'h3b560c82),
	.w4(32'hbba8e1b0),
	.w5(32'hbb95b1db),
	.w6(32'hbb58ee8c),
	.w7(32'hbbb1ac79),
	.w8(32'hba2a70e5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9376c3),
	.w1(32'h38e5055b),
	.w2(32'hbac3afaf),
	.w3(32'h3b5de4c8),
	.w4(32'h3af8b981),
	.w5(32'hba85e52e),
	.w6(32'h3ace45dd),
	.w7(32'h3b95d5e1),
	.w8(32'hbb469a6b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39d0b6),
	.w1(32'hbc0660dd),
	.w2(32'hba625ea5),
	.w3(32'h39d5e6f5),
	.w4(32'hbb1fd5d6),
	.w5(32'h3bca5f59),
	.w6(32'h3bbbe808),
	.w7(32'h3b454b7c),
	.w8(32'h3b3d078f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4cbd2),
	.w1(32'h3b913cea),
	.w2(32'hbb1e978f),
	.w3(32'h3cc51861),
	.w4(32'h3ba94de1),
	.w5(32'h3a0ae469),
	.w6(32'h3b55728e),
	.w7(32'hbab8f95e),
	.w8(32'hbb53cca5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb166b),
	.w1(32'hbae39878),
	.w2(32'h3a078616),
	.w3(32'h3b65b117),
	.w4(32'h3b40fa87),
	.w5(32'hbc3897aa),
	.w6(32'h3a8ac125),
	.w7(32'h3b371b55),
	.w8(32'hbc064ea3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b1fd),
	.w1(32'hbbf8a45b),
	.w2(32'hbbc43a9f),
	.w3(32'hbb8de1b6),
	.w4(32'h3a052e3d),
	.w5(32'hbb8b68f0),
	.w6(32'hbb7c940a),
	.w7(32'h3bb63a40),
	.w8(32'h3af7e8ad),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba673ca3),
	.w1(32'h3ac48693),
	.w2(32'hbbb9b9ec),
	.w3(32'hba9eb990),
	.w4(32'hbaef63a4),
	.w5(32'hbb2dfc21),
	.w6(32'h3c4bcb72),
	.w7(32'h3aebbf4d),
	.w8(32'h3b389311),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95c978),
	.w1(32'h3b2fd77e),
	.w2(32'h3b05e46e),
	.w3(32'hbbc97c8e),
	.w4(32'hba8d8e74),
	.w5(32'hb8940d5b),
	.w6(32'hbbadc9c4),
	.w7(32'hbaea9126),
	.w8(32'hbb148986),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a934a4f),
	.w1(32'hbb73f671),
	.w2(32'h3c15a7a3),
	.w3(32'hb73e7b47),
	.w4(32'h3a9d5ecf),
	.w5(32'hbb65f204),
	.w6(32'hb9753442),
	.w7(32'h397fe6a9),
	.w8(32'hb911f112),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc096072),
	.w1(32'h3b1eaab0),
	.w2(32'hbbc07265),
	.w3(32'h3bbaf330),
	.w4(32'h3be431f7),
	.w5(32'hbb142c9d),
	.w6(32'h3bbcfe39),
	.w7(32'h3badd2d9),
	.w8(32'h3a94cffd),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ca265),
	.w1(32'h3bedad72),
	.w2(32'h3c2ed8b2),
	.w3(32'hbbcc9b76),
	.w4(32'hba117a6f),
	.w5(32'h3bd21a3c),
	.w6(32'hbc153ffd),
	.w7(32'h3c804dc9),
	.w8(32'h3b554c24),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f944),
	.w1(32'h3be253da),
	.w2(32'h3a0c1c03),
	.w3(32'h3bab4c85),
	.w4(32'hbb201864),
	.w5(32'hbb2bda6a),
	.w6(32'h3ac4afdc),
	.w7(32'h3b3beb48),
	.w8(32'h3b57837e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88f4f),
	.w1(32'hbb49893b),
	.w2(32'hb8edb74b),
	.w3(32'h3c261fa9),
	.w4(32'hbbbf066d),
	.w5(32'hbbbb0113),
	.w6(32'h3a713557),
	.w7(32'h3bc7dd4b),
	.w8(32'h3b6bbc21),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcc822),
	.w1(32'hbc13f355),
	.w2(32'hbb98bc8a),
	.w3(32'h3991163e),
	.w4(32'hbbad682c),
	.w5(32'hbbb8f624),
	.w6(32'hbad7a413),
	.w7(32'h3b1e559b),
	.w8(32'h3baca6bd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba281045),
	.w1(32'hbad17c9a),
	.w2(32'hbaa690e2),
	.w3(32'hba727f06),
	.w4(32'h3ab625fb),
	.w5(32'hbb954ffe),
	.w6(32'h3b099931),
	.w7(32'hbba1071b),
	.w8(32'h3af9851b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf78890),
	.w1(32'hb7b7b14f),
	.w2(32'hbb57f20f),
	.w3(32'hba064caa),
	.w4(32'h3992cbbc),
	.w5(32'hba6ac25a),
	.w6(32'hbaae1827),
	.w7(32'hb938aea3),
	.w8(32'h3b835dbf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c26a5),
	.w1(32'hba97041b),
	.w2(32'h3b0192fe),
	.w3(32'hba8b9e80),
	.w4(32'h3b48a0ff),
	.w5(32'h3d08d1c1),
	.w6(32'h3ac2106b),
	.w7(32'h39f37281),
	.w8(32'hbae332e1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af26e27),
	.w1(32'h3c70aa72),
	.w2(32'h3be4c590),
	.w3(32'hbb9b9575),
	.w4(32'hbad8f58e),
	.w5(32'h3be66349),
	.w6(32'h3b957e3d),
	.w7(32'h3ba5e481),
	.w8(32'h3bbae378),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ec39a),
	.w1(32'h3b9ae941),
	.w2(32'hbb6a2031),
	.w3(32'h3bf1dba5),
	.w4(32'h3c01b52a),
	.w5(32'hbb5a4eaa),
	.w6(32'h3b8177ca),
	.w7(32'h3b95f6a7),
	.w8(32'hbad2bc9a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fd835),
	.w1(32'hbb17d327),
	.w2(32'h3c726ac5),
	.w3(32'hb87fb8da),
	.w4(32'hbb54da09),
	.w5(32'h3b01c9fc),
	.w6(32'h3aa85e20),
	.w7(32'h3a16d8ad),
	.w8(32'hba549613),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4f196),
	.w1(32'hbae7761f),
	.w2(32'hba9a0710),
	.w3(32'h3c9b56c7),
	.w4(32'hbba0eb49),
	.w5(32'hba863d0e),
	.w6(32'h3ac40169),
	.w7(32'hbbdbaf16),
	.w8(32'h3b8639ad),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b9d89),
	.w1(32'h3c11894c),
	.w2(32'h3a8dd051),
	.w3(32'hbc1f3102),
	.w4(32'hba8b38d4),
	.w5(32'h3c97b8e0),
	.w6(32'hba9bd319),
	.w7(32'h3ac4093b),
	.w8(32'hbb871b4d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef18c5),
	.w1(32'hbb8667ee),
	.w2(32'h39c9daf4),
	.w3(32'hbb8b9684),
	.w4(32'h396dfdbe),
	.w5(32'h3a011dab),
	.w6(32'h3ac311cc),
	.w7(32'hb9972055),
	.w8(32'hbb39d92d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2e705),
	.w1(32'hbb2003af),
	.w2(32'hbc00edfe),
	.w3(32'h3b966a14),
	.w4(32'hbafa7be3),
	.w5(32'hb91cf605),
	.w6(32'h3af3987a),
	.w7(32'h3bd22dff),
	.w8(32'hbb865ccb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e3bd1),
	.w1(32'h3b62d778),
	.w2(32'h3abe5d2b),
	.w3(32'hba60dd28),
	.w4(32'h38d627b8),
	.w5(32'h3c62ee1f),
	.w6(32'h3c367c38),
	.w7(32'h3bd3fdc5),
	.w8(32'h3aab4987),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba821634),
	.w1(32'h39e8b268),
	.w2(32'hb9e3a55f),
	.w3(32'h3ba658e2),
	.w4(32'hbb21c693),
	.w5(32'hbb9535d9),
	.w6(32'h3b51ec72),
	.w7(32'h3a133812),
	.w8(32'h3ac81778),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa46419),
	.w1(32'h38aa6386),
	.w2(32'hbbb806e0),
	.w3(32'h3ab7e0ec),
	.w4(32'hbbcecaa5),
	.w5(32'hba25bb14),
	.w6(32'h3b439332),
	.w7(32'hbbd0909a),
	.w8(32'hbb81303f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb72f6b),
	.w1(32'h3b0aca68),
	.w2(32'hbbabd63c),
	.w3(32'h3bdc4993),
	.w4(32'h3be0e8ad),
	.w5(32'h3a702f09),
	.w6(32'h3bc86080),
	.w7(32'h3bce16cb),
	.w8(32'hbb55e605),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa18e7),
	.w1(32'h3ac44634),
	.w2(32'hbc175b41),
	.w3(32'hbb21cf32),
	.w4(32'h3c294b60),
	.w5(32'hbbd0d5f0),
	.w6(32'hb9aa541c),
	.w7(32'h38a7ccdf),
	.w8(32'hbc18c007),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fd7ba),
	.w1(32'h3b63ee2c),
	.w2(32'h3a71fedb),
	.w3(32'h3b28ec7b),
	.w4(32'h3b5038e0),
	.w5(32'h3bf5a713),
	.w6(32'h3ca0fcba),
	.w7(32'hbb9aeeb7),
	.w8(32'h3ac94c12),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dbd17),
	.w1(32'h3a8dc1ae),
	.w2(32'hb9e05b7b),
	.w3(32'hb9b40c0d),
	.w4(32'h3b56e6cd),
	.w5(32'hbb0d115b),
	.w6(32'h3b929d78),
	.w7(32'h3b06653d),
	.w8(32'h3a8a2874),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d5bf),
	.w1(32'hb9098715),
	.w2(32'hbb658450),
	.w3(32'h3b8243e5),
	.w4(32'hbab52c32),
	.w5(32'hbc0717dc),
	.w6(32'h3bff096c),
	.w7(32'h3cda1a59),
	.w8(32'hbb9a6c2d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf86d6a),
	.w1(32'hb9f64796),
	.w2(32'hb894cc31),
	.w3(32'h3a6797e3),
	.w4(32'hbcd4dc97),
	.w5(32'hbacfea5a),
	.w6(32'h3ab2b9bc),
	.w7(32'h3b681477),
	.w8(32'h3a4cceab),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b193026),
	.w1(32'hb9aba951),
	.w2(32'hba9c56da),
	.w3(32'h3a95f299),
	.w4(32'hba32fa89),
	.w5(32'hbac10f91),
	.w6(32'hbccc4c72),
	.w7(32'h3b06a508),
	.w8(32'h3aad10a1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2e08e),
	.w1(32'h3afeb867),
	.w2(32'h397ac40e),
	.w3(32'h3ae1f047),
	.w4(32'h3addda0c),
	.w5(32'hba2367fe),
	.w6(32'h3a9a8675),
	.w7(32'hbae5cdad),
	.w8(32'hbaf62e48),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad29927),
	.w1(32'h39bbb02e),
	.w2(32'h3b232dd2),
	.w3(32'hba8571b6),
	.w4(32'h39a4b90a),
	.w5(32'hbb31eb1c),
	.w6(32'hba49609c),
	.w7(32'h3a5d235b),
	.w8(32'h3b061b69),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34154f),
	.w1(32'hbaf2ef32),
	.w2(32'hbb959a63),
	.w3(32'h3b28aa3d),
	.w4(32'hbb1adb79),
	.w5(32'hbac2f37a),
	.w6(32'h3b87b8f7),
	.w7(32'hba998964),
	.w8(32'hbad80870),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85f2e5),
	.w1(32'h3bfafdaa),
	.w2(32'hbaba2d47),
	.w3(32'hbbc4b7c6),
	.w4(32'h39f6e6fb),
	.w5(32'hbb07e5ba),
	.w6(32'h3c245994),
	.w7(32'h3c1af00f),
	.w8(32'hb981ad6a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81404a),
	.w1(32'h3b38c76e),
	.w2(32'h3bd90c3d),
	.w3(32'h38150d42),
	.w4(32'hbacdc55b),
	.w5(32'hb98c5d26),
	.w6(32'h3ac1fc39),
	.w7(32'h3a31e8eb),
	.w8(32'hba2d8f54),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7cc6b),
	.w1(32'h3818c538),
	.w2(32'hbb6799d0),
	.w3(32'h3c97b818),
	.w4(32'h3a987aa8),
	.w5(32'h3a911427),
	.w6(32'h3c101e75),
	.w7(32'h3c19152d),
	.w8(32'hbba00c86),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e0408),
	.w1(32'h3bc1276b),
	.w2(32'hbadec40b),
	.w3(32'h3b30ed1d),
	.w4(32'h3b854fea),
	.w5(32'hbb49bae6),
	.w6(32'hbb93ba92),
	.w7(32'h3c47fdb2),
	.w8(32'hbbae327b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3433c),
	.w1(32'h3b7153c7),
	.w2(32'hbac302a9),
	.w3(32'h3b11ce83),
	.w4(32'h3b86c9fb),
	.w5(32'h3ab13839),
	.w6(32'hba6f5c38),
	.w7(32'h3b38eb28),
	.w8(32'h3abee114),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7c7be),
	.w1(32'h3b594be2),
	.w2(32'h3c0cd9a3),
	.w3(32'h3c3c0642),
	.w4(32'h3bf4d562),
	.w5(32'hbacd17fe),
	.w6(32'h3c26fdf1),
	.w7(32'h3bdbba61),
	.w8(32'hb5b824b0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0dc5c1),
	.w1(32'h3aada508),
	.w2(32'h3b09cf04),
	.w3(32'h362b574e),
	.w4(32'h3968b571),
	.w5(32'h3948ba3b),
	.w6(32'hbcbd3cb6),
	.w7(32'h39fd2774),
	.w8(32'hbbd7ac93),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b100c1),
	.w1(32'h3ace5ae8),
	.w2(32'hb96e3734),
	.w3(32'h3ade01dc),
	.w4(32'h3b04b302),
	.w5(32'h3b6c3b3e),
	.w6(32'hb8d565a5),
	.w7(32'hba61d9a3),
	.w8(32'h3aad0890),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf72de3),
	.w1(32'h399557e9),
	.w2(32'h3bea60a5),
	.w3(32'hbb0b9b07),
	.w4(32'hbaf0a708),
	.w5(32'h3ce3e743),
	.w6(32'h3cb09ce2),
	.w7(32'hbba7131a),
	.w8(32'h39863d46),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba646afb),
	.w1(32'hbb6e8c2c),
	.w2(32'hbb15c005),
	.w3(32'hba781f90),
	.w4(32'hbb3ce171),
	.w5(32'hba865cc8),
	.w6(32'hbaffd52e),
	.w7(32'hbb500191),
	.w8(32'hbb010d02),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc02b8),
	.w1(32'hbb9fe3e2),
	.w2(32'hb9dd7878),
	.w3(32'hbb0b2198),
	.w4(32'hbb0bb5de),
	.w5(32'hbab48501),
	.w6(32'hbb1de0bf),
	.w7(32'hba99079a),
	.w8(32'h39da5945),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26d6a8),
	.w1(32'hba3cf763),
	.w2(32'hba61459f),
	.w3(32'h3c8524f4),
	.w4(32'hba5ae280),
	.w5(32'h37cdbf75),
	.w6(32'h3a90253a),
	.w7(32'h3cd34f33),
	.w8(32'h3a5180b5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03d4ae),
	.w1(32'hbaaa9238),
	.w2(32'h39cbd324),
	.w3(32'h3a4f4362),
	.w4(32'h3a6e043b),
	.w5(32'hbc30490e),
	.w6(32'hbb1f5eaa),
	.w7(32'hbceaccca),
	.w8(32'hbc8471d7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b209379),
	.w1(32'h3aad8e80),
	.w2(32'hbb0a133e),
	.w3(32'h3a5a2a44),
	.w4(32'hba147cb6),
	.w5(32'h3b13aef0),
	.w6(32'h3be55e73),
	.w7(32'hbc88942c),
	.w8(32'hbb64c6ad),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85aa36),
	.w1(32'h3a841ee7),
	.w2(32'h3bbcae8c),
	.w3(32'h397d7b0a),
	.w4(32'hb8a2bae5),
	.w5(32'hbabf8966),
	.w6(32'hbcde52ae),
	.w7(32'hba9f751d),
	.w8(32'h3b6cfe43),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f2c95),
	.w1(32'h3a5077b7),
	.w2(32'hb861bca1),
	.w3(32'h3af7ad10),
	.w4(32'hbbcc727e),
	.w5(32'h394b80ce),
	.w6(32'h3bbe4834),
	.w7(32'h3b442b44),
	.w8(32'h3bd72653),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac21f53),
	.w1(32'hb9b37a35),
	.w2(32'hb943fa86),
	.w3(32'h3b582f97),
	.w4(32'hbab88387),
	.w5(32'hb9c474ee),
	.w6(32'h3c1168e5),
	.w7(32'h3ade7258),
	.w8(32'h39653182),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31415d),
	.w1(32'h3b8d4c40),
	.w2(32'hba94be33),
	.w3(32'h3b3524ea),
	.w4(32'h3b70e80b),
	.w5(32'h3aa501fc),
	.w6(32'h3b461cfd),
	.w7(32'h3b61f334),
	.w8(32'hbb1e1b9d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc262c43),
	.w1(32'hba580b59),
	.w2(32'hb9d93d5a),
	.w3(32'h3a8c2840),
	.w4(32'hbb0b5818),
	.w5(32'hba63424f),
	.w6(32'hba58eaa4),
	.w7(32'h3abc275a),
	.w8(32'hbabc53c5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae63a7),
	.w1(32'h39e1560b),
	.w2(32'h3b9df00f),
	.w3(32'hba3d9f4d),
	.w4(32'hba122d80),
	.w5(32'h3adbe8e7),
	.w6(32'hba08e69b),
	.w7(32'hbacd2caf),
	.w8(32'h3a31a247),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a798f5),
	.w1(32'hbbb3826f),
	.w2(32'h3b88d2fd),
	.w3(32'h3a6d0b4f),
	.w4(32'h3b7fe852),
	.w5(32'hbaa2f9df),
	.w6(32'h3ab1ed11),
	.w7(32'hba1ec080),
	.w8(32'h3af28f7d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5d35f),
	.w1(32'hbbdca817),
	.w2(32'hbc372e20),
	.w3(32'h3b9b9327),
	.w4(32'h3ab80a6b),
	.w5(32'hbb4da91b),
	.w6(32'h3ba7cd2e),
	.w7(32'h3b6fde42),
	.w8(32'hbba0b369),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e6b24),
	.w1(32'hbb3baaff),
	.w2(32'h3b2895b8),
	.w3(32'h3a840a77),
	.w4(32'h3b90ab15),
	.w5(32'h3d8333fc),
	.w6(32'hbc7b49d2),
	.w7(32'hbc360fb8),
	.w8(32'h388de416),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9fb7f),
	.w1(32'h399ca218),
	.w2(32'h3a5aab44),
	.w3(32'hbb9084f2),
	.w4(32'hbc45962c),
	.w5(32'hbbe457c3),
	.w6(32'h3bf5c60d),
	.w7(32'h38ef8c41),
	.w8(32'h3c74ffe3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba074e5),
	.w1(32'hbc03bedf),
	.w2(32'h3c594e72),
	.w3(32'hbaaf9ddf),
	.w4(32'h3af140b3),
	.w5(32'hbb97c975),
	.w6(32'h3baca7a1),
	.w7(32'hbb9ce533),
	.w8(32'hbb21ffb0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3127f9),
	.w1(32'hbb0b5a48),
	.w2(32'h3ba27243),
	.w3(32'h3b490634),
	.w4(32'h3bc8cdbb),
	.w5(32'hbab87b13),
	.w6(32'h3c36003a),
	.w7(32'hbb03200c),
	.w8(32'hbc138731),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d078),
	.w1(32'h3b45a9f0),
	.w2(32'hba9b918e),
	.w3(32'h3b74e931),
	.w4(32'hbb6cd69c),
	.w5(32'h3bfeaafd),
	.w6(32'h3ba1be9e),
	.w7(32'h3b04fba2),
	.w8(32'hbb8555ec),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a74c6),
	.w1(32'h3b4c4f83),
	.w2(32'hbbde83d8),
	.w3(32'h3c116dcc),
	.w4(32'h3c15c21d),
	.w5(32'hbb8cf572),
	.w6(32'h3bd1b938),
	.w7(32'hbb4b594c),
	.w8(32'hbadc6c57),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba240da),
	.w1(32'h3aa9ff05),
	.w2(32'hbbf77ce2),
	.w3(32'hbb52fd40),
	.w4(32'hbad782d2),
	.w5(32'h3bdbd09b),
	.w6(32'h3b3dcaca),
	.w7(32'h3c2f4d75),
	.w8(32'hbc023f80),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d72f1),
	.w1(32'hb95cf4a2),
	.w2(32'hbb2b6db1),
	.w3(32'hba217e4a),
	.w4(32'hbb163039),
	.w5(32'h3c246d37),
	.w6(32'h3af4edc2),
	.w7(32'hba4203c0),
	.w8(32'hbac88018),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b543),
	.w1(32'h3c48ebab),
	.w2(32'hbb840f64),
	.w3(32'hbd29295f),
	.w4(32'hbd50f8d3),
	.w5(32'hbb95bba3),
	.w6(32'hbaac9d37),
	.w7(32'h3c5d40f2),
	.w8(32'h392768b6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58da0e),
	.w1(32'h3c273329),
	.w2(32'h3b78c77e),
	.w3(32'h3abc760f),
	.w4(32'hbaaa0b4d),
	.w5(32'hbb6f0bfe),
	.w6(32'hbb0e5d77),
	.w7(32'h3c574adf),
	.w8(32'hbc932aa4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0620bb),
	.w1(32'h3b8556d1),
	.w2(32'hbbd5c154),
	.w3(32'hbb8739ed),
	.w4(32'hb9e41822),
	.w5(32'h3a9dacb2),
	.w6(32'h3a92ca6a),
	.w7(32'h393c6ccb),
	.w8(32'hbc74dc92),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ce2a9),
	.w1(32'hbc4bf0be),
	.w2(32'h390f6218),
	.w3(32'h3ab61ab3),
	.w4(32'h3b11e94c),
	.w5(32'hb99837b2),
	.w6(32'h3cd66407),
	.w7(32'hbc2d3cf4),
	.w8(32'hb7aaf1b4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978487),
	.w1(32'h3bae1023),
	.w2(32'h3c2f14d2),
	.w3(32'h3c2bc702),
	.w4(32'h3c9347b1),
	.w5(32'hbbc44ec4),
	.w6(32'h3af7fc45),
	.w7(32'hb95bb32e),
	.w8(32'h3a5e578f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b193dd8),
	.w1(32'hbb245380),
	.w2(32'h3c4e8b47),
	.w3(32'h3a8d9a7f),
	.w4(32'hb95a734a),
	.w5(32'hba1031cb),
	.w6(32'h3739040c),
	.w7(32'hb9d0b8ac),
	.w8(32'h3ab6fe4d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10d527),
	.w1(32'hbaba09cc),
	.w2(32'hbccf5c96),
	.w3(32'h3bd43f61),
	.w4(32'hbb45a2c0),
	.w5(32'h3a96c0e8),
	.w6(32'h3b0e2a6c),
	.w7(32'hb9ff9ad0),
	.w8(32'hbc0b5144),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa9bf9),
	.w1(32'h3be0ccd3),
	.w2(32'h39a3c279),
	.w3(32'hbbe5104d),
	.w4(32'hb9787759),
	.w5(32'h3b4dc7aa),
	.w6(32'hbbc38b8f),
	.w7(32'h3baadd92),
	.w8(32'hbac3dc81),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a92d0),
	.w1(32'h3b3e83bd),
	.w2(32'h3bb29ee2),
	.w3(32'h3c28402f),
	.w4(32'hbaf75b27),
	.w5(32'hbd26e59e),
	.w6(32'h3bc6a473),
	.w7(32'hbc3ae44d),
	.w8(32'h3b8cd070),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18b373),
	.w1(32'hbb3d0456),
	.w2(32'h3af42c7b),
	.w3(32'hbb1a4219),
	.w4(32'h3c16e894),
	.w5(32'h3b77b437),
	.w6(32'hb9314da7),
	.w7(32'hbc91d756),
	.w8(32'h3b247a5e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dff64),
	.w1(32'hba350e01),
	.w2(32'hbafcd94b),
	.w3(32'h3c17a5b4),
	.w4(32'h3d1fcf40),
	.w5(32'h3b8b21c1),
	.w6(32'h3bf0e262),
	.w7(32'h3c88ee9e),
	.w8(32'hbc1cf721),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718265),
	.w1(32'h3c4af6ab),
	.w2(32'hbb539f66),
	.w3(32'hbb71c878),
	.w4(32'hbbd56f85),
	.w5(32'hbc4c110d),
	.w6(32'h3caeaf1a),
	.w7(32'hbc045778),
	.w8(32'hbc2f49f3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf83b6),
	.w1(32'h3b913f85),
	.w2(32'hbb954c8c),
	.w3(32'h3bcce1d9),
	.w4(32'h3bb263c1),
	.w5(32'h3baee519),
	.w6(32'h3b7029d2),
	.w7(32'hbabb4cd6),
	.w8(32'h3b64a177),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3951b986),
	.w1(32'hbc0cea37),
	.w2(32'h3a600fd1),
	.w3(32'hbc3e1f74),
	.w4(32'h3bde7e5b),
	.w5(32'hbc092ced),
	.w6(32'hbadcb8c7),
	.w7(32'hbb330588),
	.w8(32'hbce37405),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ada51),
	.w1(32'hbc794a9d),
	.w2(32'h3c9504c1),
	.w3(32'h3ba8d2b1),
	.w4(32'hbb49c321),
	.w5(32'hbabd5c08),
	.w6(32'hbac32c30),
	.w7(32'h3a8109ad),
	.w8(32'hbb881499),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a32f3),
	.w1(32'h3942b3bf),
	.w2(32'hbb4e5800),
	.w3(32'hbb1061ef),
	.w4(32'h3a78642a),
	.w5(32'hb95b5615),
	.w6(32'h39fb456d),
	.w7(32'h3c05ae11),
	.w8(32'hbaca9fbf),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b7ff9),
	.w1(32'h3d1da4e3),
	.w2(32'h3a1c244b),
	.w3(32'h3a8f0327),
	.w4(32'hbc4e914a),
	.w5(32'h3b7623b8),
	.w6(32'h3b6927d2),
	.w7(32'hbbfe2da2),
	.w8(32'hbbf5a670),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aabbe),
	.w1(32'h3bcb49dc),
	.w2(32'h3a34dd88),
	.w3(32'h3ad8e760),
	.w4(32'h3b8bac7d),
	.w5(32'hba582366),
	.w6(32'h3b7ef8bb),
	.w7(32'h3c3079a5),
	.w8(32'hbb5e4301),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba758a3),
	.w1(32'h3b97538c),
	.w2(32'h3aaf8ab2),
	.w3(32'h3c291fdb),
	.w4(32'h3bd12d69),
	.w5(32'hbc1b7864),
	.w6(32'h3c5a4cb2),
	.w7(32'h3b19cb0a),
	.w8(32'h3b59ec30),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a089b68),
	.w1(32'h3b76c834),
	.w2(32'hbb006760),
	.w3(32'hbb8b0240),
	.w4(32'h3adb45e9),
	.w5(32'h39a6032f),
	.w6(32'hba3c170c),
	.w7(32'hbb847a86),
	.w8(32'hb837261b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24fdba),
	.w1(32'h3bbd220c),
	.w2(32'hbaa7d1cf),
	.w3(32'hbb9a689b),
	.w4(32'h3bc3d8f5),
	.w5(32'h3b12e1fc),
	.w6(32'h3b4a50d7),
	.w7(32'h3be012e5),
	.w8(32'hba65f5e4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd30b36),
	.w1(32'h3bf2d311),
	.w2(32'h3b4097ce),
	.w3(32'h3b09d6d9),
	.w4(32'h3c434fb6),
	.w5(32'hbb6e3502),
	.w6(32'hbc6146f5),
	.w7(32'hb993f67c),
	.w8(32'h3c17578e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab40b9),
	.w1(32'hbc4cbed3),
	.w2(32'h3bd69c60),
	.w3(32'h3a7fb6b0),
	.w4(32'hbb911b0d),
	.w5(32'h3aa322bd),
	.w6(32'hbb096de0),
	.w7(32'h3b0cc321),
	.w8(32'hbb7548cb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a412f01),
	.w1(32'h3c25c1f8),
	.w2(32'h3b501ace),
	.w3(32'h3b46cb4d),
	.w4(32'hbb01f598),
	.w5(32'h3ac50e45),
	.w6(32'hb97ec1e7),
	.w7(32'h3b0099ed),
	.w8(32'hbae339cd),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5582),
	.w1(32'hbc154729),
	.w2(32'h3b7cdc78),
	.w3(32'h3aeec567),
	.w4(32'hbadb5947),
	.w5(32'h3bbd1974),
	.w6(32'hba88d6e5),
	.w7(32'h3bd57e83),
	.w8(32'hb9e7ab34),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cac21),
	.w1(32'h3bbd9fe5),
	.w2(32'h3b5de882),
	.w3(32'hbae7842c),
	.w4(32'h3b98066a),
	.w5(32'h3bad53fd),
	.w6(32'h3aa69ca7),
	.w7(32'h3c69f33c),
	.w8(32'hb984e546),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5f1e),
	.w1(32'hba426272),
	.w2(32'hba8501ac),
	.w3(32'hbb38b6eb),
	.w4(32'hbc1943fe),
	.w5(32'hbb51294b),
	.w6(32'h3b6d929d),
	.w7(32'hbb7786cf),
	.w8(32'h3a61b9d8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3e2b0),
	.w1(32'hbb83b0f5),
	.w2(32'hbad3bdf2),
	.w3(32'h3aaf77ba),
	.w4(32'hbb3b8bfe),
	.w5(32'hbbad6053),
	.w6(32'h3ac0532c),
	.w7(32'h3bad0309),
	.w8(32'hbb210b53),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a763d38),
	.w1(32'hbaf9d8d5),
	.w2(32'hbc228e8f),
	.w3(32'hbb0036da),
	.w4(32'hbba350c2),
	.w5(32'hbb4166fd),
	.w6(32'hbb794bd0),
	.w7(32'hbcccdc64),
	.w8(32'h3d06c133),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09d87e),
	.w1(32'h3ba93380),
	.w2(32'hbb67ee88),
	.w3(32'hbbc3f6f5),
	.w4(32'hbb0fe577),
	.w5(32'hbc17e609),
	.w6(32'h3bf94ca9),
	.w7(32'h3b1aa373),
	.w8(32'hbb862962),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03eb67),
	.w1(32'h3baa23e7),
	.w2(32'hbb763dab),
	.w3(32'hb9c1d0f3),
	.w4(32'h3c813714),
	.w5(32'hb90c279e),
	.w6(32'h3b07bedd),
	.w7(32'h3b52c474),
	.w8(32'hbb2416b4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27ad35),
	.w1(32'h3c0784b7),
	.w2(32'hbc8fe26d),
	.w3(32'h3c8a6f0e),
	.w4(32'h3c449712),
	.w5(32'hbbd9a1b5),
	.w6(32'h3c29f1b6),
	.w7(32'h3be76e67),
	.w8(32'hba3e2cba),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cb01c),
	.w1(32'hbb804074),
	.w2(32'h3aa77378),
	.w3(32'h3b80ba49),
	.w4(32'h3a8cc7ef),
	.w5(32'hbaa5ff5f),
	.w6(32'h3a40a607),
	.w7(32'hb93651e8),
	.w8(32'hbbd964a3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85740e),
	.w1(32'h3af3da1f),
	.w2(32'hb937052c),
	.w3(32'hbb74206d),
	.w4(32'h3b9b4550),
	.w5(32'h3c8505ed),
	.w6(32'hba1da731),
	.w7(32'h3ac0126a),
	.w8(32'hb86eaae1),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd983f),
	.w1(32'h3b3b2011),
	.w2(32'hbb9fbddf),
	.w3(32'h3b91b61b),
	.w4(32'h3a8cb72f),
	.w5(32'hbae3c683),
	.w6(32'h3b99cc29),
	.w7(32'h3b9bf06a),
	.w8(32'h3b45307a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc16b46),
	.w1(32'h3b4b7094),
	.w2(32'hbb34209b),
	.w3(32'h3cc7ee61),
	.w4(32'h3b9816f0),
	.w5(32'hbbd55e5f),
	.w6(32'h3c15f052),
	.w7(32'hbc821b2b),
	.w8(32'hbbf2e73b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb217a47),
	.w1(32'h3bacee08),
	.w2(32'hba3f9d2a),
	.w3(32'h3b6d48b1),
	.w4(32'h3b4d18ad),
	.w5(32'hbb9c6b90),
	.w6(32'h3be3cfa1),
	.w7(32'h3ba2da6b),
	.w8(32'hbb259975),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba25a40),
	.w1(32'hbb05d6ea),
	.w2(32'hba00316c),
	.w3(32'hba497598),
	.w4(32'h396062c9),
	.w5(32'h3acaa1ef),
	.w6(32'h3ce668d3),
	.w7(32'hb9b044b8),
	.w8(32'h3a55ac9f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cbed1),
	.w1(32'h3ad801c5),
	.w2(32'h37dbc7d5),
	.w3(32'h3a9eb66d),
	.w4(32'h3c5afec3),
	.w5(32'h39f6ec57),
	.w6(32'hbb09d9fd),
	.w7(32'h38bb5e8b),
	.w8(32'hbc9b422f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a4f7e),
	.w1(32'h3b0cdef0),
	.w2(32'h3cb5f426),
	.w3(32'hba339fbe),
	.w4(32'hbbbca644),
	.w5(32'hbb607028),
	.w6(32'h3afc29af),
	.w7(32'hbb47915e),
	.w8(32'h395d0a3d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67a28f),
	.w1(32'h3ad686a7),
	.w2(32'hbb84f8ad),
	.w3(32'h3bad7ac5),
	.w4(32'h3b324a40),
	.w5(32'h3bd12b2d),
	.w6(32'h3b92a0ca),
	.w7(32'h3b4678fb),
	.w8(32'h3b907797),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3abe19),
	.w1(32'h3bb72fee),
	.w2(32'h3baf7689),
	.w3(32'h3b6b685b),
	.w4(32'h3bc06450),
	.w5(32'h3a38f619),
	.w6(32'h3bd71076),
	.w7(32'hbb866236),
	.w8(32'h3ba45c0c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293637),
	.w1(32'h3c77d79e),
	.w2(32'h39f091a5),
	.w3(32'hbb088c68),
	.w4(32'hbb3e73a9),
	.w5(32'hbc6036a6),
	.w6(32'h3ba55372),
	.w7(32'hb913ea1e),
	.w8(32'hba512758),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1decb),
	.w1(32'h3a2926d0),
	.w2(32'hbac08291),
	.w3(32'hbc5fcc94),
	.w4(32'hbb217953),
	.w5(32'hba8e1c99),
	.w6(32'h3b3044f7),
	.w7(32'h38a0d5fc),
	.w8(32'hba4f2886),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbcb13),
	.w1(32'hbae5dd64),
	.w2(32'h3b3bc7f1),
	.w3(32'h3be86089),
	.w4(32'hba23d210),
	.w5(32'hbc4e7c0b),
	.w6(32'h3bbb0e9a),
	.w7(32'h3a021145),
	.w8(32'hbc01b996),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c9fdc),
	.w1(32'hbb1343ce),
	.w2(32'h3b5a8891),
	.w3(32'hbada5280),
	.w4(32'hbb285a7c),
	.w5(32'h3b53e501),
	.w6(32'hbb96e887),
	.w7(32'hbaa18c61),
	.w8(32'h39503b1b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcbfe5),
	.w1(32'h3b266f6b),
	.w2(32'h3b78b02b),
	.w3(32'h3935ec12),
	.w4(32'hbbd24023),
	.w5(32'h3b8623be),
	.w6(32'hbbc626d1),
	.w7(32'hbb6875d4),
	.w8(32'hb9e252a3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e4674),
	.w1(32'hbb6976fd),
	.w2(32'hbae97bf6),
	.w3(32'hba320c24),
	.w4(32'h3a8ba6e6),
	.w5(32'hbac74b72),
	.w6(32'hb9ac6d69),
	.w7(32'hbc75d87a),
	.w8(32'hb999211a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47ae8e),
	.w1(32'hba82d350),
	.w2(32'hbb499d74),
	.w3(32'hbb9c38fe),
	.w4(32'h3a9fd04f),
	.w5(32'h3c19fe62),
	.w6(32'h3a7beeac),
	.w7(32'h3af67cd9),
	.w8(32'hbb0fdeab),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020027),
	.w1(32'hb886c149),
	.w2(32'hbb01c1b9),
	.w3(32'hbb99b5ca),
	.w4(32'h39eedd7a),
	.w5(32'hbc3aff77),
	.w6(32'hbc1346ae),
	.w7(32'h3b52f2a2),
	.w8(32'hbc30df3f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34a1a5),
	.w1(32'h3c2c0b88),
	.w2(32'h3aff2050),
	.w3(32'hba05d77b),
	.w4(32'h3bdf5ed8),
	.w5(32'h3c2ee536),
	.w6(32'h3b30e999),
	.w7(32'h3c153b43),
	.w8(32'h3aebc123),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5175f8),
	.w1(32'h3b88f230),
	.w2(32'h39f90cdf),
	.w3(32'h3ba8d326),
	.w4(32'hbbbf1efc),
	.w5(32'hbb837e4a),
	.w6(32'hba060ca0),
	.w7(32'h3c0b0e89),
	.w8(32'hbc5aaa28),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03201d),
	.w1(32'hbac9d37d),
	.w2(32'hbb796f52),
	.w3(32'h3a2b1d09),
	.w4(32'h38cf897e),
	.w5(32'h3bde3263),
	.w6(32'hbab4a1e9),
	.w7(32'h3b955f29),
	.w8(32'h39228c34),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8bba5),
	.w1(32'h3c5aaa38),
	.w2(32'h3bbf3501),
	.w3(32'hbb993a39),
	.w4(32'hbae7ec62),
	.w5(32'hbc397f49),
	.w6(32'h3bf8f1f3),
	.w7(32'h3bd5ddc3),
	.w8(32'hbc7415a5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2c954),
	.w1(32'h3bdee39b),
	.w2(32'h3c360da0),
	.w3(32'hbb9bd1fa),
	.w4(32'h3bd1314d),
	.w5(32'hbaf960f1),
	.w6(32'h3b3572a2),
	.w7(32'h3c0f26d3),
	.w8(32'h3b555601),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf757c),
	.w1(32'h3a6838f8),
	.w2(32'h3bdca126),
	.w3(32'h3c11172a),
	.w4(32'h3d544353),
	.w5(32'hbb9ef761),
	.w6(32'hbb461092),
	.w7(32'hbaac7044),
	.w8(32'h3b2288a1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8620be),
	.w1(32'h3b8d61ba),
	.w2(32'hbc47b4e2),
	.w3(32'hbadd4b4c),
	.w4(32'hbb83859c),
	.w5(32'h3bf99a50),
	.w6(32'hba819f7e),
	.w7(32'hba1395d3),
	.w8(32'h3bdc6e4a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda311c6),
	.w1(32'h3b2a5d80),
	.w2(32'h3c564e93),
	.w3(32'h3ba36d61),
	.w4(32'h3bf6cbd3),
	.w5(32'hbadda1b4),
	.w6(32'h3c16a7b9),
	.w7(32'h3b175d57),
	.w8(32'h398de2fa),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39237d),
	.w1(32'h3a991369),
	.w2(32'hba3faae7),
	.w3(32'h3b3c9274),
	.w4(32'hbb21cde5),
	.w5(32'hbac210c7),
	.w6(32'hbbb78756),
	.w7(32'hbbf47b80),
	.w8(32'h39ddc82f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3ccf8),
	.w1(32'h3b507f92),
	.w2(32'h3bb233c1),
	.w3(32'hbb67ee24),
	.w4(32'hb4142f16),
	.w5(32'hbc71bbd7),
	.w6(32'h3bf7bbb5),
	.w7(32'hbc75de2e),
	.w8(32'h389499df),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950aa1b),
	.w1(32'hbb569f58),
	.w2(32'hbbe683ed),
	.w3(32'hbc373e69),
	.w4(32'hbbc0d86c),
	.w5(32'h3bb250a4),
	.w6(32'hbc710269),
	.w7(32'h3ab609c1),
	.w8(32'h3b3097ce),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bf2d4),
	.w1(32'h3b31c142),
	.w2(32'hba5e7977),
	.w3(32'hbba20d9b),
	.w4(32'h3a1f4d25),
	.w5(32'hbb438449),
	.w6(32'h3bc3b2cf),
	.w7(32'h3b746a6f),
	.w8(32'h39026779),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d7125),
	.w1(32'h3b6f8030),
	.w2(32'hbc07951a),
	.w3(32'h3c09ee56),
	.w4(32'h3c2100de),
	.w5(32'h3b76988b),
	.w6(32'h3b9bb46f),
	.w7(32'h3bdfac2f),
	.w8(32'hbb8c3420),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac32b81),
	.w1(32'h3b74a089),
	.w2(32'h39f4f353),
	.w3(32'h39ce4c85),
	.w4(32'h3be0b207),
	.w5(32'h3c4101c3),
	.w6(32'h3a8f967b),
	.w7(32'h3bad0f00),
	.w8(32'h3bf32330),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52ab06),
	.w1(32'h3c34902c),
	.w2(32'h3b33d7f0),
	.w3(32'h3c050061),
	.w4(32'h3c0660a3),
	.w5(32'h3bb3eca3),
	.w6(32'h3b42c05f),
	.w7(32'h3a9f435f),
	.w8(32'hbb6e3b16),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaaa49),
	.w1(32'h3a4b56fd),
	.w2(32'hbc4bad19),
	.w3(32'h3bd4fabb),
	.w4(32'hbb170fd0),
	.w5(32'hbbc852f9),
	.w6(32'hbaf5b933),
	.w7(32'hbbb0c874),
	.w8(32'h3a85fbd6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3b19e),
	.w1(32'hbc54b7d2),
	.w2(32'hbb58cd7c),
	.w3(32'hbb153553),
	.w4(32'h3d03d42d),
	.w5(32'h39c753be),
	.w6(32'hbbbe3f00),
	.w7(32'hbb9587b1),
	.w8(32'h3aece896),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6069537),
	.w1(32'h3ac568f3),
	.w2(32'h3bb93a16),
	.w3(32'hbb626c09),
	.w4(32'hbadcf95f),
	.w5(32'hbba67050),
	.w6(32'h3b2ed649),
	.w7(32'hbb61feff),
	.w8(32'hbcd8de0d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc57c),
	.w1(32'hba59bd46),
	.w2(32'h3a0e6aff),
	.w3(32'h3d48c0ad),
	.w4(32'hbb230df5),
	.w5(32'hbbb4d5e3),
	.w6(32'hbba95ccc),
	.w7(32'hbb84d8c4),
	.w8(32'hbca7ff73),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb4576),
	.w1(32'hba14b03a),
	.w2(32'h3c0b90d6),
	.w3(32'h3c4f5684),
	.w4(32'hbbbb683e),
	.w5(32'h3b2dbb23),
	.w6(32'h3c4f0ac7),
	.w7(32'h3a899b03),
	.w8(32'h3b6d5aea),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4cd5e0),
	.w1(32'h3a5c01b2),
	.w2(32'h3bf9ecfc),
	.w3(32'h3c07c6e3),
	.w4(32'h39c2be82),
	.w5(32'hbbf8d905),
	.w6(32'hbbe44ae8),
	.w7(32'h3ba19d71),
	.w8(32'hb9b50b27),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba2002),
	.w1(32'h3c208090),
	.w2(32'hbb0f02d2),
	.w3(32'hbbf72635),
	.w4(32'h3c2b99a6),
	.w5(32'hbaa28eef),
	.w6(32'hbd4ac926),
	.w7(32'hbcd10a7c),
	.w8(32'hbb00d96d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd2f8e),
	.w1(32'h3ab3663f),
	.w2(32'hb9db386f),
	.w3(32'h39e78671),
	.w4(32'hba7cf49e),
	.w5(32'hb7a7eed0),
	.w6(32'hbb668ae8),
	.w7(32'hbb340ed0),
	.w8(32'h39be3791),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e7a11),
	.w1(32'hba770f22),
	.w2(32'h3b26ca75),
	.w3(32'hbc395faa),
	.w4(32'h3c12d57a),
	.w5(32'h3b09152d),
	.w6(32'h3d969b47),
	.w7(32'hbc184125),
	.w8(32'hbbcd7175),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5156c0),
	.w1(32'hbafa4730),
	.w2(32'h3c29c0c5),
	.w3(32'hbc16f788),
	.w4(32'hbc21b395),
	.w5(32'h3b6fc76e),
	.w6(32'h3b858bd4),
	.w7(32'hbc0ee65f),
	.w8(32'hbb259a44),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d9c36),
	.w1(32'hbc879a30),
	.w2(32'h3a480333),
	.w3(32'hbb784600),
	.w4(32'hbcaf3bd4),
	.w5(32'h3bfa6932),
	.w6(32'hbb3866ba),
	.w7(32'hbc351384),
	.w8(32'h3baa3cf4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f72af),
	.w1(32'h3b66ba13),
	.w2(32'h3bd25a5e),
	.w3(32'h3b90c8f1),
	.w4(32'h3bbccc99),
	.w5(32'hba6cecbc),
	.w6(32'h3c1faf71),
	.w7(32'h39d602d0),
	.w8(32'h3bb6da4f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefc8a9),
	.w1(32'h3b70c80a),
	.w2(32'h3a9b6af5),
	.w3(32'hba210e4e),
	.w4(32'h3b43e57f),
	.w5(32'hba7b628c),
	.w6(32'h3a9c3c05),
	.w7(32'hb8266b0c),
	.w8(32'hbbf5ebd2),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c19d),
	.w1(32'h3bcf9c86),
	.w2(32'hbb693aa6),
	.w3(32'hbc80a8dc),
	.w4(32'hbb98d4bc),
	.w5(32'h3b1942b1),
	.w6(32'h3b811669),
	.w7(32'h3aedb676),
	.w8(32'h3b5d3952),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule