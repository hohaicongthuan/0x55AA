module layer_10_featuremap_324(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c6291),
	.w1(32'h3bba45ed),
	.w2(32'h3b41949e),
	.w3(32'h3bf9f654),
	.w4(32'h3ba2b758),
	.w5(32'h3bd5f539),
	.w6(32'h3c36a644),
	.w7(32'h3bc27843),
	.w8(32'h3baa5c28),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08ebe6),
	.w1(32'h3c244959),
	.w2(32'h3ccd275c),
	.w3(32'h39dd3e6b),
	.w4(32'hbaf3e22a),
	.w5(32'hba1d421c),
	.w6(32'h3ad892a4),
	.w7(32'h3a9bd292),
	.w8(32'hbae8abb3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2a690),
	.w1(32'hbab5c42b),
	.w2(32'hbb4d9e21),
	.w3(32'hba6149ac),
	.w4(32'hb981b767),
	.w5(32'hbb9fb417),
	.w6(32'hbb0a3d31),
	.w7(32'hbb4a0a5b),
	.w8(32'hbb9fb456),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f9040),
	.w1(32'hbb000b2f),
	.w2(32'hb9cd324d),
	.w3(32'hbb4067c8),
	.w4(32'hb997e824),
	.w5(32'hbb591fe8),
	.w6(32'hbb567f93),
	.w7(32'hbab9d235),
	.w8(32'hbbc91c47),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32ad90),
	.w1(32'hbbaa6106),
	.w2(32'hbb9763bf),
	.w3(32'hbc2292ae),
	.w4(32'hbc22ff36),
	.w5(32'hbb2362bd),
	.w6(32'hbc29a01f),
	.w7(32'hbc3d7611),
	.w8(32'hb9c495a5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf12643),
	.w1(32'hbad46fe7),
	.w2(32'hbb237dc7),
	.w3(32'hb9d7f1e5),
	.w4(32'hbb03945b),
	.w5(32'hba87dca5),
	.w6(32'h3b145f51),
	.w7(32'hbaae6db1),
	.w8(32'hbb0e814c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c061ddf),
	.w1(32'h3b513e8d),
	.w2(32'h3b117e45),
	.w3(32'h392206a2),
	.w4(32'h3adfdbc7),
	.w5(32'hbb3c457e),
	.w6(32'h3bb60703),
	.w7(32'h3a035fce),
	.w8(32'hbc3a181a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dd725),
	.w1(32'hbc69598b),
	.w2(32'hbcbd3f9e),
	.w3(32'hba934c33),
	.w4(32'h3aca8c57),
	.w5(32'h3a4f0656),
	.w6(32'hbbb19545),
	.w7(32'hba63fac8),
	.w8(32'h3bc0507d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c292243),
	.w1(32'h3ba60adc),
	.w2(32'h3b59af56),
	.w3(32'h3bb7df94),
	.w4(32'h3b9a2170),
	.w5(32'hbbb79473),
	.w6(32'h3b8cde1a),
	.w7(32'h3b46351b),
	.w8(32'hbb872394),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb952a1d),
	.w1(32'hbbbb0148),
	.w2(32'hbc16884b),
	.w3(32'h3aa14f25),
	.w4(32'hb9e2fe1d),
	.w5(32'hbc0bba0d),
	.w6(32'h3bc25afe),
	.w7(32'h3ac92de2),
	.w8(32'hbbfa19ac),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49b357),
	.w1(32'hbb7c2cb6),
	.w2(32'hbbc77722),
	.w3(32'hbaf3da8c),
	.w4(32'hbb2706cd),
	.w5(32'h39f0e913),
	.w6(32'hbaa2f2fc),
	.w7(32'hbb80f789),
	.w8(32'hbad48bc4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c519c1e),
	.w1(32'h3c0bf9b8),
	.w2(32'hbba91465),
	.w3(32'h3b7406b4),
	.w4(32'h3bee5a9e),
	.w5(32'hbbc3c5b1),
	.w6(32'h3c0fc789),
	.w7(32'h3b8508a0),
	.w8(32'hbc39389b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f763d),
	.w1(32'hbc5c0850),
	.w2(32'hbc8b2fc1),
	.w3(32'hbb683e96),
	.w4(32'hbb7d6995),
	.w5(32'hbb02f0ab),
	.w6(32'hba235c4c),
	.w7(32'hbbe5236b),
	.w8(32'hbbdb5e76),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2da22),
	.w1(32'hbbdd9626),
	.w2(32'hbc026255),
	.w3(32'hbb0a3a0a),
	.w4(32'hbc09ba6c),
	.w5(32'hbc1ab5be),
	.w6(32'hbb2d50d5),
	.w7(32'hbc1e4f89),
	.w8(32'hbc248279),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0f8ec),
	.w1(32'hbbbfd276),
	.w2(32'hbc07899e),
	.w3(32'hbb37d05f),
	.w4(32'hba42569b),
	.w5(32'h3c04f84b),
	.w6(32'hbbdc5bf7),
	.w7(32'hbbe8c5c5),
	.w8(32'h3b0a3887),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0349c3),
	.w1(32'hbbe7a462),
	.w2(32'hbba1b61b),
	.w3(32'h3bdb1499),
	.w4(32'h3b9e467c),
	.w5(32'hbafdf188),
	.w6(32'h37e51a78),
	.w7(32'h3b32571d),
	.w8(32'h393bd9e6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00cbce),
	.w1(32'h3a9d18eb),
	.w2(32'h3b1376f5),
	.w3(32'h3abfc63d),
	.w4(32'h3a46aa8e),
	.w5(32'h3a1ec99c),
	.w6(32'h3b57c228),
	.w7(32'hba8aed1d),
	.w8(32'hba7e7eb5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3174f),
	.w1(32'hbc034be3),
	.w2(32'hbc8ecdec),
	.w3(32'h3bd0a747),
	.w4(32'h3a5c8b81),
	.w5(32'hbc3b0abe),
	.w6(32'h3b8a8f4e),
	.w7(32'h3a0b7378),
	.w8(32'hbc452ea4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a288f),
	.w1(32'hbc07ac6a),
	.w2(32'hbc4c7802),
	.w3(32'h3b877a6e),
	.w4(32'h3b073edc),
	.w5(32'hbb9f804b),
	.w6(32'h3ab62f20),
	.w7(32'hbaf9375b),
	.w8(32'hbbe2fe38),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152503),
	.w1(32'h3b0f0a82),
	.w2(32'h3b12e744),
	.w3(32'h3b2cf7d3),
	.w4(32'h3aa8dad0),
	.w5(32'h3b86c308),
	.w6(32'h3b1a246d),
	.w7(32'h3aba4394),
	.w8(32'h3b1efb4b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301512),
	.w1(32'h3b1c5eae),
	.w2(32'h3be1785c),
	.w3(32'h3ba5c42f),
	.w4(32'h3c160d8d),
	.w5(32'hbb07c020),
	.w6(32'h3b3a8a49),
	.w7(32'h3be62417),
	.w8(32'hbaef92c8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9934ef9),
	.w1(32'h3b0d9d80),
	.w2(32'h3b068b2d),
	.w3(32'h3a92734c),
	.w4(32'h3b04e730),
	.w5(32'h3b270185),
	.w6(32'hbac598bb),
	.w7(32'hbab9001c),
	.w8(32'h3b13d2ed),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94009e),
	.w1(32'hbc5c8a30),
	.w2(32'hbc5f4fb7),
	.w3(32'h3ae49200),
	.w4(32'h3c4495fd),
	.w5(32'hbb69c8d0),
	.w6(32'h3bcaf118),
	.w7(32'h3c0bafd3),
	.w8(32'hbc3bae9c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9e63e),
	.w1(32'h3ba53197),
	.w2(32'h3bfa01c1),
	.w3(32'h3c133153),
	.w4(32'h3c5185a3),
	.w5(32'hba84f622),
	.w6(32'h3c1fbd46),
	.w7(32'h3c33fb01),
	.w8(32'hbb2772d3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba123aa),
	.w1(32'h3bbc2d20),
	.w2(32'h3c384c28),
	.w3(32'hbb3d941f),
	.w4(32'hba94f3cd),
	.w5(32'hba5485ac),
	.w6(32'hbc1b3643),
	.w7(32'hbc21e015),
	.w8(32'hbbd24255),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bead6),
	.w1(32'hbb5b09ca),
	.w2(32'hbb973958),
	.w3(32'hbb30dc05),
	.w4(32'hba209dc2),
	.w5(32'h38edec67),
	.w6(32'hbaff05f7),
	.w7(32'hbaa61f60),
	.w8(32'h39ef1a64),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c7641),
	.w1(32'h39908031),
	.w2(32'hbb3d8b36),
	.w3(32'h385326c7),
	.w4(32'hbabed0c6),
	.w5(32'h3bb42994),
	.w6(32'hb9a35ee0),
	.w7(32'hbb20ae79),
	.w8(32'h3bc72ec2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb80e6),
	.w1(32'h3903b428),
	.w2(32'h3bf13b78),
	.w3(32'h3aecb54a),
	.w4(32'hbbd541d2),
	.w5(32'hbbddb451),
	.w6(32'hba162a0d),
	.w7(32'hbb3835b0),
	.w8(32'hbc0b4622),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadb859),
	.w1(32'h3b9c8e45),
	.w2(32'h3ba8b843),
	.w3(32'h3b981ef9),
	.w4(32'hbab7889e),
	.w5(32'h3a58ddf3),
	.w6(32'h3b852890),
	.w7(32'h3b2423e1),
	.w8(32'h3ac6628b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe158f),
	.w1(32'h3b6e216c),
	.w2(32'h3c74a7a7),
	.w3(32'hbb7f03bb),
	.w4(32'hba160f67),
	.w5(32'hba15cab5),
	.w6(32'hbb50b7c5),
	.w7(32'hb8885b66),
	.w8(32'hbb521da9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0366ff),
	.w1(32'hb914acbc),
	.w2(32'h3a341dca),
	.w3(32'h3b811877),
	.w4(32'h3af3dd6d),
	.w5(32'h3b9e8ab5),
	.w6(32'h3b9c3d79),
	.w7(32'h3bb1ef52),
	.w8(32'h3bfe55d1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89c110),
	.w1(32'h3bb4df98),
	.w2(32'h3bdf0feb),
	.w3(32'h3b3a08aa),
	.w4(32'h3b0a2696),
	.w5(32'hbb4611aa),
	.w6(32'h3bc748ad),
	.w7(32'h3b136623),
	.w8(32'hba0f9788),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac28d5d),
	.w1(32'hbb6d7e7d),
	.w2(32'hbbd35b04),
	.w3(32'h3b90fd82),
	.w4(32'h3b3cd0d3),
	.w5(32'hb8cbf6e5),
	.w6(32'h3b8343bc),
	.w7(32'h3a5828fd),
	.w8(32'hbb586849),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bc686),
	.w1(32'h3bab2e97),
	.w2(32'h3c0aadec),
	.w3(32'h3aa8d0b4),
	.w4(32'h39c41492),
	.w5(32'h3aa082ae),
	.w6(32'h3abbaaf9),
	.w7(32'h39d165f6),
	.w8(32'h3afc80f4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b931b83),
	.w1(32'h3aeccc1a),
	.w2(32'h3a01533b),
	.w3(32'hb7238814),
	.w4(32'h3ab25ffb),
	.w5(32'hba5f37ec),
	.w6(32'h3b1240f9),
	.w7(32'h3a50c349),
	.w8(32'hb99b6d84),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5a426),
	.w1(32'h3b212878),
	.w2(32'hbaaefb74),
	.w3(32'hbaace50f),
	.w4(32'hba4b5913),
	.w5(32'hbb5140d8),
	.w6(32'h3b02e782),
	.w7(32'hba5b45c5),
	.w8(32'hbaae8fb8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2e3af),
	.w1(32'h3c5d78d6),
	.w2(32'hbb9a25a7),
	.w3(32'hbc01edde),
	.w4(32'h3c9c1144),
	.w5(32'h3c72f897),
	.w6(32'hbb9dfa9d),
	.w7(32'h3c95a323),
	.w8(32'h3c124794),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c3e7),
	.w1(32'h3b51e60d),
	.w2(32'h3c563f85),
	.w3(32'hbbd74011),
	.w4(32'hbbddf4a4),
	.w5(32'h3c7169e4),
	.w6(32'hbc2b80bb),
	.w7(32'hbc295030),
	.w8(32'h3c3dda14),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a355d),
	.w1(32'h3c233c02),
	.w2(32'h3cb52c8c),
	.w3(32'h3bcdcd78),
	.w4(32'hbaeaa2ab),
	.w5(32'h3916e48f),
	.w6(32'h3c2303e7),
	.w7(32'h3a8962a0),
	.w8(32'hbb639fc2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f77da),
	.w1(32'hba63d9a0),
	.w2(32'h3aa05943),
	.w3(32'h3ae9e2a9),
	.w4(32'h3919cef9),
	.w5(32'h3b0ff93f),
	.w6(32'hbb277105),
	.w7(32'hbb0ad284),
	.w8(32'h3b086fef),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0488c9),
	.w1(32'hb93be183),
	.w2(32'h38d3929f),
	.w3(32'h3acbc4f4),
	.w4(32'h3729ea55),
	.w5(32'hbc161183),
	.w6(32'h39217876),
	.w7(32'h39000f98),
	.w8(32'hbbc7c1e5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd78174),
	.w1(32'hbb3e75dc),
	.w2(32'hbb6ce593),
	.w3(32'hbbaec20f),
	.w4(32'hbb966801),
	.w5(32'hbb7460fa),
	.w6(32'hbb2ca528),
	.w7(32'hbb519d3e),
	.w8(32'hbb5af6bb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e73524),
	.w1(32'h3b157511),
	.w2(32'h3b723f42),
	.w3(32'hbb59cb7b),
	.w4(32'h3ad92a2f),
	.w5(32'h38111a36),
	.w6(32'hbb36e216),
	.w7(32'h3b529e0c),
	.w8(32'hbb9cc14f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35b9da),
	.w1(32'hbc54c157),
	.w2(32'hbc504d31),
	.w3(32'hba805dc6),
	.w4(32'hbb8b42d3),
	.w5(32'hbbfe8d60),
	.w6(32'hbb8769c4),
	.w7(32'hbb8c0610),
	.w8(32'hbc0db57b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1d62),
	.w1(32'h3bb51c91),
	.w2(32'h3bfcfe0a),
	.w3(32'h3bb0b0b9),
	.w4(32'h3b9620a1),
	.w5(32'h3b4ae34d),
	.w6(32'h3bae3018),
	.w7(32'h3ba826e9),
	.w8(32'h3b2fa793),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a93e6),
	.w1(32'h3a911ec2),
	.w2(32'h3bb361ff),
	.w3(32'h3aaefdc1),
	.w4(32'h3c073ad0),
	.w5(32'h3b9278ef),
	.w6(32'h3c17a5cb),
	.w7(32'h3c59f2c2),
	.w8(32'h3c0034ef),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce1007),
	.w1(32'h39b94ff1),
	.w2(32'h3a4afc68),
	.w3(32'h3b9f2cf0),
	.w4(32'h3b183372),
	.w5(32'h3bbc14f4),
	.w6(32'h3aed0e59),
	.w7(32'h3b402b7e),
	.w8(32'h3bcf0a99),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99aba6),
	.w1(32'hbaec79d0),
	.w2(32'hbc6bcc40),
	.w3(32'h3c421233),
	.w4(32'h3c24f9df),
	.w5(32'hbc6c1618),
	.w6(32'h3bf8fa2a),
	.w7(32'h3bef0d4c),
	.w8(32'hbc2a00d1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb838467),
	.w1(32'hbb61a92d),
	.w2(32'hbba51c4c),
	.w3(32'hb8059110),
	.w4(32'hbad754e3),
	.w5(32'h3ba738be),
	.w6(32'h3b93fa00),
	.w7(32'hbab3c536),
	.w8(32'h3b8b1746),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac224f8),
	.w1(32'hbb0111d8),
	.w2(32'hba18e525),
	.w3(32'h3a2512ac),
	.w4(32'h3b466dbc),
	.w5(32'hba22890b),
	.w6(32'hbabde7fd),
	.w7(32'hb8f784d9),
	.w8(32'hbaa93906),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a20e1),
	.w1(32'h39ed8d64),
	.w2(32'h3b358ade),
	.w3(32'h3aad4c48),
	.w4(32'h3b5a151d),
	.w5(32'h3852c609),
	.w6(32'h39bdd616),
	.w7(32'h3b322020),
	.w8(32'h3979478e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8efb3),
	.w1(32'hbb3d2baf),
	.w2(32'h3b005af0),
	.w3(32'hbb9f3420),
	.w4(32'hbb66f072),
	.w5(32'hb98e9815),
	.w6(32'hba913e09),
	.w7(32'hb9c7eeee),
	.w8(32'hbb2137c5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5078ee),
	.w1(32'h3b33b0e8),
	.w2(32'hbbbd0a6d),
	.w3(32'h3b8d3bab),
	.w4(32'h3adb2a47),
	.w5(32'hba83e97e),
	.w6(32'h3bab6f19),
	.w7(32'h39951f8f),
	.w8(32'hbb305853),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a16b7),
	.w1(32'hbc7964c9),
	.w2(32'hbcb05553),
	.w3(32'h3b37e3eb),
	.w4(32'h3a117915),
	.w5(32'hbc332ff1),
	.w6(32'h3b5a4985),
	.w7(32'h3bc72f50),
	.w8(32'hbc233cb7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1640e9),
	.w1(32'hbae97a67),
	.w2(32'hbbaabe36),
	.w3(32'hbb1891a8),
	.w4(32'hbb0e8bde),
	.w5(32'hba135d76),
	.w6(32'hbb006f3c),
	.w7(32'hbb64fcb8),
	.w8(32'h3a862e3f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1713d),
	.w1(32'h3b4fc3e3),
	.w2(32'h3bec11ad),
	.w3(32'hba81ace6),
	.w4(32'hbb00eb98),
	.w5(32'h3ae14881),
	.w6(32'h3b1304f8),
	.w7(32'h3b2079ea),
	.w8(32'h3b21cef2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ce6c9),
	.w1(32'h3adc80ad),
	.w2(32'hba56ab5e),
	.w3(32'h3a9db51c),
	.w4(32'hbabc547f),
	.w5(32'h3abb2b81),
	.w6(32'hb98137b2),
	.w7(32'hbaa11943),
	.w8(32'h3aee6165),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab22419),
	.w1(32'hba6f4b27),
	.w2(32'h3b5ad9eb),
	.w3(32'h3aa3bd85),
	.w4(32'hb81f9877),
	.w5(32'h3ba10f07),
	.w6(32'h3a5cac2f),
	.w7(32'h3a72d9d7),
	.w8(32'h3b7ee12e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef3552),
	.w1(32'h3b49d12b),
	.w2(32'h3adba9d4),
	.w3(32'h3b29fac7),
	.w4(32'h3b664537),
	.w5(32'hba8429b2),
	.w6(32'hba46f863),
	.w7(32'h3aa5c780),
	.w8(32'h3b237e20),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ae064),
	.w1(32'hb98c05ca),
	.w2(32'hba8ed35f),
	.w3(32'hbba800cc),
	.w4(32'h39622139),
	.w5(32'h3bacab3d),
	.w6(32'hbadbac29),
	.w7(32'hb9ee4b86),
	.w8(32'h3b96daa7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5c245),
	.w1(32'h3a5b997f),
	.w2(32'hbb276495),
	.w3(32'h3b496256),
	.w4(32'h3b8c3b5d),
	.w5(32'hbab7b02a),
	.w6(32'h3bc0f869),
	.w7(32'h3b797ab1),
	.w8(32'hbb8771c8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eaf97),
	.w1(32'hbc5f0dd3),
	.w2(32'hbb298b42),
	.w3(32'hbb4b282c),
	.w4(32'hbbbdf1a3),
	.w5(32'hbbb96fe0),
	.w6(32'hbb3d6bb6),
	.w7(32'hbb9d9b4e),
	.w8(32'hbbfbbd14),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad766ad),
	.w1(32'hb985d098),
	.w2(32'hbad903ba),
	.w3(32'hbb8092c0),
	.w4(32'hbac01d5e),
	.w5(32'hbabddbd9),
	.w6(32'hbb3b03e2),
	.w7(32'hbb41fbaf),
	.w8(32'hbb130486),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dfedf),
	.w1(32'hba8b7e59),
	.w2(32'h3ac2fac4),
	.w3(32'h398f4597),
	.w4(32'h3a22dcdc),
	.w5(32'hbb6abdc3),
	.w6(32'hba029926),
	.w7(32'h3a031852),
	.w8(32'hbb4dc947),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8bd05),
	.w1(32'hba7934ae),
	.w2(32'h3ad7ffe6),
	.w3(32'hbb112350),
	.w4(32'h3af972bf),
	.w5(32'h3bb1b629),
	.w6(32'hba144e18),
	.w7(32'h3acc83c4),
	.w8(32'h3a60bb92),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9aa59),
	.w1(32'h3ba7c151),
	.w2(32'h3ad60025),
	.w3(32'h3b2f5c85),
	.w4(32'h3b413386),
	.w5(32'h3a87f6de),
	.w6(32'h399a0d48),
	.w7(32'hba7602f9),
	.w8(32'hba7c6651),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac78b5),
	.w1(32'hbc89a954),
	.w2(32'hbcef06b2),
	.w3(32'h3c0aecf9),
	.w4(32'h397d0d3b),
	.w5(32'hbca9173c),
	.w6(32'h3bb95c05),
	.w7(32'hb99d4533),
	.w8(32'hbc677351),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b5b52),
	.w1(32'hbb3db421),
	.w2(32'hbc927981),
	.w3(32'hbb910c7a),
	.w4(32'hbba558ce),
	.w5(32'hbbb90db4),
	.w6(32'hb95bf746),
	.w7(32'hbbd0c647),
	.w8(32'h3b209f68),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe503fb),
	.w1(32'hbc2e3210),
	.w2(32'hbc0a8018),
	.w3(32'hba836813),
	.w4(32'h3b5fdc7c),
	.w5(32'hba09d9aa),
	.w6(32'hbb7848e7),
	.w7(32'hbae68e3d),
	.w8(32'hbb3c7148),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2743),
	.w1(32'h3c18215d),
	.w2(32'h3c8ff100),
	.w3(32'hba5e555d),
	.w4(32'h3a6959d1),
	.w5(32'h3bcb7cd7),
	.w6(32'hbbfc2c83),
	.w7(32'hbc3510e8),
	.w8(32'hbaec784e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3733ab),
	.w1(32'hbb073ef9),
	.w2(32'hbb6304cd),
	.w3(32'hbad8b82e),
	.w4(32'hba991d8a),
	.w5(32'h3b26b9a6),
	.w6(32'hbae9b437),
	.w7(32'hbaf93df6),
	.w8(32'h3a9afaef),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45996),
	.w1(32'h3b7c8e65),
	.w2(32'h3b61072b),
	.w3(32'h3bedc466),
	.w4(32'h3c0e8bf2),
	.w5(32'h3b81b948),
	.w6(32'h3bb3ea60),
	.w7(32'h3bbbfa4f),
	.w8(32'h3ba9db42),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1062ec),
	.w1(32'h3c174ebf),
	.w2(32'h3baf30c7),
	.w3(32'h3b394e39),
	.w4(32'h3b27f7fb),
	.w5(32'hbbd49640),
	.w6(32'h3b865901),
	.w7(32'h3ba117ed),
	.w8(32'hbbc1d03d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cf492),
	.w1(32'hbabb40ac),
	.w2(32'h3b322797),
	.w3(32'hbb808e76),
	.w4(32'hbbc7d9de),
	.w5(32'h3b7bef39),
	.w6(32'hbb43043f),
	.w7(32'hbb01e5c7),
	.w8(32'h3aa48aa6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b488c08),
	.w1(32'h3b14ea20),
	.w2(32'h3a088bab),
	.w3(32'h3bce3bac),
	.w4(32'h3ba09ddf),
	.w5(32'hbbb779be),
	.w6(32'h3b872128),
	.w7(32'h3b093e90),
	.w8(32'hbb96bc77),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86ad75),
	.w1(32'hbbba7a9d),
	.w2(32'hbc25b871),
	.w3(32'hbaf19fb9),
	.w4(32'hbb33bbbb),
	.w5(32'h3ab4cedc),
	.w6(32'hba4e413f),
	.w7(32'hba8b7985),
	.w8(32'h3a9d839e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47762f),
	.w1(32'hbb493e25),
	.w2(32'hbc81a246),
	.w3(32'h3b11ea95),
	.w4(32'hbaa25f81),
	.w5(32'hba7ee303),
	.w6(32'h3aac902a),
	.w7(32'hbb0b062d),
	.w8(32'hbb032c56),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b58f),
	.w1(32'h3c13e71f),
	.w2(32'h3c64678d),
	.w3(32'h3bde5256),
	.w4(32'h3ba1aa3f),
	.w5(32'h3b0806a5),
	.w6(32'h3bfaea4b),
	.w7(32'h3bd416dd),
	.w8(32'hba7abf20),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0dc34),
	.w1(32'hbbbc4f2b),
	.w2(32'hbc24248b),
	.w3(32'h3b892491),
	.w4(32'h3b261e22),
	.w5(32'h3b27d359),
	.w6(32'hbaaee159),
	.w7(32'hbb23d5fc),
	.w8(32'hb950e29f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c381d2b),
	.w1(32'hbb4f98df),
	.w2(32'hbbd4ea68),
	.w3(32'h3b3c5f6a),
	.w4(32'hbab28b6a),
	.w5(32'hbc0c3a0b),
	.w6(32'h3b9e12d1),
	.w7(32'h38d2c9ae),
	.w8(32'hbc1f7c34),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4f698),
	.w1(32'hbbc885a7),
	.w2(32'hbbcc2a82),
	.w3(32'hbac41231),
	.w4(32'h3aac8413),
	.w5(32'hbabaea6d),
	.w6(32'hbc11d506),
	.w7(32'hbb80bf1d),
	.w8(32'hbb13a3ae),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fe970),
	.w1(32'hbb9efc8d),
	.w2(32'hbbe06dfc),
	.w3(32'h3ba1afb0),
	.w4(32'h3b3f342d),
	.w5(32'hbad76172),
	.w6(32'h3b37bf1e),
	.w7(32'h3b0dcdde),
	.w8(32'hbaeea40b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bb8f8),
	.w1(32'hba9c5a4c),
	.w2(32'h3b173ad7),
	.w3(32'h3b15d328),
	.w4(32'h3b8dfb96),
	.w5(32'hbc6c00e9),
	.w6(32'h3a79612d),
	.w7(32'h3a2e4da4),
	.w8(32'hbc893f86),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bb6f0),
	.w1(32'hbc518fb3),
	.w2(32'hbc656d72),
	.w3(32'hbc2d258a),
	.w4(32'hbc2c9bc4),
	.w5(32'hbb31be0f),
	.w6(32'hbc5e64b4),
	.w7(32'hbc4c3c36),
	.w8(32'hba34a9b7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a6b1e),
	.w1(32'h3ae18564),
	.w2(32'h3b38fa85),
	.w3(32'hbb221224),
	.w4(32'hbb196ce5),
	.w5(32'h3b85397a),
	.w6(32'hb888280e),
	.w7(32'hbaae8309),
	.w8(32'h3b8cf731),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baff3b4),
	.w1(32'h3b80157d),
	.w2(32'h3babd7da),
	.w3(32'h3b84da5d),
	.w4(32'h3bb5f4bf),
	.w5(32'hba0557a4),
	.w6(32'h3bd4b4e2),
	.w7(32'h3bdbb7a3),
	.w8(32'hb9d70365),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ed6c9),
	.w1(32'hba34b69f),
	.w2(32'h39ae9371),
	.w3(32'hbacafea6),
	.w4(32'hbb26ff25),
	.w5(32'hb78060d4),
	.w6(32'hbb53c653),
	.w7(32'hbb2eb0d2),
	.w8(32'h38c513eb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ff1c5),
	.w1(32'hba5aa8f7),
	.w2(32'h3b140358),
	.w3(32'hbb09e2ac),
	.w4(32'hbb1575f3),
	.w5(32'h3b2a37a3),
	.w6(32'hbaa91f52),
	.w7(32'hba2abda1),
	.w8(32'h3852d2e5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98cc00),
	.w1(32'hbbaed82a),
	.w2(32'hbb91e24a),
	.w3(32'hbb3cf7da),
	.w4(32'hbb567512),
	.w5(32'h3ade1005),
	.w6(32'hbb12613f),
	.w7(32'hbb2822a1),
	.w8(32'h3be10bdb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9cbb0),
	.w1(32'hbb5a60d3),
	.w2(32'hbbee7730),
	.w3(32'h3b478296),
	.w4(32'h3a8863fd),
	.w5(32'hbbbd42c3),
	.w6(32'hb9c41357),
	.w7(32'hba145983),
	.w8(32'hbbc5cc23),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f7573),
	.w1(32'h3c31fade),
	.w2(32'h3c487c7a),
	.w3(32'hb88e24ef),
	.w4(32'h3b2fdd01),
	.w5(32'h3bb1c50f),
	.w6(32'h3b7a13ff),
	.w7(32'h3b6b5413),
	.w8(32'h3ba87702),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeadce),
	.w1(32'hbb6a0ebd),
	.w2(32'hbc0c44d6),
	.w3(32'h3bec8c39),
	.w4(32'h3c4a4e95),
	.w5(32'hbc26f5bf),
	.w6(32'h3bddff4c),
	.w7(32'h3c3a0a47),
	.w8(32'hbc14ab60),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd35bb),
	.w1(32'hbb0e7de2),
	.w2(32'h3b226486),
	.w3(32'hbbe5a9dc),
	.w4(32'hbbe09a4e),
	.w5(32'hbad015f2),
	.w6(32'hbbdc4dd9),
	.w7(32'hbc046a27),
	.w8(32'hbb951a66),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe391f7),
	.w1(32'hbc87c226),
	.w2(32'hbc980203),
	.w3(32'h3b1de302),
	.w4(32'hbb230a3c),
	.w5(32'hbb09aa0d),
	.w6(32'hbb0999c2),
	.w7(32'hbb98a445),
	.w8(32'hba364e11),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b157c86),
	.w1(32'h3ac79982),
	.w2(32'hbb11a65f),
	.w3(32'h3bce6be6),
	.w4(32'h3ba91229),
	.w5(32'hbb2111a0),
	.w6(32'h3bed3a11),
	.w7(32'h3bd9af4b),
	.w8(32'h3b89082a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba45c49),
	.w1(32'h3c244682),
	.w2(32'h3c3b73d7),
	.w3(32'hbbaa5df4),
	.w4(32'hbb9b752b),
	.w5(32'hba1eb894),
	.w6(32'h3956a00f),
	.w7(32'hbb30d79f),
	.w8(32'h392580f8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c0036),
	.w1(32'h3b457f10),
	.w2(32'h3b4fe4f0),
	.w3(32'hbb3aa5d4),
	.w4(32'hbb13fda8),
	.w5(32'h39bab758),
	.w6(32'hbb3c78dd),
	.w7(32'hba9d76e7),
	.w8(32'h3afc7a98),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248d9d),
	.w1(32'hbc063b97),
	.w2(32'hbc743495),
	.w3(32'h3bc7d7a4),
	.w4(32'h3b92ec3c),
	.w5(32'hbba43848),
	.w6(32'h3be9cb52),
	.w7(32'h3b36716d),
	.w8(32'hbbc4e86f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f9e5a),
	.w1(32'hbbebefe7),
	.w2(32'hbc000a3f),
	.w3(32'h39f33ba4),
	.w4(32'h3b151c37),
	.w5(32'hbbd0ca1d),
	.w6(32'h3b63a143),
	.w7(32'h3bb03ebc),
	.w8(32'hbbb447f8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc072e13),
	.w1(32'hbb153311),
	.w2(32'h3a129c3d),
	.w3(32'hbc3e2270),
	.w4(32'h3b386fd4),
	.w5(32'h3c659f31),
	.w6(32'hbbc8dc46),
	.w7(32'hb7cd28ee),
	.w8(32'h3c4d3e01),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78821e),
	.w1(32'h3bd39c14),
	.w2(32'h3c0d9276),
	.w3(32'hba1ad77e),
	.w4(32'h3b9c6dc9),
	.w5(32'h3c1f35cb),
	.w6(32'h3b8afe19),
	.w7(32'h3bc5e378),
	.w8(32'h3c3212df),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6c1d6),
	.w1(32'h3ae58129),
	.w2(32'h3bee6a98),
	.w3(32'hbac1d69c),
	.w4(32'hbaf34cc6),
	.w5(32'h3b2f5f1e),
	.w6(32'hba9c0f43),
	.w7(32'hba9eb9f4),
	.w8(32'h3a7b8070),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13a7e8),
	.w1(32'h3a1dab75),
	.w2(32'hbc0a052c),
	.w3(32'hba154f71),
	.w4(32'h3c81c636),
	.w5(32'h3ba60110),
	.w6(32'h3bb19783),
	.w7(32'h3c758ba3),
	.w8(32'hb982ce76),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c8c2c),
	.w1(32'h3a81ea2d),
	.w2(32'h39ebf316),
	.w3(32'h3a421a7b),
	.w4(32'h3a8787af),
	.w5(32'h3b5fa6d6),
	.w6(32'h3a3abba5),
	.w7(32'h3aaefb8d),
	.w8(32'h3b5b35fd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66f332),
	.w1(32'hbc373993),
	.w2(32'hbb866e4f),
	.w3(32'hbc4516b5),
	.w4(32'hbb642bc8),
	.w5(32'h3b62a6d2),
	.w6(32'hbb717f36),
	.w7(32'h3ad10064),
	.w8(32'h3bb45324),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af35641),
	.w1(32'hbb185e9c),
	.w2(32'hbbbc2c0d),
	.w3(32'h3af324c8),
	.w4(32'hba851eab),
	.w5(32'h3ad4816a),
	.w6(32'h3a90e676),
	.w7(32'hba851150),
	.w8(32'hbb6c5d82),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c5d79),
	.w1(32'h3b8453d0),
	.w2(32'h3b893627),
	.w3(32'hbb752b82),
	.w4(32'h3b85500e),
	.w5(32'h3acca939),
	.w6(32'h3b424c85),
	.w7(32'h3bb53d29),
	.w8(32'h3b282345),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af206b8),
	.w1(32'h3b755907),
	.w2(32'hb9678b88),
	.w3(32'h3bf6aea3),
	.w4(32'h3a1a5119),
	.w5(32'hba605d22),
	.w6(32'h3bd2030a),
	.w7(32'h3aacae04),
	.w8(32'hbb49b8f7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb7052),
	.w1(32'hbb6140c3),
	.w2(32'hbbf4e98e),
	.w3(32'h3bb35149),
	.w4(32'h3b4d3bac),
	.w5(32'h3b056bd7),
	.w6(32'h3b2cc6be),
	.w7(32'h38dd702d),
	.w8(32'h3b39eba3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d2dee),
	.w1(32'h3b7f01aa),
	.w2(32'h3b8ab700),
	.w3(32'h3b809f81),
	.w4(32'h3ab23549),
	.w5(32'hbaead83d),
	.w6(32'h3b98cd22),
	.w7(32'hba896e21),
	.w8(32'hbb6fcc48),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a3c17),
	.w1(32'hbc113209),
	.w2(32'hbba9bb1e),
	.w3(32'hbb21d75a),
	.w4(32'hbc13199f),
	.w5(32'hbb58b537),
	.w6(32'hbb63cff9),
	.w7(32'hbc2e678b),
	.w8(32'hbb3e8153),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688b1e),
	.w1(32'hb9fd25f4),
	.w2(32'h3a5bc6df),
	.w3(32'hba77275b),
	.w4(32'hba4f23ab),
	.w5(32'hba6d6673),
	.w6(32'h3b1ea617),
	.w7(32'hbac43d07),
	.w8(32'hb9ba2ff9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a310b6f),
	.w1(32'h3c5e8c73),
	.w2(32'h3c435b30),
	.w3(32'hbb230ff8),
	.w4(32'h3c196ac1),
	.w5(32'h3a8fd00d),
	.w6(32'h3bf9220b),
	.w7(32'h3c24610b),
	.w8(32'h3bb89a00),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc729c),
	.w1(32'hbc255bc6),
	.w2(32'hbc09653c),
	.w3(32'hbacb9fe6),
	.w4(32'hbb69794a),
	.w5(32'hbbe84103),
	.w6(32'h39a2d743),
	.w7(32'h3b2b5dcb),
	.w8(32'hbba6c69a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf1092),
	.w1(32'hbb40a19f),
	.w2(32'hbb4f616b),
	.w3(32'h3b72505f),
	.w4(32'hba889466),
	.w5(32'h3a0a41a2),
	.w6(32'h3b4a142a),
	.w7(32'hbababc4e),
	.w8(32'h389f2ebb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba972d23),
	.w1(32'hbac5e2d2),
	.w2(32'hba2a39ca),
	.w3(32'hbb1b4bee),
	.w4(32'hbaf3b458),
	.w5(32'h3b4bea2a),
	.w6(32'hba535b0d),
	.w7(32'hb987c5a2),
	.w8(32'h3a00d242),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a503a82),
	.w1(32'hbb860158),
	.w2(32'hbaf98ec3),
	.w3(32'hba940764),
	.w4(32'hbb18fc7e),
	.w5(32'hbae997af),
	.w6(32'hbb9140f0),
	.w7(32'hba71061c),
	.w8(32'h3b027613),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b621e6d),
	.w1(32'h38864b1a),
	.w2(32'hb8ba48b5),
	.w3(32'h3a284f67),
	.w4(32'hbaf7f74f),
	.w5(32'hbb076722),
	.w6(32'h3990cc26),
	.w7(32'hbb8b4454),
	.w8(32'hba00f892),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e8160),
	.w1(32'h3934283d),
	.w2(32'h3abed37b),
	.w3(32'hba9a8f8c),
	.w4(32'h3b0d14b2),
	.w5(32'h38616917),
	.w6(32'h3a939351),
	.w7(32'h3b36b26a),
	.w8(32'h38046518),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba009819),
	.w1(32'hb987f04b),
	.w2(32'hbba90726),
	.w3(32'hbaf31d1b),
	.w4(32'hbb181b22),
	.w5(32'h3bc1754b),
	.w6(32'hba8876d6),
	.w7(32'hbacd6c79),
	.w8(32'h3b98cada),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b3d1f),
	.w1(32'hba685f5d),
	.w2(32'hbb634b0c),
	.w3(32'h3b68fe75),
	.w4(32'h3af03f2f),
	.w5(32'h3a588720),
	.w6(32'h3b198e45),
	.w7(32'hba43e6fb),
	.w8(32'hbabe3ce2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0059fb),
	.w1(32'hbb81539f),
	.w2(32'hbb896c85),
	.w3(32'hbb832aa9),
	.w4(32'h3bd52ccc),
	.w5(32'hbb6b5346),
	.w6(32'hbb356bef),
	.w7(32'h3b825905),
	.w8(32'hbbb08f36),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadac9a),
	.w1(32'h3b147b06),
	.w2(32'h3c4d2aa1),
	.w3(32'hbb218c08),
	.w4(32'hbb923372),
	.w5(32'hba99d6ef),
	.w6(32'hbb9e520e),
	.w7(32'hbb73235c),
	.w8(32'h3a20ddff),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34e0b0),
	.w1(32'hba5b8f02),
	.w2(32'hb944daba),
	.w3(32'hba4fb073),
	.w4(32'h3afc842d),
	.w5(32'hbaa63765),
	.w6(32'hba5efa93),
	.w7(32'h3ae5c97b),
	.w8(32'hbb4f0848),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b469),
	.w1(32'hbb256841),
	.w2(32'h37e2d8e8),
	.w3(32'hbb0dcace),
	.w4(32'hbb638a07),
	.w5(32'h3b40c986),
	.w6(32'hbb5dc74b),
	.w7(32'hbb7f948a),
	.w8(32'h3b8752fe),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89e1b1),
	.w1(32'hbacebd6c),
	.w2(32'hbaf9654d),
	.w3(32'h3ad81900),
	.w4(32'hbb2085c1),
	.w5(32'h3ac38675),
	.w6(32'hba0dd2a0),
	.w7(32'hbb0dc8d8),
	.w8(32'h3b2d7864),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2842fd),
	.w1(32'h3a463aa7),
	.w2(32'hba0ec504),
	.w3(32'h3b520c5a),
	.w4(32'hbafcb319),
	.w5(32'h3b083ec8),
	.w6(32'h3b559d3d),
	.w7(32'hba924349),
	.w8(32'hba30c6dd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56a94b),
	.w1(32'h39393d80),
	.w2(32'hbbab6a36),
	.w3(32'hbb4eec14),
	.w4(32'hbac61a35),
	.w5(32'hbba56725),
	.w6(32'h3bdae07e),
	.w7(32'hb963f41c),
	.w8(32'hbb3c196e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6e754),
	.w1(32'hbb753802),
	.w2(32'hbc84960d),
	.w3(32'h3b7689e5),
	.w4(32'hb905b3eb),
	.w5(32'hbc05b02f),
	.w6(32'h3be3e954),
	.w7(32'hbb2a91dd),
	.w8(32'hbc00b114),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b26760),
	.w1(32'hbb22f229),
	.w2(32'hbba335a7),
	.w3(32'hbaf3f4d9),
	.w4(32'hbb8db726),
	.w5(32'h39fc8651),
	.w6(32'hbaa859a8),
	.w7(32'hbb1755e8),
	.w8(32'h3aa10f25),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b0927),
	.w1(32'h3b44582c),
	.w2(32'hbb9d1c00),
	.w3(32'hbb5bc292),
	.w4(32'hbb6aff9b),
	.w5(32'hba039dc8),
	.w6(32'hba1e49bf),
	.w7(32'hbb0fa8bd),
	.w8(32'h3a33e0ed),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ed4c),
	.w1(32'h3a8e5ea8),
	.w2(32'h3907b46d),
	.w3(32'hbad9d72f),
	.w4(32'hbb1b419f),
	.w5(32'hb9865e29),
	.w6(32'hbaaf6310),
	.w7(32'hbb0c433e),
	.w8(32'h3b5217fa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04fb93),
	.w1(32'hbbcdab62),
	.w2(32'hbba44c46),
	.w3(32'h3ab9c182),
	.w4(32'hbbbd4a90),
	.w5(32'h3ab4623a),
	.w6(32'h3a943cea),
	.w7(32'hbb1387e7),
	.w8(32'h3b47c40d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d1bf0),
	.w1(32'hbaf0cffe),
	.w2(32'hbaf793c2),
	.w3(32'h3ac4b5d8),
	.w4(32'hbbac0a5b),
	.w5(32'h3992b3ce),
	.w6(32'h3b4ed45e),
	.w7(32'hba9abeb9),
	.w8(32'hbb8583f2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c8a0f),
	.w1(32'hbc36a572),
	.w2(32'hbc9aff60),
	.w3(32'hba8080eb),
	.w4(32'h3ab2564c),
	.w5(32'hbb9debd5),
	.w6(32'hba485366),
	.w7(32'hba9b5ec3),
	.w8(32'hbbbd6d5a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc824e),
	.w1(32'h3c623b4a),
	.w2(32'h3c1c72a5),
	.w3(32'h3a8a1e20),
	.w4(32'h3b7bdc8d),
	.w5(32'h3b1f03b2),
	.w6(32'h3c0c233d),
	.w7(32'h3b4bf1b9),
	.w8(32'h3b44b6f0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8cd89),
	.w1(32'hbb76b9d7),
	.w2(32'hbbd8a814),
	.w3(32'h3a5a83df),
	.w4(32'h3a69f65f),
	.w5(32'h3b1a251d),
	.w6(32'h3b8bafab),
	.w7(32'h3a94316e),
	.w8(32'h3ad252d8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef7109),
	.w1(32'hba13864f),
	.w2(32'hbc390680),
	.w3(32'h3bad4c75),
	.w4(32'h3ba3d40e),
	.w5(32'hbb66cee0),
	.w6(32'h3c2c18e8),
	.w7(32'h3bea3bbf),
	.w8(32'hbba4d029),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb039fbd),
	.w1(32'h3b5f60fc),
	.w2(32'h3a9ba791),
	.w3(32'hbac3e5e7),
	.w4(32'hbab4e2ef),
	.w5(32'h3af58ad9),
	.w6(32'hb9c11808),
	.w7(32'hbb3a97a9),
	.w8(32'h3bb5fd4f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f297d9),
	.w1(32'hba3945ee),
	.w2(32'hbbc66a22),
	.w3(32'h39a9924c),
	.w4(32'h3bc7097e),
	.w5(32'hbc4e7581),
	.w6(32'h3bc632c1),
	.w7(32'h3b63d935),
	.w8(32'hbbf5b329),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8009b5),
	.w1(32'h3bb7c6b1),
	.w2(32'h3ad083b2),
	.w3(32'h3b00ade1),
	.w4(32'h3be3df89),
	.w5(32'hbb71640c),
	.w6(32'h3b655a2b),
	.w7(32'h3ba7920b),
	.w8(32'h3a028d2b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c98bd),
	.w1(32'hbb1dda67),
	.w2(32'h3c033402),
	.w3(32'h3b83f7a6),
	.w4(32'hbbc5c10a),
	.w5(32'hbb4f4396),
	.w6(32'h3be93652),
	.w7(32'hbba94c55),
	.w8(32'hbbd836ab),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb872bfc),
	.w1(32'hbab72d30),
	.w2(32'hbaf3c096),
	.w3(32'hbad7d151),
	.w4(32'hbb248854),
	.w5(32'hbc00d7f5),
	.w6(32'hbb28fc8f),
	.w7(32'hbb70061a),
	.w8(32'hbb815ee7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f68d5),
	.w1(32'h3b4d7c10),
	.w2(32'hbbc3aed5),
	.w3(32'h3aecb05e),
	.w4(32'hbb485d66),
	.w5(32'h3ab55da6),
	.w6(32'h3b87d576),
	.w7(32'hbbc8b984),
	.w8(32'h3b7a408d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af63076),
	.w1(32'h3b6754c0),
	.w2(32'h3a5cab10),
	.w3(32'h3bb2347a),
	.w4(32'h3ac68866),
	.w5(32'h3b4e5bab),
	.w6(32'h3bb768dc),
	.w7(32'hb8a43f14),
	.w8(32'h3a46ce97),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b730060),
	.w1(32'h38ed455b),
	.w2(32'hb9bc2489),
	.w3(32'h3afe69d6),
	.w4(32'hbaa88d8d),
	.w5(32'h3a06327e),
	.w6(32'h39ad1904),
	.w7(32'hba67f910),
	.w8(32'h39c03c97),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf1ff3),
	.w1(32'h3b686ee4),
	.w2(32'h3b1d2604),
	.w3(32'hbb10d0eb),
	.w4(32'hbb09aaab),
	.w5(32'h3bb6e523),
	.w6(32'hbbc294d9),
	.w7(32'hbb7b0192),
	.w8(32'h3ba2b569),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5fedf),
	.w1(32'hbbe31bbc),
	.w2(32'hbac1a9e1),
	.w3(32'h3b1913c1),
	.w4(32'h3a73ee5f),
	.w5(32'hbbfaeb8d),
	.w6(32'h3bafafbe),
	.w7(32'h3a78794e),
	.w8(32'hbb9ebaa3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e84a),
	.w1(32'h3bb9535b),
	.w2(32'hbb7b0c28),
	.w3(32'h3b181c09),
	.w4(32'h3a0072b1),
	.w5(32'h3ab90c45),
	.w6(32'h3bbcc79f),
	.w7(32'hbb0d4878),
	.w8(32'hbab6dd1e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec738),
	.w1(32'hbc001198),
	.w2(32'hbbdeb893),
	.w3(32'h3adeb2d3),
	.w4(32'h3ae9502d),
	.w5(32'hbb773aa9),
	.w6(32'hba20b7f9),
	.w7(32'h39336a86),
	.w8(32'hbb4d5ea5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641f89),
	.w1(32'h3b3ff16a),
	.w2(32'h3b83c822),
	.w3(32'h3a80d2ea),
	.w4(32'h3b8196e9),
	.w5(32'hbc0d17bd),
	.w6(32'h3b7fe257),
	.w7(32'h3b93727a),
	.w8(32'hbb32f2f2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65c8de),
	.w1(32'hba95925f),
	.w2(32'hbc7ba6d5),
	.w3(32'h3cad3763),
	.w4(32'h3a459e7a),
	.w5(32'hbb810a0a),
	.w6(32'h3c72cbce),
	.w7(32'hbb5ee11c),
	.w8(32'h393b96b1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03ee90),
	.w1(32'hbbea54ed),
	.w2(32'h3b841f70),
	.w3(32'h3ac57e0f),
	.w4(32'hbba96d5e),
	.w5(32'hbb89155c),
	.w6(32'hbbea7ba1),
	.w7(32'hbb9d2d3a),
	.w8(32'hbbf91108),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0262a),
	.w1(32'hb79986b3),
	.w2(32'h3a467097),
	.w3(32'hb97279d4),
	.w4(32'hbb554d2d),
	.w5(32'h3b427695),
	.w6(32'hbaa4db20),
	.w7(32'hbb6065bb),
	.w8(32'h3a8d4925),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80f6c9),
	.w1(32'hb9e7a18c),
	.w2(32'h3b56a327),
	.w3(32'hba690e3f),
	.w4(32'h3aa7920d),
	.w5(32'h3b9feeb9),
	.w6(32'hba14aad4),
	.w7(32'h3a9a723b),
	.w8(32'h3c096293),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b207a9c),
	.w1(32'hb9ffb62b),
	.w2(32'hbb03ff88),
	.w3(32'h3b3c6f64),
	.w4(32'hba423d19),
	.w5(32'h3af6516d),
	.w6(32'h3b0d7567),
	.w7(32'hbaef2903),
	.w8(32'h3b7af323),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a964c3b),
	.w1(32'hbb101fab),
	.w2(32'h3b44762d),
	.w3(32'hba50713d),
	.w4(32'hba7f73c2),
	.w5(32'hbb7d5e06),
	.w6(32'h3b2f8eec),
	.w7(32'h3af012bc),
	.w8(32'hbb58c7df),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb672d46),
	.w1(32'h3b833938),
	.w2(32'h3bdd1228),
	.w3(32'hbb8e7bac),
	.w4(32'h3baaca08),
	.w5(32'h3b9d5fb3),
	.w6(32'hb922c6b5),
	.w7(32'h3bb32fb1),
	.w8(32'h3bb3a111),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45a70e),
	.w1(32'hbb304af8),
	.w2(32'hbafd62ca),
	.w3(32'h3ba9a43d),
	.w4(32'hbbdf0615),
	.w5(32'hb5dfec92),
	.w6(32'h3b525621),
	.w7(32'hbbc43043),
	.w8(32'hba024ff9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff3f40),
	.w1(32'hbb25461f),
	.w2(32'hbb5b3135),
	.w3(32'h3b37617b),
	.w4(32'hbb311f97),
	.w5(32'h3b788489),
	.w6(32'h3a5b1f19),
	.w7(32'h3a2748dd),
	.w8(32'h3b40aa94),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb54d31),
	.w1(32'hbc14d2d8),
	.w2(32'hbbef2c33),
	.w3(32'hbbbc12f7),
	.w4(32'hbb8ea742),
	.w5(32'h3a1e32eb),
	.w6(32'hba3db6c8),
	.w7(32'hba89fd63),
	.w8(32'hb8b5f6bd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba09b72),
	.w1(32'hb7e37a44),
	.w2(32'hbb37e1f3),
	.w3(32'h3ba6890e),
	.w4(32'h39f6693f),
	.w5(32'h382260a5),
	.w6(32'h3b5f385a),
	.w7(32'hbaee0fd5),
	.w8(32'h3b500968),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd14cf),
	.w1(32'h3b4130d0),
	.w2(32'h3a3ce7d0),
	.w3(32'hbb5b120a),
	.w4(32'hbab9b887),
	.w5(32'hbbd929db),
	.w6(32'hba1a49d0),
	.w7(32'hba4224f4),
	.w8(32'hbb1efc86),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b97a4),
	.w1(32'h3a88757c),
	.w2(32'hbad0668f),
	.w3(32'h3b66ca8b),
	.w4(32'h39e77161),
	.w5(32'h3b24ad2d),
	.w6(32'h3b7adcb7),
	.w7(32'hbb412003),
	.w8(32'h3bb5cae6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c556035),
	.w1(32'h3b48df5f),
	.w2(32'hba6bec7a),
	.w3(32'h3b308352),
	.w4(32'hba9d91dd),
	.w5(32'h3b7c9a14),
	.w6(32'h3b54ac69),
	.w7(32'hbbe6b4f6),
	.w8(32'hba251890),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e833b),
	.w1(32'hbafb4fca),
	.w2(32'hbb1c3300),
	.w3(32'hba47f93a),
	.w4(32'hbb628fec),
	.w5(32'h3b8c8a61),
	.w6(32'hb9aa0040),
	.w7(32'hbb4df819),
	.w8(32'h3ab09aaf),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8731ca),
	.w1(32'hba009687),
	.w2(32'hba94230a),
	.w3(32'h3b464cc4),
	.w4(32'hb905120c),
	.w5(32'h3b2ec6ef),
	.w6(32'hbab1536c),
	.w7(32'hbba9f63b),
	.w8(32'h3a4657bb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06c543),
	.w1(32'h3b8c5ebc),
	.w2(32'h3a735dbc),
	.w3(32'h3b8191d4),
	.w4(32'h3bda4936),
	.w5(32'hbab185d9),
	.w6(32'h3b9ae16e),
	.w7(32'h3b90f1dc),
	.w8(32'hbb4f31ba),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b396b4d),
	.w1(32'h3b815e4d),
	.w2(32'hbb9101f8),
	.w3(32'hbae3ffde),
	.w4(32'h3be2366c),
	.w5(32'h3a667d97),
	.w6(32'h3b5783f7),
	.w7(32'h3bd825a3),
	.w8(32'hb96e85d6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b999300),
	.w1(32'h3b96c2c3),
	.w2(32'h392eaea5),
	.w3(32'h3b19f059),
	.w4(32'h3a612fde),
	.w5(32'h3babc9d0),
	.w6(32'h3b680bab),
	.w7(32'h3835c309),
	.w8(32'h3b75090e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c5a69),
	.w1(32'h3b3bc5d9),
	.w2(32'h3bb5e69d),
	.w3(32'hba56d112),
	.w4(32'hba607487),
	.w5(32'h3a07712b),
	.w6(32'h3a8bfdf4),
	.w7(32'h3ad0c25e),
	.w8(32'hba479f6c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95e901),
	.w1(32'hbb07f3b5),
	.w2(32'hba8c6a75),
	.w3(32'hb8757e66),
	.w4(32'hbb8e8b58),
	.w5(32'hb9944c11),
	.w6(32'hbb0e5034),
	.w7(32'hbb1edd4c),
	.w8(32'h3aabc387),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2437ac),
	.w1(32'hbbd0404d),
	.w2(32'hbc1bbe8f),
	.w3(32'hba66aab0),
	.w4(32'hb95c1b52),
	.w5(32'hbbafa470),
	.w6(32'hbb1dc728),
	.w7(32'hba9d7cf9),
	.w8(32'hbbac42bf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a676e4d),
	.w1(32'hba9a33a7),
	.w2(32'hbba1f60d),
	.w3(32'h3c15d57b),
	.w4(32'h3b33d941),
	.w5(32'hbabd1bc6),
	.w6(32'h3bd7d959),
	.w7(32'h3ad1e476),
	.w8(32'hbabb7146),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c8f1b),
	.w1(32'hbc1e381c),
	.w2(32'hbc67442b),
	.w3(32'h3b019f48),
	.w4(32'hbb02e5c2),
	.w5(32'hbbdd3146),
	.w6(32'h3a5be02b),
	.w7(32'hbaed3134),
	.w8(32'hbb8c6b01),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d336c8),
	.w1(32'h3a776431),
	.w2(32'h3b88c085),
	.w3(32'h3958a442),
	.w4(32'h3b0b4a89),
	.w5(32'hbacbb86d),
	.w6(32'h3a946b8e),
	.w7(32'h3b59163c),
	.w8(32'h3a895b17),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa937a),
	.w1(32'h3b66103d),
	.w2(32'hbb6213f0),
	.w3(32'h3bb12bcb),
	.w4(32'h3ae40ea7),
	.w5(32'hba924fe1),
	.w6(32'h3bfebd94),
	.w7(32'h3b00fcd5),
	.w8(32'hbb5159f1),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0c3fe),
	.w1(32'hbb558934),
	.w2(32'hb7bc776d),
	.w3(32'hbb9c079a),
	.w4(32'hba431b68),
	.w5(32'h3ae3eba0),
	.w6(32'hbb8895f8),
	.w7(32'hb841cdd5),
	.w8(32'h3b65b157),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1c39c),
	.w1(32'hbbcd83ea),
	.w2(32'h3b056853),
	.w3(32'hb889e7ea),
	.w4(32'hbaa93641),
	.w5(32'h3ac6e249),
	.w6(32'hbb8acc9d),
	.w7(32'h3a12c19f),
	.w8(32'h3aa1e23d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bace87b),
	.w1(32'h3a1ca782),
	.w2(32'h3973cc32),
	.w3(32'h3b1a1d03),
	.w4(32'hb99034b6),
	.w5(32'hb9e647ad),
	.w6(32'hb9927571),
	.w7(32'hbb3c7d66),
	.w8(32'hba4748fa),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8518f1),
	.w1(32'hbb88191c),
	.w2(32'hbbcda857),
	.w3(32'h3aeaadb0),
	.w4(32'hbab1021d),
	.w5(32'hbba5d0e4),
	.w6(32'h3a85f340),
	.w7(32'hbb20aaa4),
	.w8(32'hb8f042e0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae88eba),
	.w1(32'h3b996bd6),
	.w2(32'h3c153d21),
	.w3(32'hbb30d882),
	.w4(32'h3c6a9dba),
	.w5(32'hb9376daa),
	.w6(32'h3b1d478c),
	.w7(32'h3c3d6cc2),
	.w8(32'h391015e8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb017b93),
	.w1(32'hbb62e662),
	.w2(32'hb9583911),
	.w3(32'hb9932425),
	.w4(32'hbaba1f7e),
	.w5(32'hbb8ed1eb),
	.w6(32'h39c6d6e4),
	.w7(32'hba44a3c6),
	.w8(32'hba48bf3a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56a523),
	.w1(32'hbb049981),
	.w2(32'hba42f660),
	.w3(32'hbac3b346),
	.w4(32'hbb1ae830),
	.w5(32'hbba12981),
	.w6(32'hbaca8ef7),
	.w7(32'hbab6b85c),
	.w8(32'hbb3eef38),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6478bc),
	.w1(32'hba708299),
	.w2(32'hbbe374da),
	.w3(32'h3a20838b),
	.w4(32'h3bdd2f3c),
	.w5(32'h3b6d0840),
	.w6(32'h3b39bdf6),
	.w7(32'h3bcb8f60),
	.w8(32'hba8d10dc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39333a89),
	.w1(32'h3b8db097),
	.w2(32'h3bcf1d64),
	.w3(32'hbbf51b24),
	.w4(32'h3c0f13c5),
	.w5(32'h3be3a540),
	.w6(32'h390f1480),
	.w7(32'h3c13ca14),
	.w8(32'h3ba01780),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc2d16),
	.w1(32'hbbbacadb),
	.w2(32'hbb1c04db),
	.w3(32'hbbbd86f7),
	.w4(32'hbb2e5771),
	.w5(32'h3a9ab5ac),
	.w6(32'hbbc449ab),
	.w7(32'hbafba064),
	.w8(32'h3b49d621),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13eed2),
	.w1(32'hbc8a687f),
	.w2(32'hbc71d4bb),
	.w3(32'h3b817b99),
	.w4(32'hbb765a6e),
	.w5(32'hbbda7931),
	.w6(32'hba31caf7),
	.w7(32'hb9810e55),
	.w8(32'hbc276742),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb2031),
	.w1(32'hbbc32fb3),
	.w2(32'h35d4e070),
	.w3(32'h3bdf73b9),
	.w4(32'hbaf4629b),
	.w5(32'hbc065dce),
	.w6(32'h3b468de6),
	.w7(32'hbb98b677),
	.w8(32'hbb5a9059),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ed0a7),
	.w1(32'hba9ae286),
	.w2(32'hbb865761),
	.w3(32'h3a9ce04b),
	.w4(32'hbb38f9ca),
	.w5(32'h3ae07b99),
	.w6(32'h3b38ed33),
	.w7(32'hbb94a6d1),
	.w8(32'h3b9c3a10),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dd547),
	.w1(32'h3a168c22),
	.w2(32'hbaa86972),
	.w3(32'h3b06cb6f),
	.w4(32'hbb17d13e),
	.w5(32'hbaadff78),
	.w6(32'h3a31cd45),
	.w7(32'hbb015421),
	.w8(32'h3af2dd04),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991697d),
	.w1(32'h3b8cb3f9),
	.w2(32'h384d4749),
	.w3(32'hb854f2c4),
	.w4(32'h3b3dc91a),
	.w5(32'h3ad91246),
	.w6(32'h3b805102),
	.w7(32'h3b30330a),
	.w8(32'h3ba20e42),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b596ddf),
	.w1(32'h3a0902bb),
	.w2(32'hbacd6b6c),
	.w3(32'hbb40e546),
	.w4(32'hbb22a311),
	.w5(32'h38d7c2a4),
	.w6(32'h3a909678),
	.w7(32'hba72cabc),
	.w8(32'h3ab0f5da),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b671c74),
	.w1(32'h3b25d3a5),
	.w2(32'hb9720f28),
	.w3(32'hbabb570d),
	.w4(32'hbad33c1c),
	.w5(32'hbb77bd17),
	.w6(32'h3b16ed3a),
	.w7(32'hba117065),
	.w8(32'hbb9772f8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dd3d7),
	.w1(32'h3c32d259),
	.w2(32'h3b4e0ef8),
	.w3(32'h39e90be6),
	.w4(32'h3be985b2),
	.w5(32'hbaac6cf6),
	.w6(32'h3c1ee736),
	.w7(32'h3b7b1193),
	.w8(32'h3ad6322f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a920a7b),
	.w1(32'h3c512ce4),
	.w2(32'h3ca5c584),
	.w3(32'h3b8e9c9e),
	.w4(32'h3c39c7d0),
	.w5(32'h3b8ce0d1),
	.w6(32'h3ba68e4e),
	.w7(32'h3c0dfae9),
	.w8(32'hb9925eee),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b234874),
	.w1(32'hbb2ed00c),
	.w2(32'hba49d793),
	.w3(32'hbb6a6083),
	.w4(32'hbb45f24a),
	.w5(32'h3a60b69f),
	.w6(32'hbb239bb4),
	.w7(32'hba70a755),
	.w8(32'h3912f23f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a7627),
	.w1(32'hbaa91bf1),
	.w2(32'hbbf3d476),
	.w3(32'h3a020736),
	.w4(32'h3b806f88),
	.w5(32'hbabe4c49),
	.w6(32'h3b88c66e),
	.w7(32'h3b0edbb2),
	.w8(32'hbb4a9017),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56202c),
	.w1(32'h3a8b255c),
	.w2(32'h39a7183e),
	.w3(32'hbb0186b7),
	.w4(32'h3a4c8a97),
	.w5(32'h395e3399),
	.w6(32'hbafbaf25),
	.w7(32'h3a09de2d),
	.w8(32'hb96c46b8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeed9a),
	.w1(32'h3ca10819),
	.w2(32'h3b0995c0),
	.w3(32'h3c37d9af),
	.w4(32'h3c4e1bc7),
	.w5(32'h3b49c1c2),
	.w6(32'h3ca0cfa1),
	.w7(32'h3b30b606),
	.w8(32'h3bce1c91),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0408ec),
	.w1(32'hbb8eb1d0),
	.w2(32'hbad82b02),
	.w3(32'hbac9508f),
	.w4(32'hbba12a73),
	.w5(32'h3ab808bf),
	.w6(32'h3a3e2649),
	.w7(32'hbbaea9e8),
	.w8(32'h3bb9ecc7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93269a),
	.w1(32'hb9966efb),
	.w2(32'hb8d723cf),
	.w3(32'hbb421a5b),
	.w4(32'h3b341386),
	.w5(32'h3b71beb9),
	.w6(32'hbaebb0a9),
	.w7(32'hba058bb7),
	.w8(32'h3b2a28f4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27c806),
	.w1(32'h3be1e539),
	.w2(32'h3a27b7ce),
	.w3(32'h3acee624),
	.w4(32'h3bc5dbd3),
	.w5(32'hbb9d2fdc),
	.w6(32'h3bd757f8),
	.w7(32'h3b44dbb8),
	.w8(32'hbb62787f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5b671),
	.w1(32'h3b29e6a4),
	.w2(32'h3b9767f9),
	.w3(32'h3b586508),
	.w4(32'hbab3f3a5),
	.w5(32'h3ab0029d),
	.w6(32'hb982bf4c),
	.w7(32'hbb363f97),
	.w8(32'hbb19780d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf33ccd),
	.w1(32'h3b2fa60e),
	.w2(32'h3b3cea06),
	.w3(32'hbab4bbe0),
	.w4(32'h3a7a9da9),
	.w5(32'h3aabc374),
	.w6(32'h3a1b3241),
	.w7(32'h3ac30d97),
	.w8(32'h3a352980),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0aed1),
	.w1(32'hb9960b95),
	.w2(32'hba771216),
	.w3(32'h3b26bbab),
	.w4(32'hbae66f1d),
	.w5(32'hba803262),
	.w6(32'hb97f1b50),
	.w7(32'hbb6325c6),
	.w8(32'hbaea6e3d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6abde2),
	.w1(32'h3b99b83e),
	.w2(32'h3bac0a32),
	.w3(32'hbb2a7d28),
	.w4(32'h3ac13026),
	.w5(32'h3a4577ce),
	.w6(32'h3b6b2cf9),
	.w7(32'h3a86f92c),
	.w8(32'h3b8bf178),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fb684),
	.w1(32'h3b461aa8),
	.w2(32'hbb5148e6),
	.w3(32'h3b958e7e),
	.w4(32'h3b0ba5f3),
	.w5(32'hbbb695ce),
	.w6(32'h3c2fb0a4),
	.w7(32'h3a82dccf),
	.w8(32'hbbde71c1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a94bf),
	.w1(32'hb9da8eb4),
	.w2(32'h3b6a9d32),
	.w3(32'h3ac4cd1f),
	.w4(32'h3bbf4ad1),
	.w5(32'hba7e268d),
	.w6(32'h3be0d7e9),
	.w7(32'h3be6ce2f),
	.w8(32'hbb2491c1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b65411),
	.w1(32'h3a486f43),
	.w2(32'hb9331848),
	.w3(32'hba36824e),
	.w4(32'hb9cbc6e8),
	.w5(32'hb998eb2d),
	.w6(32'hb96ae858),
	.w7(32'hb83c42f9),
	.w8(32'hbb179cc0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba975462),
	.w1(32'hbaeef329),
	.w2(32'hbaa3c47d),
	.w3(32'hbbb2d0b4),
	.w4(32'hbb85b555),
	.w5(32'hbaff4fc9),
	.w6(32'hbb927dbc),
	.w7(32'h38f88641),
	.w8(32'h39ac76fa),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe4a01),
	.w1(32'h3c2dbcd9),
	.w2(32'h3c24dcc4),
	.w3(32'h3c0f55ec),
	.w4(32'h3c581358),
	.w5(32'hba17d078),
	.w6(32'h3c7741ec),
	.w7(32'h3c39eb20),
	.w8(32'h3bb94022),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7f3e5),
	.w1(32'h3a638bc3),
	.w2(32'hbba97764),
	.w3(32'h398f123f),
	.w4(32'h3bbb3924),
	.w5(32'hbb4fe69a),
	.w6(32'hb9cb4897),
	.w7(32'h3ba7ae79),
	.w8(32'hbb7d96da),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8df3b),
	.w1(32'h3adc4551),
	.w2(32'h3b81da30),
	.w3(32'h3bfc36f7),
	.w4(32'hbb2fb78a),
	.w5(32'h3b289cd3),
	.w6(32'h3b215813),
	.w7(32'h371600c2),
	.w8(32'h3af0a369),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c243835),
	.w1(32'h3995079a),
	.w2(32'hbc05fd84),
	.w3(32'hbb338d78),
	.w4(32'h3b838218),
	.w5(32'h3b8acc13),
	.w6(32'h3bb92921),
	.w7(32'h3b9d8d1c),
	.w8(32'h3b2d7381),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a979b68),
	.w1(32'hba77b28e),
	.w2(32'hba067260),
	.w3(32'h3b15d25d),
	.w4(32'hbac2fff6),
	.w5(32'h3aa3d399),
	.w6(32'h3a2c2f8b),
	.w7(32'hbb3ea8a6),
	.w8(32'h38d30151),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4f743),
	.w1(32'hbb8c0d73),
	.w2(32'hbb70f8df),
	.w3(32'hba8ef75e),
	.w4(32'hbbaf4ce0),
	.w5(32'hbc2a10a8),
	.w6(32'h3983f8de),
	.w7(32'hbb5e95a0),
	.w8(32'hbc1a9134),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe946b),
	.w1(32'h3c359205),
	.w2(32'hbbbfb5bd),
	.w3(32'hbc3af3a8),
	.w4(32'h3be717a6),
	.w5(32'hba235dc2),
	.w6(32'h3b170e5a),
	.w7(32'h3c0afa5b),
	.w8(32'h3abc4516),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdc6d0),
	.w1(32'hbc428436),
	.w2(32'hbc52a2bd),
	.w3(32'h3ba6a50d),
	.w4(32'hbba961c8),
	.w5(32'hbc0c00a6),
	.w6(32'h3b36722b),
	.w7(32'hbbc02ad3),
	.w8(32'hbc1d3738),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee518b),
	.w1(32'hbab7770f),
	.w2(32'h3a378432),
	.w3(32'hb9ca95b0),
	.w4(32'h3c1597ba),
	.w5(32'h3ba1e426),
	.w6(32'h39c6cedd),
	.w7(32'h3c4767a7),
	.w8(32'h3b4d2b66),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20702e),
	.w1(32'hba9f87c9),
	.w2(32'h37ba318c),
	.w3(32'hbbc504a3),
	.w4(32'hbbb20ad2),
	.w5(32'h3b863c14),
	.w6(32'hbc0437f7),
	.w7(32'hbbb9ffc5),
	.w8(32'h3ba1d9d5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92c130),
	.w1(32'hbb8ada9d),
	.w2(32'h3bf97c5a),
	.w3(32'hbb9a79d8),
	.w4(32'hbb149402),
	.w5(32'h3b438062),
	.w6(32'hbb962d64),
	.w7(32'hb8c791f5),
	.w8(32'h3a40870d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9819723),
	.w1(32'h3b79fcb3),
	.w2(32'hbb3caf38),
	.w3(32'h3acbc828),
	.w4(32'hb9853179),
	.w5(32'h3bbc3b1e),
	.w6(32'h3b83700b),
	.w7(32'hbb190f8e),
	.w8(32'h3b5172f2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a73875),
	.w1(32'hb9ba5523),
	.w2(32'hb99a1ce9),
	.w3(32'h38c9eb16),
	.w4(32'hbae8d9ee),
	.w5(32'h3a41fcef),
	.w6(32'hbb0751fd),
	.w7(32'h3a5bbe76),
	.w8(32'h3ae749c7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54ee7),
	.w1(32'hbb21c7f5),
	.w2(32'hb9cf079b),
	.w3(32'hb9f7ed33),
	.w4(32'hbb872667),
	.w5(32'h3af7f9c0),
	.w6(32'hb98b0665),
	.w7(32'hbb3961ad),
	.w8(32'h3b3f9c46),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9de75),
	.w1(32'hbb89ef4e),
	.w2(32'hbb73409d),
	.w3(32'h3a91e95d),
	.w4(32'hbc0158cd),
	.w5(32'h3b1d731a),
	.w6(32'hbb00f73f),
	.w7(32'hbb86d3e9),
	.w8(32'h3b0c0c4e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2efd9),
	.w1(32'h3abc9c79),
	.w2(32'hba9b1d8e),
	.w3(32'h3a42d079),
	.w4(32'hba8101e1),
	.w5(32'hbbab24b2),
	.w6(32'h3b143509),
	.w7(32'hb9c8f38e),
	.w8(32'hbb497368),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac21f9e),
	.w1(32'hbb4c41d9),
	.w2(32'hbbec1f50),
	.w3(32'h3b1ce4e4),
	.w4(32'h3b4f49f5),
	.w5(32'hbae54d5b),
	.w6(32'h3b08f1a1),
	.w7(32'h3af58c54),
	.w8(32'hbae78ffa),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881114),
	.w1(32'h3b2b174e),
	.w2(32'h3aa532b6),
	.w3(32'h3a9fed30),
	.w4(32'h3ac957ab),
	.w5(32'h3a0ac433),
	.w6(32'h3b37017f),
	.w7(32'hba5489b4),
	.w8(32'hbb17d86f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7b359),
	.w1(32'h3ae8bcec),
	.w2(32'h3b30e0b2),
	.w3(32'hb98c23c4),
	.w4(32'h3a994f53),
	.w5(32'h3ac6151a),
	.w6(32'hbad75cbe),
	.w7(32'h38508c69),
	.w8(32'h3abe730c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bd2ea),
	.w1(32'hba86963b),
	.w2(32'hbc158cf3),
	.w3(32'h3954a876),
	.w4(32'h3c02e7eb),
	.w5(32'h3bae69ed),
	.w6(32'h3b41d3b6),
	.w7(32'h3c0370a8),
	.w8(32'h3b11cdab),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83d17c),
	.w1(32'h3a3c8315),
	.w2(32'hb9ff1d26),
	.w3(32'h3b6e45bb),
	.w4(32'h3acaf77f),
	.w5(32'hb97abada),
	.w6(32'h3b8cddb0),
	.w7(32'h3b062d54),
	.w8(32'hbb0ddd91),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eade0),
	.w1(32'h3b2a1564),
	.w2(32'h3b2bc31f),
	.w3(32'h3afec7f6),
	.w4(32'h3af77ef3),
	.w5(32'hbb3335d0),
	.w6(32'h3a2cc81b),
	.w7(32'h3aad334e),
	.w8(32'hbb875f7f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba276bb2),
	.w1(32'hbbec418d),
	.w2(32'hbc0e57b6),
	.w3(32'hbaa4691f),
	.w4(32'hbae35d8f),
	.w5(32'hbadb65df),
	.w6(32'hbace6233),
	.w7(32'hbb2cffca),
	.w8(32'hbb2cbcbb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aa2eb),
	.w1(32'h37bb7b1e),
	.w2(32'hbb1120c6),
	.w3(32'h39ba7e98),
	.w4(32'hbb074fa3),
	.w5(32'h3b5155a1),
	.w6(32'hb91fa899),
	.w7(32'hbb093ad2),
	.w8(32'h3b51adb9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81f1ff),
	.w1(32'h3b35cf67),
	.w2(32'h3a721605),
	.w3(32'h3b4d7d3f),
	.w4(32'h3af1ba92),
	.w5(32'h3b44378a),
	.w6(32'h3b2cbce1),
	.w7(32'h3ae002ee),
	.w8(32'h3b2a2de4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bea11),
	.w1(32'h39ddf84d),
	.w2(32'h3a19c2e1),
	.w3(32'h3b0809db),
	.w4(32'h3ab89826),
	.w5(32'h3ba1b549),
	.w6(32'h392e8a06),
	.w7(32'h3a736898),
	.w8(32'h3b9d0663),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9d078),
	.w1(32'h3b1d59c5),
	.w2(32'h3a10ae2f),
	.w3(32'h3b0fe28b),
	.w4(32'hb9e97cd6),
	.w5(32'hbb248925),
	.w6(32'h3ae37c2b),
	.w7(32'hba9dc9c8),
	.w8(32'hbabd2eee),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94b64f),
	.w1(32'h3a853f8a),
	.w2(32'h3b39a4bc),
	.w3(32'hbb5b6588),
	.w4(32'hb9a54db9),
	.w5(32'hbac18c13),
	.w6(32'hbb33cc43),
	.w7(32'hbaf4f43a),
	.w8(32'hb9c43ab0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d9c9b),
	.w1(32'hbbdb14d5),
	.w2(32'hbc53f82b),
	.w3(32'h3b19f92b),
	.w4(32'hba146897),
	.w5(32'hbbf29895),
	.w6(32'h39c94ec0),
	.w7(32'h39a19080),
	.w8(32'hbc08bcc7),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ef008),
	.w1(32'hbbf26c13),
	.w2(32'hbc270b62),
	.w3(32'h3aceaed4),
	.w4(32'h3a373b9d),
	.w5(32'hbb9c91ce),
	.w6(32'h3b0110a8),
	.w7(32'h3a993e67),
	.w8(32'hbb998634),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e3989),
	.w1(32'hbbadad26),
	.w2(32'hbc269875),
	.w3(32'hba269818),
	.w4(32'h3b05f6e7),
	.w5(32'hbbf3fd86),
	.w6(32'h3a61e038),
	.w7(32'h3a864815),
	.w8(32'hbc00895c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf591df),
	.w1(32'hba35ee46),
	.w2(32'hba1b55a3),
	.w3(32'hbad8946f),
	.w4(32'hb9c4c5e9),
	.w5(32'hba5bdc7e),
	.w6(32'hbb3382db),
	.w7(32'hba890e1c),
	.w8(32'h3a9a8c1b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae756db),
	.w1(32'hba884194),
	.w2(32'hb9ba67ee),
	.w3(32'hbb5b44de),
	.w4(32'hbb264ab8),
	.w5(32'hbb083211),
	.w6(32'hba2365ea),
	.w7(32'hba445261),
	.w8(32'hba96bef9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d2157),
	.w1(32'hb92fb12e),
	.w2(32'hbac37382),
	.w3(32'hb92f7db6),
	.w4(32'hba82f454),
	.w5(32'h39af4c1c),
	.w6(32'h39d3f7ff),
	.w7(32'hba151eee),
	.w8(32'h3a084500),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c4973),
	.w1(32'hba1f824f),
	.w2(32'hba0aba05),
	.w3(32'hb701067a),
	.w4(32'hba861d0d),
	.w5(32'hbac91baa),
	.w6(32'hbadc2259),
	.w7(32'hba5e0f03),
	.w8(32'hbb32afbe),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1eadc),
	.w1(32'hbbf9e145),
	.w2(32'hbc277dde),
	.w3(32'hba5647f5),
	.w4(32'hbb8e6c7d),
	.w5(32'hbbeea412),
	.w6(32'h39801bc5),
	.w7(32'hbb59b93b),
	.w8(32'hbb7a016e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2af0da),
	.w1(32'h3a21affb),
	.w2(32'hba93d6c6),
	.w3(32'hba8ba65c),
	.w4(32'hb9ca12f5),
	.w5(32'hbb497276),
	.w6(32'hbabbc98c),
	.w7(32'hbaf678d2),
	.w8(32'hbb0719a7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3dd20),
	.w1(32'hba2e0ecc),
	.w2(32'hbac28df3),
	.w3(32'hb981b9b3),
	.w4(32'hbaebd144),
	.w5(32'hba29eff2),
	.w6(32'hba090c6b),
	.w7(32'hbb352381),
	.w8(32'hbaa68e70),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74044e),
	.w1(32'hbb465d84),
	.w2(32'hbb16ebb9),
	.w3(32'hbb8253f6),
	.w4(32'hbb5a97d0),
	.w5(32'hbafd0b69),
	.w6(32'hbb38de00),
	.w7(32'hba4fa07c),
	.w8(32'h39d87c5a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24497a),
	.w1(32'hbb597afd),
	.w2(32'hbab3166e),
	.w3(32'hba9de81c),
	.w4(32'hb7ef8d47),
	.w5(32'h38f09df8),
	.w6(32'hbaed8619),
	.w7(32'hbac4a635),
	.w8(32'hb9707137),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a804e04),
	.w1(32'hba9dd88c),
	.w2(32'hbb058c21),
	.w3(32'h3acf51d6),
	.w4(32'h3a365c05),
	.w5(32'hbacc630a),
	.w6(32'h39f56fca),
	.w7(32'h394ea860),
	.w8(32'hbae57c62),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3937e361),
	.w1(32'hba348200),
	.w2(32'hba3767a6),
	.w3(32'hba1c2a16),
	.w4(32'h39a28815),
	.w5(32'hba4ffa0f),
	.w6(32'hbac96f47),
	.w7(32'hb9e66a66),
	.w8(32'hba8a96fd),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cdb0f),
	.w1(32'hbc76f625),
	.w2(32'hbc66bc4d),
	.w3(32'h3b8d988f),
	.w4(32'hbbd1b6a4),
	.w5(32'hbc02ee20),
	.w6(32'h3985f531),
	.w7(32'hbb8568ff),
	.w8(32'hbbbbce04),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa09e),
	.w1(32'h3a82d301),
	.w2(32'hb8293274),
	.w3(32'h3b43caac),
	.w4(32'h394d6eb2),
	.w5(32'hbaef1a2a),
	.w6(32'h3b0a82e6),
	.w7(32'hb9a864c6),
	.w8(32'hbb39f849),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb38515),
	.w1(32'h3a2be436),
	.w2(32'h3b35b44c),
	.w3(32'hb924ef58),
	.w4(32'h3b944b48),
	.w5(32'h3ba19c20),
	.w6(32'hb9a21887),
	.w7(32'h3b5383b2),
	.w8(32'h3c02758e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule