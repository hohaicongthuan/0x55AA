module layer_10_featuremap_129(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7403a8e),
	.w1(32'h38bc6c1a),
	.w2(32'h3a27c491),
	.w3(32'hb8f925d2),
	.w4(32'h3a34b16a),
	.w5(32'h3a1d97a3),
	.w6(32'hb998c051),
	.w7(32'h3ad99ac9),
	.w8(32'h3aafa41e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa60daa),
	.w1(32'h3a1cbf1c),
	.w2(32'h3a62ec99),
	.w3(32'h3acbdbf3),
	.w4(32'h3a067d4a),
	.w5(32'h3a2632f4),
	.w6(32'h3a39b156),
	.w7(32'hb9a14b71),
	.w8(32'h3a35bd15),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a563eed),
	.w1(32'h399449ce),
	.w2(32'hb978c2e1),
	.w3(32'h3a1e97ac),
	.w4(32'h397915c6),
	.w5(32'h37e78006),
	.w6(32'h392c16ae),
	.w7(32'hb93bf95c),
	.w8(32'h38c1de53),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eec67d),
	.w1(32'h38e9b667),
	.w2(32'hbab02746),
	.w3(32'hb94372f6),
	.w4(32'hba219672),
	.w5(32'hba51d8d5),
	.w6(32'hba909385),
	.w7(32'hbaa488a5),
	.w8(32'hbac51f17),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab520f7),
	.w1(32'h38a404b9),
	.w2(32'h3a09df4b),
	.w3(32'hba9e09ae),
	.w4(32'h3a08ff90),
	.w5(32'hb8e15f31),
	.w6(32'hb934fd89),
	.w7(32'hb981db55),
	.w8(32'hb95dc24b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370e7ab6),
	.w1(32'h399a2d33),
	.w2(32'hb92dc6e6),
	.w3(32'hb99a4c8f),
	.w4(32'hb770e9a3),
	.w5(32'hb9aadd39),
	.w6(32'h396c0aca),
	.w7(32'hb83a37e2),
	.w8(32'hb81902ca),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce097a),
	.w1(32'h3a9dc4ff),
	.w2(32'h3acc39b3),
	.w3(32'hb9018caf),
	.w4(32'h3aff14ce),
	.w5(32'h3b1a5133),
	.w6(32'h3a3c94fa),
	.w7(32'h3a9ab50a),
	.w8(32'h3b151f5a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eb6ef),
	.w1(32'h3ab51520),
	.w2(32'h3a4e68ee),
	.w3(32'h3b80be52),
	.w4(32'h3b0c2ea6),
	.w5(32'h39bc17cb),
	.w6(32'h3b4c5d65),
	.w7(32'h3a89cc1a),
	.w8(32'h3a1a405a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997ce70),
	.w1(32'hb8633739),
	.w2(32'h34561c18),
	.w3(32'h3a0fc5ad),
	.w4(32'h3a0a1b6f),
	.w5(32'hb90a251e),
	.w6(32'h395ad56f),
	.w7(32'h3a039428),
	.w8(32'hb8aeeb50),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b909923),
	.w1(32'h3b342bd8),
	.w2(32'h3b5e1127),
	.w3(32'h3b872964),
	.w4(32'h3b0be9ed),
	.w5(32'h3b4012b3),
	.w6(32'h3b3e647e),
	.w7(32'h3a3b4122),
	.w8(32'h3b1f6dbc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba028f2c),
	.w1(32'h391e6e33),
	.w2(32'hba5d7afc),
	.w3(32'hb98b961b),
	.w4(32'hb9bb981c),
	.w5(32'hba17de69),
	.w6(32'hba575155),
	.w7(32'hba1d1735),
	.w8(32'hba9ebdd9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cdcaf2),
	.w1(32'hba460960),
	.w2(32'hbae018dc),
	.w3(32'hb8df9b53),
	.w4(32'hba858b84),
	.w5(32'h396242b0),
	.w6(32'h39289ba7),
	.w7(32'hbaccced8),
	.w8(32'hb814a5c1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1edd02),
	.w1(32'h3a0fedde),
	.w2(32'h3ac2a8f9),
	.w3(32'h3b2bc3e2),
	.w4(32'h394580b7),
	.w5(32'h3a8155c8),
	.w6(32'h3acc202d),
	.w7(32'h39d28234),
	.w8(32'h3a833d03),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a9684),
	.w1(32'h3a526b15),
	.w2(32'h3a98d03d),
	.w3(32'hba1ae626),
	.w4(32'h3a5120ac),
	.w5(32'h3aaab857),
	.w6(32'h39bdee8b),
	.w7(32'h3a526342),
	.w8(32'h3a93b5bf),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac66e0b),
	.w1(32'h3acb2b67),
	.w2(32'h3a90bab1),
	.w3(32'h3abbe96e),
	.w4(32'h39075337),
	.w5(32'h3ae8a9e8),
	.w6(32'h3974481f),
	.w7(32'hba162442),
	.w8(32'h3a2cf8aa),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2574d7),
	.w1(32'h3a7fa48b),
	.w2(32'h3aadd5bb),
	.w3(32'h3b234975),
	.w4(32'h3a1c2b59),
	.w5(32'h3889b12a),
	.w6(32'h3b0b68f8),
	.w7(32'h399924e6),
	.w8(32'h38e57c55),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68dd792),
	.w1(32'hb94face4),
	.w2(32'hba3da5cc),
	.w3(32'h39554a75),
	.w4(32'hb9359c53),
	.w5(32'hba412abd),
	.w6(32'hb8fe1009),
	.w7(32'hb93ff62e),
	.w8(32'h381c9908),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9486),
	.w1(32'h3a9ccedb),
	.w2(32'h3ae56f51),
	.w3(32'h3ac18038),
	.w4(32'h3ab30b80),
	.w5(32'h3ad7681d),
	.w6(32'h3b03cbc9),
	.w7(32'h39977b6a),
	.w8(32'h3a427bfd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b361a97),
	.w1(32'h3a87e1cf),
	.w2(32'h3ab16ffc),
	.w3(32'h3b02ad3b),
	.w4(32'h3ac7f926),
	.w5(32'h3ac33c9a),
	.w6(32'h3a9ec9ec),
	.w7(32'h3a39e329),
	.w8(32'h3aac7040),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39413a1b),
	.w1(32'hb97ea908),
	.w2(32'hb8d03de2),
	.w3(32'h37c9a369),
	.w4(32'hb8a02ddc),
	.w5(32'hb9519250),
	.w6(32'hb97624bb),
	.w7(32'hb99a2cb4),
	.w8(32'h390c4276),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a894c),
	.w1(32'hba055a77),
	.w2(32'hba63d6ba),
	.w3(32'h387ab148),
	.w4(32'hba02d195),
	.w5(32'hb9fbd2c4),
	.w6(32'hba3a0c3a),
	.w7(32'hba5f4202),
	.w8(32'hb9ecdf4f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f2218),
	.w1(32'hb9932607),
	.w2(32'hbaf7dba6),
	.w3(32'h385cdf9c),
	.w4(32'hb9d0b4f6),
	.w5(32'hb9224ff2),
	.w6(32'hb9fa0e6a),
	.w7(32'hba540eda),
	.w8(32'hb8a081a0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f8fc7),
	.w1(32'hba8e9af9),
	.w2(32'h3a564e35),
	.w3(32'h3b0484b0),
	.w4(32'hb939aea9),
	.w5(32'h3a1144f2),
	.w6(32'hb987e311),
	.w7(32'hba84dce3),
	.w8(32'h39d250ad),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407d2b),
	.w1(32'h3ac68045),
	.w2(32'h3b367662),
	.w3(32'h3b24794c),
	.w4(32'h3a4f5d31),
	.w5(32'h3ad8c38a),
	.w6(32'h3b049d1b),
	.w7(32'hb99b10d1),
	.w8(32'h3a6994f7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b531532),
	.w1(32'hba3d34ae),
	.w2(32'h3a137535),
	.w3(32'h3b56317e),
	.w4(32'hb990b842),
	.w5(32'h388e0dd3),
	.w6(32'h3b067ae5),
	.w7(32'hbad9755c),
	.w8(32'hb9b97753),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92626c5),
	.w1(32'h39dacbc6),
	.w2(32'h36b385d4),
	.w3(32'hb9bf5c81),
	.w4(32'h39e38189),
	.w5(32'h398fdcbe),
	.w6(32'hb7b7d97c),
	.w7(32'h3a130d19),
	.w8(32'h3a0ae2bd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10ddd3),
	.w1(32'hb8b237e3),
	.w2(32'hb958e442),
	.w3(32'hb9ddc678),
	.w4(32'h37136b4c),
	.w5(32'hb94a4552),
	.w6(32'hb966e12f),
	.w7(32'hb98e2f0f),
	.w8(32'h38df7238),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eaa0ee),
	.w1(32'hbabaf1ba),
	.w2(32'hb8cbf70b),
	.w3(32'h3a334517),
	.w4(32'hba62bc08),
	.w5(32'hba389070),
	.w6(32'h393252df),
	.w7(32'hbb0d72c2),
	.w8(32'hbad2cf36),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c5230),
	.w1(32'hbaffef3c),
	.w2(32'hbb21aca9),
	.w3(32'h3a0c33f0),
	.w4(32'hba85f2d1),
	.w5(32'hbae2d061),
	.w6(32'hb9a1eda2),
	.w7(32'hbb2e0ed6),
	.w8(32'hbada2bcf),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7b158),
	.w1(32'hba5d216f),
	.w2(32'h3ae4e0dc),
	.w3(32'h3af9f0b0),
	.w4(32'hba31e490),
	.w5(32'h3ab4a9c1),
	.w6(32'h3a1752c6),
	.w7(32'hbada135b),
	.w8(32'h3a0ca3bf),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89847ff),
	.w1(32'hb9668591),
	.w2(32'hb9ec309f),
	.w3(32'hb9904f49),
	.w4(32'hb9702338),
	.w5(32'hb984493e),
	.w6(32'hb9923cc1),
	.w7(32'hb9e25dad),
	.w8(32'hb950ff36),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f29fa),
	.w1(32'hb8827965),
	.w2(32'hb9920162),
	.w3(32'h388d4b2a),
	.w4(32'hb92256fb),
	.w5(32'hb9d8b2b1),
	.w6(32'hb88602cc),
	.w7(32'hb93d21b6),
	.w8(32'hb8a71c74),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5ccb5),
	.w1(32'h39036100),
	.w2(32'h3b24edc8),
	.w3(32'h3aa20d2e),
	.w4(32'h3a05053c),
	.w5(32'h3ae377e4),
	.w6(32'h3a091fa0),
	.w7(32'h3a5a63f7),
	.w8(32'h3a505eed),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11c3b5),
	.w1(32'h39c7b4e9),
	.w2(32'hb95dbc94),
	.w3(32'h3b23c563),
	.w4(32'h39ff7242),
	.w5(32'hbac19a00),
	.w6(32'h3aba6d31),
	.w7(32'hba7a98d6),
	.w8(32'hba56cc6a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb6146),
	.w1(32'h3a90ef24),
	.w2(32'hb8162370),
	.w3(32'hb6d16429),
	.w4(32'h3a91dc6f),
	.w5(32'h390eca4e),
	.w6(32'h3aa794a0),
	.w7(32'h3a098197),
	.w8(32'h39b9e36c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a315970),
	.w1(32'h39b2e9d7),
	.w2(32'h3976bdfe),
	.w3(32'h39f79a94),
	.w4(32'h39daabd9),
	.w5(32'h39adec19),
	.w6(32'hb8dbae58),
	.w7(32'h398b02ac),
	.w8(32'h3a24610e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b058258),
	.w1(32'h3a121315),
	.w2(32'h3a761490),
	.w3(32'h3ae99d0c),
	.w4(32'hb9e70c78),
	.w5(32'hb88511d7),
	.w6(32'hba65d1b7),
	.w7(32'hbb04fbad),
	.w8(32'h3936fc32),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65e73f),
	.w1(32'hbb404ffc),
	.w2(32'hba8b49f4),
	.w3(32'h3b3bca56),
	.w4(32'hbb5e7aeb),
	.w5(32'hba491ed4),
	.w6(32'h3ab9d699),
	.w7(32'hbbaab389),
	.w8(32'hbaf48329),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d138d),
	.w1(32'hbba9a2d4),
	.w2(32'hbb75ca62),
	.w3(32'h3b0dd3c0),
	.w4(32'hbb8c15c5),
	.w5(32'hbb11a5a7),
	.w6(32'h3a1656d9),
	.w7(32'hbb95dd5b),
	.w8(32'hbb05abda),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a957684),
	.w1(32'h3a5dd692),
	.w2(32'h3a772d04),
	.w3(32'h3a6a0675),
	.w4(32'h3a6b98fd),
	.w5(32'h3a65b6ef),
	.w6(32'h3aa8a2f5),
	.w7(32'h39df1d25),
	.w8(32'h3a3ab649),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34ee32),
	.w1(32'h38d737e1),
	.w2(32'h39bca683),
	.w3(32'h3a35b95f),
	.w4(32'h3814070b),
	.w5(32'h38c9e680),
	.w6(32'h3902dca4),
	.w7(32'h396963b4),
	.w8(32'hb96e8d06),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d41b16),
	.w1(32'hb82d3888),
	.w2(32'hba227182),
	.w3(32'hba23b948),
	.w4(32'hb9774376),
	.w5(32'hb990096d),
	.w6(32'h37af4150),
	.w7(32'hb9c266e2),
	.w8(32'hb938e235),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d60e9),
	.w1(32'h39293f1c),
	.w2(32'h37f37a5c),
	.w3(32'h3a027d1c),
	.w4(32'hb8b1d025),
	.w5(32'hb9feefc4),
	.w6(32'h391eaad5),
	.w7(32'h38fe02bb),
	.w8(32'h3982b0eb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82c129),
	.w1(32'h3b0af83c),
	.w2(32'h3acc9047),
	.w3(32'h3b60a7b8),
	.w4(32'h3b1100b7),
	.w5(32'h3ab865db),
	.w6(32'h3b80593a),
	.w7(32'h3a5a138b),
	.w8(32'h3a25dcbe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b323587),
	.w1(32'h3a85762c),
	.w2(32'h3b28a2a1),
	.w3(32'h3b0aa909),
	.w4(32'h3a31cbff),
	.w5(32'h3af590ef),
	.w6(32'h3ae7d077),
	.w7(32'hb93a8e0e),
	.w8(32'h3a33f284),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bd1f2),
	.w1(32'h3a53fb2e),
	.w2(32'h3b184dff),
	.w3(32'h3b489bbe),
	.w4(32'h3a88a573),
	.w5(32'h3aa598ce),
	.w6(32'h3b289c5b),
	.w7(32'hba18d745),
	.w8(32'h3a2a81de),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b6c45),
	.w1(32'h3a983476),
	.w2(32'h3a4f8483),
	.w3(32'h3b6459e7),
	.w4(32'h3affaca2),
	.w5(32'h3b3b525e),
	.w6(32'h3b130b7f),
	.w7(32'hb9a988c5),
	.w8(32'h3942edba),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395293e4),
	.w1(32'hb98f4cb2),
	.w2(32'hb955bda3),
	.w3(32'h3b006418),
	.w4(32'h3a97bb77),
	.w5(32'h3a98fd97),
	.w6(32'hba2a20f7),
	.w7(32'h388e004d),
	.w8(32'h3a93a934),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d4f1),
	.w1(32'hb9856015),
	.w2(32'hb8cb980b),
	.w3(32'hba344f03),
	.w4(32'hb974ae4a),
	.w5(32'hb9fa8ab5),
	.w6(32'hb9a25a3c),
	.w7(32'hb91ac203),
	.w8(32'h38818896),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a57f4),
	.w1(32'h3a22b754),
	.w2(32'h3a93014e),
	.w3(32'h39868ad1),
	.w4(32'h3a699c9e),
	.w5(32'h3a66f25b),
	.w6(32'h3a56441e),
	.w7(32'h3a87b784),
	.w8(32'h3a863c0f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f61eaf),
	.w1(32'hb98c0e7a),
	.w2(32'hb981882f),
	.w3(32'hb8824919),
	.w4(32'h391a169f),
	.w5(32'hb7c9678a),
	.w6(32'h38b45110),
	.w7(32'hb9ac5a51),
	.w8(32'hb75d12b1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfe6e5),
	.w1(32'h3732fdb8),
	.w2(32'h3b4c42f2),
	.w3(32'h3ab3d9ed),
	.w4(32'h39ee4d35),
	.w5(32'h3b02f226),
	.w6(32'h3ab13831),
	.w7(32'h3948ab36),
	.w8(32'h39ec7f45),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7b8e3),
	.w1(32'h3968d806),
	.w2(32'hb991f628),
	.w3(32'h3afda939),
	.w4(32'h39ce8228),
	.w5(32'h38bf1578),
	.w6(32'h3a1389ee),
	.w7(32'hb945c89e),
	.w8(32'hb90d4e92),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f4481),
	.w1(32'h3aa71ab2),
	.w2(32'h3b0b354f),
	.w3(32'h3ae25aaa),
	.w4(32'h3ad2fcce),
	.w5(32'h3b0a9f3a),
	.w6(32'h3a954957),
	.w7(32'hb8e8e1cf),
	.w8(32'h3a791c75),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39237acc),
	.w1(32'hb947929a),
	.w2(32'hb99281ea),
	.w3(32'h395311bf),
	.w4(32'hb91d5195),
	.w5(32'hb9ef5155),
	.w6(32'h3a02bf7e),
	.w7(32'hb98886a7),
	.w8(32'hb998d49e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6ca1c),
	.w1(32'hb7ebef62),
	.w2(32'h398fc315),
	.w3(32'hba39d284),
	.w4(32'hb97b0308),
	.w5(32'hb9d33491),
	.w6(32'hba2201f2),
	.w7(32'hb5b0cfec),
	.w8(32'hb9a007bb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396741d1),
	.w1(32'h3a09cd04),
	.w2(32'h389e2aa1),
	.w3(32'h39039a2d),
	.w4(32'h39dae14a),
	.w5(32'h3a079277),
	.w6(32'h39d65a7b),
	.w7(32'hb95658e3),
	.w8(32'h391e31d1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36d289),
	.w1(32'h3a1cea1c),
	.w2(32'h3aba469c),
	.w3(32'h3a100de3),
	.w4(32'h3a688750),
	.w5(32'hb97c6c20),
	.w6(32'h3a8b4a72),
	.w7(32'h39632f6f),
	.w8(32'h3a1eb109),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2750e),
	.w1(32'h39a64ee1),
	.w2(32'hb990a327),
	.w3(32'hb9103bbb),
	.w4(32'h3a434692),
	.w5(32'h3a128107),
	.w6(32'h3a9eb569),
	.w7(32'h39dfd10c),
	.w8(32'h3a2fe14b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d52a3),
	.w1(32'h39d0d282),
	.w2(32'h3905dab5),
	.w3(32'h3a3e0a1a),
	.w4(32'h398ea1a3),
	.w5(32'h390537bc),
	.w6(32'h36803ecd),
	.w7(32'h37a29852),
	.w8(32'h392d70db),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ceeab),
	.w1(32'h3aa6c201),
	.w2(32'h3a7da9c3),
	.w3(32'h3b0c6c83),
	.w4(32'h3adc2216),
	.w5(32'h3a8df080),
	.w6(32'h3b148cf6),
	.w7(32'h3aa69dfe),
	.w8(32'h39200f95),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09bc78),
	.w1(32'h398bc5e0),
	.w2(32'h39e1fc98),
	.w3(32'h3aae0d3b),
	.w4(32'h39a3ed04),
	.w5(32'hb525ba2b),
	.w6(32'h3a93c13f),
	.w7(32'h39b48d6f),
	.w8(32'h38abecc4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10f894),
	.w1(32'hb7f38338),
	.w2(32'h3b865798),
	.w3(32'h39e614b5),
	.w4(32'hb7c8ce21),
	.w5(32'h3b2e02b1),
	.w6(32'h3943794b),
	.w7(32'h3b4b4333),
	.w8(32'h3ae79d40),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4c620),
	.w1(32'h3a037448),
	.w2(32'hb956bbfd),
	.w3(32'h3aa0c303),
	.w4(32'h3a20f297),
	.w5(32'h385adac3),
	.w6(32'h3a1f193d),
	.w7(32'hb689793f),
	.w8(32'h398289e4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94344c4),
	.w1(32'hb7a61615),
	.w2(32'h39592a59),
	.w3(32'hb9a5e2f7),
	.w4(32'h39d05c6d),
	.w5(32'h3949b29a),
	.w6(32'hb81ea50a),
	.w7(32'h3989b1ef),
	.w8(32'h3a06831a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2fc91),
	.w1(32'h3976423e),
	.w2(32'h3a574655),
	.w3(32'h38ea71af),
	.w4(32'h37bfc00b),
	.w5(32'hba1cbdd0),
	.w6(32'h3a2307be),
	.w7(32'hb90e764e),
	.w8(32'hb60908dc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b153578),
	.w1(32'h395c685c),
	.w2(32'h395276ee),
	.w3(32'h3b05d2a7),
	.w4(32'h39e9926d),
	.w5(32'h38ebb2d9),
	.w6(32'h3a86bd1d),
	.w7(32'h39a1d4c4),
	.w8(32'hba5224bb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b6507),
	.w1(32'hb9bfc629),
	.w2(32'h3a4cef0a),
	.w3(32'h3b0f007d),
	.w4(32'h3927de0e),
	.w5(32'h3a2b1af5),
	.w6(32'h3a994332),
	.w7(32'hbab52016),
	.w8(32'hba53b4fb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad582b1),
	.w1(32'hbaf92a98),
	.w2(32'hbae0121a),
	.w3(32'h3a2ca128),
	.w4(32'hbb0847e9),
	.w5(32'hbae05100),
	.w6(32'h3a7ee345),
	.w7(32'hbb57028c),
	.w8(32'hbb288c16),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e0267),
	.w1(32'hbaa99a70),
	.w2(32'h3b28d60e),
	.w3(32'h3b3809b6),
	.w4(32'hbacd76a7),
	.w5(32'h395f4f2a),
	.w6(32'h3b013c2c),
	.w7(32'hbb5cb0d4),
	.w8(32'h38fc9c8a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865707e),
	.w1(32'h3a3b9a50),
	.w2(32'h39a51eb8),
	.w3(32'hb78efaa3),
	.w4(32'h3a3eef5d),
	.w5(32'h39a06777),
	.w6(32'h3a46f941),
	.w7(32'h3a3f7227),
	.w8(32'h3a314dde),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a264847),
	.w1(32'h39a68fcd),
	.w2(32'h39087be5),
	.w3(32'h398a09d0),
	.w4(32'h39237874),
	.w5(32'h390563bc),
	.w6(32'h391f7dc4),
	.w7(32'h37f4365a),
	.w8(32'h36dfde53),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a5016),
	.w1(32'h393c0b1c),
	.w2(32'h38729e3f),
	.w3(32'h37cd3ea3),
	.w4(32'h391afba1),
	.w5(32'h383b867f),
	.w6(32'h38a036c3),
	.w7(32'hb8081aef),
	.w8(32'h38c0d7b5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa26ebc),
	.w1(32'h3809906a),
	.w2(32'hba37ec1b),
	.w3(32'h3a7174e7),
	.w4(32'hb7c2b322),
	.w5(32'hba1c9e9b),
	.w6(32'h3a058032),
	.w7(32'hb9a48951),
	.w8(32'hb97a35b3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963763d),
	.w1(32'h3a8b659e),
	.w2(32'h39e59c2d),
	.w3(32'h3303cbf5),
	.w4(32'h3ab02686),
	.w5(32'h3a899723),
	.w6(32'h3a80a9ec),
	.w7(32'h3a3c7757),
	.w8(32'h3a8468f4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac56895),
	.w1(32'h3a675401),
	.w2(32'h397dd215),
	.w3(32'h3aebf7ef),
	.w4(32'h3a886b9f),
	.w5(32'h3acf3042),
	.w6(32'h3a29af29),
	.w7(32'h3a3640a4),
	.w8(32'hba2fe6a9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aec55),
	.w1(32'h3ae22e14),
	.w2(32'h3a8cb28c),
	.w3(32'h3b666176),
	.w4(32'h3a6953f3),
	.w5(32'h39e752c6),
	.w6(32'h3b012a99),
	.w7(32'h3aa73b38),
	.w8(32'h3a13d76e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17ed41),
	.w1(32'h3aa46936),
	.w2(32'h3b105020),
	.w3(32'h3b06f036),
	.w4(32'h3aa12b8d),
	.w5(32'h3b078095),
	.w6(32'h3ac1ec8c),
	.w7(32'h3a6b3118),
	.w8(32'h3aa1d348),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d872c),
	.w1(32'h39b9a1ef),
	.w2(32'h3a3fa799),
	.w3(32'h3a6d5f5b),
	.w4(32'hb9cc9973),
	.w5(32'hba0e7aca),
	.w6(32'h3ad9351b),
	.w7(32'h39d03278),
	.w8(32'h386ca8ed),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c3bfc),
	.w1(32'hb9233eb8),
	.w2(32'hb7647eff),
	.w3(32'h3a96395f),
	.w4(32'h399dc2d6),
	.w5(32'h39fa3aa8),
	.w6(32'hb9ab3906),
	.w7(32'hb9d97fac),
	.w8(32'h39b10ca0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa64cce),
	.w1(32'hb9c21a6a),
	.w2(32'hb9b6e2a7),
	.w3(32'h3a79ff5e),
	.w4(32'hba0d5e13),
	.w5(32'hba41a409),
	.w6(32'h3a15782d),
	.w7(32'hbab12ccf),
	.w8(32'hba902862),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc3b6f),
	.w1(32'h3a201671),
	.w2(32'h37ab8a57),
	.w3(32'hb8e05921),
	.w4(32'h3a688f24),
	.w5(32'h3aa5ca49),
	.w6(32'h39e96a1a),
	.w7(32'hba00663b),
	.w8(32'h3994e9a4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1035de),
	.w1(32'hba16f60b),
	.w2(32'hb9fab2cc),
	.w3(32'h3a255849),
	.w4(32'hb9a3d33f),
	.w5(32'hb9b6fee7),
	.w6(32'hb9c38a7b),
	.w7(32'hb9469384),
	.w8(32'hb90ffc35),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f8364),
	.w1(32'h3a6a5ec6),
	.w2(32'h3a101147),
	.w3(32'hb9677d5e),
	.w4(32'h3a94d000),
	.w5(32'h3aa9c3ad),
	.w6(32'h3a57a486),
	.w7(32'h3a339869),
	.w8(32'h3a723cd0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53d6ea),
	.w1(32'h38e04b56),
	.w2(32'hba28c139),
	.w3(32'h3a74d696),
	.w4(32'h39ec16a3),
	.w5(32'hb96a96a8),
	.w6(32'h39424033),
	.w7(32'hb88f51c0),
	.w8(32'hb9a789af),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90db057),
	.w1(32'hb97e13a8),
	.w2(32'hb8374c94),
	.w3(32'h38e8f9d8),
	.w4(32'hb9578d77),
	.w5(32'h39999855),
	.w6(32'hb9b712ab),
	.w7(32'hb9da1114),
	.w8(32'hb934728e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b49ce),
	.w1(32'hba22654a),
	.w2(32'h3a3c7be6),
	.w3(32'h3b1047b9),
	.w4(32'hb97f3833),
	.w5(32'h38f4c5bf),
	.w6(32'h3aa8baa9),
	.w7(32'hba4ead19),
	.w8(32'hba31705b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974cfb1),
	.w1(32'hb9ad436a),
	.w2(32'hba10b49b),
	.w3(32'h39d23054),
	.w4(32'hb9861ec3),
	.w5(32'hb9bd6929),
	.w6(32'hb92d13fc),
	.w7(32'hb9ab1503),
	.w8(32'hb9a5a8e7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f75154),
	.w1(32'h3979876d),
	.w2(32'h3a627ce7),
	.w3(32'h3a2d8a96),
	.w4(32'h3979364d),
	.w5(32'h3a46d9df),
	.w6(32'h39093d49),
	.w7(32'hba10ce84),
	.w8(32'h38b19268),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd2ee3),
	.w1(32'hb90dbdb6),
	.w2(32'hb9c98153),
	.w3(32'h3ab4dfa4),
	.w4(32'hb998ed4c),
	.w5(32'hb9e6d166),
	.w6(32'h3aae80ae),
	.w7(32'hba5693ab),
	.w8(32'hbaa39527),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398934ac),
	.w1(32'hbadd9947),
	.w2(32'hba9d8b55),
	.w3(32'h39e4b200),
	.w4(32'hbad7e063),
	.w5(32'hba3ef206),
	.w6(32'hb9fbef37),
	.w7(32'hbb1d2d54),
	.w8(32'hba9b7ac4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb945832d),
	.w1(32'hba8d3b57),
	.w2(32'hba13a86c),
	.w3(32'h3aad269a),
	.w4(32'h3a13c090),
	.w5(32'h3a5aefae),
	.w6(32'h3a313764),
	.w7(32'h39ace770),
	.w8(32'h39ce2eb0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c723a),
	.w1(32'h39fbf0c3),
	.w2(32'h398ca133),
	.w3(32'h37b59878),
	.w4(32'h39d8a0b2),
	.w5(32'h3a0ed7f1),
	.w6(32'hb7378194),
	.w7(32'hba323d03),
	.w8(32'hb88f49fc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d78c),
	.w1(32'h3a1c174e),
	.w2(32'h3ae124a2),
	.w3(32'h3b03c548),
	.w4(32'hb8654717),
	.w5(32'h3a57e385),
	.w6(32'h3a90ba52),
	.w7(32'hba8b6424),
	.w8(32'hb89512bd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf0234),
	.w1(32'h3894fb44),
	.w2(32'h3a783eca),
	.w3(32'h3a1d545c),
	.w4(32'h39203027),
	.w5(32'h3a24eae9),
	.w6(32'h39b09ba9),
	.w7(32'hba0c61a0),
	.w8(32'h394328d0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae96868),
	.w1(32'hb9e21359),
	.w2(32'h3a0f5291),
	.w3(32'h3abc7586),
	.w4(32'hba32a358),
	.w5(32'h3a8c6045),
	.w6(32'h3aab6e81),
	.w7(32'hbaa95e00),
	.w8(32'hb881b906),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2b153),
	.w1(32'hbab409b1),
	.w2(32'hba53aac6),
	.w3(32'hba2af7c5),
	.w4(32'hbadcbfa0),
	.w5(32'hbb0a1f7b),
	.w6(32'hbacb27ed),
	.w7(32'hbaad67b0),
	.w8(32'hbae001fd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7165f),
	.w1(32'hb7837c4f),
	.w2(32'h3b3f36df),
	.w3(32'h3a82d89e),
	.w4(32'h391a4152),
	.w5(32'h3aa5de56),
	.w6(32'h3ac1d802),
	.w7(32'h3a78bfc1),
	.w8(32'h3aecfb78),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9392af),
	.w1(32'hba6ebd73),
	.w2(32'hbac285b7),
	.w3(32'h3b2addfa),
	.w4(32'hb78ca966),
	.w5(32'hb8f7c765),
	.w6(32'h3b0914d4),
	.w7(32'h399d0035),
	.w8(32'h3a215440),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11de89),
	.w1(32'hba2f15e6),
	.w2(32'hbab4e686),
	.w3(32'h3aa7f5db),
	.w4(32'hba4cedc2),
	.w5(32'hba81524f),
	.w6(32'hba209bf5),
	.w7(32'hbaf14da9),
	.w8(32'hbae97315),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b3951),
	.w1(32'hbb454360),
	.w2(32'h3b0e2f38),
	.w3(32'h3b111d38),
	.w4(32'hbb0b8dce),
	.w5(32'h395ba689),
	.w6(32'h3b4c2738),
	.w7(32'hbb3f4ef8),
	.w8(32'hb90ee107),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b379106),
	.w1(32'h3b196239),
	.w2(32'h3b9b3ce6),
	.w3(32'h3b305486),
	.w4(32'h3af2c813),
	.w5(32'h3b1ebfb6),
	.w6(32'h3af33d8a),
	.w7(32'h3997ce8e),
	.w8(32'h3aff3345),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58f960),
	.w1(32'hb8fc8ada),
	.w2(32'hb99afdbf),
	.w3(32'h3a106908),
	.w4(32'hba5c89fd),
	.w5(32'hba1efadb),
	.w6(32'hbab40acc),
	.w7(32'hbab1b474),
	.w8(32'hb9839d77),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1abb09),
	.w1(32'hba1e0348),
	.w2(32'hba233ff1),
	.w3(32'h38d47f80),
	.w4(32'hb9932093),
	.w5(32'hba44faed),
	.w6(32'hb9d7d547),
	.w7(32'hba1472fe),
	.w8(32'hba96a78f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aa4c6),
	.w1(32'h3a60e8d6),
	.w2(32'h39a26d4b),
	.w3(32'h3b2fc0cb),
	.w4(32'hba1d0415),
	.w5(32'hb844eec2),
	.w6(32'h390326b9),
	.w7(32'hbac6d2e6),
	.w8(32'hbabbaf67),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae060a7),
	.w1(32'h39548857),
	.w2(32'h3a1a7804),
	.w3(32'h3abf70c1),
	.w4(32'h39f8d6ce),
	.w5(32'h3a428a6c),
	.w6(32'h39b450e5),
	.w7(32'hb7e634a6),
	.w8(32'h3a177dc7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39802104),
	.w1(32'h3a50eee5),
	.w2(32'h397825a0),
	.w3(32'h38ee7f31),
	.w4(32'h3a430b05),
	.w5(32'h3a0d68ba),
	.w6(32'h3a4d5dbd),
	.w7(32'h3a106e36),
	.w8(32'h39ccd6a7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a546111),
	.w1(32'hba41428a),
	.w2(32'hba264810),
	.w3(32'h394d9713),
	.w4(32'hba2b8c9e),
	.w5(32'hb9c5d21d),
	.w6(32'hb993a2c8),
	.w7(32'hba46f27e),
	.w8(32'hb9d4738d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae35386),
	.w1(32'h3a424de4),
	.w2(32'h3aa96a51),
	.w3(32'h3ace673d),
	.w4(32'h3a52a0f7),
	.w5(32'h3a82fc3b),
	.w6(32'h3ace74ef),
	.w7(32'h3a8c833b),
	.w8(32'h3ad408f4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e3009),
	.w1(32'h3a8484f1),
	.w2(32'h3b44335c),
	.w3(32'h3a328b2f),
	.w4(32'h3aae5965),
	.w5(32'h3b1160fa),
	.w6(32'h3a6c3270),
	.w7(32'h3a309b38),
	.w8(32'h3b06a535),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0e917),
	.w1(32'h39528d55),
	.w2(32'h3a9e305a),
	.w3(32'h3b0a808c),
	.w4(32'h388d082a),
	.w5(32'h3a62136d),
	.w6(32'h39e6bcf6),
	.w7(32'hba35ba5e),
	.w8(32'h3a9dbd3a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b6cfe),
	.w1(32'hb91ccb69),
	.w2(32'h3b7db29c),
	.w3(32'h3a4ae551),
	.w4(32'hb96b0df0),
	.w5(32'h3af8aba4),
	.w6(32'h39bc8f2b),
	.w7(32'h3a9588b1),
	.w8(32'h3aa3ead5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a141158),
	.w1(32'hba90fba1),
	.w2(32'hbab07073),
	.w3(32'h3a913362),
	.w4(32'hba2a24bb),
	.w5(32'hb9b8d493),
	.w6(32'hb8405ac6),
	.w7(32'hbad6b6d6),
	.w8(32'hba8fda05),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac68873),
	.w1(32'h3ad6740d),
	.w2(32'h3adfb727),
	.w3(32'h3a9901cf),
	.w4(32'h3a8320d0),
	.w5(32'h3a51608c),
	.w6(32'h3add53e7),
	.w7(32'h39e87f9c),
	.w8(32'hb815ddb0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9282a),
	.w1(32'h399f85fe),
	.w2(32'h3a9d614a),
	.w3(32'h3abecb23),
	.w4(32'h3a0d3936),
	.w5(32'h3a1d952e),
	.w6(32'h3a513631),
	.w7(32'h399c9ffb),
	.w8(32'h39fc9d9a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ac73c),
	.w1(32'h39c9b3e5),
	.w2(32'h3990cd53),
	.w3(32'h3996ee1c),
	.w4(32'h34cdce3c),
	.w5(32'hb93ec908),
	.w6(32'h392edceb),
	.w7(32'h380eb41f),
	.w8(32'hb822ddd7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a05845),
	.w1(32'h398e1d48),
	.w2(32'h3947848d),
	.w3(32'hb754a0fc),
	.w4(32'hb8bc25a5),
	.w5(32'hb992cbbc),
	.w6(32'h39a15940),
	.w7(32'hb7b2ece4),
	.w8(32'hb92fbe79),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39940dc3),
	.w1(32'h399c463a),
	.w2(32'h38ac60d9),
	.w3(32'h3850e565),
	.w4(32'hb854e1c6),
	.w5(32'hb99de5d5),
	.w6(32'h39992bdc),
	.w7(32'hb740ba73),
	.w8(32'hb8f5e133),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370f4edb),
	.w1(32'h39974cae),
	.w2(32'hba071b0b),
	.w3(32'hb987b4eb),
	.w4(32'h39e83dca),
	.w5(32'h39ccb444),
	.w6(32'hb86c81e8),
	.w7(32'h394495a4),
	.w8(32'hb99a852e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc24ed),
	.w1(32'h3975a9dd),
	.w2(32'h3ab30201),
	.w3(32'h3aca42cf),
	.w4(32'h3a1022ff),
	.w5(32'hb8da3b04),
	.w6(32'h3a33b799),
	.w7(32'hba7d3220),
	.w8(32'h3963cbc8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383a8c07),
	.w1(32'hba26f1c0),
	.w2(32'hbab26465),
	.w3(32'hb9ffb844),
	.w4(32'hba247ead),
	.w5(32'hba7aa105),
	.w6(32'hba1f9843),
	.w7(32'hba6fcced),
	.w8(32'hba4aaa0f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d60ad),
	.w1(32'h39979c5d),
	.w2(32'hb74ad2da),
	.w3(32'h39b1ac39),
	.w4(32'h3a259d99),
	.w5(32'h397e86a3),
	.w6(32'hb9a048b4),
	.w7(32'hb68c20c5),
	.w8(32'h38dfefb7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf5b7e),
	.w1(32'h39a82001),
	.w2(32'h3abd8524),
	.w3(32'h3abba074),
	.w4(32'hb98a2753),
	.w5(32'h3a214dc7),
	.w6(32'h3acbe2c2),
	.w7(32'hba8ba7cf),
	.w8(32'h3a073c52),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e876c9),
	.w1(32'h39ca0dec),
	.w2(32'hba9df759),
	.w3(32'h3992b592),
	.w4(32'h3a084057),
	.w5(32'h3a665c2d),
	.w6(32'hb9b6f87a),
	.w7(32'hb8427e02),
	.w8(32'h398a0543),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba455d49),
	.w1(32'hb9c6ede4),
	.w2(32'hbaab45d5),
	.w3(32'h39defa11),
	.w4(32'hba0f3433),
	.w5(32'hba66a0f4),
	.w6(32'hb98ccae4),
	.w7(32'hb9f65903),
	.w8(32'hba16e445),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2451b0),
	.w1(32'hba217c44),
	.w2(32'hba3a56c5),
	.w3(32'hba6b91dc),
	.w4(32'hb9e07e0e),
	.w5(32'hba0037fb),
	.w6(32'hba193b93),
	.w7(32'hba3c8523),
	.w8(32'hb980738c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b631ed),
	.w1(32'h396bc6de),
	.w2(32'h39caa4fd),
	.w3(32'h397a7e32),
	.w4(32'h396ba074),
	.w5(32'h39a9ec4f),
	.w6(32'h38ea18a2),
	.w7(32'h39c846fe),
	.w8(32'h39ff77f3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a4903),
	.w1(32'h3a133a9e),
	.w2(32'h3a82b011),
	.w3(32'h3a6d7e69),
	.w4(32'h3ab3b88b),
	.w5(32'h3a9cc464),
	.w6(32'h38607903),
	.w7(32'h3983aeed),
	.w8(32'hb9f057ae),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae92eac),
	.w1(32'h3af70d36),
	.w2(32'h3b3e2a64),
	.w3(32'h3ad2685f),
	.w4(32'h3abd527f),
	.w5(32'h3b09ae20),
	.w6(32'h3a224881),
	.w7(32'h3a716b31),
	.w8(32'h3ab37b4d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39213af7),
	.w1(32'h38c5b8f7),
	.w2(32'hb73ec939),
	.w3(32'h38f852d3),
	.w4(32'h38bcbd71),
	.w5(32'hb7bbedb5),
	.w6(32'hb8c0d044),
	.w7(32'hb8c7c0a3),
	.w8(32'hb911cd00),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22331e),
	.w1(32'h392c7e3e),
	.w2(32'h39dcb673),
	.w3(32'h3a627fce),
	.w4(32'h39ac95e4),
	.w5(32'h39df9ead),
	.w6(32'h3a752569),
	.w7(32'h397abe45),
	.w8(32'h39811cbb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc4ee5),
	.w1(32'hb91ad885),
	.w2(32'h38c366dd),
	.w3(32'h3a01a9dc),
	.w4(32'hb7fb5cfa),
	.w5(32'h38a99888),
	.w6(32'h3956e19d),
	.w7(32'hb9dd4c64),
	.w8(32'hb907a2fa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69a56d),
	.w1(32'h388564c6),
	.w2(32'h39f59b22),
	.w3(32'h3a3df704),
	.w4(32'hb7e063ab),
	.w5(32'h38e194a2),
	.w6(32'h3a25289a),
	.w7(32'hb80b0cb3),
	.w8(32'h38ee201e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c8ed5),
	.w1(32'h39dcfa98),
	.w2(32'h3a5c456e),
	.w3(32'h3a85728c),
	.w4(32'h3973a267),
	.w5(32'hb7b56f0d),
	.w6(32'h39f7f3ae),
	.w7(32'hb9f4ee15),
	.w8(32'hba6109d5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed112a),
	.w1(32'h3a20fb04),
	.w2(32'h3a95b263),
	.w3(32'h3ae35942),
	.w4(32'h3a25a3bd),
	.w5(32'h3ab735c9),
	.w6(32'h3a679bc5),
	.w7(32'h38bd9159),
	.w8(32'h39ee0d2c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a33ca),
	.w1(32'h38cf2249),
	.w2(32'h3a452361),
	.w3(32'h3a8134ac),
	.w4(32'hb90f4a30),
	.w5(32'h3a24997b),
	.w6(32'h3a0cab37),
	.w7(32'hb9f28cf7),
	.w8(32'h39fec54f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c6c3a),
	.w1(32'h38991cae),
	.w2(32'h3a641033),
	.w3(32'h3a1f4c19),
	.w4(32'hb9bb43a8),
	.w5(32'h377b15c7),
	.w6(32'hb99f83c6),
	.w7(32'hba72b741),
	.w8(32'hb802ccbd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1e4dc),
	.w1(32'hb7994f71),
	.w2(32'h37b25b42),
	.w3(32'h3a87b06b),
	.w4(32'hb9139111),
	.w5(32'h3a307525),
	.w6(32'h3985f5e1),
	.w7(32'hba1af179),
	.w8(32'h38f8acb1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a830b28),
	.w1(32'hb9e5e13e),
	.w2(32'hb9e99f37),
	.w3(32'h3a91eec1),
	.w4(32'hb959f574),
	.w5(32'hba1e601b),
	.w6(32'h3a065c6a),
	.w7(32'hba761cfb),
	.w8(32'hba74642d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac90bcf),
	.w1(32'h3a9aab13),
	.w2(32'h3af23401),
	.w3(32'h3ae0e548),
	.w4(32'h3a65b4e7),
	.w5(32'h3ab22331),
	.w6(32'h3a1efced),
	.w7(32'h39dee029),
	.w8(32'h3a9b7cf6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00ef0b),
	.w1(32'hb83acdd9),
	.w2(32'h38be5590),
	.w3(32'h39ccedd5),
	.w4(32'hb8f39eb0),
	.w5(32'hb6c939b7),
	.w6(32'h39b053b2),
	.w7(32'hb900fe6f),
	.w8(32'h36bcc0a6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdbf5f),
	.w1(32'hba6f2f76),
	.w2(32'h3b0ecdb8),
	.w3(32'h3b2d84f1),
	.w4(32'hba798967),
	.w5(32'h3afabcbe),
	.w6(32'h3aabeaf8),
	.w7(32'hbae65f8c),
	.w8(32'h3ac55ba9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959a408),
	.w1(32'hb9b4f520),
	.w2(32'h38dc73f7),
	.w3(32'h3a009937),
	.w4(32'hb9a0b9d4),
	.w5(32'hb99c87e7),
	.w6(32'h39cd3d03),
	.w7(32'hba2292a2),
	.w8(32'hb9bd8169),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e81973),
	.w1(32'hb7a02a3c),
	.w2(32'h376ba0da),
	.w3(32'h3808cadb),
	.w4(32'h3715ffe3),
	.w5(32'h38059243),
	.w6(32'h37522bf7),
	.w7(32'h367ac6e3),
	.w8(32'h35488db4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb590ee1f),
	.w1(32'hb794dfe7),
	.w2(32'h36fc6b2b),
	.w3(32'h37703fbb),
	.w4(32'hb5c252d3),
	.w5(32'h37afc746),
	.w6(32'h3629b57c),
	.w7(32'h37170fd5),
	.w8(32'h3837ce6d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d6a72),
	.w1(32'h385c5a0a),
	.w2(32'h38522795),
	.w3(32'h3a58c81f),
	.w4(32'h38d7ae1b),
	.w5(32'hb8ca501e),
	.w6(32'h39ba5cb1),
	.w7(32'h39161f44),
	.w8(32'hb6b678ac),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cfe49),
	.w1(32'h39ca1bb0),
	.w2(32'h3ae236d8),
	.w3(32'h3a96b2b5),
	.w4(32'hb8a6e3d4),
	.w5(32'h3aee31db),
	.w6(32'h3962d666),
	.w7(32'hba443d05),
	.w8(32'h3a7fb503),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b146ae5),
	.w1(32'h39797710),
	.w2(32'h3a2db61d),
	.w3(32'h3b23912a),
	.w4(32'h38bb8c8b),
	.w5(32'h3a16a63e),
	.w6(32'h3b022ba9),
	.w7(32'h399fb73e),
	.w8(32'h3a74146e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35418fd1),
	.w1(32'hb7a9823c),
	.w2(32'h3736369e),
	.w3(32'h36a3cbb8),
	.w4(32'hb4943144),
	.w5(32'h37ab817e),
	.w6(32'hb7c63d53),
	.w7(32'h380419df),
	.w8(32'h36f33987),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b162e9e),
	.w1(32'h3ab14158),
	.w2(32'h3b056d08),
	.w3(32'h3b1e06fd),
	.w4(32'h3a8146a7),
	.w5(32'h3ab64150),
	.w6(32'h3af8aecf),
	.w7(32'h3a25040a),
	.w8(32'h3a94c073),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3d17d),
	.w1(32'h3a8e16e8),
	.w2(32'h3afcffa8),
	.w3(32'h3ad43c75),
	.w4(32'h3a8f8e7a),
	.w5(32'h3aab2af8),
	.w6(32'h3a40ca12),
	.w7(32'h3a53f24f),
	.w8(32'h3aa01d33),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae73bbc),
	.w1(32'h3b00128b),
	.w2(32'h3b0ea099),
	.w3(32'h3ace0ec9),
	.w4(32'h3ab8b2cf),
	.w5(32'h3b039887),
	.w6(32'h39315f93),
	.w7(32'h3a63dc4f),
	.w8(32'h3a954a73),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a127a37),
	.w1(32'hbaae8eb5),
	.w2(32'h3a84167f),
	.w3(32'h3a824c2d),
	.w4(32'hbaf031de),
	.w5(32'h3a18147f),
	.w6(32'h39f23820),
	.w7(32'hbb2522da),
	.w8(32'hb9ba4784),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba207189),
	.w1(32'hbabff1cf),
	.w2(32'hba109b92),
	.w3(32'hba2c340e),
	.w4(32'hba98a8ff),
	.w5(32'hba15cb79),
	.w6(32'hb99eb99e),
	.w7(32'hbaaa40ab),
	.w8(32'hb8f1da6a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d6d11),
	.w1(32'hba6a0ec9),
	.w2(32'hb9a71ef1),
	.w3(32'hbaa133d7),
	.w4(32'hbabc8caa),
	.w5(32'hba8e6d9a),
	.w6(32'hba9f3464),
	.w7(32'hbaad44eb),
	.w8(32'hba908cc3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd69b1),
	.w1(32'h397458a6),
	.w2(32'h3a0b5512),
	.w3(32'h3b112b43),
	.w4(32'h393004b0),
	.w5(32'h3a284270),
	.w6(32'h3aea5fc6),
	.w7(32'hb9902c82),
	.w8(32'h39df983f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42e0a2),
	.w1(32'hbaeb2d19),
	.w2(32'hb88446e6),
	.w3(32'h3a0caebd),
	.w4(32'hbafabac1),
	.w5(32'hb906b0ee),
	.w6(32'h398c9c8b),
	.w7(32'hbaf4f1a0),
	.w8(32'hb9a4b270),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb67f3),
	.w1(32'hba95cde2),
	.w2(32'hba1cc82e),
	.w3(32'h3a35d84a),
	.w4(32'hba86da35),
	.w5(32'hba0d5033),
	.w6(32'h3a20a879),
	.w7(32'hba9b4db7),
	.w8(32'hba29ff4c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a89331),
	.w1(32'h383ef0f4),
	.w2(32'hb8e6c3e8),
	.w3(32'h39e61885),
	.w4(32'h3988a490),
	.w5(32'h391bfe94),
	.w6(32'h39213006),
	.w7(32'h3846358a),
	.w8(32'hb88269d5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383ad14d),
	.w1(32'h370a0e46),
	.w2(32'h3890d135),
	.w3(32'h3711fdf4),
	.w4(32'hb70454a4),
	.w5(32'h382499b4),
	.w6(32'h3793d851),
	.w7(32'h3825ecca),
	.w8(32'h38de51a0),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8a38a),
	.w1(32'h3a8eee78),
	.w2(32'h3aca16bd),
	.w3(32'h3ab81640),
	.w4(32'h3a36cbbd),
	.w5(32'h3aa09979),
	.w6(32'h3a697d8d),
	.w7(32'h3a0c9c22),
	.w8(32'h3a45249e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386d3578),
	.w1(32'h382aeb46),
	.w2(32'h390be804),
	.w3(32'h38524d8e),
	.w4(32'h37b507e8),
	.w5(32'h3970f2b3),
	.w6(32'hb91fd763),
	.w7(32'h36f81f90),
	.w8(32'h3916a7b7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cc85b),
	.w1(32'hb9c5a7c7),
	.w2(32'h39ba2666),
	.w3(32'h3a992eed),
	.w4(32'h386a0f13),
	.w5(32'h372cfb89),
	.w6(32'h3a2de2c9),
	.w7(32'hba234b67),
	.w8(32'hb9ab45f3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9388cdc),
	.w1(32'hb9218d6c),
	.w2(32'hb927e2d3),
	.w3(32'hb8f82ba2),
	.w4(32'hb9662b51),
	.w5(32'hb8083a83),
	.w6(32'hb851c6b0),
	.w7(32'hb9413c3e),
	.w8(32'h38172f05),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac62cb0),
	.w1(32'h395e2a93),
	.w2(32'hb8a63d57),
	.w3(32'h3af34a81),
	.w4(32'h3a81d7b6),
	.w5(32'h39d222a3),
	.w6(32'h3a8e6718),
	.w7(32'h39d4cb9b),
	.w8(32'hb96b7246),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fde0af),
	.w1(32'hb9342557),
	.w2(32'hb95a6471),
	.w3(32'hb8f97deb),
	.w4(32'hb95b3b35),
	.w5(32'hb95aecd9),
	.w6(32'hb966454d),
	.w7(32'hb9ccb6bf),
	.w8(32'hb9bb0301),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb887f38a),
	.w1(32'hb8288e7d),
	.w2(32'hb9339b4a),
	.w3(32'hb9371a00),
	.w4(32'hb9045e70),
	.w5(32'hb92d77f6),
	.w6(32'hb8e87c44),
	.w7(32'hb89807f6),
	.w8(32'hb922b221),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39878442),
	.w1(32'h386f71fc),
	.w2(32'h3ad74542),
	.w3(32'h398b19de),
	.w4(32'hb94781fa),
	.w5(32'h3aad3007),
	.w6(32'hb98d98c7),
	.w7(32'hba0dd51a),
	.w8(32'h3a870d0f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8119ab),
	.w1(32'h3b3020a9),
	.w2(32'h3b7bb86b),
	.w3(32'h3ba245ab),
	.w4(32'h3b44a98a),
	.w5(32'h3b787350),
	.w6(32'h3b2f789a),
	.w7(32'h3a9676a7),
	.w8(32'h3a854662),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3937647e),
	.w1(32'hba80632b),
	.w2(32'hba8ecdb7),
	.w3(32'h398a3fda),
	.w4(32'hba298b76),
	.w5(32'hba3618d2),
	.w6(32'h39c3d008),
	.w7(32'hba7d0d66),
	.w8(32'hba906688),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a1c93),
	.w1(32'hb9a65516),
	.w2(32'h3a8d621f),
	.w3(32'h39abffd4),
	.w4(32'hba51eb73),
	.w5(32'h3a19e804),
	.w6(32'h3939bfb5),
	.w7(32'hba2b9af6),
	.w8(32'h39067907),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a6926),
	.w1(32'hb98d5a19),
	.w2(32'h399a5a84),
	.w3(32'h398d718a),
	.w4(32'hb996c777),
	.w5(32'h39004984),
	.w6(32'h391923f5),
	.w7(32'hb9ce665b),
	.w8(32'hb89dc910),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a8b50),
	.w1(32'h39a29eeb),
	.w2(32'h3ad913c1),
	.w3(32'h3b827963),
	.w4(32'h39845f14),
	.w5(32'h3af58212),
	.w6(32'h3b78a267),
	.w7(32'h39c8aa8e),
	.w8(32'h3ae6dbd9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf14b9),
	.w1(32'hb99742b7),
	.w2(32'h37e69d32),
	.w3(32'h3ac9e1c8),
	.w4(32'hb9ef5a29),
	.w5(32'hb95f2077),
	.w6(32'h3a86a8d9),
	.w7(32'hba7254e7),
	.w8(32'hba2a46fb),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cc27e),
	.w1(32'h3a745082),
	.w2(32'h3b066587),
	.w3(32'h3b0cb8b3),
	.w4(32'h3a8ec757),
	.w5(32'h3af6f752),
	.w6(32'h3ab989c3),
	.w7(32'h39ac3755),
	.w8(32'h3a8100a3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c28df7),
	.w1(32'hb9a3522b),
	.w2(32'h37cee28f),
	.w3(32'hb99bff63),
	.w4(32'hba0a2907),
	.w5(32'hb9bee863),
	.w6(32'hba12d8b8),
	.w7(32'hba2f13a8),
	.w8(32'hb9cd292e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a968169),
	.w1(32'h3a575b0f),
	.w2(32'h3ad90744),
	.w3(32'h3aac8cdf),
	.w4(32'h3a3ee3fb),
	.w5(32'h3a95b05d),
	.w6(32'h3a1aeb31),
	.w7(32'h3919b374),
	.w8(32'h39871f0f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c2da41),
	.w1(32'h3688ee15),
	.w2(32'h367dd1fa),
	.w3(32'hb78e2c7c),
	.w4(32'h3770fefd),
	.w5(32'h369d5494),
	.w6(32'hb7a8f85b),
	.w7(32'h377958b0),
	.w8(32'hb75526cf),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cc85c),
	.w1(32'h3a158ce4),
	.w2(32'h3a2f3c7c),
	.w3(32'h3a04820a),
	.w4(32'h39cd4aeb),
	.w5(32'h39d9961c),
	.w6(32'h39fc75b1),
	.w7(32'h39b3a1bb),
	.w8(32'h39966905),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982f100),
	.w1(32'hb914384e),
	.w2(32'h38733005),
	.w3(32'h3977681b),
	.w4(32'hb8664d71),
	.w5(32'h37950bff),
	.w6(32'h3925a8a2),
	.w7(32'hb926000f),
	.w8(32'h37a37951),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2d42d),
	.w1(32'h3874735d),
	.w2(32'h3a7fd0b3),
	.w3(32'h3afd442c),
	.w4(32'h39248aa9),
	.w5(32'h39d3416c),
	.w6(32'h3b031c6a),
	.w7(32'h39be9155),
	.w8(32'h3a11e976),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b2fe6b),
	.w1(32'hb524be62),
	.w2(32'h365502e4),
	.w3(32'h36a0581b),
	.w4(32'hb6d6fe2d),
	.w5(32'h36864c35),
	.w6(32'h370ac569),
	.w7(32'h37546d43),
	.w8(32'hb5e0e41b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ace3fe),
	.w1(32'hb867325a),
	.w2(32'h383dec68),
	.w3(32'hb82373b6),
	.w4(32'hb85a8b86),
	.w5(32'h37c1079a),
	.w6(32'hb8673d7e),
	.w7(32'h35d884c0),
	.w8(32'h387f1652),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d30f8),
	.w1(32'hba015a1b),
	.w2(32'hb9743c82),
	.w3(32'h3a2c99f3),
	.w4(32'hba0dab78),
	.w5(32'hba05f71d),
	.w6(32'h39abbf70),
	.w7(32'hba37b69b),
	.w8(32'hba11293a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c62842),
	.w1(32'hbaa2b986),
	.w2(32'hba1349d7),
	.w3(32'h3a2f6570),
	.w4(32'hba09ef3a),
	.w5(32'hb9b247b5),
	.w6(32'h39b9b8c1),
	.w7(32'hba337c22),
	.w8(32'hb9842afa),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a300dde),
	.w1(32'h3a319453),
	.w2(32'h38642886),
	.w3(32'h3a7357ef),
	.w4(32'h3998b1f5),
	.w5(32'h387b9d38),
	.w6(32'hb8fe3d72),
	.w7(32'hb99b1d30),
	.w8(32'h37cefb95),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968d618),
	.w1(32'hb9f0757f),
	.w2(32'hb9ca3a41),
	.w3(32'hb7f822d7),
	.w4(32'hb8c76e52),
	.w5(32'hb91e3096),
	.w6(32'hb88acb76),
	.w7(32'hb9b330e0),
	.w8(32'hb973ec77),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e8ee1),
	.w1(32'h3b1a49f2),
	.w2(32'h3b922534),
	.w3(32'h3b7df487),
	.w4(32'h3acecc45),
	.w5(32'h3b3fbff0),
	.w6(32'h3add4592),
	.w7(32'h3a0004d1),
	.w8(32'h3a636ec1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77d39d),
	.w1(32'hba5b9af5),
	.w2(32'h3a4358bd),
	.w3(32'h3b4ebf61),
	.w4(32'hbaca718d),
	.w5(32'hba0091b3),
	.w6(32'h3ad6aa54),
	.w7(32'hbb4954dd),
	.w8(32'hbabeeb79),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ff399),
	.w1(32'h3887ac95),
	.w2(32'h389cbc59),
	.w3(32'h38a83471),
	.w4(32'hb86ac5f1),
	.w5(32'h39152a0a),
	.w6(32'hb98cec69),
	.w7(32'hb90d8f55),
	.w8(32'h387a227f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37404baf),
	.w1(32'hb76f6459),
	.w2(32'hb8289173),
	.w3(32'h36234c88),
	.w4(32'h3686436b),
	.w5(32'hb8183dad),
	.w6(32'h36fe27b0),
	.w7(32'hb72ad5e3),
	.w8(32'h38896245),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb852a832),
	.w1(32'hb6d0281a),
	.w2(32'h3905d3fa),
	.w3(32'h376375ba),
	.w4(32'h37a23f02),
	.w5(32'hb74016ec),
	.w6(32'h38646f04),
	.w7(32'h39315b70),
	.w8(32'h392dc142),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1d36b),
	.w1(32'hb7795d01),
	.w2(32'hb7584337),
	.w3(32'hb824c4de),
	.w4(32'hb79dd0af),
	.w5(32'hb75e094e),
	.w6(32'hb7dcaaf2),
	.w7(32'h371254d1),
	.w8(32'h372116cd),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92cad6e),
	.w1(32'h39ad90b6),
	.w2(32'h3a5dc150),
	.w3(32'h38e2d6e1),
	.w4(32'h3a090bfe),
	.w5(32'h3a97a47d),
	.w6(32'hb94ed828),
	.w7(32'h3a06be0e),
	.w8(32'h3a8a897a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33add0),
	.w1(32'h3842aefc),
	.w2(32'h3a4f3948),
	.w3(32'h3a887425),
	.w4(32'hb9be5291),
	.w5(32'h39ae913b),
	.w6(32'h39992dae),
	.w7(32'hba374148),
	.w8(32'h3a1e4e8c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b461fb1),
	.w1(32'h3acaf3f6),
	.w2(32'h3b135c7a),
	.w3(32'h3b324f55),
	.w4(32'h3a8c5ec7),
	.w5(32'h3ad5525f),
	.w6(32'h3b022d48),
	.w7(32'h3a489952),
	.w8(32'h3a87302e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a563b95),
	.w1(32'h37798b33),
	.w2(32'hb86b0a3d),
	.w3(32'h3a8c42b6),
	.w4(32'h393edc56),
	.w5(32'hb80a1e0d),
	.w6(32'h39dc1b90),
	.w7(32'hb830da36),
	.w8(32'hb975fe4b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9b38),
	.w1(32'h39eec45b),
	.w2(32'h3a98a577),
	.w3(32'h3ad563fd),
	.w4(32'h3a442eaa),
	.w5(32'h3ab37933),
	.w6(32'h3abebb59),
	.w7(32'h3a54c4e8),
	.w8(32'h3ac71560),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7f0d2),
	.w1(32'h37578a6e),
	.w2(32'h38fe45ff),
	.w3(32'h39d052c4),
	.w4(32'h38d0c7ae),
	.w5(32'h388c3c8a),
	.w6(32'h390a839f),
	.w7(32'h382891bd),
	.w8(32'hb936e895),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7611621),
	.w1(32'hb751802d),
	.w2(32'h3679bdc6),
	.w3(32'hb78f6242),
	.w4(32'hb669f15b),
	.w5(32'h374cce81),
	.w6(32'hb7f72877),
	.w7(32'h36818663),
	.w8(32'hb613fc6a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d08dc2),
	.w1(32'h394761ed),
	.w2(32'hb91b0605),
	.w3(32'h39869423),
	.w4(32'hb7e07d89),
	.w5(32'hb99ddd75),
	.w6(32'h37dd2178),
	.w7(32'hb91fa1c4),
	.w8(32'hba0c2d0f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84aa60d),
	.w1(32'h3615353f),
	.w2(32'h3793eaa9),
	.w3(32'hb85ca08e),
	.w4(32'h36dfb82d),
	.w5(32'h37828437),
	.w6(32'hb88d72c0),
	.w7(32'h3769bb98),
	.w8(32'hb718e69b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adccda4),
	.w1(32'hb8f7eace),
	.w2(32'h3889e713),
	.w3(32'h3a9929a3),
	.w4(32'hb7bd3f28),
	.w5(32'hb9d4f8d6),
	.w6(32'h3a313129),
	.w7(32'hb977be6b),
	.w8(32'hb9cc7d37),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c464f),
	.w1(32'hb8a8e334),
	.w2(32'h39b23f0f),
	.w3(32'h3b0756cf),
	.w4(32'hba648bc8),
	.w5(32'hba3c6709),
	.w6(32'h3adc5035),
	.w7(32'hbaa69701),
	.w8(32'hba8bd30d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a574805),
	.w1(32'hb8aa0728),
	.w2(32'h3a159fed),
	.w3(32'h3a1c1b0b),
	.w4(32'hb9eb02ae),
	.w5(32'h39347743),
	.w6(32'h391185b1),
	.w7(32'hba5a7c0a),
	.w8(32'hb9096ce3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4f365),
	.w1(32'hba778fa2),
	.w2(32'hbaa16e5e),
	.w3(32'hb99a833f),
	.w4(32'hba41d366),
	.w5(32'hba7ce749),
	.w6(32'hb99f907c),
	.w7(32'hba49bcfe),
	.w8(32'hba6ea64c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0a5b5),
	.w1(32'hb98f58b6),
	.w2(32'h3a9a5062),
	.w3(32'h3ab64bff),
	.w4(32'hba179a5d),
	.w5(32'h3a2f47c1),
	.w6(32'h3a2f097e),
	.w7(32'hba6ee0ac),
	.w8(32'h396b8b26),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ae8b),
	.w1(32'h3a1fe17d),
	.w2(32'h3aa75b2d),
	.w3(32'h3aa44023),
	.w4(32'h39eafca6),
	.w5(32'h3a4b2c8b),
	.w6(32'h3a4b5ac0),
	.w7(32'h39f79ccf),
	.w8(32'h3a3c75f4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90228f),
	.w1(32'h3a516e6a),
	.w2(32'h3a986f26),
	.w3(32'h3ba80968),
	.w4(32'h3a84abf8),
	.w5(32'h3ab12f92),
	.w6(32'h3b7175b5),
	.w7(32'h3a777e45),
	.w8(32'h3a85623a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a3bc2),
	.w1(32'h37dd4727),
	.w2(32'h37622bb0),
	.w3(32'h38c4a380),
	.w4(32'h3758b16e),
	.w5(32'hb6061ec8),
	.w6(32'h35292c08),
	.w7(32'hb5572db0),
	.w8(32'h36d25deb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816cab8),
	.w1(32'hb8b33b66),
	.w2(32'hb7c02651),
	.w3(32'hb6178d6f),
	.w4(32'hb7a2b58f),
	.w5(32'h375d4e28),
	.w6(32'hb70a4100),
	.w7(32'hb7a6f731),
	.w8(32'h37373b6c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea6b33),
	.w1(32'hb8bc6c99),
	.w2(32'h398f20ef),
	.w3(32'h3ae90284),
	.w4(32'h394b004b),
	.w5(32'h39a036aa),
	.w6(32'h3a85aa6f),
	.w7(32'hb9fbdc7f),
	.w8(32'hb9aae076),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3707ea),
	.w1(32'h3aaa55de),
	.w2(32'h3b2694f9),
	.w3(32'h3b3cce2e),
	.w4(32'h3aabceb5),
	.w5(32'h3b0ba032),
	.w6(32'h3ae232e5),
	.w7(32'hb788df40),
	.w8(32'h398d4b2c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2370c2),
	.w1(32'h3aae4a44),
	.w2(32'h3b020c0d),
	.w3(32'h3b18482e),
	.w4(32'h3a24b646),
	.w5(32'h3a8a700f),
	.w6(32'h3aa831d2),
	.w7(32'hb9573f2d),
	.w8(32'h3a20be72),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982c1d3),
	.w1(32'h38dc90cf),
	.w2(32'hb970a215),
	.w3(32'h3aa213c5),
	.w4(32'h3a6686bf),
	.w5(32'h3a0bb92d),
	.w6(32'hb9e69119),
	.w7(32'h388f57a5),
	.w8(32'h39690b36),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38972906),
	.w1(32'h377069a2),
	.w2(32'h388a0455),
	.w3(32'h388c5bb5),
	.w4(32'h389d9626),
	.w5(32'h384d22e4),
	.w6(32'h382cc121),
	.w7(32'h38bf1acb),
	.w8(32'h37bd16b0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395fa7bb),
	.w1(32'h399b68d8),
	.w2(32'h394cc1ea),
	.w3(32'h39a0c194),
	.w4(32'h39c774b3),
	.w5(32'h396c384d),
	.w6(32'h39c07f3e),
	.w7(32'h3998b8dd),
	.w8(32'h38ed73f9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52e924),
	.w1(32'h3a0f9511),
	.w2(32'h3a3aef4e),
	.w3(32'h3a891cd2),
	.w4(32'h3aa69ba9),
	.w5(32'h3ae61063),
	.w6(32'hb99ac2a9),
	.w7(32'h3a029a8b),
	.w8(32'h3a824608),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a1d7d),
	.w1(32'h3b05bcd3),
	.w2(32'h3aa19fe4),
	.w3(32'h3b61e31b),
	.w4(32'h3ae267ff),
	.w5(32'h3b084cb7),
	.w6(32'h3b446127),
	.w7(32'h3aa1f693),
	.w8(32'h3a7ad5ec),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a1765),
	.w1(32'h3a3d2105),
	.w2(32'h3a4e23fe),
	.w3(32'h3a875d62),
	.w4(32'h3a7e9ad6),
	.w5(32'h3a99d49f),
	.w6(32'hb8cd714a),
	.w7(32'h39c61a04),
	.w8(32'h39b7faa2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a283f60),
	.w1(32'hbab3f4f7),
	.w2(32'hba15d4b9),
	.w3(32'h3a86f5dc),
	.w4(32'hbaa415b6),
	.w5(32'hb9ef93c8),
	.w6(32'h3a37bbbb),
	.w7(32'hbacaf3ba),
	.w8(32'hba15f45a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e8c58),
	.w1(32'h39800c77),
	.w2(32'h3ad67778),
	.w3(32'h3aef7fc7),
	.w4(32'hba2dc8d8),
	.w5(32'h39e3b73e),
	.w6(32'h3a683bc3),
	.w7(32'hbabbe234),
	.w8(32'hba05c7db),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384d028d),
	.w1(32'hb636b4ee),
	.w2(32'hb7179d14),
	.w3(32'h3871c846),
	.w4(32'hb7229723),
	.w5(32'hb734280a),
	.w6(32'hb753f09c),
	.w7(32'hb77be6c3),
	.w8(32'hb723e10c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35cfd595),
	.w1(32'h36813a1c),
	.w2(32'h36a4f39c),
	.w3(32'hb448aa2c),
	.w4(32'h372517b2),
	.w5(32'h379535a6),
	.w6(32'hb74d0ac1),
	.w7(32'hb6845c58),
	.w8(32'hb6ce49c5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7f169),
	.w1(32'hb96ca6cc),
	.w2(32'hb84e10a3),
	.w3(32'hb8d33680),
	.w4(32'hb8977575),
	.w5(32'h394e1353),
	.w6(32'hb98414f9),
	.w7(32'h3733c218),
	.w8(32'h38b82648),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ef1fb8),
	.w1(32'hb7e15ade),
	.w2(32'hb788795d),
	.w3(32'h38303143),
	.w4(32'hb7963bab),
	.w5(32'hb769a6a9),
	.w6(32'hb8568a0b),
	.w7(32'hb68efc26),
	.w8(32'h37b1f1f2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ad87b),
	.w1(32'h37c7b09d),
	.w2(32'hb7d10223),
	.w3(32'h39140c20),
	.w4(32'h3868c229),
	.w5(32'h392ef506),
	.w6(32'h3911e992),
	.w7(32'h385084d0),
	.w8(32'h392f0d9f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9d5c),
	.w1(32'h3a62b10f),
	.w2(32'h3b1aff81),
	.w3(32'h3b061fca),
	.w4(32'h3ab4745e),
	.w5(32'h3af52977),
	.w6(32'h3a925704),
	.w7(32'h3a09ef00),
	.w8(32'h3aa321dd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dac80),
	.w1(32'h39f2f575),
	.w2(32'h3a87b28d),
	.w3(32'h3ae5e4b3),
	.w4(32'h3a283878),
	.w5(32'h3a87e8f4),
	.w6(32'h3a3eeb3e),
	.w7(32'h39a8d471),
	.w8(32'h3a32c64a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e53f5c),
	.w1(32'hb7f6639f),
	.w2(32'hb7f419ca),
	.w3(32'h380c569b),
	.w4(32'hb811a25f),
	.w5(32'hb830992d),
	.w6(32'h366d9d13),
	.w7(32'hb7b3e21b),
	.w8(32'hb863d0cf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d65a5),
	.w1(32'h3ad04406),
	.w2(32'h3a8ddd8f),
	.w3(32'h3b04c8be),
	.w4(32'h3ac44bf6),
	.w5(32'h3af0517e),
	.w6(32'h39f88209),
	.w7(32'h3a254fc9),
	.w8(32'h3a85db00),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9674ac),
	.w1(32'h3a37809a),
	.w2(32'h3a10ac9b),
	.w3(32'h3a7fb96e),
	.w4(32'h3a11570d),
	.w5(32'h39f16f48),
	.w6(32'h3a256e09),
	.w7(32'h39cb4266),
	.w8(32'h39263b75),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bfa31a),
	.w1(32'h391ffb10),
	.w2(32'h38f86e28),
	.w3(32'hb8869dbf),
	.w4(32'h39078acf),
	.w5(32'h392b0e87),
	.w6(32'hb8e888a6),
	.w7(32'h38b4d2a8),
	.w8(32'h390ea19d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7500d),
	.w1(32'hb8cf3a7c),
	.w2(32'hb980ff44),
	.w3(32'h39ebdf4e),
	.w4(32'h3900b143),
	.w5(32'h388f0315),
	.w6(32'h3987a4d2),
	.w7(32'h37a7106d),
	.w8(32'hb892e1a9),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f45d5),
	.w1(32'hb8f452b5),
	.w2(32'hb84340b4),
	.w3(32'hb9336662),
	.w4(32'hb91ac056),
	.w5(32'hb8e84d77),
	.w6(32'hb92269e1),
	.w7(32'hb9007b32),
	.w8(32'hb870c3ac),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376145f3),
	.w1(32'hb8989383),
	.w2(32'hb89fd3d3),
	.w3(32'h3961bd80),
	.w4(32'h3971a47c),
	.w5(32'h38c7a75f),
	.w6(32'h3903a45e),
	.w7(32'h38ebaf31),
	.w8(32'hb7953035),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d84188),
	.w1(32'hb8127ab3),
	.w2(32'hb78445d6),
	.w3(32'hb499dc83),
	.w4(32'hb64a8b32),
	.w5(32'hb6ca85bd),
	.w6(32'hb7989a55),
	.w7(32'h378ad284),
	.w8(32'hb6a71a6d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0375e),
	.w1(32'hb5f59ea9),
	.w2(32'hb720f65f),
	.w3(32'hb7c73f3c),
	.w4(32'hb77ed711),
	.w5(32'hb7249cf2),
	.w6(32'hb7b00735),
	.w7(32'hb7abc153),
	.w8(32'h36259865),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aea9d8),
	.w1(32'hba6a0816),
	.w2(32'hba2a6878),
	.w3(32'h3937d878),
	.w4(32'hb9e0eda6),
	.w5(32'hb45c1c7c),
	.w6(32'h39c17cdd),
	.w7(32'hba000f34),
	.w8(32'h3887beda),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ed311),
	.w1(32'h3a8af915),
	.w2(32'h3b239dc5),
	.w3(32'h3b0fa3e2),
	.w4(32'h3a41a217),
	.w5(32'h3ae26599),
	.w6(32'h3a99f98d),
	.w7(32'h390ea321),
	.w8(32'h3a5fb852),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac99960),
	.w1(32'h3a200843),
	.w2(32'h3a80f23c),
	.w3(32'h3a84d525),
	.w4(32'hb79c43ee),
	.w5(32'h3a20b317),
	.w6(32'h39a2ded5),
	.w7(32'hba006896),
	.w8(32'hb7dd7a6e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a648d),
	.w1(32'h3ac161be),
	.w2(32'h3b179d41),
	.w3(32'h3b254d5a),
	.w4(32'h3aab2730),
	.w5(32'h3b0aaa1c),
	.w6(32'h3ac35517),
	.w7(32'h3a8aab03),
	.w8(32'h3a914be5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809af47),
	.w1(32'hb85007be),
	.w2(32'hb959354b),
	.w3(32'h38983741),
	.w4(32'h3817885a),
	.w5(32'hb8a2b6a6),
	.w6(32'h36ff09d0),
	.w7(32'hb7912893),
	.w8(32'hb908c5bf),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e9a9b),
	.w1(32'h38349ef9),
	.w2(32'h36c5e146),
	.w3(32'h3858d699),
	.w4(32'h3849b24c),
	.w5(32'hb7acc3b5),
	.w6(32'h37a65803),
	.w7(32'h387b3d04),
	.w8(32'hb88835b1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83c6757),
	.w1(32'hb7bacf43),
	.w2(32'h36c8c63d),
	.w3(32'hb7b70d4f),
	.w4(32'hb672fb95),
	.w5(32'h3756acdc),
	.w6(32'h37460f5c),
	.w7(32'h378d77c2),
	.w8(32'h37fa4b53),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cda47c),
	.w1(32'h364b4b3f),
	.w2(32'h3644df3c),
	.w3(32'hb70b3e5b),
	.w4(32'h378a3024),
	.w5(32'h3710751d),
	.w6(32'h3793a603),
	.w7(32'h38011de9),
	.w8(32'hb77dbc64),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acab6d1),
	.w1(32'h3a250e3f),
	.w2(32'h3ab38939),
	.w3(32'h3a88c624),
	.w4(32'h39e3bef3),
	.w5(32'h3a7e44ff),
	.w6(32'h3a67dce6),
	.w7(32'h358582b4),
	.w8(32'h38c9c179),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b191af),
	.w1(32'h394c83a4),
	.w2(32'h39aca464),
	.w3(32'h3976e5e4),
	.w4(32'h39d58e98),
	.w5(32'h39d1d972),
	.w6(32'h39e87461),
	.w7(32'h3a1379f4),
	.w8(32'h39fe67e8),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79b44bc),
	.w1(32'hb9cd752d),
	.w2(32'hba7f23c7),
	.w3(32'hb6c50733),
	.w4(32'hb95496c2),
	.w5(32'hba7d577c),
	.w6(32'hb9ce54e9),
	.w7(32'hba112b7e),
	.w8(32'hba922c28),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2c360),
	.w1(32'hb9e10743),
	.w2(32'hb9dd5fe8),
	.w3(32'h3995645a),
	.w4(32'hb96bdaef),
	.w5(32'hb9d99f0b),
	.w6(32'h393fcef1),
	.w7(32'hb9dd79e7),
	.w8(32'hba1504fc),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88106b9),
	.w1(32'h3802b54f),
	.w2(32'h38004800),
	.w3(32'hb84d2905),
	.w4(32'h38106abd),
	.w5(32'h373023d6),
	.w6(32'hb708c98f),
	.w7(32'h388facbb),
	.w8(32'h37c48ba9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19c3cd),
	.w1(32'h399d3142),
	.w2(32'h393ac762),
	.w3(32'h3a20b29f),
	.w4(32'h39aee4b4),
	.w5(32'h39bf6123),
	.w6(32'h395c71c9),
	.w7(32'h3982e9e9),
	.w8(32'h3981539f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900993c),
	.w1(32'h38c85ff8),
	.w2(32'h386f553a),
	.w3(32'h38bcef04),
	.w4(32'h38aa7ff9),
	.w5(32'h3715df71),
	.w6(32'h387ea50d),
	.w7(32'h38b6de89),
	.w8(32'hb8471fb5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a790478),
	.w1(32'hba09bc66),
	.w2(32'h3a3b83cf),
	.w3(32'h3a6545b0),
	.w4(32'hb95ae4a1),
	.w5(32'hb79cdfaa),
	.w6(32'h3a4e8468),
	.w7(32'hba7e3d85),
	.w8(32'hbaacf56c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37678cd5),
	.w1(32'hb99988b8),
	.w2(32'hbbd2f12a),
	.w3(32'hb70a8e8f),
	.w4(32'h3a2aca5a),
	.w5(32'hbbee5ad2),
	.w6(32'hba4eee2d),
	.w7(32'hbbfde320),
	.w8(32'hbaeb46d7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84bf6a),
	.w1(32'h3aef48f2),
	.w2(32'h3adbaded),
	.w3(32'hba49eed9),
	.w4(32'h3b4836b0),
	.w5(32'hb8a69653),
	.w6(32'h3ba17b40),
	.w7(32'h3b22045a),
	.w8(32'hbad8a182),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule