module layer_10_featuremap_212(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae20e00),
	.w1(32'hbbd6d03a),
	.w2(32'hba82f7cf),
	.w3(32'h3a41b477),
	.w4(32'hbb0a0604),
	.w5(32'h3a653bdc),
	.w6(32'hbb0245f5),
	.w7(32'hb9a0a543),
	.w8(32'h3a071c4c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64a2d3),
	.w1(32'hba98f286),
	.w2(32'hbaab8fff),
	.w3(32'hb7b346ed),
	.w4(32'h3a7b9e34),
	.w5(32'h39dae998),
	.w6(32'hba9be603),
	.w7(32'h38cbd388),
	.w8(32'hbabf7b89),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae22ca7),
	.w1(32'h37f86a94),
	.w2(32'h3b39384f),
	.w3(32'h3ade7e0e),
	.w4(32'h3898e522),
	.w5(32'h399c0471),
	.w6(32'hba933dc2),
	.w7(32'hb9a0cd90),
	.w8(32'h3a9d3f00),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25611a),
	.w1(32'hba9f3718),
	.w2(32'h3bf2797a),
	.w3(32'h3b1b4cb9),
	.w4(32'hbb4b204a),
	.w5(32'h3a85b778),
	.w6(32'h3b1b62fd),
	.w7(32'h3bef8a1a),
	.w8(32'h3b676ee4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f48d35),
	.w1(32'hbacee7ca),
	.w2(32'hbab799e1),
	.w3(32'hbb0ed51c),
	.w4(32'hba0aa6c3),
	.w5(32'h3b4467a0),
	.w6(32'hbb845d31),
	.w7(32'hbb0d79ba),
	.w8(32'hbb4321ed),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadba59),
	.w1(32'hbb0b1819),
	.w2(32'h3a3ed281),
	.w3(32'h3a345b97),
	.w4(32'hba5ae1e7),
	.w5(32'h3ab75b7e),
	.w6(32'hbb441aa0),
	.w7(32'hbac8d665),
	.w8(32'hba3656ff),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d72d9),
	.w1(32'hb9ab8605),
	.w2(32'hbaa02627),
	.w3(32'h3b914967),
	.w4(32'hbb04cad2),
	.w5(32'hbaea9202),
	.w6(32'h39169e7a),
	.w7(32'hb8970ccd),
	.w8(32'hba5ab151),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4fa0b),
	.w1(32'hbbe48198),
	.w2(32'hbbc8c753),
	.w3(32'hbbb3583b),
	.w4(32'hbb8c2d6a),
	.w5(32'hba7035b2),
	.w6(32'hbc0f49db),
	.w7(32'hbb2d32ce),
	.w8(32'h3ae0fc35),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dcf0b),
	.w1(32'hbb08ff1e),
	.w2(32'h3a6eb7a3),
	.w3(32'hba5dcc23),
	.w4(32'hbb21bac3),
	.w5(32'h3a53506e),
	.w6(32'hbb4d7f22),
	.w7(32'hbadfa710),
	.w8(32'hba8f38ea),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ceae3),
	.w1(32'hbbc79ed7),
	.w2(32'hbbb63dde),
	.w3(32'hbb1c771f),
	.w4(32'hbbcb42ec),
	.w5(32'hbbc2acfb),
	.w6(32'hbbf128a1),
	.w7(32'hbbaae58a),
	.w8(32'hbc0597e2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1abeb4),
	.w1(32'hbba9dc00),
	.w2(32'hbb9a27b9),
	.w3(32'h39c2a206),
	.w4(32'hbb08be83),
	.w5(32'h390d0540),
	.w6(32'hbaeed654),
	.w7(32'hbb5815a0),
	.w8(32'hbaecad4f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60ce0),
	.w1(32'hb90e882c),
	.w2(32'hbb4fd8a9),
	.w3(32'h3c519e41),
	.w4(32'h3b6b4fb0),
	.w5(32'h3b600063),
	.w6(32'h39479989),
	.w7(32'hbadde698),
	.w8(32'h3b297a18),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a008d87),
	.w1(32'hbae93662),
	.w2(32'hbb8524a7),
	.w3(32'h3b9c3efb),
	.w4(32'hba889c54),
	.w5(32'hbab3e747),
	.w6(32'hbb634d79),
	.w7(32'hbb27c00e),
	.w8(32'hbb5b7842),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd5135),
	.w1(32'hba440afe),
	.w2(32'hbab97cd0),
	.w3(32'h3a659d16),
	.w4(32'h3a8a80f9),
	.w5(32'hb9abb351),
	.w6(32'h391fb16f),
	.w7(32'hb9f39ee5),
	.w8(32'hb8438489),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a28cb),
	.w1(32'hbadcec54),
	.w2(32'hbbe66336),
	.w3(32'h3b1918a7),
	.w4(32'hb885a382),
	.w5(32'h3ae0e16c),
	.w6(32'h383a58db),
	.w7(32'h3ae36e08),
	.w8(32'h3912c434),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7802d4),
	.w1(32'hbbfc7cb8),
	.w2(32'hbb994783),
	.w3(32'hbab86ad0),
	.w4(32'hbba3bb33),
	.w5(32'hbb3180ac),
	.w6(32'hbbf2f2ec),
	.w7(32'hbb8cc864),
	.w8(32'hbb8c89e5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7cf4c),
	.w1(32'hbb13cf64),
	.w2(32'h3b29ffa3),
	.w3(32'h3b11f923),
	.w4(32'h3abe52a1),
	.w5(32'hba575cb8),
	.w6(32'hbc2d147f),
	.w7(32'hbbbe0389),
	.w8(32'hbbed2551),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32bc64),
	.w1(32'hbb9ed031),
	.w2(32'h3a287407),
	.w3(32'hbc3d2e52),
	.w4(32'hbb618b77),
	.w5(32'hba804961),
	.w6(32'hbbd9df93),
	.w7(32'hbb24ffa1),
	.w8(32'hbaec1579),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cccf9),
	.w1(32'hbac35fdd),
	.w2(32'h3a6018cf),
	.w3(32'hbae3f8a8),
	.w4(32'hbab530f7),
	.w5(32'h37c3055a),
	.w6(32'hbb25bcca),
	.w7(32'hba918d3f),
	.w8(32'hba80e442),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89fd5f),
	.w1(32'hba5025d7),
	.w2(32'h3af9996f),
	.w3(32'h3ab11aa1),
	.w4(32'hba86b457),
	.w5(32'h3b023e36),
	.w6(32'hba4f8b90),
	.w7(32'h3a22fc6d),
	.w8(32'h3aae1f1f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920d364),
	.w1(32'h39a80e11),
	.w2(32'h3b036f18),
	.w3(32'h3acbef64),
	.w4(32'hbae4b2c8),
	.w5(32'hb826464c),
	.w6(32'hbaf70ee7),
	.w7(32'h39f905f6),
	.w8(32'h3a56b348),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9a70c),
	.w1(32'hba83c743),
	.w2(32'h3b210bf3),
	.w3(32'hbae3a4a7),
	.w4(32'hbc1b9589),
	.w5(32'hbc173842),
	.w6(32'h3b53aa36),
	.w7(32'h3b9dee08),
	.w8(32'h3bf71196),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba115f26),
	.w1(32'h3bfee348),
	.w2(32'h3bea3c23),
	.w3(32'hbb8c7a21),
	.w4(32'hbb7ef25e),
	.w5(32'hbbacd1c9),
	.w6(32'hbc83755b),
	.w7(32'hbc2ba6f7),
	.w8(32'hbc75f175),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933055),
	.w1(32'hbb3b6d1a),
	.w2(32'hbbd20ca4),
	.w3(32'hbc541cc1),
	.w4(32'hba9cb4f6),
	.w5(32'hbb5fd4bb),
	.w6(32'hbb4fde90),
	.w7(32'hbad9523d),
	.w8(32'hbb9dfd5d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae554e),
	.w1(32'hb898b3da),
	.w2(32'hbb49ab05),
	.w3(32'hba70ff2a),
	.w4(32'hb9c864a6),
	.w5(32'hbb827e3f),
	.w6(32'hbb2b3ae9),
	.w7(32'hbb3e063f),
	.w8(32'hbbce91ed),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39619c44),
	.w1(32'hba0207f4),
	.w2(32'h3b1a99e8),
	.w3(32'hb952d47f),
	.w4(32'hbb7ffb86),
	.w5(32'hbb8cdedc),
	.w6(32'hbc14d0ca),
	.w7(32'hbba18d0c),
	.w8(32'hbb9324fd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa73ba2),
	.w1(32'hba34fb87),
	.w2(32'h3a792986),
	.w3(32'hbbb165ff),
	.w4(32'hba56c1e9),
	.w5(32'h3ae15184),
	.w6(32'hba8f89fd),
	.w7(32'h3a46cfdb),
	.w8(32'h3aaf4c51),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3489c0),
	.w1(32'hbb282673),
	.w2(32'hba655cf1),
	.w3(32'h3b78a24b),
	.w4(32'hbb9f398d),
	.w5(32'hbbafd611),
	.w6(32'h3abfb3b3),
	.w7(32'hbaa21679),
	.w8(32'hbac7147a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19db21),
	.w1(32'hb934c1b7),
	.w2(32'h3bb72d4c),
	.w3(32'hba64bf32),
	.w4(32'hbb0b3f21),
	.w5(32'h3b7b318e),
	.w6(32'hbba0af76),
	.w7(32'h3b91a947),
	.w8(32'hbb3b3764),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c12ad),
	.w1(32'hba6373ca),
	.w2(32'hbc469f7c),
	.w3(32'hbbeaeb18),
	.w4(32'h3b9aabf1),
	.w5(32'hbc3309b0),
	.w6(32'h3b14acc8),
	.w7(32'hbbfa7458),
	.w8(32'hbb7bdd4b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f06e0),
	.w1(32'hb99affc3),
	.w2(32'h3a065003),
	.w3(32'hbbb17d2d),
	.w4(32'hb977a0fc),
	.w5(32'h3a3cbee3),
	.w6(32'hba876d94),
	.w7(32'h3a10ff02),
	.w8(32'h3970f98c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc08ee),
	.w1(32'h3ab3f2ee),
	.w2(32'h3afc6c8a),
	.w3(32'hb9503c9a),
	.w4(32'h38215373),
	.w5(32'h3b0d924b),
	.w6(32'hba83f27e),
	.w7(32'h3a207faf),
	.w8(32'h3a5f6f7a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eaefc1),
	.w1(32'hbbd5bcf1),
	.w2(32'hba854ffa),
	.w3(32'h3a41104f),
	.w4(32'hbaee5cdb),
	.w5(32'h3a2ee754),
	.w6(32'hbb9fc084),
	.w7(32'h3a336981),
	.w8(32'h3b03c885),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396dca71),
	.w1(32'hbbe84cef),
	.w2(32'hbb46287e),
	.w3(32'h3b0ff4c4),
	.w4(32'hbc197b82),
	.w5(32'h3bf08756),
	.w6(32'hbc15e7c7),
	.w7(32'h3a8a4424),
	.w8(32'hbc2e859a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02da8a),
	.w1(32'hbb953a9c),
	.w2(32'hb94f8e1f),
	.w3(32'hba25d53e),
	.w4(32'hbba3bfef),
	.w5(32'hbaf83cc2),
	.w6(32'hbb9a3fe7),
	.w7(32'hbb50821f),
	.w8(32'hbb727f16),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13e5d6),
	.w1(32'h3a98a0f2),
	.w2(32'h3a488c72),
	.w3(32'hba428a42),
	.w4(32'h387db858),
	.w5(32'h3a3b5f45),
	.w6(32'hba60cbf0),
	.w7(32'h3acc320d),
	.w8(32'h3afb2f44),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaff5d6),
	.w1(32'hbb7d3257),
	.w2(32'hbc0182eb),
	.w3(32'hba214dbf),
	.w4(32'hb9efb4c5),
	.w5(32'hbb0b1cdb),
	.w6(32'hbba4129b),
	.w7(32'hbafdcd19),
	.w8(32'hbbc195d3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1d9aa),
	.w1(32'h3bcd9e27),
	.w2(32'h3bd8cec1),
	.w3(32'hbb808fa6),
	.w4(32'h3bba34ee),
	.w5(32'h3bbf65a5),
	.w6(32'hbaff3000),
	.w7(32'h3b5daa10),
	.w8(32'hba8692b3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8c13),
	.w1(32'h3bd22cf8),
	.w2(32'h3bb9589f),
	.w3(32'h3bc02850),
	.w4(32'h3910c79a),
	.w5(32'hb971f444),
	.w6(32'h3b4c0871),
	.w7(32'hba654ae1),
	.w8(32'hbbaab145),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e07b5),
	.w1(32'h3a6f9ed1),
	.w2(32'hb91f60b5),
	.w3(32'h3b1ee3c1),
	.w4(32'h3ab28fb5),
	.w5(32'h3a801316),
	.w6(32'hba6dadac),
	.w7(32'h38ea4308),
	.w8(32'hba67fb6f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a6535),
	.w1(32'h3b896ba4),
	.w2(32'hbc869d20),
	.w3(32'h3acb059d),
	.w4(32'h3c22644d),
	.w5(32'hbc5b05b3),
	.w6(32'h3c4e4e48),
	.w7(32'hbb1c00ef),
	.w8(32'h3be48ada),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75c8c6),
	.w1(32'hba8cd5b4),
	.w2(32'hba31280f),
	.w3(32'hbc40bbfb),
	.w4(32'hba4fc194),
	.w5(32'h3b0f1bb5),
	.w6(32'hb90675be),
	.w7(32'hb8fa9c7a),
	.w8(32'h39d933f9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00e161),
	.w1(32'hba40d786),
	.w2(32'hba13ab0a),
	.w3(32'h3b63f22d),
	.w4(32'hba75b4a0),
	.w5(32'h386fa951),
	.w6(32'hbb23c348),
	.w7(32'hbab23323),
	.w8(32'hba7da969),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad7d53),
	.w1(32'hbc103775),
	.w2(32'hbb960505),
	.w3(32'hbb0511ef),
	.w4(32'hbc00bad8),
	.w5(32'hbbf81a6c),
	.w6(32'hbbec789b),
	.w7(32'hbbf61460),
	.w8(32'hbc200107),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab3a59),
	.w1(32'hbb73ae46),
	.w2(32'hbb1684c7),
	.w3(32'hbb4111f7),
	.w4(32'hbb4b70c6),
	.w5(32'hbb9fcbf7),
	.w6(32'hbbb3c406),
	.w7(32'hbb2db8f3),
	.w8(32'hbb9d5148),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1870f),
	.w1(32'hbb356eaa),
	.w2(32'hbbe8daf5),
	.w3(32'hbb32daa5),
	.w4(32'hbbbaa28d),
	.w5(32'hbbf33230),
	.w6(32'hbbad6d1f),
	.w7(32'hbb277a3c),
	.w8(32'hbbe464f5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe154d9),
	.w1(32'hbbc466d6),
	.w2(32'hbc1ec44e),
	.w3(32'hbb8f4601),
	.w4(32'hbaea912f),
	.w5(32'hbb8e3c63),
	.w6(32'hbb505cb8),
	.w7(32'hb9c08a50),
	.w8(32'hbb8d6603),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba748625),
	.w1(32'hbb684bc6),
	.w2(32'h3bf3ed40),
	.w3(32'h3a198b9e),
	.w4(32'hbb993f75),
	.w5(32'h3c1e3606),
	.w6(32'hbc447c12),
	.w7(32'h38d7d861),
	.w8(32'hbc3f9efc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c35c9),
	.w1(32'hba24073a),
	.w2(32'hb9de0b08),
	.w3(32'hbb23b06a),
	.w4(32'hbaf2eece),
	.w5(32'hb914ee67),
	.w6(32'hba977970),
	.w7(32'hb9ab3990),
	.w8(32'hba61cba3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa332f9),
	.w1(32'hb9a1de31),
	.w2(32'hbb41d40a),
	.w3(32'h3a8a3cec),
	.w4(32'h3a281790),
	.w5(32'hbac1d5b7),
	.w6(32'hba3874a8),
	.w7(32'hbae4ad8e),
	.w8(32'hbb4abd66),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c66c7),
	.w1(32'h3ae12856),
	.w2(32'h3afe7314),
	.w3(32'h3b7fbedb),
	.w4(32'h3b05cf15),
	.w5(32'h3ac762c9),
	.w6(32'hb8078b4a),
	.w7(32'h3a3c7f75),
	.w8(32'h3a89960c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f3c0d6),
	.w1(32'hbb234008),
	.w2(32'hbb8838d7),
	.w3(32'hb9ec969d),
	.w4(32'hbbc46a35),
	.w5(32'hbb8cd1e8),
	.w6(32'hba8f99a0),
	.w7(32'hbb84f9e8),
	.w8(32'hbac116f4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9856ba9),
	.w1(32'h39a49677),
	.w2(32'h3aa693b7),
	.w3(32'h3b233a7a),
	.w4(32'hb9984694),
	.w5(32'hb9ed108f),
	.w6(32'hb9ad8f66),
	.w7(32'hb8241f2c),
	.w8(32'h3a77c8d7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf4dad),
	.w1(32'hbbd5e15b),
	.w2(32'hbbb19e0a),
	.w3(32'h3ac125ae),
	.w4(32'hbb8a05ab),
	.w5(32'hbab495d2),
	.w6(32'hbbb61644),
	.w7(32'hbaba3ec8),
	.w8(32'hb9b649f7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b4787),
	.w1(32'hbb2d09b4),
	.w2(32'hba8e439d),
	.w3(32'h3b107ac8),
	.w4(32'hbaa49b0c),
	.w5(32'hbb31087a),
	.w6(32'hbbbcdf98),
	.w7(32'hbb8baa28),
	.w8(32'hbb90b6bd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6fd0),
	.w1(32'h3afe7a1e),
	.w2(32'hbc5bcb8b),
	.w3(32'hbb6456f4),
	.w4(32'h3bf2f4f0),
	.w5(32'hbc4b7ce9),
	.w6(32'h3cb69461),
	.w7(32'h3bbe3387),
	.w8(32'h3c869776),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2b3c9),
	.w1(32'hba9d37e0),
	.w2(32'hbba9badc),
	.w3(32'hbc2423ce),
	.w4(32'hbabcfd15),
	.w5(32'hbbda0050),
	.w6(32'hbb1a6f58),
	.w7(32'hbb58672c),
	.w8(32'hbb06a89a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52b287),
	.w1(32'h3ae92339),
	.w2(32'hbb963cc6),
	.w3(32'hbb75576e),
	.w4(32'h3bc2fe27),
	.w5(32'h3b5c94e8),
	.w6(32'hbaa1bb5c),
	.w7(32'hba27d17b),
	.w8(32'hbadb31d2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25e5d4),
	.w1(32'h3aaf88b8),
	.w2(32'h3ae567c9),
	.w3(32'h3aa42396),
	.w4(32'h3a9dac7b),
	.w5(32'h3ab2f7ce),
	.w6(32'hba11405c),
	.w7(32'hb9a210f2),
	.w8(32'h3a23662f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28de84),
	.w1(32'hba1d4d86),
	.w2(32'h3882e106),
	.w3(32'h3b318ead),
	.w4(32'h38addde9),
	.w5(32'h3aa5e1a3),
	.w6(32'hb979f3d5),
	.w7(32'h399839be),
	.w8(32'hb96d3e41),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb220c54),
	.w1(32'hbb0a4f28),
	.w2(32'hbb05c98e),
	.w3(32'h3a83525f),
	.w4(32'h38e53437),
	.w5(32'hbb05ffe7),
	.w6(32'hbb4ae2a5),
	.w7(32'hbac1a47c),
	.w8(32'h38d572ab),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad75f7f),
	.w1(32'hbb1f1f33),
	.w2(32'hb920fe59),
	.w3(32'hbad349e2),
	.w4(32'hbab1cbee),
	.w5(32'hbb17365f),
	.w6(32'hba4a8af2),
	.w7(32'h3a9c019c),
	.w8(32'h3a750e1f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9514d78),
	.w1(32'hba05f922),
	.w2(32'h3b4223f1),
	.w3(32'hb8860425),
	.w4(32'h3ae4256d),
	.w5(32'h3b5037d8),
	.w6(32'hbadc4ace),
	.w7(32'hb9b8a136),
	.w8(32'h3b850d9c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad74151),
	.w1(32'hbb26655f),
	.w2(32'h3a7cd1c7),
	.w3(32'h39ce1ec9),
	.w4(32'hbb7c50fb),
	.w5(32'hbab50534),
	.w6(32'hbb218d0e),
	.w7(32'hbb6d2f21),
	.w8(32'hbb587622),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcafba),
	.w1(32'hbaf1b438),
	.w2(32'h39b8777a),
	.w3(32'h3931d9bc),
	.w4(32'hba914ce3),
	.w5(32'hb94597cc),
	.w6(32'hba7778a6),
	.w7(32'h3ae95360),
	.w8(32'h3a148b7b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9d765),
	.w1(32'h39eef7f9),
	.w2(32'hbb8c6460),
	.w3(32'hba979ffe),
	.w4(32'hba15c3a2),
	.w5(32'h390541e0),
	.w6(32'hbaad21a4),
	.w7(32'hb9e96b70),
	.w8(32'hbb8b2464),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc294ff9),
	.w1(32'h3c3d1cf6),
	.w2(32'hbb88a60d),
	.w3(32'hbb05785c),
	.w4(32'h3c9370eb),
	.w5(32'hbb177332),
	.w6(32'h3ca3cc79),
	.w7(32'h3bcb4156),
	.w8(32'h3be8384f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51f92c),
	.w1(32'h3c6ba22f),
	.w2(32'h3c2a3a7c),
	.w3(32'hbaf504ef),
	.w4(32'hbb056d76),
	.w5(32'hbb016e35),
	.w6(32'hbc0b4965),
	.w7(32'h3aaa1001),
	.w8(32'hbbe72e21),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa7d2d),
	.w1(32'hb9d4e986),
	.w2(32'hbadfd2fb),
	.w3(32'hbc48b00e),
	.w4(32'h3ab17441),
	.w5(32'hbb11fafc),
	.w6(32'hbb90fb79),
	.w7(32'hba913434),
	.w8(32'hbac4c97c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a153c77),
	.w1(32'hbb277d1a),
	.w2(32'hbbd40740),
	.w3(32'hba9a4093),
	.w4(32'hbb80750d),
	.w5(32'hbb632dc0),
	.w6(32'hbc053e6d),
	.w7(32'hbb929382),
	.w8(32'hbc28f128),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26989),
	.w1(32'hba5dc197),
	.w2(32'h3a74ead8),
	.w3(32'hbaad7c41),
	.w4(32'hbaa63c98),
	.w5(32'h3980f632),
	.w6(32'hba9da64d),
	.w7(32'hba60d989),
	.w8(32'hbb0008aa),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989706a),
	.w1(32'hb923efe1),
	.w2(32'hb9c3db1e),
	.w3(32'hb90045eb),
	.w4(32'h3a1db342),
	.w5(32'h39c41c71),
	.w6(32'hba3232cb),
	.w7(32'hb9615804),
	.w8(32'hba187804),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bc1df),
	.w1(32'hb9af329f),
	.w2(32'h3a15ac9c),
	.w3(32'h3a8503ca),
	.w4(32'h37ac27b3),
	.w5(32'h3aa95c3f),
	.w6(32'hb9a73221),
	.w7(32'h39362d41),
	.w8(32'hb9642b1e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66cba8),
	.w1(32'h3b3d6333),
	.w2(32'h3b89f1da),
	.w3(32'h3afc2245),
	.w4(32'h3a9147ac),
	.w5(32'h3b48c874),
	.w6(32'hbae07c98),
	.w7(32'h3b00829d),
	.w8(32'h3a532a71),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1d82a),
	.w1(32'hba032bad),
	.w2(32'hb79db85e),
	.w3(32'h3b141a32),
	.w4(32'hb91f106c),
	.w5(32'hb9d5051d),
	.w6(32'h38b099a9),
	.w7(32'hb9dbea43),
	.w8(32'hbac812a8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba265345),
	.w1(32'hbc0660c3),
	.w2(32'hbc29f32a),
	.w3(32'hba1c2ff2),
	.w4(32'hbbeb48b6),
	.w5(32'hbb68baba),
	.w6(32'hbb54b2f4),
	.w7(32'hbb95f58a),
	.w8(32'hba49625d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fd8b3),
	.w1(32'hbb60bbcf),
	.w2(32'hbb9111e1),
	.w3(32'hbb822304),
	.w4(32'hbb69087b),
	.w5(32'hbb544a2b),
	.w6(32'hbbbfd5a9),
	.w7(32'hbb884a9c),
	.w8(32'hbb6eeec9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac6433),
	.w1(32'hbb34bb46),
	.w2(32'hbac38b8a),
	.w3(32'hbb67e216),
	.w4(32'hbb218db5),
	.w5(32'hba8c4d86),
	.w6(32'hbb92ac73),
	.w7(32'hbb96d273),
	.w8(32'hbb4b8214),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28c5ec),
	.w1(32'hbbbdd0a6),
	.w2(32'h3a9c22d1),
	.w3(32'hba788ba0),
	.w4(32'hbbcb2e3a),
	.w5(32'hbb5c70e7),
	.w6(32'hbc670ca0),
	.w7(32'hbbcb7886),
	.w8(32'hbc19f242),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9db9e2),
	.w1(32'hbb1cb3e5),
	.w2(32'hba6cfdea),
	.w3(32'hbbe71d96),
	.w4(32'hbb4a27ee),
	.w5(32'hbaa9a158),
	.w6(32'hbb443ff0),
	.w7(32'h396c74f8),
	.w8(32'hbb305f47),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9335aa),
	.w1(32'h3c1c26d4),
	.w2(32'h3b048486),
	.w3(32'hbb616772),
	.w4(32'hba899c73),
	.w5(32'hbb4915bc),
	.w6(32'h3c154492),
	.w7(32'h3c3bb183),
	.w8(32'h3b485292),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8485d),
	.w1(32'hba9e1aa6),
	.w2(32'hbaec8c79),
	.w3(32'hbc6362cd),
	.w4(32'hbafe28d9),
	.w5(32'hbaec54fd),
	.w6(32'hbaac0706),
	.w7(32'hba16b97d),
	.w8(32'h3987bf1c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904394b),
	.w1(32'hba1842f8),
	.w2(32'hbac15db6),
	.w3(32'hba407938),
	.w4(32'h3a6160c3),
	.w5(32'hbae393f3),
	.w6(32'h3b564bc9),
	.w7(32'h3a6b18e7),
	.w8(32'h3b3dcf58),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6eef7),
	.w1(32'hb87e5067),
	.w2(32'hba08df86),
	.w3(32'hb7e7a6c6),
	.w4(32'h39b9837c),
	.w5(32'hba370323),
	.w6(32'h388a7c81),
	.w7(32'h3980369f),
	.w8(32'h3993df58),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a412f76),
	.w1(32'h3c8e6287),
	.w2(32'h3d05e3aa),
	.w3(32'h3aa710b4),
	.w4(32'hbbb9bab9),
	.w5(32'h3d020bed),
	.w6(32'hbc220a55),
	.w7(32'h3c53232a),
	.w8(32'hbc9d5863),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bfed5),
	.w1(32'h3b124f63),
	.w2(32'h3aa000b6),
	.w3(32'h3a19022d),
	.w4(32'h3afddfdb),
	.w5(32'hb842857e),
	.w6(32'h3b0ad89b),
	.w7(32'h3a06b371),
	.w8(32'h38f31a82),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba084896),
	.w1(32'hba90f9bc),
	.w2(32'hbb03d54d),
	.w3(32'hba6991e5),
	.w4(32'hba417440),
	.w5(32'hba64a8b2),
	.w6(32'hbb13cda7),
	.w7(32'hba8a7fb7),
	.w8(32'hbaff919e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6cb7b),
	.w1(32'h3977faf3),
	.w2(32'h3a8ffc90),
	.w3(32'hbad0a31f),
	.w4(32'hb8cc7651),
	.w5(32'h39fffb32),
	.w6(32'hbaa1719b),
	.w7(32'h3a0b1b77),
	.w8(32'hb8054d1d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47d29e),
	.w1(32'hbadbcd81),
	.w2(32'hbb0b1608),
	.w3(32'hbaa01691),
	.w4(32'hba19d394),
	.w5(32'hbb27819f),
	.w6(32'hbba2ae5e),
	.w7(32'hbb7c08bc),
	.w8(32'hbb7bba63),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35f8a0),
	.w1(32'hba8586aa),
	.w2(32'h3aa841d6),
	.w3(32'hbb26315c),
	.w4(32'hb9cdee49),
	.w5(32'h3a1606e3),
	.w6(32'hbbde84ff),
	.w7(32'hba4f95ed),
	.w8(32'hb964ec95),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adcfd6),
	.w1(32'h3bacb61f),
	.w2(32'h3bb063d4),
	.w3(32'hb92cb938),
	.w4(32'h3ab414cf),
	.w5(32'h3adffaec),
	.w6(32'h3b23e515),
	.w7(32'h3a6ea9a9),
	.w8(32'hbaa00a1b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e798c),
	.w1(32'hbb7c2bdd),
	.w2(32'hb9c0ac3c),
	.w3(32'h3ac8d65c),
	.w4(32'hbb65dbf6),
	.w5(32'hbb406315),
	.w6(32'hbbd0b705),
	.w7(32'hbbc4ad58),
	.w8(32'hbbdd5d40),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba69bb4),
	.w1(32'h3a26e0a2),
	.w2(32'hba303dcb),
	.w3(32'h3ac614dc),
	.w4(32'hbb015c7d),
	.w5(32'hbba0edbc),
	.w6(32'hba9b06f8),
	.w7(32'hbb141260),
	.w8(32'hbb48dd7d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51e04c),
	.w1(32'h3b9c9e08),
	.w2(32'hbbd21019),
	.w3(32'hbbbc342a),
	.w4(32'hbb90f1bd),
	.w5(32'hbc6bf9fb),
	.w6(32'h3b99fa90),
	.w7(32'h3b939ce3),
	.w8(32'h3b096faf),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8771d1),
	.w1(32'hba2d8833),
	.w2(32'hb9e3a947),
	.w3(32'hbc7b52fc),
	.w4(32'hb8eaba30),
	.w5(32'hbb0f0825),
	.w6(32'hb986c6fd),
	.w7(32'hb9986dfc),
	.w8(32'hbab2cacd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4288be),
	.w1(32'hbb8246f6),
	.w2(32'hbbb9b8c6),
	.w3(32'h3a25ee60),
	.w4(32'hbb43ce27),
	.w5(32'hbb87fa45),
	.w6(32'hbb952d77),
	.w7(32'hbb8b7bc8),
	.w8(32'hbb31bda7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cd6bd),
	.w1(32'h3b4ca76f),
	.w2(32'h3bd8321e),
	.w3(32'h39b8b3e2),
	.w4(32'hbae34a2a),
	.w5(32'h3c030c5b),
	.w6(32'hbc1ad6e8),
	.w7(32'hbb7c1101),
	.w8(32'hbc106732),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e8f3c),
	.w1(32'h3a9ed942),
	.w2(32'hbc4c6c75),
	.w3(32'hbc02df08),
	.w4(32'h3afa81df),
	.w5(32'hbc02121e),
	.w6(32'hbb3278b7),
	.w7(32'hbc007adb),
	.w8(32'hbc12eece),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd667a),
	.w1(32'h3ae89654),
	.w2(32'hba9c0ed7),
	.w3(32'h3b9d19fd),
	.w4(32'h3977ac0d),
	.w5(32'hbb07e740),
	.w6(32'hbb20ed37),
	.w7(32'hbb508991),
	.w8(32'hbbae4dea),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb494c2b),
	.w1(32'hbb4de270),
	.w2(32'hbb379ead),
	.w3(32'hbb306f56),
	.w4(32'hba65f8d4),
	.w5(32'hb9c90b58),
	.w6(32'hbb8bde82),
	.w7(32'hb8f2d9e3),
	.w8(32'hb9caae07),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad5276),
	.w1(32'h3b908697),
	.w2(32'hbc024679),
	.w3(32'hbbdca9b1),
	.w4(32'h3be3d4bb),
	.w5(32'h35671268),
	.w6(32'hbbd06eec),
	.w7(32'hbb2bcc95),
	.w8(32'hbb140146),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37958756),
	.w1(32'hbbe4e763),
	.w2(32'hbc749969),
	.w3(32'h3a902a07),
	.w4(32'hbbf127b3),
	.w5(32'hbc214829),
	.w6(32'hbb9f6df2),
	.w7(32'hbba97761),
	.w8(32'hbba96554),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade88c1),
	.w1(32'hbae16d58),
	.w2(32'hbb8124c7),
	.w3(32'hbba6ce15),
	.w4(32'hb91b341e),
	.w5(32'h38283762),
	.w6(32'hbb761167),
	.w7(32'hbb3829f7),
	.w8(32'hbbc66c59),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebb2cd),
	.w1(32'h389f59fa),
	.w2(32'hbb14b05d),
	.w3(32'hba036d5d),
	.w4(32'h3a3a0294),
	.w5(32'h3a013297),
	.w6(32'hbae29c56),
	.w7(32'hbacb4e2d),
	.w8(32'hbb3cb7e2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3829c),
	.w1(32'hbb5e19f6),
	.w2(32'hbbcbcc39),
	.w3(32'hbb1062b4),
	.w4(32'hbaac6d48),
	.w5(32'hb8b869fe),
	.w6(32'hbb4e35a7),
	.w7(32'hbb1bdd19),
	.w8(32'hbba75092),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cd9aa),
	.w1(32'hbb43f3c1),
	.w2(32'hbb515a8d),
	.w3(32'hba36aaba),
	.w4(32'hbb809c7f),
	.w5(32'hbb47738c),
	.w6(32'hb9e2b260),
	.w7(32'hbae7c3bc),
	.w8(32'hbaeedd4d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c79691),
	.w1(32'hba538fac),
	.w2(32'h3b13a53f),
	.w3(32'h395efe41),
	.w4(32'hbafe3d97),
	.w5(32'hbaaa08b3),
	.w6(32'hbaa74765),
	.w7(32'hba92723c),
	.w8(32'hba49555d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01885c),
	.w1(32'h3b188735),
	.w2(32'h3b42011b),
	.w3(32'hbb0c5521),
	.w4(32'h3aae2ec1),
	.w5(32'h3a8fd1c9),
	.w6(32'hba7fa6a8),
	.w7(32'h390bfc9b),
	.w8(32'hba34df59),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38488717),
	.w1(32'hbafe331a),
	.w2(32'hbb80a173),
	.w3(32'h3adbca74),
	.w4(32'hbb179061),
	.w5(32'hbba4a68d),
	.w6(32'hbb696c94),
	.w7(32'hbbce5c81),
	.w8(32'hbc0a48ac),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368ade10),
	.w1(32'h3935cea1),
	.w2(32'hbb2bd823),
	.w3(32'h3ac6398d),
	.w4(32'hbad88348),
	.w5(32'hbbb9e3d9),
	.w6(32'h390e50ee),
	.w7(32'hba5de686),
	.w8(32'hbb76e018),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b281fc0),
	.w1(32'hb914215d),
	.w2(32'hba1016c4),
	.w3(32'hbaa7d45e),
	.w4(32'hba7c6eeb),
	.w5(32'hba7accc4),
	.w6(32'hb950a078),
	.w7(32'hbab83bea),
	.w8(32'hbb8c8c1d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5a007),
	.w1(32'hbad862d4),
	.w2(32'hbb1e84e7),
	.w3(32'h3b104c44),
	.w4(32'hbab63f3e),
	.w5(32'h38ed3390),
	.w6(32'hb967f3d7),
	.w7(32'hba4f832a),
	.w8(32'h3a86de9a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5dd9a5),
	.w1(32'h3a626fd7),
	.w2(32'h3b5539f6),
	.w3(32'h3a14c31b),
	.w4(32'hba5652be),
	.w5(32'h3b03f55e),
	.w6(32'hbbb1a9f3),
	.w7(32'hbab4c834),
	.w8(32'hb9fdb6fd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5f0f0),
	.w1(32'hbbc4585d),
	.w2(32'hbba1a661),
	.w3(32'hbaf03a95),
	.w4(32'hbba024c9),
	.w5(32'hbb6b006b),
	.w6(32'hbb81434d),
	.w7(32'hbae1ff56),
	.w8(32'hba1532c9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd541),
	.w1(32'hbb7ac9d5),
	.w2(32'hbb8559c8),
	.w3(32'h38ed73da),
	.w4(32'hbb91b5ae),
	.w5(32'hbbc91d0f),
	.w6(32'hbb8c653b),
	.w7(32'hbbad876c),
	.w8(32'hbbde2185),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69c6c0),
	.w1(32'hbae29c96),
	.w2(32'hba1e531c),
	.w3(32'hbb93ae06),
	.w4(32'hbb08fe5c),
	.w5(32'hba6c282f),
	.w6(32'hbb0adb8d),
	.w7(32'hbb50ff87),
	.w8(32'hbb88fa48),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ef0b2),
	.w1(32'hbab3aec0),
	.w2(32'hbad6b5ba),
	.w3(32'hbaad1bfc),
	.w4(32'hba5a3a2f),
	.w5(32'hba08bb26),
	.w6(32'hbabe8c41),
	.w7(32'hbabba8e2),
	.w8(32'hbb11646c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbb8cf),
	.w1(32'hbace206a),
	.w2(32'hbab18d15),
	.w3(32'hb94c1a4d),
	.w4(32'hbab3d41d),
	.w5(32'hba301d4b),
	.w6(32'hbad6f834),
	.w7(32'hbb019e41),
	.w8(32'hbb499d36),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e2982),
	.w1(32'h3ae41b2e),
	.w2(32'h3acd8a8a),
	.w3(32'hba79bf34),
	.w4(32'hb8b403a5),
	.w5(32'hba25c3dd),
	.w6(32'h3b36c1a3),
	.w7(32'h3b1a44e7),
	.w8(32'h3b6642df),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a6342),
	.w1(32'hb9384b63),
	.w2(32'h3ae6b40f),
	.w3(32'h3af45e73),
	.w4(32'h3942b4de),
	.w5(32'h3ac7f68f),
	.w6(32'hbb2ea40d),
	.w7(32'h3b62b62f),
	.w8(32'hbbbf8257),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74470),
	.w1(32'hb736ee40),
	.w2(32'h3acfb832),
	.w3(32'hbb3b78ab),
	.w4(32'hba86de9e),
	.w5(32'h3ad8bc91),
	.w6(32'hbb3eca7f),
	.w7(32'h39f96259),
	.w8(32'hbac01272),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac72750),
	.w1(32'hbae04094),
	.w2(32'h390b5f05),
	.w3(32'h386fc870),
	.w4(32'hbb202709),
	.w5(32'hb9614b1e),
	.w6(32'hbb25d027),
	.w7(32'hba99edf0),
	.w8(32'hbaee1411),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b34d6),
	.w1(32'hbb087045),
	.w2(32'hbb2f99fe),
	.w3(32'hbaf828b4),
	.w4(32'hbaa3cec2),
	.w5(32'hba9b46c7),
	.w6(32'hbb676423),
	.w7(32'hbb642f1c),
	.w8(32'hbbab8c6e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14acfc),
	.w1(32'hbbb5567f),
	.w2(32'hbba5fcb1),
	.w3(32'h3b00920d),
	.w4(32'hb9993075),
	.w5(32'hbb0d4550),
	.w6(32'hbb58f98d),
	.w7(32'h3ad0f581),
	.w8(32'h3a05c1a7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4402af),
	.w1(32'h3957e97a),
	.w2(32'h3b5962e6),
	.w3(32'hbaa16213),
	.w4(32'hba6c0315),
	.w5(32'h39e160d3),
	.w6(32'hbaf5f3ff),
	.w7(32'hb94063d6),
	.w8(32'hbaa3398d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1ba53),
	.w1(32'h3af0beb9),
	.w2(32'h3bbeef4d),
	.w3(32'hba7396c1),
	.w4(32'h38f17ba2),
	.w5(32'h3b87f40a),
	.w6(32'hb9671a4a),
	.w7(32'h3b880cfb),
	.w8(32'h3a6a470b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa13777),
	.w1(32'hb991e511),
	.w2(32'hba17a82a),
	.w3(32'h39884520),
	.w4(32'hb7f21632),
	.w5(32'hb8f54512),
	.w6(32'hb93f0fb0),
	.w7(32'hba093aae),
	.w8(32'hb93478d8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b742139),
	.w1(32'hb9f64db8),
	.w2(32'hbb29686b),
	.w3(32'h3a879092),
	.w4(32'hbb67240e),
	.w5(32'hbba89c15),
	.w6(32'hbb67f6d4),
	.w7(32'hbb4694f4),
	.w8(32'hbae60ee2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c2ea4),
	.w1(32'hbb6522e9),
	.w2(32'hbba03ea6),
	.w3(32'hb94759c6),
	.w4(32'hbb02603d),
	.w5(32'hbb6dc9eb),
	.w6(32'hba1715d6),
	.w7(32'hbaac0b30),
	.w8(32'hbb33d50c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32ff3a),
	.w1(32'h3950fd1c),
	.w2(32'h39a2284c),
	.w3(32'h391e90fd),
	.w4(32'h39a49efb),
	.w5(32'h39f40fa5),
	.w6(32'h391f8515),
	.w7(32'h39399c0a),
	.w8(32'h39aa9d50),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba23d4),
	.w1(32'hba5fd154),
	.w2(32'hbace674f),
	.w3(32'hbaa305b1),
	.w4(32'hb94a9923),
	.w5(32'hb9e0fa50),
	.w6(32'hbacba279),
	.w7(32'hba0e91d3),
	.w8(32'h38adb05b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39729166),
	.w1(32'hb982f7d1),
	.w2(32'hba1cd3bc),
	.w3(32'h3913eb03),
	.w4(32'h390a6f6a),
	.w5(32'h38f94797),
	.w6(32'hba03bc80),
	.w7(32'hb9bc5225),
	.w8(32'hba9da8a3),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf4ec),
	.w1(32'hba600a64),
	.w2(32'hbad86a54),
	.w3(32'hba68cb01),
	.w4(32'hb841e1bf),
	.w5(32'hba93b5c5),
	.w6(32'hbabe4f51),
	.w7(32'hba03190e),
	.w8(32'hba488a32),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11dfcb),
	.w1(32'hbb0807ba),
	.w2(32'hbb0b9b1c),
	.w3(32'hbaca21eb),
	.w4(32'hb90fc4cf),
	.w5(32'hba15b672),
	.w6(32'hb9851ada),
	.w7(32'h397e2235),
	.w8(32'hb98976ba),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba464953),
	.w1(32'hbb33331f),
	.w2(32'hbb81dc4c),
	.w3(32'h38a0a72c),
	.w4(32'hbaa0a5d6),
	.w5(32'hbb5f260e),
	.w6(32'hbb05a9ca),
	.w7(32'hbb4981da),
	.w8(32'hbb3d09ea),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6b6b5),
	.w1(32'hba12fa8f),
	.w2(32'hbaf96ff8),
	.w3(32'hba1ffc88),
	.w4(32'hb9b12a22),
	.w5(32'hbabbcda6),
	.w6(32'hba8bce54),
	.w7(32'hba8f2c70),
	.w8(32'hbb30aedc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1a980),
	.w1(32'hb9bb6f2b),
	.w2(32'hbb351d17),
	.w3(32'h39972e22),
	.w4(32'h38e8fed3),
	.w5(32'hba5fb0b5),
	.w6(32'hbaaff8b0),
	.w7(32'h39b12227),
	.w8(32'hbabd2c5a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b63df),
	.w1(32'hba9ff520),
	.w2(32'hbac9a473),
	.w3(32'h38b0955b),
	.w4(32'h39ae6863),
	.w5(32'hba9553b7),
	.w6(32'hbacfa314),
	.w7(32'hba9d79fe),
	.w8(32'hb7aa275b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b50a7),
	.w1(32'h3a0139c0),
	.w2(32'h38a47c2c),
	.w3(32'hbab21193),
	.w4(32'h38ce7a37),
	.w5(32'h3a8ba0a2),
	.w6(32'hbb5a954b),
	.w7(32'hba6bc629),
	.w8(32'hbaae1337),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba512906),
	.w1(32'hbb579f4b),
	.w2(32'hbbb24638),
	.w3(32'h391c25bd),
	.w4(32'hbb116ae3),
	.w5(32'hbb813a83),
	.w6(32'hbae284ff),
	.w7(32'hbb133923),
	.w8(32'hbb6a7ae5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a63366),
	.w1(32'hb995c8db),
	.w2(32'hba113adf),
	.w3(32'hba076dd2),
	.w4(32'hb8647b10),
	.w5(32'hb9b67ded),
	.w6(32'hba7800df),
	.w7(32'hb9e97a24),
	.w8(32'hba34290d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b001822),
	.w1(32'hba6c76c4),
	.w2(32'hbacf9ff7),
	.w3(32'h39b8b4e6),
	.w4(32'hbb1e4b58),
	.w5(32'hbb842534),
	.w6(32'h3a27ef1c),
	.w7(32'hbb484f4a),
	.w8(32'hbbc9613d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a651d6f),
	.w1(32'h3a10a72a),
	.w2(32'hb988ff67),
	.w3(32'h3a8eaac1),
	.w4(32'h3ab788e9),
	.w5(32'h3a21cfb9),
	.w6(32'hb9a4ddfd),
	.w7(32'hb95ca458),
	.w8(32'hb937c510),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb73a2),
	.w1(32'h39537e9a),
	.w2(32'h37ac16be),
	.w3(32'hb9069038),
	.w4(32'h396fa50e),
	.w5(32'h38722917),
	.w6(32'h394ae239),
	.w7(32'h3942a434),
	.w8(32'h39c73995),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989bbec),
	.w1(32'h39ed3d2c),
	.w2(32'h3a1b7bbb),
	.w3(32'h39fa1035),
	.w4(32'h38c0241c),
	.w5(32'h39e9bc26),
	.w6(32'h39b12b03),
	.w7(32'h3a0e903a),
	.w8(32'h39fd12ab),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67a3f3),
	.w1(32'hb98a91e8),
	.w2(32'hba248695),
	.w3(32'hb95d9cee),
	.w4(32'h389a7700),
	.w5(32'hb9c6a79c),
	.w6(32'hb99b581b),
	.w7(32'hba144c55),
	.w8(32'hba101be3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b7378),
	.w1(32'hb8d0cd6e),
	.w2(32'hbad959e3),
	.w3(32'h3a66d414),
	.w4(32'h3b026af7),
	.w5(32'hb922cfad),
	.w6(32'hb92757bf),
	.w7(32'h39af22f6),
	.w8(32'hbb4cbdd7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e55d8),
	.w1(32'hba279885),
	.w2(32'hba728837),
	.w3(32'hbaa2b46a),
	.w4(32'hb9b4bf45),
	.w5(32'hbac17a31),
	.w6(32'hbb4661d5),
	.w7(32'hbac73739),
	.w8(32'hbad36ac0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380b7041),
	.w1(32'h39acbec3),
	.w2(32'h392afd64),
	.w3(32'h39623b3f),
	.w4(32'h39a4623c),
	.w5(32'h39cabaf7),
	.w6(32'h399a4872),
	.w7(32'h394fcc82),
	.w8(32'h3a4777b4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d1971),
	.w1(32'hbb401471),
	.w2(32'hbbba379e),
	.w3(32'h38da7a76),
	.w4(32'hba86d1ee),
	.w5(32'hbb3506fb),
	.w6(32'hbb788d41),
	.w7(32'hbb813f5c),
	.w8(32'hbba1bb96),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117658),
	.w1(32'hba0ecf21),
	.w2(32'hbb828b29),
	.w3(32'h3b121457),
	.w4(32'hbabf248b),
	.w5(32'hbb929f78),
	.w6(32'hb8fff7a6),
	.w7(32'hbb1674b7),
	.w8(32'hbba34427),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3421e0),
	.w1(32'hbb89e1e7),
	.w2(32'hbbba47e3),
	.w3(32'hbae31574),
	.w4(32'hbb1e9e6a),
	.w5(32'hbb268958),
	.w6(32'hbb9be6ea),
	.w7(32'hbb876c8c),
	.w8(32'hbb5cfb36),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac51099),
	.w1(32'h390c50d6),
	.w2(32'hb8ec5ec5),
	.w3(32'h3a712082),
	.w4(32'hb9c00176),
	.w5(32'hbab2d14c),
	.w6(32'h3a9d8cfb),
	.w7(32'hb9fa07ac),
	.w8(32'hbb7b76eb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7db13),
	.w1(32'h3b0d99a0),
	.w2(32'h3a288af5),
	.w3(32'h3b00b05a),
	.w4(32'h3abfd0af),
	.w5(32'hb9885837),
	.w6(32'h39dc25a5),
	.w7(32'h3978b0b0),
	.w8(32'hbaafac43),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af022d0),
	.w1(32'h3a329687),
	.w2(32'hbaa2e4fc),
	.w3(32'h3b4daedd),
	.w4(32'h3b8f90cf),
	.w5(32'h3ae0198d),
	.w6(32'h3b25db04),
	.w7(32'h3adf2219),
	.w8(32'h3a2b650f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf79ad3),
	.w1(32'hba8d7bd4),
	.w2(32'hbb409dbe),
	.w3(32'hbad4b488),
	.w4(32'hba1f9b80),
	.w5(32'hbb0e403e),
	.w6(32'hbaee12e0),
	.w7(32'h3974db9c),
	.w8(32'hbb22a5fd),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d7535),
	.w1(32'h3b26255f),
	.w2(32'h3a315eb0),
	.w3(32'h384ba4ba),
	.w4(32'h3b406e71),
	.w5(32'h3aa1aa0c),
	.w6(32'h3a668804),
	.w7(32'h3b1a606c),
	.w8(32'hb9b45524),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c523e1),
	.w1(32'h3b010584),
	.w2(32'h3b02b946),
	.w3(32'hb932190c),
	.w4(32'h3a859152),
	.w5(32'h3acf9d69),
	.w6(32'h38f86761),
	.w7(32'h3a6c05e7),
	.w8(32'h39f00424),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba005d67),
	.w1(32'h38aced6e),
	.w2(32'h37547031),
	.w3(32'hb8ad3d51),
	.w4(32'hb903e725),
	.w5(32'h3986e57c),
	.w6(32'hba3140cb),
	.w7(32'hb9c620fc),
	.w8(32'h38bb3b0e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905b433),
	.w1(32'hb9053947),
	.w2(32'hb995fd9c),
	.w3(32'h39795cfc),
	.w4(32'h38e62de2),
	.w5(32'hb83e0214),
	.w6(32'hb9457165),
	.w7(32'hb96fc950),
	.w8(32'hb83ef0cf),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aab0cd),
	.w1(32'hbafb2238),
	.w2(32'hbb6b9682),
	.w3(32'h3980e02a),
	.w4(32'hba934e0b),
	.w5(32'hbb1467a2),
	.w6(32'hbaba4f7a),
	.w7(32'hbafe72e9),
	.w8(32'hbb054015),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe9b98),
	.w1(32'h3a465263),
	.w2(32'h37b42d76),
	.w3(32'h3a3f6d7a),
	.w4(32'h3a780c51),
	.w5(32'h38d882b8),
	.w6(32'h3a7629ab),
	.w7(32'h39549b80),
	.w8(32'hb8e17e5d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898de71),
	.w1(32'hb7a60987),
	.w2(32'hb9940116),
	.w3(32'hbaa35574),
	.w4(32'hbaace2aa),
	.w5(32'hba8f4744),
	.w6(32'hba184ae8),
	.w7(32'h3799158b),
	.w8(32'h3875ec3c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4e020),
	.w1(32'h39d890d5),
	.w2(32'h38ce3685),
	.w3(32'h3a77d2e8),
	.w4(32'h3a2eb21a),
	.w5(32'h39bd333e),
	.w6(32'h3940c6a8),
	.w7(32'h3a97d90d),
	.w8(32'h3a86a2ba),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e1b52),
	.w1(32'h390cb06c),
	.w2(32'h3a474d78),
	.w3(32'hb98a0b0e),
	.w4(32'hbaad4eb1),
	.w5(32'hba627c56),
	.w6(32'hba1b51d9),
	.w7(32'hbad28594),
	.w8(32'hb9eba406),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f43538),
	.w1(32'h39ee0211),
	.w2(32'h3a212ff7),
	.w3(32'h39f24a05),
	.w4(32'h3a37e03f),
	.w5(32'h3a6683de),
	.w6(32'h3a2ba389),
	.w7(32'h3a575633),
	.w8(32'h3a5831ad),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a345697),
	.w1(32'h3877dc18),
	.w2(32'hb93d0529),
	.w3(32'h3a8bb688),
	.w4(32'h397a8f0b),
	.w5(32'h35b5c299),
	.w6(32'h39534bac),
	.w7(32'h361e8383),
	.w8(32'h390f61b2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba633676),
	.w1(32'hb85e73d6),
	.w2(32'hbb2d70e4),
	.w3(32'hb8e049fe),
	.w4(32'h3a75433d),
	.w5(32'hba798ffa),
	.w6(32'h370dbd4f),
	.w7(32'hb8858a33),
	.w8(32'hbb124fa6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8ee4b),
	.w1(32'hb9597bda),
	.w2(32'hbb7554a8),
	.w3(32'hbb25fd68),
	.w4(32'hba8194fd),
	.w5(32'hbba82c81),
	.w6(32'hbb90936e),
	.w7(32'hba88d7dd),
	.w8(32'hbb4d75b8),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f1384),
	.w1(32'h3ad52b74),
	.w2(32'h3a8d2456),
	.w3(32'h3a69bf36),
	.w4(32'h3a4b0b42),
	.w5(32'h3a38d42c),
	.w6(32'h3ac08365),
	.w7(32'h3aacea3b),
	.w8(32'h3ab1c7c9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69fa66),
	.w1(32'h38c4417e),
	.w2(32'hba161e42),
	.w3(32'h3a441aa5),
	.w4(32'h3abfe437),
	.w5(32'hb981de19),
	.w6(32'hb9a3f4a7),
	.w7(32'hb847a6d4),
	.w8(32'hbae23d45),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b5d38),
	.w1(32'h3a24c48e),
	.w2(32'h3901fc7b),
	.w3(32'h3aa10c67),
	.w4(32'h3a362f06),
	.w5(32'hba2cef94),
	.w6(32'h3abe7a2c),
	.w7(32'h3a3ffa75),
	.w8(32'h38445775),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86207d),
	.w1(32'hbb76f8a5),
	.w2(32'hbb661205),
	.w3(32'hbb5fc9cb),
	.w4(32'hbaecc65e),
	.w5(32'hbb3566cb),
	.w6(32'hbb7e6df2),
	.w7(32'hba950782),
	.w8(32'hbb285406),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba7e2b),
	.w1(32'hbab6aa2c),
	.w2(32'hbb79ddfe),
	.w3(32'hb9875150),
	.w4(32'hba0c70ed),
	.w5(32'hbaf8124b),
	.w6(32'hbb13fa5d),
	.w7(32'hba69d3cb),
	.w8(32'hbad9a06b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fff9d),
	.w1(32'hbb67e371),
	.w2(32'hbbafeba9),
	.w3(32'hbaae557e),
	.w4(32'hbacd1943),
	.w5(32'hbb7251f4),
	.w6(32'hbb54c2f3),
	.w7(32'hbb0c5c2a),
	.w8(32'hbb586cd4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a994ccb),
	.w1(32'h3a8c005b),
	.w2(32'h3944fced),
	.w3(32'h3a3f824b),
	.w4(32'h3ad5c11b),
	.w5(32'h3a8dee13),
	.w6(32'h3ad824e3),
	.w7(32'h3b1f8f0e),
	.w8(32'h3a9fdedf),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a3b9),
	.w1(32'hbb26aa7e),
	.w2(32'hbb42e585),
	.w3(32'hbac593ca),
	.w4(32'hba2e6e6a),
	.w5(32'hbaa1d030),
	.w6(32'hba9dd0bd),
	.w7(32'hb9cb684e),
	.w8(32'hba09d669),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3f1e6),
	.w1(32'hb85cf1e4),
	.w2(32'h38213d85),
	.w3(32'h3a070fb8),
	.w4(32'hb9053894),
	.w5(32'hb8750f5f),
	.w6(32'hb8dc8929),
	.w7(32'hb8ae4c65),
	.w8(32'hb8863f64),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45259b),
	.w1(32'hb9b7b456),
	.w2(32'h3991906b),
	.w3(32'hb9e9fa44),
	.w4(32'hb906737b),
	.w5(32'h39c4ed39),
	.w6(32'hba5b3574),
	.w7(32'hba209030),
	.w8(32'h39350d79),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caed3f),
	.w1(32'h3a0f40c3),
	.w2(32'hb819e1db),
	.w3(32'h390f6672),
	.w4(32'h382e0a39),
	.w5(32'hb9e52ea4),
	.w6(32'h39fbb7a7),
	.w7(32'hb8030eec),
	.w8(32'hba5e71db),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f424f),
	.w1(32'hbb6fde9d),
	.w2(32'hbb71ff46),
	.w3(32'hbb78a498),
	.w4(32'hbb259b55),
	.w5(32'hbb2488ad),
	.w6(32'hbb603b80),
	.w7(32'hbb1f50f4),
	.w8(32'hbb2c9fae),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f51e75),
	.w1(32'hba066d17),
	.w2(32'h398f48f1),
	.w3(32'h3a268947),
	.w4(32'hba10d0da),
	.w5(32'hb927aaa1),
	.w6(32'hba02fc20),
	.w7(32'hb9375c89),
	.w8(32'hb46b160f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb803a3be),
	.w1(32'h39a643d1),
	.w2(32'h3a125a80),
	.w3(32'h390e1b2b),
	.w4(32'h39f75edc),
	.w5(32'h3a0507e8),
	.w6(32'h39fc5120),
	.w7(32'h3a3bdcd3),
	.w8(32'h3a0f1aa0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fe17b),
	.w1(32'h3a540dce),
	.w2(32'h3a825325),
	.w3(32'h399f78d0),
	.w4(32'h3954aac8),
	.w5(32'h3a2c34e7),
	.w6(32'hb9f89d58),
	.w7(32'hb981c728),
	.w8(32'hbaae2e3a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94871e3),
	.w1(32'h38bf265d),
	.w2(32'hbb2e4ed8),
	.w3(32'h391a3403),
	.w4(32'hba2690ae),
	.w5(32'hbb01dd1a),
	.w6(32'hba9a1832),
	.w7(32'hbaaf90ae),
	.w8(32'hbb6aecd3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043161),
	.w1(32'hba693825),
	.w2(32'hba30f9cd),
	.w3(32'hba222b73),
	.w4(32'h38cac0c9),
	.w5(32'h39fd4b23),
	.w6(32'hb9893955),
	.w7(32'hba5ca6bd),
	.w8(32'hba150cf8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb838ba2b),
	.w1(32'h3a2b52bc),
	.w2(32'h3a88c4a7),
	.w3(32'hb877d823),
	.w4(32'h3a1f192f),
	.w5(32'h3a4c797a),
	.w6(32'h3a02be23),
	.w7(32'h3a2faeaf),
	.w8(32'h3a830840),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60dd71),
	.w1(32'hbbae775b),
	.w2(32'hbc116273),
	.w3(32'hb85be249),
	.w4(32'hbab7a1b0),
	.w5(32'hbbe6e07b),
	.w6(32'hbb866107),
	.w7(32'hba648739),
	.w8(32'hbae63ea2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4561c7),
	.w1(32'hb9bc5dad),
	.w2(32'hbaaaaee5),
	.w3(32'hb96e28a2),
	.w4(32'h3acd83a8),
	.w5(32'hba67a8b5),
	.w6(32'h3a4de5e7),
	.w7(32'h3ab9a4a7),
	.w8(32'hbb9d27ec),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f896c),
	.w1(32'hb947e33f),
	.w2(32'hba947cdb),
	.w3(32'h3af1b6b6),
	.w4(32'h3948aa28),
	.w5(32'hba53fd88),
	.w6(32'h3a10d1c4),
	.w7(32'hb9061d64),
	.w8(32'hba06c104),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d3a1e0),
	.w1(32'h3a676340),
	.w2(32'h3a5e6c2e),
	.w3(32'h390031c8),
	.w4(32'h3a5ddac6),
	.w5(32'h39655790),
	.w6(32'h39efff3a),
	.w7(32'h39b15467),
	.w8(32'hb62ebb38),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22e08e),
	.w1(32'h39f6c664),
	.w2(32'hb82838d7),
	.w3(32'h397ad5b5),
	.w4(32'h3a4b6e75),
	.w5(32'h39246039),
	.w6(32'h3a2d1f8a),
	.w7(32'h39042ab5),
	.w8(32'h38b93e6f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d51d35),
	.w1(32'h38da3e79),
	.w2(32'h3919de28),
	.w3(32'h39b6819a),
	.w4(32'h38f3d145),
	.w5(32'h38f8a5c6),
	.w6(32'h38d82eea),
	.w7(32'hb8ad4e00),
	.w8(32'h3883a242),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1da9f4),
	.w1(32'h3a73eaa4),
	.w2(32'hbaadd408),
	.w3(32'h3b0413df),
	.w4(32'h389e0792),
	.w5(32'hbab83652),
	.w6(32'h39ab71e0),
	.w7(32'hba0fb3bb),
	.w8(32'hba3317b4),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7244a5),
	.w1(32'h3a5e398f),
	.w2(32'hbabf4bd0),
	.w3(32'h3b224050),
	.w4(32'h3a32b5db),
	.w5(32'hba0e4656),
	.w6(32'hba64cb2e),
	.w7(32'h39cea303),
	.w8(32'hbae8a786),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e908),
	.w1(32'hbb0fd7bd),
	.w2(32'hbb1624e0),
	.w3(32'hbb2dbe9c),
	.w4(32'hba6fc244),
	.w5(32'hba82f68b),
	.w6(32'hbb115ea1),
	.w7(32'hba5c4f3a),
	.w8(32'hbb3a0917),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adef42),
	.w1(32'h39af5d73),
	.w2(32'h3a47e455),
	.w3(32'hb9a8969f),
	.w4(32'hb8b72c20),
	.w5(32'h383c1779),
	.w6(32'hb9ac831d),
	.w7(32'hb868c516),
	.w8(32'h38c3db67),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a021dfb),
	.w1(32'hba7d0c2e),
	.w2(32'hbb849430),
	.w3(32'h3aa7639d),
	.w4(32'hba67b810),
	.w5(32'hbb4b7d6f),
	.w6(32'hbb30ca0d),
	.w7(32'hbb386381),
	.w8(32'hbb718f41),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3743b),
	.w1(32'hb986a74d),
	.w2(32'hba967f8d),
	.w3(32'h399e2b10),
	.w4(32'hb9b8548f),
	.w5(32'hba4d84e8),
	.w6(32'hb9741acb),
	.w7(32'hb97b83df),
	.w8(32'hba0da2a3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03b471),
	.w1(32'hb7b4f9f7),
	.w2(32'h381b4a63),
	.w3(32'h3a191be5),
	.w4(32'h38431a32),
	.w5(32'h38a94797),
	.w6(32'hb8db393e),
	.w7(32'hb832052f),
	.w8(32'h38dbeaa1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacef2fc),
	.w1(32'hbaed887e),
	.w2(32'hbac40a14),
	.w3(32'hb9b4d032),
	.w4(32'hbaa543ba),
	.w5(32'hba0e8b3a),
	.w6(32'hb9a09801),
	.w7(32'hb90ee674),
	.w8(32'h399bf347),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357da75b),
	.w1(32'h37f5a512),
	.w2(32'h38eee8f0),
	.w3(32'h3920bbe6),
	.w4(32'h38b9fb76),
	.w5(32'h394425ab),
	.w6(32'h3936c2a7),
	.w7(32'h38c4568f),
	.w8(32'h3a007fde),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a845887),
	.w1(32'h3a7415f9),
	.w2(32'hba282d3e),
	.w3(32'h3aa80163),
	.w4(32'h388ab558),
	.w5(32'hba886cb3),
	.w6(32'hba3ff70e),
	.w7(32'hba393685),
	.w8(32'hbacb8270),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d368),
	.w1(32'h3aaeed60),
	.w2(32'h37e1ccff),
	.w3(32'hbaeaa802),
	.w4(32'h3aecf28b),
	.w5(32'h39a328f4),
	.w6(32'hba8e996a),
	.w7(32'h3a302727),
	.w8(32'hbb02814e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f1842),
	.w1(32'hb97d8cc7),
	.w2(32'hbad960e8),
	.w3(32'hb94460a4),
	.w4(32'hb812db15),
	.w5(32'hbab87274),
	.w6(32'hba97d133),
	.w7(32'hba63eae3),
	.w8(32'hbb2c8561),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39058109),
	.w1(32'h3abb044a),
	.w2(32'h3a990629),
	.w3(32'h3920b9d0),
	.w4(32'h3a72ca30),
	.w5(32'h3a6e8029),
	.w6(32'h3a00d47c),
	.w7(32'h3a45dfdc),
	.w8(32'h398f35bd),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb971d),
	.w1(32'hba69140d),
	.w2(32'hb9ac3173),
	.w3(32'hbaaf246d),
	.w4(32'h38d0e560),
	.w5(32'hba3bbc03),
	.w6(32'hba9f2141),
	.w7(32'h39294118),
	.w8(32'hbb13a916),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e4941),
	.w1(32'hbaa72721),
	.w2(32'hbb3997e7),
	.w3(32'h3a9d683c),
	.w4(32'hb9cb4945),
	.w5(32'hbaa719eb),
	.w6(32'hba7f4d4a),
	.w7(32'hb9fb2d6a),
	.w8(32'hba295331),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a18f3),
	.w1(32'hbb5ae73d),
	.w2(32'hbb755d55),
	.w3(32'hbb4bc689),
	.w4(32'hbb04e086),
	.w5(32'hbb23f47b),
	.w6(32'hbbb0fcce),
	.w7(32'hbb4cc598),
	.w8(32'hbb9070e0),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c21bb5),
	.w1(32'h3a5f38e1),
	.w2(32'h3a3faaea),
	.w3(32'h38c868e3),
	.w4(32'h3a1e2c09),
	.w5(32'h3a14c29d),
	.w6(32'h3a636dc5),
	.w7(32'h3a44054e),
	.w8(32'h3a23538e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e708c8),
	.w1(32'h39d28f84),
	.w2(32'h390bbd30),
	.w3(32'h39e166d0),
	.w4(32'h392dbbc3),
	.w5(32'hb8b04d5c),
	.w6(32'h3a2ec8a4),
	.w7(32'h39e83850),
	.w8(32'h39108c32),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f0b39),
	.w1(32'h3ab69859),
	.w2(32'hbb1c1470),
	.w3(32'hba543fa9),
	.w4(32'hb9d3e360),
	.w5(32'hbb143ee9),
	.w6(32'hbb585911),
	.w7(32'hbaa93227),
	.w8(32'hbb544f7d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a201400),
	.w1(32'hba852adf),
	.w2(32'hbb5da521),
	.w3(32'hb804ed6f),
	.w4(32'hbab2e6d1),
	.w5(32'hbbb421e9),
	.w6(32'hbb4a2f69),
	.w7(32'hba915128),
	.w8(32'hbb5d297c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac63472),
	.w1(32'hbad3a45a),
	.w2(32'hbb991384),
	.w3(32'hbb05fa13),
	.w4(32'hbaf35ec3),
	.w5(32'hbb5d492a),
	.w6(32'hbb17f224),
	.w7(32'hbb11400d),
	.w8(32'hbba7b46b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84aebc),
	.w1(32'hbb137010),
	.w2(32'hb993bd07),
	.w3(32'h3ad9674a),
	.w4(32'hba71f0a1),
	.w5(32'hbab61430),
	.w6(32'h3ae4d571),
	.w7(32'h388de4e0),
	.w8(32'hba2845dc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f250d7),
	.w1(32'hb922f8e5),
	.w2(32'hb9c489b9),
	.w3(32'h397929aa),
	.w4(32'hb8c0e14f),
	.w5(32'h36af37aa),
	.w6(32'hb8e81b7f),
	.w7(32'hb9559d56),
	.w8(32'h3a054da1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb938ad18),
	.w1(32'hba34cf95),
	.w2(32'hb9c24aa7),
	.w3(32'h3979c3d3),
	.w4(32'hb8890047),
	.w5(32'h3903c5e9),
	.w6(32'hb9966fa3),
	.w7(32'h3a027e03),
	.w8(32'h3a80da00),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4200fc),
	.w1(32'h3acd469b),
	.w2(32'hbb154adb),
	.w3(32'h3a925d9f),
	.w4(32'hbab70c37),
	.w5(32'hbb20e5e0),
	.w6(32'hbafd14f7),
	.w7(32'hbaf19295),
	.w8(32'hbaac6252),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95c9e5),
	.w1(32'hbb8a3486),
	.w2(32'hbb18e232),
	.w3(32'hbb314ae1),
	.w4(32'hbb1bdaea),
	.w5(32'hbb42e53a),
	.w6(32'hbbd7869b),
	.w7(32'hbb16dfe0),
	.w8(32'hba5c887f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a627213),
	.w1(32'hb9ee4985),
	.w2(32'hbb255acc),
	.w3(32'h3abb2d21),
	.w4(32'h3a82edd5),
	.w5(32'hb9a7e76a),
	.w6(32'hbacefda3),
	.w7(32'hbaa43cee),
	.w8(32'hba7adea6),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefd38d),
	.w1(32'h3b308df0),
	.w2(32'h3afd9364),
	.w3(32'h39981a12),
	.w4(32'h3ac0384a),
	.w5(32'h3a4290e1),
	.w6(32'h393afb5e),
	.w7(32'h3a09f79e),
	.w8(32'hba3db378),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a9b7d),
	.w1(32'hba92851b),
	.w2(32'hbb3bbd09),
	.w3(32'hbb145205),
	.w4(32'hb92eabf1),
	.w5(32'hbaf17501),
	.w6(32'hbab636c9),
	.w7(32'hba6a9fda),
	.w8(32'hbb7956dd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b83119),
	.w1(32'h39fd9c05),
	.w2(32'h3a111f24),
	.w3(32'h39428db4),
	.w4(32'h39d9a7da),
	.w5(32'h3a132f02),
	.w6(32'h39b01874),
	.w7(32'h39bf2daf),
	.w8(32'h39ab8308),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ad2b4),
	.w1(32'hb9fb18b5),
	.w2(32'hb9e929cd),
	.w3(32'h3a119a33),
	.w4(32'hb8f460f5),
	.w5(32'hb73d478f),
	.w6(32'hb9c12733),
	.w7(32'hb8c53dbf),
	.w8(32'h38ed3344),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89e167),
	.w1(32'h39bda441),
	.w2(32'h39990d76),
	.w3(32'h3a93a215),
	.w4(32'h3918591a),
	.w5(32'hba0e1dc8),
	.w6(32'h3a14440f),
	.w7(32'h3850d0c9),
	.w8(32'h39c37e3c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab9d2a),
	.w1(32'h39b52432),
	.w2(32'h36b9544d),
	.w3(32'h38a1dce4),
	.w4(32'h39bc7e91),
	.w5(32'hb93fabe8),
	.w6(32'h39ee7631),
	.w7(32'h3591bde3),
	.w8(32'hb98db534),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21f24a),
	.w1(32'h38b25497),
	.w2(32'hba88126b),
	.w3(32'h39a1b662),
	.w4(32'hb9a2cc22),
	.w5(32'hbaaf49f9),
	.w6(32'hb9467344),
	.w7(32'hb91403d2),
	.w8(32'hb9d21eea),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a676e),
	.w1(32'hbb1ae41d),
	.w2(32'hbba43ed7),
	.w3(32'hbaae4dae),
	.w4(32'hbb5c5e81),
	.w5(32'hbbb53b06),
	.w6(32'hbb70541c),
	.w7(32'hbb53e46f),
	.w8(32'hbb81e8e4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b921d8),
	.w1(32'hb9c1da12),
	.w2(32'hbaf045a2),
	.w3(32'hba9a7432),
	.w4(32'hba77fbd7),
	.w5(32'hbb2576d6),
	.w6(32'hbad9d92c),
	.w7(32'hbb0b91bd),
	.w8(32'hbb334ba7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b967f3),
	.w1(32'h3a8cdcd0),
	.w2(32'h395b6ec2),
	.w3(32'h3a0cfe1b),
	.w4(32'hb8f70c82),
	.w5(32'hb9fb56ed),
	.w6(32'h3a43153b),
	.w7(32'h39f9ae77),
	.w8(32'h39de657c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb554277),
	.w1(32'hbb3f24b9),
	.w2(32'hbb926e2b),
	.w3(32'hb9666f01),
	.w4(32'hba602319),
	.w5(32'hbae27876),
	.w6(32'hbb995d75),
	.w7(32'hbb3dc6dc),
	.w8(32'hba54b79b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6472d7),
	.w1(32'hbad59467),
	.w2(32'hbacc4aca),
	.w3(32'hb8b4c205),
	.w4(32'hba6dd930),
	.w5(32'hba9ed8d6),
	.w6(32'hbad31a81),
	.w7(32'hbaadabc5),
	.w8(32'hba281379),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fd26b2),
	.w1(32'hb8a915a4),
	.w2(32'hb8d486e2),
	.w3(32'h3985c35b),
	.w4(32'hb8421d45),
	.w5(32'hb8779462),
	.w6(32'hb8167bc8),
	.w7(32'hb891aa0e),
	.w8(32'h38c481be),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fede6),
	.w1(32'hba3e496a),
	.w2(32'hba840c27),
	.w3(32'h38c08b03),
	.w4(32'hb9f741db),
	.w5(32'hb9d4a2bc),
	.w6(32'hbab4baa0),
	.w7(32'hba8c6909),
	.w8(32'h39814c00),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a212fc6),
	.w1(32'h3a99332f),
	.w2(32'h3a5b39e9),
	.w3(32'h3a6410a0),
	.w4(32'h3a9c23de),
	.w5(32'h3a83e66c),
	.w6(32'h3a563b42),
	.w7(32'h3a3c39c1),
	.w8(32'h39b8ba7a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9313d),
	.w1(32'hb92ee225),
	.w2(32'hb9e216af),
	.w3(32'h39b33bc7),
	.w4(32'h38b1d3a1),
	.w5(32'h382b5dfa),
	.w6(32'hb7d5b6f1),
	.w7(32'hb746f6e9),
	.w8(32'h3980199d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e24d44),
	.w1(32'h382be7b0),
	.w2(32'h380a581e),
	.w3(32'h3a0f07c4),
	.w4(32'h36a2e7fa),
	.w5(32'h3864ad36),
	.w6(32'hb8ad843c),
	.w7(32'hb885470a),
	.w8(32'h38a50e75),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956953c),
	.w1(32'h398aebb3),
	.w2(32'h3a4ab1c9),
	.w3(32'h39a0d9f9),
	.w4(32'h39b16ec0),
	.w5(32'h39f012fe),
	.w6(32'h394d8f1b),
	.w7(32'h39acd2f8),
	.w8(32'hb902c152),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5966e8),
	.w1(32'h3aa8f707),
	.w2(32'h39f1c343),
	.w3(32'hb88ed6ed),
	.w4(32'h39f71e26),
	.w5(32'hb985d55b),
	.w6(32'hb89c404d),
	.w7(32'hb8c6b6c2),
	.w8(32'hba3c45c9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1722bf),
	.w1(32'hbb75c39e),
	.w2(32'hbb9eb50d),
	.w3(32'hbb0c5808),
	.w4(32'hbb2e49b1),
	.w5(32'hbb994701),
	.w6(32'hbb275e4c),
	.w7(32'hbaef7c66),
	.w8(32'hbba39bbd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb28a5),
	.w1(32'hbb179d04),
	.w2(32'hbb8316d2),
	.w3(32'hba51a1b9),
	.w4(32'hbac4552f),
	.w5(32'hbb281380),
	.w6(32'hba89a3c5),
	.w7(32'hba32d732),
	.w8(32'hba5060bf),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb317acc),
	.w1(32'hbb7b1734),
	.w2(32'hbb980367),
	.w3(32'hbb003b8d),
	.w4(32'hbb059b24),
	.w5(32'hbb4ffc78),
	.w6(32'hbb1d1977),
	.w7(32'hbb0d78ab),
	.w8(32'hbb2c6e8c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a424f7c),
	.w1(32'h393953c0),
	.w2(32'h3a2a84e8),
	.w3(32'h3a4d9a92),
	.w4(32'h39c5d7e5),
	.w5(32'h3a19180b),
	.w6(32'hb810bf6e),
	.w7(32'h39bd03da),
	.w8(32'h3a07f674),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87abf0f),
	.w1(32'hb9b1fe41),
	.w2(32'hb9967ee0),
	.w3(32'h39d1b6df),
	.w4(32'hb8decc26),
	.w5(32'hb886ed51),
	.w6(32'hb9345f1c),
	.w7(32'hb8f48247),
	.w8(32'h3923b6f7),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c7e8de),
	.w1(32'hb89045df),
	.w2(32'hb7b9e2a4),
	.w3(32'h39845006),
	.w4(32'hb5e4fcd4),
	.w5(32'h3878d6fe),
	.w6(32'hb9007cf6),
	.w7(32'hb8bb80dd),
	.w8(32'h38ab598a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a254cb),
	.w1(32'hb823fc00),
	.w2(32'hb8c51667),
	.w3(32'h39629b8a),
	.w4(32'hb81615ab),
	.w5(32'hb867550c),
	.w6(32'hb8856344),
	.w7(32'hb8bbc8a5),
	.w8(32'h383b7f0d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb309412),
	.w1(32'hbbaafee1),
	.w2(32'hbbab2846),
	.w3(32'hba8f4ffa),
	.w4(32'hbb0f7485),
	.w5(32'hbb2c8afa),
	.w6(32'hbb4e5859),
	.w7(32'hbb0438f0),
	.w8(32'hbb27c668),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80203f),
	.w1(32'hba1f3130),
	.w2(32'hba3c98ac),
	.w3(32'h39541844),
	.w4(32'hb9b6a9d8),
	.w5(32'hba0ba0a8),
	.w6(32'hba281a81),
	.w7(32'hba2e98f0),
	.w8(32'hba6183bf),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5cc4a),
	.w1(32'h39ba6340),
	.w2(32'h3a44ef7c),
	.w3(32'h3a568888),
	.w4(32'h39c63dc3),
	.w5(32'h3a7558ac),
	.w6(32'h3a5f7b81),
	.w7(32'h3a31405e),
	.w8(32'h3a979ba7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a717e),
	.w1(32'hb947a2ef),
	.w2(32'h37bf1f69),
	.w3(32'hba032427),
	.w4(32'hb9968e67),
	.w5(32'hb97989a9),
	.w6(32'h39acf6a2),
	.w7(32'h3a1a545b),
	.w8(32'h3a4f9699),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39374b6e),
	.w1(32'hb8805859),
	.w2(32'hb8f54689),
	.w3(32'h39f17a9d),
	.w4(32'h37f88959),
	.w5(32'hb8875f9e),
	.w6(32'hb81492e4),
	.w7(32'hb902e433),
	.w8(32'hb873bc3c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e814d7),
	.w1(32'hba92d98d),
	.w2(32'hbb0a425a),
	.w3(32'h396443a4),
	.w4(32'hb8bdfa44),
	.w5(32'hba0459bf),
	.w6(32'hbaa64a78),
	.w7(32'hbaa1cb27),
	.w8(32'hbadf409f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3183dd),
	.w1(32'h37bb9faf),
	.w2(32'hb7b9f461),
	.w3(32'h3a072961),
	.w4(32'h39ca826e),
	.w5(32'h39853fd6),
	.w6(32'h399444dc),
	.w7(32'h39c88df0),
	.w8(32'h3a0a4d4f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5df71a),
	.w1(32'hbbb2f25c),
	.w2(32'hbb9cb223),
	.w3(32'hbb4cb9f7),
	.w4(32'hbb08d4a1),
	.w5(32'hbb0051b1),
	.w6(32'hbb849f6c),
	.w7(32'hb99f74ab),
	.w8(32'hba1407a6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5cae4),
	.w1(32'h3b2412b2),
	.w2(32'hbacb2cb1),
	.w3(32'h3a1dd7ea),
	.w4(32'h3aca76a8),
	.w5(32'h3a01e3ff),
	.w6(32'h3b3fd77c),
	.w7(32'hbad915bd),
	.w8(32'h395f39cb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396adfe8),
	.w1(32'hbb1da448),
	.w2(32'h3afe2f70),
	.w3(32'h3aa898f8),
	.w4(32'hbbaac8e6),
	.w5(32'hba3534b1),
	.w6(32'hbbe513cd),
	.w7(32'h3806108c),
	.w8(32'h3b322108),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule