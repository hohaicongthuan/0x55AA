module layer_8_featuremap_167(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c818a26),
	.w1(32'hbaf4d758),
	.w2(32'h3b13934f),
	.w3(32'h3c8aa2f1),
	.w4(32'h3b454f2b),
	.w5(32'h3c0e0245),
	.w6(32'h3b2270de),
	.w7(32'h3bc7dc09),
	.w8(32'h3bf82805),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a4d5),
	.w1(32'h3b2985c2),
	.w2(32'h3bb696e6),
	.w3(32'h3c32de36),
	.w4(32'h3b23fec6),
	.w5(32'h3c0372cb),
	.w6(32'h37a45e0c),
	.w7(32'h3a7bf6fa),
	.w8(32'hbb2f845e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae005a),
	.w1(32'h3c259c24),
	.w2(32'h3babb4d7),
	.w3(32'h3c51617d),
	.w4(32'h3b90b1f8),
	.w5(32'hba171cf0),
	.w6(32'h3c6641d3),
	.w7(32'h3bfda428),
	.w8(32'hb9dfbd4c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc922e1),
	.w1(32'h3b64cb19),
	.w2(32'h3c031b08),
	.w3(32'h3aec724d),
	.w4(32'h3abefb82),
	.w5(32'hba9a9712),
	.w6(32'h3c1789e1),
	.w7(32'h3c116914),
	.w8(32'h3c19a7bb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf507f6),
	.w1(32'h3c947c0c),
	.w2(32'h3bc1043c),
	.w3(32'h3c3e54cc),
	.w4(32'h3c9b0692),
	.w5(32'h3c38e356),
	.w6(32'h3bf57df1),
	.w7(32'h3ae95f06),
	.w8(32'hbc1a419d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b48f0),
	.w1(32'h3a6e2344),
	.w2(32'h3a9907b5),
	.w3(32'hbbace554),
	.w4(32'h3b0af4c5),
	.w5(32'h39f9de63),
	.w6(32'h3bc4dff9),
	.w7(32'h3ba61d3c),
	.w8(32'h3b1468a0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3df53),
	.w1(32'h3b500785),
	.w2(32'hbb61fa99),
	.w3(32'hba9f2fba),
	.w4(32'h3a406206),
	.w5(32'hbbd07d88),
	.w6(32'h3b73c03a),
	.w7(32'h3a2c389d),
	.w8(32'h39dbffbf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf55938),
	.w1(32'h3b78b608),
	.w2(32'h3bff833c),
	.w3(32'hba7e83ae),
	.w4(32'hba2bddd5),
	.w5(32'hba20b789),
	.w6(32'h3c0adc8c),
	.w7(32'h3c0edfc5),
	.w8(32'h3c46e3b5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90ea7c),
	.w1(32'h3d2fcc02),
	.w2(32'h3b898ec3),
	.w3(32'h3c0b14d9),
	.w4(32'h3d2623b7),
	.w5(32'h3c00748e),
	.w6(32'h3cee5d5b),
	.w7(32'h3b8101b3),
	.w8(32'hbce29f3b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd279857),
	.w1(32'hbb867fd8),
	.w2(32'hbbe22c3c),
	.w3(32'hbcb671f3),
	.w4(32'hbbc5cfda),
	.w5(32'hbbaa86a9),
	.w6(32'hbb08ed30),
	.w7(32'hbbefc19e),
	.w8(32'hbb2b7571),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a987825),
	.w1(32'h3b44a192),
	.w2(32'h3b4be667),
	.w3(32'h3824e0d7),
	.w4(32'hbac75b6d),
	.w5(32'hbc4c3833),
	.w6(32'h3c586975),
	.w7(32'h3ba974f9),
	.w8(32'h3b466c31),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9c716),
	.w1(32'hbb1e1d0c),
	.w2(32'hbbfe36ad),
	.w3(32'hbbb09a0f),
	.w4(32'hbb42e95b),
	.w5(32'hbbfd7893),
	.w6(32'h3b0b6ecc),
	.w7(32'hbb10a58a),
	.w8(32'h3ba8ef9d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7618b9),
	.w1(32'h3c1bf9f4),
	.w2(32'h3c1fc988),
	.w3(32'h3bb6000b),
	.w4(32'h3ae478d5),
	.w5(32'h3bcbc274),
	.w6(32'h3c704655),
	.w7(32'h3baa633b),
	.w8(32'h3b27ca14),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2fe28),
	.w1(32'h3b4338a6),
	.w2(32'hbb189369),
	.w3(32'h3b95ca3d),
	.w4(32'hb9aa600c),
	.w5(32'h3a7e742e),
	.w6(32'h3aa0ed28),
	.w7(32'h3bb9a597),
	.w8(32'h3b81642d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba13fa5),
	.w1(32'h3c5a0358),
	.w2(32'hb9fc10dc),
	.w3(32'hbb1be34c),
	.w4(32'h3c4a2db0),
	.w5(32'hbaa16ca4),
	.w6(32'h3c4b98f0),
	.w7(32'h3b2166e1),
	.w8(32'hbbdf3a59),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc027c55),
	.w1(32'hbb524a81),
	.w2(32'hbc9996b5),
	.w3(32'hbc287e2e),
	.w4(32'hb9f83227),
	.w5(32'hbc89e08e),
	.w6(32'h3b7c1202),
	.w7(32'hbc04fde6),
	.w8(32'hba8f4151),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83dff4),
	.w1(32'hbc083b73),
	.w2(32'h3b870172),
	.w3(32'hbc66f0c1),
	.w4(32'hb8eb3eec),
	.w5(32'h3af443ce),
	.w6(32'h3b52f3a8),
	.w7(32'h3c36fb54),
	.w8(32'h3ba67800),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c442e0f),
	.w1(32'hbc30e9af),
	.w2(32'hba4202a3),
	.w3(32'h3c23619d),
	.w4(32'hbbeda36f),
	.w5(32'hbbcbed27),
	.w6(32'hbba05835),
	.w7(32'hbbe49d1e),
	.w8(32'hbb147708),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56cec),
	.w1(32'hbcbc6d6e),
	.w2(32'hbc77555d),
	.w3(32'h3c0b583d),
	.w4(32'hbbc46234),
	.w5(32'hbc03880d),
	.w6(32'hbbfd26e0),
	.w7(32'hbb472729),
	.w8(32'hbbdff20f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79ec76),
	.w1(32'h3c016663),
	.w2(32'h3bb26c50),
	.w3(32'h3b8a80da),
	.w4(32'h3c1b915e),
	.w5(32'h3b09a591),
	.w6(32'h3c034b9d),
	.w7(32'h3a04d09b),
	.w8(32'h3ba6d09a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dfa7f),
	.w1(32'h3cc87ea3),
	.w2(32'h3c88d930),
	.w3(32'hbc07125e),
	.w4(32'h3b8f44b9),
	.w5(32'h3caa7c1f),
	.w6(32'h3ca0d507),
	.w7(32'h3c86884d),
	.w8(32'h3c10968b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0d004),
	.w1(32'h38a01344),
	.w2(32'h3bf394a2),
	.w3(32'h3c93c0c9),
	.w4(32'h3a62219c),
	.w5(32'hb936b0fc),
	.w6(32'h3bb8425c),
	.w7(32'hba7b7a19),
	.w8(32'hbb76e5c7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8328b),
	.w1(32'h3be1009b),
	.w2(32'hbc74fcad),
	.w3(32'h3c3a2349),
	.w4(32'h3c2b96b2),
	.w5(32'hbaaba0e2),
	.w6(32'h3c04bef5),
	.w7(32'h3b46f217),
	.w8(32'hbc3a3d3f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccd5dd),
	.w1(32'h3c0f5d26),
	.w2(32'h3c01f6d2),
	.w3(32'h3c1e75bf),
	.w4(32'h3c0f5229),
	.w5(32'h3c60b0aa),
	.w6(32'h3b434635),
	.w7(32'h3b215724),
	.w8(32'h3aa53702),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58fe4f),
	.w1(32'hbba4a33d),
	.w2(32'hbc72d337),
	.w3(32'h3a7eed6c),
	.w4(32'h3b2a4460),
	.w5(32'h3c3d40ca),
	.w6(32'h3c15bd73),
	.w7(32'h3be4a32b),
	.w8(32'hbb1e7f0b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc483875),
	.w1(32'h3c734484),
	.w2(32'h3cad89c7),
	.w3(32'h3c9da354),
	.w4(32'h3c2b7b4b),
	.w5(32'h3caab2a1),
	.w6(32'h3c8401ff),
	.w7(32'h3c616e2a),
	.w8(32'h3c6d12d6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c234d49),
	.w1(32'hbb599147),
	.w2(32'hbbaaf29c),
	.w3(32'h3b60accc),
	.w4(32'hbb2e6cc8),
	.w5(32'hbc009a69),
	.w6(32'hba34ee1d),
	.w7(32'h3c2647ee),
	.w8(32'h3c3b45ad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c212c9f),
	.w1(32'h3c3916ea),
	.w2(32'h3cc0d24f),
	.w3(32'h3be22421),
	.w4(32'hbb56ccd4),
	.w5(32'h3c482d5d),
	.w6(32'h3cacd14c),
	.w7(32'h3c3c3311),
	.w8(32'h3c50b98b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c519e),
	.w1(32'h3c5342b9),
	.w2(32'h3d154a4f),
	.w3(32'h3c43ea8b),
	.w4(32'h3c72da3f),
	.w5(32'h3ce70e1b),
	.w6(32'h3bde40b3),
	.w7(32'h3ca86539),
	.w8(32'h3d0ac516),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d484dce),
	.w1(32'h3bac96e8),
	.w2(32'h3b9925cd),
	.w3(32'h3d16f066),
	.w4(32'h3be98eb5),
	.w5(32'h3c443751),
	.w6(32'h3af971c7),
	.w7(32'h3b97d471),
	.w8(32'h3b6ff51b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80786e),
	.w1(32'hbc82dcff),
	.w2(32'hbc0e7907),
	.w3(32'h3a67f0db),
	.w4(32'hbb3d2b68),
	.w5(32'hbbe03f1c),
	.w6(32'hbc47ed36),
	.w7(32'hbb179a43),
	.w8(32'h3c1a951f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90204d),
	.w1(32'h3c450162),
	.w2(32'h3c447909),
	.w3(32'hbc3ab374),
	.w4(32'h3c522f75),
	.w5(32'h3c2622d5),
	.w6(32'h3c762388),
	.w7(32'h3b9d2580),
	.w8(32'hbac6a9cc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99ddad),
	.w1(32'hbc078b5d),
	.w2(32'h3aeefba4),
	.w3(32'h3c00beaf),
	.w4(32'h3ad3f3e2),
	.w5(32'hba92abcf),
	.w6(32'hbaf38468),
	.w7(32'hbb9a9349),
	.w8(32'h3b3e5531),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfef5b),
	.w1(32'hbbca2a02),
	.w2(32'hbb8c820a),
	.w3(32'h3b531bdd),
	.w4(32'hbbba3577),
	.w5(32'hbbbd62af),
	.w6(32'hbb6d8a71),
	.w7(32'hbb297b9c),
	.w8(32'h3b899031),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be80e1a),
	.w1(32'hbbe7286c),
	.w2(32'hbb614626),
	.w3(32'h3b9592bc),
	.w4(32'hbc533ee7),
	.w5(32'hb9a5bd42),
	.w6(32'hbb60fb6e),
	.w7(32'h3a9f752d),
	.w8(32'h3b7e0941),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10e11e),
	.w1(32'h3c3179f0),
	.w2(32'h3b7372e6),
	.w3(32'h3b3c1601),
	.w4(32'h3bc027ca),
	.w5(32'hba22896f),
	.w6(32'h369b5ce4),
	.w7(32'h3b82affc),
	.w8(32'hb88d2cea),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9452f),
	.w1(32'h3c9f7149),
	.w2(32'h3cb39c31),
	.w3(32'h3a9b3b64),
	.w4(32'h3c6ce761),
	.w5(32'h3ca9944d),
	.w6(32'h3c9dee30),
	.w7(32'h3c8a4612),
	.w8(32'h3c4d23cd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdf04e),
	.w1(32'h3ca5418c),
	.w2(32'h3bc69342),
	.w3(32'h3cdc3185),
	.w4(32'h3c861be0),
	.w5(32'h3bcb46b2),
	.w6(32'h3c00c88f),
	.w7(32'hba96d376),
	.w8(32'hbc2e5136),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3531b5),
	.w1(32'hbb565520),
	.w2(32'hbab35fa7),
	.w3(32'hbbf7b99b),
	.w4(32'hbb77f272),
	.w5(32'hbadd3fb6),
	.w6(32'hbb392eca),
	.w7(32'hbbaaf277),
	.w8(32'h3a0ced32),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0c72d),
	.w1(32'h3bd698b1),
	.w2(32'h3b9131c1),
	.w3(32'hbbfb6e4c),
	.w4(32'h3bb00c2d),
	.w5(32'h3bb8c907),
	.w6(32'hb90a2d00),
	.w7(32'hba6a8e6d),
	.w8(32'hbad7c046),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f4fd2),
	.w1(32'hbb87a5de),
	.w2(32'hbb683f80),
	.w3(32'h3c202b0b),
	.w4(32'hbb8276db),
	.w5(32'hbb5f94c0),
	.w6(32'h3b80a051),
	.w7(32'hbb73dbf2),
	.w8(32'h3b806210),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f3955),
	.w1(32'hbd191e99),
	.w2(32'hbd7b8708),
	.w3(32'hbbaa4215),
	.w4(32'hbd0927dd),
	.w5(32'hbd49764a),
	.w6(32'hbc87f680),
	.w7(32'hbd2697cd),
	.w8(32'hbd079031),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd37d084),
	.w1(32'h3c2cb151),
	.w2(32'h3ca475a0),
	.w3(32'hbd2e1738),
	.w4(32'h3baba184),
	.w5(32'h3c79deab),
	.w6(32'h3afe8800),
	.w7(32'h3c03b9cf),
	.w8(32'h39946bcc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c790827),
	.w1(32'hbb14a2bc),
	.w2(32'hbc27a511),
	.w3(32'h3c3ba5ed),
	.w4(32'h3b16516d),
	.w5(32'hbbce309b),
	.w6(32'h3b2ace08),
	.w7(32'hbb8e8d5b),
	.w8(32'h3ac82a36),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b484c),
	.w1(32'h3c0333d1),
	.w2(32'h3c450e7c),
	.w3(32'h392edf04),
	.w4(32'h3c2305b4),
	.w5(32'h3c3eb864),
	.w6(32'h3b3c7f64),
	.w7(32'h3b37c312),
	.w8(32'h3b39b14d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b266f),
	.w1(32'hbb0bd73f),
	.w2(32'hbb875e2f),
	.w3(32'h3c14b54d),
	.w4(32'hba25b126),
	.w5(32'hbbee4d8e),
	.w6(32'h3b639023),
	.w7(32'h3a9b3c48),
	.w8(32'h3b3c0624),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e3075),
	.w1(32'hbc373d0a),
	.w2(32'hbb70294a),
	.w3(32'hbb1f41a9),
	.w4(32'hbbe37928),
	.w5(32'h3ba636f7),
	.w6(32'hbbb07632),
	.w7(32'hbac3bd75),
	.w8(32'h3a50dac4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b366371),
	.w1(32'hbacb82b5),
	.w2(32'h3b9f7ef9),
	.w3(32'h3c2b1f78),
	.w4(32'hbb6d7786),
	.w5(32'h3b2cd85e),
	.w6(32'h3bbe4646),
	.w7(32'hb9a4694e),
	.w8(32'hba0998f3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a664b2c),
	.w1(32'h3b4985a5),
	.w2(32'h3b9e0f9a),
	.w3(32'h3b51d3ff),
	.w4(32'h3b086af5),
	.w5(32'hbad389ad),
	.w6(32'h3bc47501),
	.w7(32'h3ba753f2),
	.w8(32'hbb44e03e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dbc3d),
	.w1(32'h3a38328a),
	.w2(32'hbb4ebc66),
	.w3(32'h3bb91dc9),
	.w4(32'h3ac09539),
	.w5(32'hb9bedbe8),
	.w6(32'h3ae265c6),
	.w7(32'hbb2fc68a),
	.w8(32'h3b515771),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c336a4e),
	.w1(32'h39cfd410),
	.w2(32'hbbbce77e),
	.w3(32'h3b2a2ecd),
	.w4(32'h3a90e0d5),
	.w5(32'hbbe5c2b6),
	.w6(32'h3b60e46f),
	.w7(32'hbbfe5df7),
	.w8(32'hbba8d2d4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46591d),
	.w1(32'hbcd2f6fb),
	.w2(32'hbcc0eb96),
	.w3(32'h3bf9e6e1),
	.w4(32'hbc9b280c),
	.w5(32'hbc698b04),
	.w6(32'hbbf86905),
	.w7(32'hbc421c6b),
	.w8(32'hbc18a54e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd072527),
	.w1(32'h3b3141e7),
	.w2(32'hbb82dd8f),
	.w3(32'hbc8f41da),
	.w4(32'h3b98ee93),
	.w5(32'h3b04e21c),
	.w6(32'h3b31458b),
	.w7(32'hbb98ab80),
	.w8(32'hbc1ecb7c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d49c6),
	.w1(32'h3b6dc647),
	.w2(32'h37b90a12),
	.w3(32'hbadb27a7),
	.w4(32'h3c0211cf),
	.w5(32'h3c132274),
	.w6(32'h3a9351d0),
	.w7(32'hba9a0e79),
	.w8(32'hbbdca21c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72fb90),
	.w1(32'hbc8434ad),
	.w2(32'hbc7d0b50),
	.w3(32'h3b0494db),
	.w4(32'hbc368f9e),
	.w5(32'hbaf50f7b),
	.w6(32'hbc879c4b),
	.w7(32'hbac44a94),
	.w8(32'h3bc370d9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1e299),
	.w1(32'h3bbd27b9),
	.w2(32'h3bb1d01f),
	.w3(32'h3bdc17d0),
	.w4(32'h3b5d3db8),
	.w5(32'h3bec7a96),
	.w6(32'hb95ccf12),
	.w7(32'h3aec11ff),
	.w8(32'h3c255c1b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f262b),
	.w1(32'hbc782a6d),
	.w2(32'hbbeb7e02),
	.w3(32'h3ba1d221),
	.w4(32'hbc34573f),
	.w5(32'hbc38cf00),
	.w6(32'hbb9ff267),
	.w7(32'hbbc570fb),
	.w8(32'hbae9f215),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d01c),
	.w1(32'h3cd5907f),
	.w2(32'h3d274e16),
	.w3(32'hb9a040ce),
	.w4(32'h3ca58657),
	.w5(32'h3d0b77db),
	.w6(32'h3cbdc60b),
	.w7(32'h3cd3ab03),
	.w8(32'h3c7573d9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd7af35),
	.w1(32'hbc05a45d),
	.w2(32'hbb7fda0d),
	.w3(32'h3cb6be12),
	.w4(32'hbc0e5752),
	.w5(32'hbbdb14d4),
	.w6(32'hbc1df335),
	.w7(32'hbbf7b8f0),
	.w8(32'hbb1d299e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bcee6),
	.w1(32'h3c08ffb0),
	.w2(32'h3c2e4f11),
	.w3(32'hbb24b6f3),
	.w4(32'h3c4f9bb9),
	.w5(32'h3c14668f),
	.w6(32'h3b12b9f9),
	.w7(32'h3b2df715),
	.w8(32'h3a585e0a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eba02),
	.w1(32'hbbaade20),
	.w2(32'hbbfd554b),
	.w3(32'h3bac0620),
	.w4(32'hbbef8710),
	.w5(32'hbc320892),
	.w6(32'h3ad70abc),
	.w7(32'h3b58b10f),
	.w8(32'h3b940a85),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb480c56),
	.w1(32'h3c1747b9),
	.w2(32'hbb96c936),
	.w3(32'hbc35a2c8),
	.w4(32'h3ab3d3fc),
	.w5(32'hbaac404e),
	.w6(32'h3c79629c),
	.w7(32'h3b107b53),
	.w8(32'hbc503602),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84acea),
	.w1(32'h3c704f30),
	.w2(32'h3c74e5f2),
	.w3(32'h3c048d5c),
	.w4(32'h3c8f4099),
	.w5(32'h3be2386c),
	.w6(32'h3c6ef230),
	.w7(32'h3c117f8f),
	.w8(32'h3c9ee17e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94ab6b),
	.w1(32'hbc83c066),
	.w2(32'hbc80128c),
	.w3(32'h3c79bf1f),
	.w4(32'hbc550d9f),
	.w5(32'hbc6233cc),
	.w6(32'hbc3ad4c7),
	.w7(32'hbc1d32e0),
	.w8(32'hbca7cd5b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1c429),
	.w1(32'hbc2f2340),
	.w2(32'hbb44a00e),
	.w3(32'hbcc9d41f),
	.w4(32'hbc031e06),
	.w5(32'hbb6f4fd9),
	.w6(32'hbbdaf98b),
	.w7(32'hbba662df),
	.w8(32'hb6f0e67f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1efc33),
	.w1(32'h3bd02b00),
	.w2(32'h3bfdd3f7),
	.w3(32'h3b814136),
	.w4(32'h3c47d8a7),
	.w5(32'h3c18eb70),
	.w6(32'h3b75ef31),
	.w7(32'h3b9b775e),
	.w8(32'h3b8ef4a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a9eb8),
	.w1(32'h3b7074db),
	.w2(32'h3a107b84),
	.w3(32'h3c3c81ca),
	.w4(32'h3b577140),
	.w5(32'h3c45557c),
	.w6(32'h3bece7c7),
	.w7(32'h3c8564a0),
	.w8(32'h3b3988c4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0acb20),
	.w1(32'h3c0fc982),
	.w2(32'h3c0046c8),
	.w3(32'h3b80f26f),
	.w4(32'h3c23051c),
	.w5(32'h3bda76e4),
	.w6(32'h3c32d5e0),
	.w7(32'h3c4460d4),
	.w8(32'h3c5d7765),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7bde8),
	.w1(32'h3bfa2d9d),
	.w2(32'h3c144cc1),
	.w3(32'h3c327176),
	.w4(32'h3b88fed0),
	.w5(32'h3a74640b),
	.w6(32'hba7dc1fe),
	.w7(32'h3a1a80ee),
	.w8(32'h3b6d6483),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01f682),
	.w1(32'hbb40a2c1),
	.w2(32'h3b0b9073),
	.w3(32'h3c33c850),
	.w4(32'h3bc96a71),
	.w5(32'h3bbc39ee),
	.w6(32'h3b1e2c0b),
	.w7(32'h3b96463e),
	.w8(32'h3c182050),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68abc8),
	.w1(32'hbcf4bd16),
	.w2(32'hbd669f38),
	.w3(32'hba48b9d8),
	.w4(32'hbcc1567f),
	.w5(32'hbd3499b8),
	.w6(32'hbca3f8c1),
	.w7(32'hbd13afa5),
	.w8(32'hbce0fa5c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd48e400),
	.w1(32'h3c72a0c4),
	.w2(32'h3c7ccb9c),
	.w3(32'hbd1eab6b),
	.w4(32'h3c3e1289),
	.w5(32'h3c2c2e0b),
	.w6(32'h3b07c7e7),
	.w7(32'h3c13f8b9),
	.w8(32'h3c398ca3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3ded3),
	.w1(32'hb914d30d),
	.w2(32'h3bbcd41d),
	.w3(32'h3c0f07e1),
	.w4(32'hbad2d217),
	.w5(32'h3bf34c49),
	.w6(32'h3bb2db09),
	.w7(32'h3bfc829b),
	.w8(32'h3aaf92f4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109bc4),
	.w1(32'h3b9a5f3d),
	.w2(32'h3c69ec81),
	.w3(32'h3c67549e),
	.w4(32'h3bea3399),
	.w5(32'h3c103a04),
	.w6(32'h3b2c77ec),
	.w7(32'h3c13dfa3),
	.w8(32'h3b8d26b4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc7949),
	.w1(32'hbcfab156),
	.w2(32'hbd32e5c2),
	.w3(32'h3b18d040),
	.w4(32'hbd09e4ac),
	.w5(32'hbce1e9b0),
	.w6(32'hbc4f0fe7),
	.w7(32'hbcbf404e),
	.w8(32'hbc6186c4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc84a94),
	.w1(32'hbb38fe22),
	.w2(32'hbc8c419f),
	.w3(32'hbc2d00ce),
	.w4(32'hbbd10823),
	.w5(32'hbc6f986f),
	.w6(32'hbbde9775),
	.w7(32'hbc86c120),
	.w8(32'hbc93adb2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceaaaf0),
	.w1(32'h3c0e6bc4),
	.w2(32'h3c8f5439),
	.w3(32'hbcbd3335),
	.w4(32'h3bab411e),
	.w5(32'h3c67a5d7),
	.w6(32'h3b814ca6),
	.w7(32'h3c1be2d7),
	.w8(32'h3ba6a477),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d07dc),
	.w1(32'h3caa3f4c),
	.w2(32'h3ce12f31),
	.w3(32'h3c331dca),
	.w4(32'h3c91d69a),
	.w5(32'h3ca92188),
	.w6(32'h3c524bea),
	.w7(32'h3c842407),
	.w8(32'h3c2db6ec),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f4c64),
	.w1(32'hbce5a466),
	.w2(32'hbd045cc7),
	.w3(32'h3cb5a796),
	.w4(32'hbbdcc001),
	.w5(32'hbc2d1577),
	.w6(32'hbbd650c5),
	.w7(32'hbbc17bcc),
	.w8(32'hbb8f77d4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6587e),
	.w1(32'h3c281990),
	.w2(32'h3a4494ef),
	.w3(32'hbc84577a),
	.w4(32'h3b8ef934),
	.w5(32'h3b2c24a8),
	.w6(32'h3b683d52),
	.w7(32'h3b2e4e3a),
	.w8(32'h3aa64d04),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67d28e),
	.w1(32'h3b697e03),
	.w2(32'h3b955edb),
	.w3(32'h3b8e619b),
	.w4(32'h3baf51d9),
	.w5(32'h3a0ab49d),
	.w6(32'h3c495052),
	.w7(32'h3bcf63fb),
	.w8(32'h37f5889c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d8dfb),
	.w1(32'h3c281e9a),
	.w2(32'h3bc0aa92),
	.w3(32'h3c21215e),
	.w4(32'h3b7faa51),
	.w5(32'h3a927076),
	.w6(32'h3bafaa8c),
	.w7(32'h3bc8a156),
	.w8(32'h3b7b820c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7603ac),
	.w1(32'hbb12fa0d),
	.w2(32'hbc6e054a),
	.w3(32'h3c158b97),
	.w4(32'h3b876cb2),
	.w5(32'hbbbd5399),
	.w6(32'hbb35b51b),
	.w7(32'hbbde5920),
	.w8(32'hbb882d69),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f5079),
	.w1(32'h3b8857b0),
	.w2(32'h3c9ab533),
	.w3(32'h3ad40c4a),
	.w4(32'h3bc8843a),
	.w5(32'h3c9df6ec),
	.w6(32'h3c21aa6e),
	.w7(32'h3c5fb576),
	.w8(32'h3c87ec2e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ffd40),
	.w1(32'h3ba8159c),
	.w2(32'hbb8cc5ed),
	.w3(32'h3c943eb7),
	.w4(32'h3c15ac75),
	.w5(32'h3b559280),
	.w6(32'h3c47d30f),
	.w7(32'h3b2a8280),
	.w8(32'h3c07267f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c675f),
	.w1(32'h3aae2ee7),
	.w2(32'h3b6f6ed7),
	.w3(32'hbbfe9554),
	.w4(32'h3b327f76),
	.w5(32'h3a94d044),
	.w6(32'h3c4d648e),
	.w7(32'h3c26125f),
	.w8(32'hbad95ad4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3ee76),
	.w1(32'hbc95cd3e),
	.w2(32'hbc76637c),
	.w3(32'hbbe6ea26),
	.w4(32'hbc00ea85),
	.w5(32'hbc03b812),
	.w6(32'hbc5b8827),
	.w7(32'hbc03b0f6),
	.w8(32'hba5953be),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30296b),
	.w1(32'h3ade045c),
	.w2(32'h3b6cb7ae),
	.w3(32'hbc0caa6e),
	.w4(32'hbc37934b),
	.w5(32'h3bbf4fbc),
	.w6(32'h3c85d069),
	.w7(32'h3bcb92cc),
	.w8(32'hbb7b9a17),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf99f0),
	.w1(32'hbbadd503),
	.w2(32'hbb90e2f0),
	.w3(32'h3c841e55),
	.w4(32'h3ba39e5f),
	.w5(32'h3bd35f4d),
	.w6(32'hbab530c1),
	.w7(32'h3ba17f09),
	.w8(32'h3c2e8ae2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fba07),
	.w1(32'hb984b006),
	.w2(32'h3bae0dbb),
	.w3(32'h3b85e41b),
	.w4(32'hbbe1b264),
	.w5(32'hbab1a16c),
	.w6(32'h3b018f8b),
	.w7(32'h3b4c64e4),
	.w8(32'hbb5aef04),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab23c8),
	.w1(32'h3b8f7a04),
	.w2(32'h3c89fbbf),
	.w3(32'h3ae57bad),
	.w4(32'hbab5796f),
	.w5(32'h3be8b26a),
	.w6(32'h3c319277),
	.w7(32'h3c127102),
	.w8(32'h3be41f69),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b6448),
	.w1(32'hba9053a7),
	.w2(32'h3b47c0f0),
	.w3(32'h3b059d40),
	.w4(32'h3ad8b2ab),
	.w5(32'h3b78ee19),
	.w6(32'hbb1daaef),
	.w7(32'h3b85049c),
	.w8(32'hbb74842a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe8c10),
	.w1(32'hbb9e5b64),
	.w2(32'h3ab5aebd),
	.w3(32'h38edf80c),
	.w4(32'hbb9ab85c),
	.w5(32'h39c2c842),
	.w6(32'hbb47644c),
	.w7(32'hbab279ba),
	.w8(32'h3b1613ad),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed2011),
	.w1(32'hbc3e38e9),
	.w2(32'h3b169c8a),
	.w3(32'h3b8a001a),
	.w4(32'hbc045f48),
	.w5(32'h3bd76fc9),
	.w6(32'hbbf5de9f),
	.w7(32'h3b20a4f4),
	.w8(32'h3c236c78),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20ea6f),
	.w1(32'hbb48bf7e),
	.w2(32'hbc3fe46d),
	.w3(32'h3c3097f1),
	.w4(32'hbbbafc11),
	.w5(32'hbc499d6d),
	.w6(32'hbc1c1b1f),
	.w7(32'hbc23e6eb),
	.w8(32'hbc039583),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc196e65),
	.w1(32'h3cc69297),
	.w2(32'h3cd219dc),
	.w3(32'hbc3bb054),
	.w4(32'h3cd7d643),
	.w5(32'h3cb28ddb),
	.w6(32'h3ca313df),
	.w7(32'h3c9d6c1d),
	.w8(32'h3cbb8b33),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a213f),
	.w1(32'hbacebb61),
	.w2(32'h3bbe1260),
	.w3(32'h3cfcb52e),
	.w4(32'h3ad1f666),
	.w5(32'h3a6560d5),
	.w6(32'hbbb9443e),
	.w7(32'hba964ee0),
	.w8(32'h3beaaf08),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad871ef),
	.w1(32'hbb6def0b),
	.w2(32'hbb9c7cc6),
	.w3(32'h3b64cc66),
	.w4(32'h3b6a7e33),
	.w5(32'hbb87e11f),
	.w6(32'hbbd4613d),
	.w7(32'hbba31628),
	.w8(32'h3bc8a72c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb484666),
	.w1(32'hbbc7645d),
	.w2(32'hbc2cc677),
	.w3(32'hbb83eede),
	.w4(32'h3a06ae0c),
	.w5(32'hbb88fdc7),
	.w6(32'hbb5246c4),
	.w7(32'hbc446d09),
	.w8(32'hbbd3e277),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc815a76),
	.w1(32'hbc71b4b7),
	.w2(32'hbc4748e2),
	.w3(32'hbc5b4ea6),
	.w4(32'h3a1766f1),
	.w5(32'hbbb646a8),
	.w6(32'hbb9e7a6a),
	.w7(32'hbad3bd2e),
	.w8(32'h3b45acd1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d33a06),
	.w1(32'h3c084979),
	.w2(32'h3b06d1aa),
	.w3(32'hbb834fc1),
	.w4(32'h3b3eda0f),
	.w5(32'h3b384741),
	.w6(32'h3c13f2c5),
	.w7(32'h3ab4d2c5),
	.w8(32'h3aae2cc9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe440e),
	.w1(32'h3c64172e),
	.w2(32'h3c024796),
	.w3(32'h3b6fb718),
	.w4(32'h3c81e0a7),
	.w5(32'h3b177ba5),
	.w6(32'h3c23c2f4),
	.w7(32'h39d88e9e),
	.w8(32'h3bd1eff2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b391633),
	.w1(32'h3ab4cd20),
	.w2(32'h3a949250),
	.w3(32'h3a89ce62),
	.w4(32'h3b9f1869),
	.w5(32'h3bc64992),
	.w6(32'h3b678d31),
	.w7(32'h3a9e2d5a),
	.w8(32'h37b276ff),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77c94d),
	.w1(32'h3b611aad),
	.w2(32'h3be34257),
	.w3(32'h3b847179),
	.w4(32'h3c36f067),
	.w5(32'h3bc02fc7),
	.w6(32'h3c51d01d),
	.w7(32'h3bf79cf8),
	.w8(32'h3c5405a4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf60d42),
	.w1(32'h3ba236e8),
	.w2(32'h3b016106),
	.w3(32'h3c04d209),
	.w4(32'h3b62472a),
	.w5(32'h3a83b998),
	.w6(32'h3bb9175b),
	.w7(32'h3a819c44),
	.w8(32'hbb60ed1c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7e36e),
	.w1(32'hb9cbe9a3),
	.w2(32'hbb74f3fa),
	.w3(32'h3b7cfb84),
	.w4(32'h3b587386),
	.w5(32'hbb84b88b),
	.w6(32'h3c0fa268),
	.w7(32'h3bac45c5),
	.w8(32'h3bb68103),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85a5f6),
	.w1(32'hbc08686a),
	.w2(32'hbbffe06f),
	.w3(32'hba601d9d),
	.w4(32'h3c14541b),
	.w5(32'h3b3c4867),
	.w6(32'hbb375f11),
	.w7(32'h3b8079c6),
	.w8(32'h3c5925a8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e224b),
	.w1(32'h3c17b861),
	.w2(32'h3bc52ce0),
	.w3(32'h3b285477),
	.w4(32'h3bddee23),
	.w5(32'h3c59ba57),
	.w6(32'h3bc7d12e),
	.w7(32'h3aedc4f9),
	.w8(32'hba4c1296),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f1df2),
	.w1(32'h3936d2c5),
	.w2(32'hbaa07b98),
	.w3(32'h3bf83d65),
	.w4(32'h3af77313),
	.w5(32'hba038839),
	.w6(32'h3be93636),
	.w7(32'hbac17938),
	.w8(32'hbb70bcf9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb3d5e),
	.w1(32'h3b7d2b88),
	.w2(32'h3bce5534),
	.w3(32'hba5fb739),
	.w4(32'h3b686635),
	.w5(32'h3beda156),
	.w6(32'h37a3294a),
	.w7(32'h3b52d39a),
	.w8(32'h3bc34611),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bb8bf),
	.w1(32'hba8948ba),
	.w2(32'h3a085917),
	.w3(32'h3c59e59f),
	.w4(32'h3a392edb),
	.w5(32'h3c016a9a),
	.w6(32'h3b9f887e),
	.w7(32'h3b38a50f),
	.w8(32'h3a88c425),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a3416),
	.w1(32'hbc7e9218),
	.w2(32'hbb20ea92),
	.w3(32'h3b6c59b7),
	.w4(32'hbc6a2b9c),
	.w5(32'hbbe5672d),
	.w6(32'hbc0a4733),
	.w7(32'hbb94c483),
	.w8(32'h3b9a508b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e3bd),
	.w1(32'hbc23615b),
	.w2(32'hbb96308b),
	.w3(32'hbb0d4011),
	.w4(32'hbb06ad58),
	.w5(32'hbb95c22b),
	.w6(32'hbb3ae213),
	.w7(32'h3b1c19c4),
	.w8(32'h39f8cf85),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd6894),
	.w1(32'h3bda192e),
	.w2(32'h3c23fc09),
	.w3(32'hbb1c00b1),
	.w4(32'hbab84954),
	.w5(32'h3c526569),
	.w6(32'h3b95ae32),
	.w7(32'h3b46a164),
	.w8(32'h3bfdb8a3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed54dc),
	.w1(32'hbc692fa4),
	.w2(32'hbcff825a),
	.w3(32'h3c1e7608),
	.w4(32'hbbd157f9),
	.w5(32'hbcb7ea1f),
	.w6(32'hba575f0f),
	.w7(32'hbc413efd),
	.w8(32'hbc04d67b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda631b),
	.w1(32'hbb114935),
	.w2(32'h3bd4f152),
	.w3(32'hbcb430b8),
	.w4(32'hb92275d0),
	.w5(32'h3bf5bf4e),
	.w6(32'hb9e66f3b),
	.w7(32'h3b2e379c),
	.w8(32'h3bf7f45d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c662761),
	.w1(32'hbc2dfb35),
	.w2(32'hbc8ecc9d),
	.w3(32'h3c4e7d7e),
	.w4(32'h3bf3c0ba),
	.w5(32'hbb229a35),
	.w6(32'hbbeeed05),
	.w7(32'hbc1ea41a),
	.w8(32'hbbbec0d3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b0c5e),
	.w1(32'h3ab0b4aa),
	.w2(32'hbad1a7bb),
	.w3(32'hbbcc3485),
	.w4(32'h3b94a654),
	.w5(32'h3993fa3f),
	.w6(32'h3bfc4ae7),
	.w7(32'hb9ba7ce1),
	.w8(32'hbad939ac),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e1669),
	.w1(32'h3b223ee8),
	.w2(32'hba0b9f3c),
	.w3(32'h3b6ea493),
	.w4(32'h3b8d9b24),
	.w5(32'h3c167b76),
	.w6(32'h3ba02c98),
	.w7(32'h3ae97e21),
	.w8(32'hbb3169d3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb876d9f),
	.w1(32'hbc83a402),
	.w2(32'hbcb10acf),
	.w3(32'h3bcb227e),
	.w4(32'hbc4bbefc),
	.w5(32'hbc76d217),
	.w6(32'hbba5c59a),
	.w7(32'hbc21f5e5),
	.w8(32'hbbbd9594),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc887419),
	.w1(32'h3c2121c3),
	.w2(32'h3bd93e9a),
	.w3(32'hbbf73949),
	.w4(32'h3c1c02af),
	.w5(32'h3c2ab640),
	.w6(32'h3acc256b),
	.w7(32'hba065cbc),
	.w8(32'h3ba6ffee),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb54913),
	.w1(32'h3ba5febe),
	.w2(32'hbb9f8b19),
	.w3(32'h3c611e40),
	.w4(32'h3bb4cc7c),
	.w5(32'hbb916c09),
	.w6(32'h3bc2a5a1),
	.w7(32'h3b93666f),
	.w8(32'hbc05bfb4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4aba5c),
	.w1(32'hbb7e4432),
	.w2(32'hbab7a71a),
	.w3(32'hbc5907de),
	.w4(32'hbb267c0c),
	.w5(32'h3b17906e),
	.w6(32'hbb187dea),
	.w7(32'h3a0a2807),
	.w8(32'hbb6c26ac),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc316c91),
	.w1(32'hbbb9dbb7),
	.w2(32'hb9530c83),
	.w3(32'hbbc42e34),
	.w4(32'hbb4e0440),
	.w5(32'hba069a3d),
	.w6(32'h3ac68e33),
	.w7(32'hbb980d8f),
	.w8(32'hbbbb33e3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a5688),
	.w1(32'hbb1c890a),
	.w2(32'hbbc70f1c),
	.w3(32'hbb5402ae),
	.w4(32'h3c488098),
	.w5(32'h3c3e0972),
	.w6(32'hbb313ff4),
	.w7(32'h3a455a7c),
	.w8(32'hbb511805),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb37409),
	.w1(32'h3b3129f9),
	.w2(32'hbb6ddf56),
	.w3(32'h3afc55c2),
	.w4(32'h3c0e2308),
	.w5(32'h3b14f68a),
	.w6(32'hbb1b706e),
	.w7(32'hbb64ae06),
	.w8(32'hbba184f7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bbcdc),
	.w1(32'h3c5120d2),
	.w2(32'h3d169cdd),
	.w3(32'h3b1eaa18),
	.w4(32'h3c026f6b),
	.w5(32'h3ca3e01d),
	.w6(32'h3ad390ea),
	.w7(32'h3baa4639),
	.w8(32'hbbc39bb2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b978b26),
	.w1(32'h3c3742a4),
	.w2(32'h3c8cf4e1),
	.w3(32'hba0eeebb),
	.w4(32'h3b3e3d01),
	.w5(32'h3c41ae0f),
	.w6(32'h3bf27c1b),
	.w7(32'h3c4cf82b),
	.w8(32'hbb93c79d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule