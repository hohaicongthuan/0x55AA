module layer_6_featuremap_102(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9c42e),
	.w1(32'hba39194e),
	.w2(32'hbba07eb6),
	.w3(32'hbbadbc6d),
	.w4(32'hbb81fdf4),
	.w5(32'hbb7fa1a8),
	.w6(32'h3ba03465),
	.w7(32'h3bbb34a7),
	.w8(32'h3bd804c8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2b030),
	.w1(32'hbbffab6d),
	.w2(32'hbb8ce0a7),
	.w3(32'hba9d042a),
	.w4(32'h3b0ece55),
	.w5(32'h3b70c28a),
	.w6(32'h3be48be5),
	.w7(32'h3c0ad56b),
	.w8(32'h3c00ae1d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47b14f),
	.w1(32'hbcc6afdd),
	.w2(32'hbbb2a50b),
	.w3(32'hbc9e9f75),
	.w4(32'hbb8de209),
	.w5(32'hbb0faca1),
	.w6(32'h3c4b5c35),
	.w7(32'h3c6c0e9a),
	.w8(32'h3cc2d982),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8daeb5),
	.w1(32'h3bfe3302),
	.w2(32'h3b91705c),
	.w3(32'h3bd18832),
	.w4(32'h3bbe3b1d),
	.w5(32'h3b427b39),
	.w6(32'h3b386f88),
	.w7(32'h3b018030),
	.w8(32'hbabc3892),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9244d9e),
	.w1(32'hbc98a977),
	.w2(32'hbc3bae20),
	.w3(32'hbc502d5a),
	.w4(32'hbc7ebc47),
	.w5(32'hbce2bb41),
	.w6(32'h3cd8ceed),
	.w7(32'h3d56fb7b),
	.w8(32'h3d4993cf),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca72dbb),
	.w1(32'hba404924),
	.w2(32'hbb84de78),
	.w3(32'hbae323cb),
	.w4(32'hbb034690),
	.w5(32'hbac0252f),
	.w6(32'h3b8911e3),
	.w7(32'h3ba71109),
	.w8(32'h3b90d5d0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188d2f),
	.w1(32'h3a282020),
	.w2(32'h3b4655c3),
	.w3(32'h3b10e267),
	.w4(32'h3b009eb5),
	.w5(32'h3ad935d7),
	.w6(32'hbbb453f0),
	.w7(32'hbb890fe7),
	.w8(32'hbbf3a926),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0375c0),
	.w1(32'hbc85d0b7),
	.w2(32'h3c4d9d6b),
	.w3(32'hbbbbd91c),
	.w4(32'h3b647931),
	.w5(32'h3be7db41),
	.w6(32'h3cab293b),
	.w7(32'hbb8f75f1),
	.w8(32'hbcd3b936),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b947a6b),
	.w1(32'h3d8c312a),
	.w2(32'h3dcb4856),
	.w3(32'h3cde5628),
	.w4(32'h3b1a1dbf),
	.w5(32'h3aafc359),
	.w6(32'hbd3a65ee),
	.w7(32'hbda7b218),
	.w8(32'hbd04e01e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5e616c),
	.w1(32'hbb96f056),
	.w2(32'hbbce8ad1),
	.w3(32'hbac15edd),
	.w4(32'hb89d51cd),
	.w5(32'hba98daf6),
	.w6(32'hbb16853f),
	.w7(32'hbb142af3),
	.w8(32'hbb2173ee),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f53c9),
	.w1(32'hb95ab6f7),
	.w2(32'hbb70c324),
	.w3(32'h3c0cc9ed),
	.w4(32'h3ba5418d),
	.w5(32'h3bbd2bd1),
	.w6(32'h3c54fd1f),
	.w7(32'hbc30a654),
	.w8(32'hba07ffe6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcf2ba),
	.w1(32'h3cb0a88d),
	.w2(32'h3ce55b24),
	.w3(32'hbc297023),
	.w4(32'hbc276ba8),
	.w5(32'hbc94ee98),
	.w6(32'hbbcb67c9),
	.w7(32'hbb775794),
	.w8(32'hbb92ffce),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdab05b),
	.w1(32'h3a0e1f8f),
	.w2(32'h3baffee0),
	.w3(32'h3a519c2d),
	.w4(32'h3b816e51),
	.w5(32'h3b314241),
	.w6(32'hb9e7e7c1),
	.w7(32'h3b2125f0),
	.w8(32'h3a16de5c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02c1ab),
	.w1(32'h3bd6cbe7),
	.w2(32'h3ca86c51),
	.w3(32'h3b175e6a),
	.w4(32'h3c9653de),
	.w5(32'h3c1ee189),
	.w6(32'h3d6b972a),
	.w7(32'h3dbb5fed),
	.w8(32'h3d464650),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc291298),
	.w1(32'h39b552d5),
	.w2(32'h3b3f8f67),
	.w3(32'hba88e9da),
	.w4(32'hbaba0dd6),
	.w5(32'hbbdf1863),
	.w6(32'hba732cc9),
	.w7(32'hbbe22265),
	.w8(32'hbba6c772),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4b216),
	.w1(32'h3a8f8fc3),
	.w2(32'h3b57cb2b),
	.w3(32'h3ad00961),
	.w4(32'h3a1cd338),
	.w5(32'hbb21abd6),
	.w6(32'h39e0ebc3),
	.w7(32'h3b135ed2),
	.w8(32'h39455d34),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f6386),
	.w1(32'h3b853499),
	.w2(32'hbbafb8cd),
	.w3(32'h3b82d56b),
	.w4(32'hbc18652d),
	.w5(32'hbad62561),
	.w6(32'hbc41d1d5),
	.w7(32'hbbddf8f4),
	.w8(32'hbbd76e14),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7964cc),
	.w1(32'hbb8f2d24),
	.w2(32'hbbb6d59a),
	.w3(32'h3b07e02c),
	.w4(32'h3b273f58),
	.w5(32'h3b093628),
	.w6(32'hbbb0a0ec),
	.w7(32'hbbd9e360),
	.w8(32'hbb65dfff),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b749d),
	.w1(32'hbb7101c9),
	.w2(32'hbbb2670a),
	.w3(32'h3a1db5e9),
	.w4(32'hba09f47b),
	.w5(32'hbaa0e7fe),
	.w6(32'hba460603),
	.w7(32'hba068aea),
	.w8(32'hbb4d7fa5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3d76e),
	.w1(32'hbbc00209),
	.w2(32'hbb7e1840),
	.w3(32'hbbe6da23),
	.w4(32'hbb87191f),
	.w5(32'hb9a2a2cb),
	.w6(32'hbb43224a),
	.w7(32'hbbf4876d),
	.w8(32'hbb44807d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc324e87),
	.w1(32'hbb36fffb),
	.w2(32'hbb2c5956),
	.w3(32'hb79cfc49),
	.w4(32'hb9c17d69),
	.w5(32'hb993fd37),
	.w6(32'hba94ae3f),
	.w7(32'hbb0399b4),
	.w8(32'hbadfe627),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df335b),
	.w1(32'h3b0111e7),
	.w2(32'h3ba1c026),
	.w3(32'h3b138cf0),
	.w4(32'hbb4044f8),
	.w5(32'hb91c451d),
	.w6(32'h3b11b4df),
	.w7(32'hbb1ae22b),
	.w8(32'h3b30620b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba136452),
	.w1(32'h3a95acde),
	.w2(32'hbc16cc48),
	.w3(32'hbc9cd0cd),
	.w4(32'hbbc80c3a),
	.w5(32'hbb8f2aab),
	.w6(32'h3bdf3322),
	.w7(32'hbad90737),
	.w8(32'h3bb6b8b4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4284c3),
	.w1(32'hbaf2e01f),
	.w2(32'h3c2ec1e6),
	.w3(32'hbb87abed),
	.w4(32'h3bd8ac69),
	.w5(32'h3c99612a),
	.w6(32'hbb1400b0),
	.w7(32'hbb95d753),
	.w8(32'hbc12a469),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba606c9e),
	.w1(32'hbb75b54b),
	.w2(32'h3c9b6f2a),
	.w3(32'h3b5fccff),
	.w4(32'h3cbcaf33),
	.w5(32'h3ce486b1),
	.w6(32'h3ca8e5ad),
	.w7(32'h3d2e7d3d),
	.w8(32'h3cdaaa38),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfdbc3a),
	.w1(32'h3c32c5f5),
	.w2(32'hbc4223e7),
	.w3(32'hb9d16d4f),
	.w4(32'hbc0eb797),
	.w5(32'h3ad7615e),
	.w6(32'hbbf05e90),
	.w7(32'hbc50b540),
	.w8(32'hbc32e062),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7dbb5),
	.w1(32'h3c802acb),
	.w2(32'h3c1d7ea9),
	.w3(32'h3b8b0725),
	.w4(32'hbb40b728),
	.w5(32'hbacbf078),
	.w6(32'h3c255740),
	.w7(32'h3c7fc817),
	.w8(32'h3b597ac4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c200d4f),
	.w1(32'hbb196dd2),
	.w2(32'hb9de411d),
	.w3(32'h3b5d2b68),
	.w4(32'h3bb9cc67),
	.w5(32'h3bf84f46),
	.w6(32'hba74ae64),
	.w7(32'hb88f3a3a),
	.w8(32'hbb2317ff),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d3c70),
	.w1(32'h3b675290),
	.w2(32'h3aa356f4),
	.w3(32'h3b126bf8),
	.w4(32'hba88bb4f),
	.w5(32'hba2eb516),
	.w6(32'h3bbc6b48),
	.w7(32'h3b307185),
	.w8(32'h3b933435),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebc9ef),
	.w1(32'hb9eca758),
	.w2(32'h3cad817d),
	.w3(32'h3b4e7dad),
	.w4(32'h3c6cadeb),
	.w5(32'hb963eef6),
	.w6(32'hbbe3f3bc),
	.w7(32'hbcb627e8),
	.w8(32'hbbd4ea73),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47adbf),
	.w1(32'hbc2b59a1),
	.w2(32'h3c984ccb),
	.w3(32'h3b828d7e),
	.w4(32'h3c443928),
	.w5(32'h3bc0bbbf),
	.w6(32'h3c3cd490),
	.w7(32'h3c15e110),
	.w8(32'hba3b222f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86c54b),
	.w1(32'hbbfda023),
	.w2(32'h3c23fd86),
	.w3(32'h3c559139),
	.w4(32'h3c9fbb0d),
	.w5(32'h3c43645b),
	.w6(32'hbcd6bf7b),
	.w7(32'hbd097627),
	.w8(32'hbcc38b2e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca17622),
	.w1(32'hbc699f7f),
	.w2(32'hbaec5633),
	.w3(32'h3c8c8c0c),
	.w4(32'h3c107425),
	.w5(32'h3bde4a24),
	.w6(32'hbc9c5fe9),
	.w7(32'hbd01449c),
	.w8(32'hbca17811),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06a89b),
	.w1(32'h3cbbd3e2),
	.w2(32'h3a35ba6c),
	.w3(32'h3c221440),
	.w4(32'h3b5ee15d),
	.w5(32'h3c43fe24),
	.w6(32'hbc445139),
	.w7(32'hbc067ea1),
	.w8(32'hba9e384d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e5988),
	.w1(32'hbb9aa63c),
	.w2(32'hbb696989),
	.w3(32'h3a892590),
	.w4(32'h3aa7088e),
	.w5(32'h3abe16fc),
	.w6(32'hba4a858d),
	.w7(32'hbb25f490),
	.w8(32'h3b0aad7a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a543b5c),
	.w1(32'h3be93780),
	.w2(32'h3c696902),
	.w3(32'h3a811aea),
	.w4(32'hbbd8c2c5),
	.w5(32'hbc09241a),
	.w6(32'h3b55d8d5),
	.w7(32'h3b3499d9),
	.w8(32'h3b677788),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c215a03),
	.w1(32'hba2f266f),
	.w2(32'hbbdb375e),
	.w3(32'hba9808b0),
	.w4(32'hba0435b4),
	.w5(32'h3ae7281e),
	.w6(32'h3b0b5ec2),
	.w7(32'h3bce6d03),
	.w8(32'h3b53924b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb547a1d),
	.w1(32'h3b42775e),
	.w2(32'h3930f217),
	.w3(32'h3b69a80c),
	.w4(32'h3b0b2ac4),
	.w5(32'h3b77a458),
	.w6(32'h3b133497),
	.w7(32'h3b436bb1),
	.w8(32'h3b95dbc2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a466b39),
	.w1(32'hbc21e293),
	.w2(32'hbc345a08),
	.w3(32'hbbf93759),
	.w4(32'h3b130daf),
	.w5(32'h3ca4576f),
	.w6(32'hbd0ee96b),
	.w7(32'hbd467395),
	.w8(32'hbd2fbf03),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91ece7),
	.w1(32'hbc176338),
	.w2(32'h3c1551c5),
	.w3(32'h3cd0ed6e),
	.w4(32'h3a81daeb),
	.w5(32'hbbda357b),
	.w6(32'hbca76bb0),
	.w7(32'hbc0a6b2e),
	.w8(32'h3c351615),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67793d),
	.w1(32'hbcc39ee7),
	.w2(32'hbc0e1703),
	.w3(32'h3b90617d),
	.w4(32'h3b188f21),
	.w5(32'h3c1de7e6),
	.w6(32'hbab37239),
	.w7(32'hbc2e262d),
	.w8(32'hbca14f08),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca850b),
	.w1(32'h3a0faf54),
	.w2(32'hba0a2e2a),
	.w3(32'h39b468ed),
	.w4(32'h3ac9d3dd),
	.w5(32'hbab6c2d5),
	.w6(32'hb99e6027),
	.w7(32'h3a81880f),
	.w8(32'hbafaf3d7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904ff9a),
	.w1(32'h3b21e5cf),
	.w2(32'hbaf7b233),
	.w3(32'h3b051046),
	.w4(32'h3bee49d2),
	.w5(32'h3a0a6ec2),
	.w6(32'hbb6abc87),
	.w7(32'hbbff4c33),
	.w8(32'hbbc22092),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c4dff),
	.w1(32'h3b45bec4),
	.w2(32'h3bdff1bb),
	.w3(32'hbb0f64bb),
	.w4(32'hbb227c62),
	.w5(32'hbb39192b),
	.w6(32'h3aff770e),
	.w7(32'h3c5d0844),
	.w8(32'h3c2f25ff),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1b4d3),
	.w1(32'hbb22ec2e),
	.w2(32'hbb55f079),
	.w3(32'hbb653849),
	.w4(32'hbb6f79e7),
	.w5(32'hbc10fb91),
	.w6(32'hbba1829e),
	.w7(32'hbb4901e9),
	.w8(32'hbba6a50e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff8ddf),
	.w1(32'hbc63491b),
	.w2(32'hbc42238d),
	.w3(32'hbbbc926b),
	.w4(32'hbc3ae42c),
	.w5(32'hbbe32ee3),
	.w6(32'hb99bd45f),
	.w7(32'hbc2dd64b),
	.w8(32'hbc19190d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86220b),
	.w1(32'hbc79740b),
	.w2(32'hbbce50e2),
	.w3(32'h3b715fc3),
	.w4(32'h3c31943f),
	.w5(32'h3c919d29),
	.w6(32'hbbdadfd4),
	.w7(32'hbbcf1705),
	.w8(32'hba581140),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c015d18),
	.w1(32'h3c496c0b),
	.w2(32'h3b8bff4b),
	.w3(32'h3c0bcb94),
	.w4(32'h3bd58d00),
	.w5(32'hba34dc9d),
	.w6(32'h3c0967b9),
	.w7(32'hbb2ca312),
	.w8(32'hba8df3d8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee7057),
	.w1(32'h3b921edb),
	.w2(32'h3b541146),
	.w3(32'h3aadc10f),
	.w4(32'h3a1f8f06),
	.w5(32'hb9fe0298),
	.w6(32'hb98a50f8),
	.w7(32'hbad258d1),
	.w8(32'hbb056217),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be32850),
	.w1(32'hbd9bed21),
	.w2(32'hbded8e01),
	.w3(32'hbba42cf2),
	.w4(32'hbba78364),
	.w5(32'h3ba1b352),
	.w6(32'h3d2b6fb0),
	.w7(32'h3d8a0009),
	.w8(32'h3d47770b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7fd4e8),
	.w1(32'h3aef73c2),
	.w2(32'h3b8cc390),
	.w3(32'hbaecf769),
	.w4(32'h3af9a3e9),
	.w5(32'hbb436f4c),
	.w6(32'hb9a494d9),
	.w7(32'hba0a1ace),
	.w8(32'hbbf7e6e4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa05dcc),
	.w1(32'hbb7d3fdf),
	.w2(32'hba10c4ce),
	.w3(32'hbb9c7989),
	.w4(32'hbb39a22c),
	.w5(32'h3bd92042),
	.w6(32'hbbd6d1a4),
	.w7(32'hbb0ef20e),
	.w8(32'h3b953e4f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e5bc7),
	.w1(32'hbac722da),
	.w2(32'h3a8632ad),
	.w3(32'h3b0ae3af),
	.w4(32'hba7dbff2),
	.w5(32'hb8c5835f),
	.w6(32'hbac2910a),
	.w7(32'hbb283392),
	.w8(32'hbb719193),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee6932),
	.w1(32'h3a906d7f),
	.w2(32'h3b136141),
	.w3(32'hbbc7744d),
	.w4(32'hbb85d2d6),
	.w5(32'hbb872c3c),
	.w6(32'hbbded8a7),
	.w7(32'hbbd93049),
	.w8(32'hbbe95860),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31fd46),
	.w1(32'h3b50405d),
	.w2(32'h3b37c4fc),
	.w3(32'hba9796ea),
	.w4(32'h3ab34a44),
	.w5(32'hba3ec68f),
	.w6(32'hbbc0e520),
	.w7(32'hbbfa37c5),
	.w8(32'hbc26cb6a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81fe18),
	.w1(32'hbb72fc7c),
	.w2(32'hbb9d29bf),
	.w3(32'h3b9fda75),
	.w4(32'h3b5fa3c5),
	.w5(32'hbb765e99),
	.w6(32'h3c9c9f03),
	.w7(32'h3d55761f),
	.w8(32'h3ca5868c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff97ab),
	.w1(32'hbbb249a7),
	.w2(32'hbbb2c776),
	.w3(32'hbb9df84d),
	.w4(32'hbbbf8dfc),
	.w5(32'hbbc00c82),
	.w6(32'hbc1b70f8),
	.w7(32'hbc35fa45),
	.w8(32'hbc3349ec),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f0e8b),
	.w1(32'hbc0e744c),
	.w2(32'hbc88d3b4),
	.w3(32'hbc2eed97),
	.w4(32'hbba2a0fd),
	.w5(32'h3a2422b9),
	.w6(32'hbc9b1195),
	.w7(32'hbbd7aef2),
	.w8(32'hbcafdb7a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f896d),
	.w1(32'hbbdde741),
	.w2(32'hbc0a71f2),
	.w3(32'hbc09dc27),
	.w4(32'hbc2c22b1),
	.w5(32'hbc6146f6),
	.w6(32'hbbb7eb8d),
	.w7(32'hbc07f535),
	.w8(32'hbbeb07d6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1be0d),
	.w1(32'h3cb1790c),
	.w2(32'h3af6cac2),
	.w3(32'hbb0e4f84),
	.w4(32'h3c5cdca4),
	.w5(32'h3c2f0f25),
	.w6(32'hb9bccbdb),
	.w7(32'hbc63ca58),
	.w8(32'hbccdad4b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35bd5c),
	.w1(32'h3a5acd8d),
	.w2(32'hbc31e5ca),
	.w3(32'h3c113730),
	.w4(32'hbb778978),
	.w5(32'hbc1f6d21),
	.w6(32'hbbf1e26a),
	.w7(32'hbc6bbf7f),
	.w8(32'hbc969635),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbc122),
	.w1(32'h3bbff12b),
	.w2(32'h3c107009),
	.w3(32'h3ba25744),
	.w4(32'hbb4e9538),
	.w5(32'hbbb1c559),
	.w6(32'hbbfe84d1),
	.w7(32'hbbe8b6ec),
	.w8(32'hbc4a4930),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03e6a4),
	.w1(32'h3c585b45),
	.w2(32'h3cc83b81),
	.w3(32'h3c964658),
	.w4(32'h3d3a372b),
	.w5(32'h3d2178f4),
	.w6(32'hbc76fed7),
	.w7(32'hbd42f9d2),
	.w8(32'hbd4ecd78),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc13434),
	.w1(32'hbc41bacb),
	.w2(32'hbc9e8f8e),
	.w3(32'hbbb9bc7d),
	.w4(32'hbc17a396),
	.w5(32'hbc4dcf4e),
	.w6(32'hbb4852b9),
	.w7(32'hbb0072de),
	.w8(32'hbc2a7016),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule