module layer_10_featuremap_9(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12b03c),
	.w1(32'h3ac0a32f),
	.w2(32'h3bc101ef),
	.w3(32'hbc0774d4),
	.w4(32'hbbf6d00b),
	.w5(32'h3bc1b8b6),
	.w6(32'h39809898),
	.w7(32'hbb54dca1),
	.w8(32'hba999f3c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b424ade),
	.w1(32'h3a35fd5c),
	.w2(32'h3bebe63e),
	.w3(32'hbb065be5),
	.w4(32'hb8ddc9ee),
	.w5(32'hbbb6a324),
	.w6(32'hbc9399be),
	.w7(32'hbc0cd86a),
	.w8(32'hbc3d39c3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c230849),
	.w1(32'h3bbdee0c),
	.w2(32'h3bee45f9),
	.w3(32'hbc46acef),
	.w4(32'hbc1830d3),
	.w5(32'h3b2afa13),
	.w6(32'hbc283d8b),
	.w7(32'hbb32597a),
	.w8(32'hbc05af75),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ba9b4),
	.w1(32'h39ea00d4),
	.w2(32'hbb995dc2),
	.w3(32'hb9ac6ac6),
	.w4(32'hbbae8287),
	.w5(32'hb9a386be),
	.w6(32'hbb860532),
	.w7(32'h3c543e20),
	.w8(32'h3ba89436),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6f3d8),
	.w1(32'h3b4d1d78),
	.w2(32'h3b754dad),
	.w3(32'hbb7e3c3b),
	.w4(32'hbc0508a1),
	.w5(32'hbb6f5ccc),
	.w6(32'h395464a1),
	.w7(32'h398fb400),
	.w8(32'h3aa9e1fe),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23b70d),
	.w1(32'h3b9de5de),
	.w2(32'hbc157c20),
	.w3(32'hba922bbb),
	.w4(32'h3b160d1a),
	.w5(32'hbaa10dda),
	.w6(32'hbae41d90),
	.w7(32'h3a3b05a3),
	.w8(32'h3b4f3fb2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd49ed6),
	.w1(32'hbb80f350),
	.w2(32'hbb575ab4),
	.w3(32'h3b05267d),
	.w4(32'h3b934876),
	.w5(32'hbb59c670),
	.w6(32'h3c3dc9f8),
	.w7(32'h3c02f2fa),
	.w8(32'hbc43916f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f000),
	.w1(32'hbba2cab2),
	.w2(32'hbc540982),
	.w3(32'hbba385a0),
	.w4(32'hbc2a1374),
	.w5(32'h3a85a134),
	.w6(32'hbc445e47),
	.w7(32'hbc68f982),
	.w8(32'hbb2596fc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17e70b),
	.w1(32'hbb4dab2f),
	.w2(32'hbaecd65b),
	.w3(32'h3a99ed04),
	.w4(32'h3a7b8d69),
	.w5(32'hbbaec16d),
	.w6(32'hbaf1d135),
	.w7(32'hbb1bca42),
	.w8(32'hbb634eff),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982d82),
	.w1(32'hbb20a89d),
	.w2(32'hbbbadbbd),
	.w3(32'h3bdfa020),
	.w4(32'hb9c89d78),
	.w5(32'hbb5dcfa3),
	.w6(32'h3b22005c),
	.w7(32'h3bb025e5),
	.w8(32'hbb6cabec),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387da090),
	.w1(32'h3af884f6),
	.w2(32'hbad7f1ce),
	.w3(32'h37a1326d),
	.w4(32'h3afc1b99),
	.w5(32'h3c1e82ca),
	.w6(32'h3b4d0883),
	.w7(32'h3b5862c7),
	.w8(32'hbc81654a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29d29d),
	.w1(32'h3be777d8),
	.w2(32'h3a53c4e3),
	.w3(32'h3bf0bb13),
	.w4(32'h3c1ff5f0),
	.w5(32'h3c0b29bf),
	.w6(32'hba369648),
	.w7(32'h3c96eea0),
	.w8(32'h3b898dd9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c39ee),
	.w1(32'h3bf09b79),
	.w2(32'hbb65d20d),
	.w3(32'h3c82e196),
	.w4(32'h3c19017f),
	.w5(32'h3abe7359),
	.w6(32'h3c1b4991),
	.w7(32'h3ba9c2fa),
	.w8(32'hbbc1c94f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b485941),
	.w1(32'hbb04c429),
	.w2(32'hbc5cd512),
	.w3(32'hba43b4bd),
	.w4(32'hbc06237e),
	.w5(32'h3b6bbf0b),
	.w6(32'h3b366aa7),
	.w7(32'hba2b37db),
	.w8(32'h3a1d3ea8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c217b),
	.w1(32'hbbbe7179),
	.w2(32'hbc097d98),
	.w3(32'h3b9efb32),
	.w4(32'h3adbc741),
	.w5(32'hbb777539),
	.w6(32'h3c2b4bce),
	.w7(32'h3b8d52d5),
	.w8(32'hbc05478b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a252fb3),
	.w1(32'hba7832be),
	.w2(32'hbc1c81c3),
	.w3(32'h3b5f519d),
	.w4(32'hbaff52de),
	.w5(32'hbc0b1c56),
	.w6(32'h3afedbb2),
	.w7(32'hba329b35),
	.w8(32'hbbd2bb42),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d04572),
	.w1(32'h3a36b8d4),
	.w2(32'h3b228287),
	.w3(32'hbb4d8ba1),
	.w4(32'hbb059282),
	.w5(32'hbc00aa6c),
	.w6(32'h3af4a966),
	.w7(32'h3a8692f7),
	.w8(32'hbc34f73d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0930bb),
	.w1(32'h3bfbbe33),
	.w2(32'hbc020cc9),
	.w3(32'h3c495463),
	.w4(32'h3b91ed48),
	.w5(32'h3b22f68e),
	.w6(32'h3ca5116a),
	.w7(32'h3c05cc3c),
	.w8(32'h3bb5633a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4889e),
	.w1(32'h3b75e027),
	.w2(32'hbbf70046),
	.w3(32'h3bbc6e4d),
	.w4(32'h3bb54894),
	.w5(32'h3b6cf844),
	.w6(32'h3c72dcf6),
	.w7(32'h3c3d4a8f),
	.w8(32'hb87182a6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5eed4c),
	.w1(32'hbbcfa7ce),
	.w2(32'h3b1ec61a),
	.w3(32'hbbc30cd6),
	.w4(32'hbba27e0b),
	.w5(32'h3b7ec771),
	.w6(32'hbb3682ef),
	.w7(32'h3a58f859),
	.w8(32'h3b0130b7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb0214),
	.w1(32'h3a786120),
	.w2(32'h3ba21681),
	.w3(32'h3b2d5916),
	.w4(32'h3b40c9b4),
	.w5(32'hbb893a4f),
	.w6(32'h39ba8441),
	.w7(32'hbae3dd6d),
	.w8(32'h3c8936b4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c120e17),
	.w1(32'h3c2048b7),
	.w2(32'hbbeb357b),
	.w3(32'hbc41c0d2),
	.w4(32'hbb659654),
	.w5(32'h3ba6152c),
	.w6(32'h3c6487a8),
	.w7(32'h3c04aca1),
	.w8(32'h3b395c0b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f16c3),
	.w1(32'h3a6d551d),
	.w2(32'hbc41e174),
	.w3(32'h3c3a436c),
	.w4(32'h3cb9dc68),
	.w5(32'hbb50e7de),
	.w6(32'h3cd81619),
	.w7(32'h3ca49f1e),
	.w8(32'hbbff13aa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f23b),
	.w1(32'h39b5fbef),
	.w2(32'hbbdcbd98),
	.w3(32'h3b386abb),
	.w4(32'h3b9481be),
	.w5(32'hbb38d298),
	.w6(32'hbb2b3a4a),
	.w7(32'hbc064ad7),
	.w8(32'hbb591462),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3542f6),
	.w1(32'hbb54b429),
	.w2(32'h3c8862b3),
	.w3(32'h3a6f32ee),
	.w4(32'h3b9b4bb3),
	.w5(32'hbbc46407),
	.w6(32'hba81b09f),
	.w7(32'hba8a0770),
	.w8(32'hbbadf9e8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8fe5f),
	.w1(32'h3b852503),
	.w2(32'hbbe383bc),
	.w3(32'hbc1324d6),
	.w4(32'hbb1ac77c),
	.w5(32'hbc287054),
	.w6(32'h3b8970bc),
	.w7(32'h3bd30e82),
	.w8(32'h3bf4c931),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc2ed5),
	.w1(32'h3b0beff3),
	.w2(32'h3a716ac4),
	.w3(32'hbc142da8),
	.w4(32'hbbe4f3da),
	.w5(32'h3abbafba),
	.w6(32'h3bbf66e7),
	.w7(32'hb9f2c388),
	.w8(32'h3a3f88d7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b360846),
	.w1(32'h3bfb79a2),
	.w2(32'h3b0abedd),
	.w3(32'h3b717d4c),
	.w4(32'h3b9505d6),
	.w5(32'h3c1db7ad),
	.w6(32'hba2278b1),
	.w7(32'h3a45b3b8),
	.w8(32'h3c0457bc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6ea93),
	.w1(32'h3c837be1),
	.w2(32'hba21e8ab),
	.w3(32'h3bc701df),
	.w4(32'h3a823fb2),
	.w5(32'hbc53d998),
	.w6(32'hbc60ed52),
	.w7(32'h3b9e6462),
	.w8(32'h3b416921),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc155975),
	.w1(32'hbbc2b802),
	.w2(32'hbc1720f9),
	.w3(32'hbc4defab),
	.w4(32'hbb7934bb),
	.w5(32'hbc102d36),
	.w6(32'hbc42bb6f),
	.w7(32'hbc25b73b),
	.w8(32'hbc458497),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f32eae),
	.w1(32'hbb32e34e),
	.w2(32'hbc2cb0c6),
	.w3(32'hba6c7c45),
	.w4(32'hbb0b170d),
	.w5(32'hbc3149d8),
	.w6(32'hbb81c2d1),
	.w7(32'hbb19c99d),
	.w8(32'hbc539fd2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99e515),
	.w1(32'hbc524b1a),
	.w2(32'hbc837bf2),
	.w3(32'hbce75f6d),
	.w4(32'hbca953a0),
	.w5(32'h3b484068),
	.w6(32'hbc09e100),
	.w7(32'hbb1cff44),
	.w8(32'hbc43474a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bc908),
	.w1(32'hbba38f3c),
	.w2(32'hbbc8bbb1),
	.w3(32'hbb426c24),
	.w4(32'hbc8dc970),
	.w5(32'hbb886c30),
	.w6(32'hbca42faa),
	.w7(32'hbbcfea4b),
	.w8(32'hbc35bc75),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f63d96),
	.w1(32'h3bf86b2a),
	.w2(32'h3bd951c0),
	.w3(32'h3baf3905),
	.w4(32'h3adf19a5),
	.w5(32'h3c220dcc),
	.w6(32'hbc2705f1),
	.w7(32'hbc226496),
	.w8(32'hbc3caa28),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccac641),
	.w1(32'hbbb5b054),
	.w2(32'h3ab89eaa),
	.w3(32'hbc25f417),
	.w4(32'hb9e607bb),
	.w5(32'h3b836f7a),
	.w6(32'h3c391a12),
	.w7(32'h3d205ebf),
	.w8(32'hbba11d64),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2974d7),
	.w1(32'h3bfc66f4),
	.w2(32'hbb802f5a),
	.w3(32'h3c1725c6),
	.w4(32'h3b431a8a),
	.w5(32'h3b0f7e46),
	.w6(32'h3bbd1973),
	.w7(32'h3bbf689b),
	.w8(32'h3ad61723),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac54a2),
	.w1(32'h3c0bd62b),
	.w2(32'hbc61a7b9),
	.w3(32'hbc81b552),
	.w4(32'h3c1cc673),
	.w5(32'h3a89e659),
	.w6(32'h3d4bbdf7),
	.w7(32'h3d54a07e),
	.w8(32'h3a60f452),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc004659),
	.w1(32'h3c2e5226),
	.w2(32'h3c518b13),
	.w3(32'hbb8c1450),
	.w4(32'h3b5feea1),
	.w5(32'h3c07f8bb),
	.w6(32'hbce07fbb),
	.w7(32'hba71245c),
	.w8(32'h3b869d0d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaab336),
	.w1(32'h3b398cf3),
	.w2(32'h38fecdf7),
	.w3(32'h3cc5b8b6),
	.w4(32'h3c44a6c8),
	.w5(32'h3c00d29a),
	.w6(32'hbd0a604b),
	.w7(32'hbcecefb4),
	.w8(32'h3a94956a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e9247),
	.w1(32'h3bdbf28c),
	.w2(32'hbb734eda),
	.w3(32'hbb617c2f),
	.w4(32'hbbde71c6),
	.w5(32'hbb188d21),
	.w6(32'hbc9d8050),
	.w7(32'hbc78476b),
	.w8(32'hbb873c4f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb209fe9),
	.w1(32'h3b74c416),
	.w2(32'hbbfc3e04),
	.w3(32'h3ac2429f),
	.w4(32'h3a8888f0),
	.w5(32'hbc0bd689),
	.w6(32'hbbbffb90),
	.w7(32'hbc781501),
	.w8(32'h3c6dfd60),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e27d7),
	.w1(32'hbb58b891),
	.w2(32'h3a91a0f1),
	.w3(32'h3c4a6638),
	.w4(32'h3c515301),
	.w5(32'hba87e32f),
	.w6(32'hbbdfd470),
	.w7(32'hbc8ab925),
	.w8(32'h3bd82fb4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e8e27),
	.w1(32'h3a28fad1),
	.w2(32'hbaec0134),
	.w3(32'hbb2207ad),
	.w4(32'h3beed473),
	.w5(32'h3b82d1d6),
	.w6(32'h3b13facc),
	.w7(32'h3c27617a),
	.w8(32'h3a976d8d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c61bb),
	.w1(32'hbb5b6543),
	.w2(32'h3a1d7972),
	.w3(32'h3bed3d2a),
	.w4(32'hbbc5a2aa),
	.w5(32'hbc2f7864),
	.w6(32'h3b3e9af1),
	.w7(32'hbb1ffc21),
	.w8(32'hbc15b213),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d0736),
	.w1(32'h3ac21544),
	.w2(32'hbc167ed5),
	.w3(32'h3bacc5e7),
	.w4(32'h3c773e6e),
	.w5(32'hbb88fe9c),
	.w6(32'hbb831c8d),
	.w7(32'hbbb65403),
	.w8(32'hbb2296fa),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba93c7c),
	.w1(32'h3c74a960),
	.w2(32'hbc929f11),
	.w3(32'h3d295403),
	.w4(32'hbbcd7ec0),
	.w5(32'hbc55d42f),
	.w6(32'hbc7c5c53),
	.w7(32'h3bade09a),
	.w8(32'hbca66aa4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b68aa),
	.w1(32'h3b8b8104),
	.w2(32'hb99fa6a3),
	.w3(32'hbc15176d),
	.w4(32'hbc5b5ed4),
	.w5(32'hbb47a2a9),
	.w6(32'hbc754067),
	.w7(32'h3ba62d2e),
	.w8(32'hbc8c2a6e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caff289),
	.w1(32'hbbaba731),
	.w2(32'hbbfe2127),
	.w3(32'h3b9e6d7c),
	.w4(32'hbb8e8c54),
	.w5(32'h3a6043a5),
	.w6(32'h3d27d8cf),
	.w7(32'h3d69d331),
	.w8(32'h3bd1b258),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa80a9d),
	.w1(32'hbb2894aa),
	.w2(32'h38b6f35a),
	.w3(32'hbb8531a0),
	.w4(32'hbb9fae02),
	.w5(32'h39b8c36e),
	.w6(32'hba83dba2),
	.w7(32'h3b2b28f0),
	.w8(32'hbbc2ffe8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0437e2),
	.w1(32'hbc06d9d6),
	.w2(32'hbb19aeea),
	.w3(32'h3c69576e),
	.w4(32'hbb07506f),
	.w5(32'h3aba714a),
	.w6(32'hbbd9ddd3),
	.w7(32'hbc888c70),
	.w8(32'h396523bd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29cf14),
	.w1(32'hbbc46e86),
	.w2(32'h3b405871),
	.w3(32'h3c03b7df),
	.w4(32'h3cf687b2),
	.w5(32'hbc4b3250),
	.w6(32'h3c88ceff),
	.w7(32'h3b670a5b),
	.w8(32'h3c70de38),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d9a0e),
	.w1(32'hbc0fbeb3),
	.w2(32'hbc188e8c),
	.w3(32'h3b10a0db),
	.w4(32'h3d4ee0c7),
	.w5(32'hbc82bfc7),
	.w6(32'h3d276560),
	.w7(32'hb9601ece),
	.w8(32'hbc706146),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8f1e6),
	.w1(32'hbc8402d4),
	.w2(32'h3b225c57),
	.w3(32'hbcbd7933),
	.w4(32'h3b4560f9),
	.w5(32'h3b1ce082),
	.w6(32'hbb930777),
	.w7(32'hbc6b7730),
	.w8(32'hbc1c1204),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c572fa7),
	.w1(32'h3be14ab9),
	.w2(32'h38e11ced),
	.w3(32'h3c1eca3c),
	.w4(32'h3c06976c),
	.w5(32'hbca6a90c),
	.w6(32'h3cdf3f38),
	.w7(32'h3c681c2d),
	.w8(32'h3c6cd5e8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d0253),
	.w1(32'hbc19f026),
	.w2(32'h3beebde3),
	.w3(32'h3b2964c2),
	.w4(32'h3cc15b48),
	.w5(32'h3d125779),
	.w6(32'h3c81f7e0),
	.w7(32'hba5156f0),
	.w8(32'hbc820af4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4c25b),
	.w1(32'h3c2a2d9d),
	.w2(32'h3ad8e048),
	.w3(32'h3c0ea5f2),
	.w4(32'hbc577e68),
	.w5(32'hbc1a6534),
	.w6(32'h3cc0a1bc),
	.w7(32'h3d42a69b),
	.w8(32'hbba9f8c2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdede6a),
	.w1(32'hbc51534a),
	.w2(32'h3be65b5a),
	.w3(32'hbc802f1b),
	.w4(32'hbc7029c2),
	.w5(32'h3b477f8d),
	.w6(32'hbc108dfb),
	.w7(32'h3b100589),
	.w8(32'h3b8016c3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8acace),
	.w1(32'hbc0c9b03),
	.w2(32'h3a11e8e9),
	.w3(32'hb8a17e4d),
	.w4(32'hbb88ac9c),
	.w5(32'h3a167986),
	.w6(32'hbb03ee65),
	.w7(32'hbba7c087),
	.w8(32'hba470961),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95b70e),
	.w1(32'h3ba05f1e),
	.w2(32'h3bcf1dfe),
	.w3(32'h3b8e1b30),
	.w4(32'h3baa1cf0),
	.w5(32'h3b73a4de),
	.w6(32'hb9426168),
	.w7(32'h3b03e5f1),
	.w8(32'h3b60afc0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67fa21),
	.w1(32'h3bac3e84),
	.w2(32'hb90cab89),
	.w3(32'h3bcf4bc4),
	.w4(32'h3ba6083a),
	.w5(32'hbc1aa26c),
	.w6(32'hbc0cf43d),
	.w7(32'hbcc47360),
	.w8(32'h3bb89dd0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38a7fa),
	.w1(32'hbb104e32),
	.w2(32'h3a46b18d),
	.w3(32'h3bcfe4ff),
	.w4(32'h3cbc6c8a),
	.w5(32'h3ca8bae2),
	.w6(32'h3ce156f9),
	.w7(32'h3cb1b472),
	.w8(32'hba31fe03),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67298e),
	.w1(32'h3c05161e),
	.w2(32'hbc251718),
	.w3(32'h3cb7802d),
	.w4(32'hba846d5b),
	.w5(32'h3b2bcf41),
	.w6(32'h3bed3b57),
	.w7(32'h3c2f4a8f),
	.w8(32'h3a521864),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0e95a),
	.w1(32'h3aa6b9e0),
	.w2(32'hbb86fffd),
	.w3(32'h3baa92b4),
	.w4(32'hbab6fa47),
	.w5(32'h3baa9593),
	.w6(32'hbb9eca70),
	.w7(32'h3bdd58e7),
	.w8(32'h3ac75fee),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986b3b1),
	.w1(32'h3ba17ff0),
	.w2(32'h3b74b9c2),
	.w3(32'h3c6090c1),
	.w4(32'h3c16e6bf),
	.w5(32'hbbf918e1),
	.w6(32'hb9bf1b9b),
	.w7(32'hbc1730f0),
	.w8(32'hbbeecf2f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61672c),
	.w1(32'hbc87e9d2),
	.w2(32'hbb0ab7ab),
	.w3(32'hbc9e97c0),
	.w4(32'hbcb66605),
	.w5(32'hbb4e4746),
	.w6(32'h3c2fb762),
	.w7(32'h3bfd8ecb),
	.w8(32'h3ab6c0f6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae97d6d),
	.w1(32'hbb408d60),
	.w2(32'hbb3b9159),
	.w3(32'hbb432005),
	.w4(32'hbab61592),
	.w5(32'h3bb79d28),
	.w6(32'h39ceadea),
	.w7(32'h3b783daf),
	.w8(32'h392efc31),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6e144),
	.w1(32'h38a4b5c4),
	.w2(32'hbb5b2813),
	.w3(32'h3bc53abc),
	.w4(32'hbbfa75c3),
	.w5(32'hbb9d0a06),
	.w6(32'h3bbbf8c5),
	.w7(32'h3b32dee6),
	.w8(32'hbbcb9ffd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5260),
	.w1(32'h3a74cd99),
	.w2(32'hbbacb3a2),
	.w3(32'hbc555dff),
	.w4(32'h3b64d2f2),
	.w5(32'hbb7b840c),
	.w6(32'hbb53856b),
	.w7(32'h3a09f526),
	.w8(32'hbc24429d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb00b94),
	.w1(32'hbb8f11d8),
	.w2(32'hbb25b7d9),
	.w3(32'hbb8ea7e4),
	.w4(32'h3c625d34),
	.w5(32'h3a857f23),
	.w6(32'h3c812ea3),
	.w7(32'h3bfafb2f),
	.w8(32'hb9c0826a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10b8b9),
	.w1(32'h3bef0db3),
	.w2(32'hbb118260),
	.w3(32'h39b12204),
	.w4(32'h3be96c6e),
	.w5(32'hbb36c0e5),
	.w6(32'hbbd2a62b),
	.w7(32'hbbc1436d),
	.w8(32'hbc17235f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f8a7a),
	.w1(32'h3b434281),
	.w2(32'hb94bb138),
	.w3(32'hbc06c185),
	.w4(32'h3bbfc884),
	.w5(32'hbbc6ba23),
	.w6(32'h3bacbe00),
	.w7(32'h3bad9060),
	.w8(32'hba9265cb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4ec61),
	.w1(32'hbb3f9c9e),
	.w2(32'h38fe538b),
	.w3(32'hbbfcf846),
	.w4(32'hbbad0c4e),
	.w5(32'h39d07768),
	.w6(32'hba283236),
	.w7(32'h3a56f720),
	.w8(32'hbbc4b4eb),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8cdd3),
	.w1(32'h3c5f712a),
	.w2(32'hbc032f43),
	.w3(32'h3a8bc4b1),
	.w4(32'hbaf07d86),
	.w5(32'hbc6dbe99),
	.w6(32'hbb79c304),
	.w7(32'h3c81136a),
	.w8(32'h3beaccdc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c73ab),
	.w1(32'hbbc980ce),
	.w2(32'h3b1bb4c7),
	.w3(32'hb9942dc2),
	.w4(32'hbb3c5bf8),
	.w5(32'h3b2786bd),
	.w6(32'h3c5bfc45),
	.w7(32'hbbf473b7),
	.w8(32'h3ac4e9dc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37dd95),
	.w1(32'hba943d4c),
	.w2(32'h3b53e648),
	.w3(32'hbbb13c38),
	.w4(32'hbc04a491),
	.w5(32'hbc3b88e7),
	.w6(32'hbba10d08),
	.w7(32'hba9042ca),
	.w8(32'hbc3b7d01),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbb6a0),
	.w1(32'hbbc0e7d2),
	.w2(32'h3b660e17),
	.w3(32'hbbda93f8),
	.w4(32'hbc4279d6),
	.w5(32'hbc89d400),
	.w6(32'h3c112370),
	.w7(32'h3b0acef4),
	.w8(32'h3c35dcbf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf39b3),
	.w1(32'hbc0c64a9),
	.w2(32'hbb09ae74),
	.w3(32'hbcaf4ae1),
	.w4(32'h3c761a76),
	.w5(32'hbbd8f97e),
	.w6(32'h3d0f07c2),
	.w7(32'h3c6e0845),
	.w8(32'h3ce29569),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c296e52),
	.w1(32'hbbed0b53),
	.w2(32'hba570cd7),
	.w3(32'h3c7ff297),
	.w4(32'h3d105d08),
	.w5(32'hbc2b0feb),
	.w6(32'h3d308343),
	.w7(32'h3c26f3e9),
	.w8(32'hbc41124d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e008d4),
	.w1(32'hbb6ff36b),
	.w2(32'hbb0ffb22),
	.w3(32'hbc2a4e9e),
	.w4(32'hbc796b64),
	.w5(32'hbb0cd258),
	.w6(32'hbc57ad21),
	.w7(32'hba9e8fa8),
	.w8(32'hbb0cc8c0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26994d),
	.w1(32'h3ab006b0),
	.w2(32'hbb9cf021),
	.w3(32'hbbba28a5),
	.w4(32'hbabc5ea6),
	.w5(32'hbbbbe3d1),
	.w6(32'hba4ea96b),
	.w7(32'h39fa129a),
	.w8(32'hbc25c112),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97a16b),
	.w1(32'hbc11f654),
	.w2(32'hbbcad971),
	.w3(32'hbc29403e),
	.w4(32'hbc3dd232),
	.w5(32'hbb4f2f2d),
	.w6(32'hbb4baeb6),
	.w7(32'h3b531a56),
	.w8(32'hbb9002b1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89e8eb),
	.w1(32'hba352d7a),
	.w2(32'hbae869bf),
	.w3(32'h3c013244),
	.w4(32'h3ad2c52a),
	.w5(32'h3a8e4d01),
	.w6(32'h3be88b4b),
	.w7(32'h3a0cc490),
	.w8(32'hba17d926),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe712c1),
	.w1(32'hbb972f4e),
	.w2(32'hbb3fa82e),
	.w3(32'hbc5f04ef),
	.w4(32'h3ae76813),
	.w5(32'hbba1c22b),
	.w6(32'h3a468d05),
	.w7(32'hbbe4c7b4),
	.w8(32'hbc48c9fb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41439d),
	.w1(32'h3be25d3a),
	.w2(32'hbbe4a100),
	.w3(32'h39e187a2),
	.w4(32'hbbc8d2fe),
	.w5(32'hbaa2ad16),
	.w6(32'hba5d2ecc),
	.w7(32'h3bba01d5),
	.w8(32'hbb4a6feb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedec4e),
	.w1(32'h3bdd7ef3),
	.w2(32'hbbfc1420),
	.w3(32'h3b9315ba),
	.w4(32'h395faea4),
	.w5(32'hbbfd9151),
	.w6(32'hb976c106),
	.w7(32'h3bcd0e86),
	.w8(32'h3b1f2db3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc886036),
	.w1(32'h3b9b3046),
	.w2(32'h3aaf0f43),
	.w3(32'h3c82831b),
	.w4(32'h3c5cf24d),
	.w5(32'h3b73642e),
	.w6(32'hbc21f9b1),
	.w7(32'hbcd0c36c),
	.w8(32'h3be51308),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75f4c0),
	.w1(32'h3a4d4369),
	.w2(32'hba626c1d),
	.w3(32'hbc0861eb),
	.w4(32'hba037690),
	.w5(32'hbb867f93),
	.w6(32'hbc736c79),
	.w7(32'hbbbebb8d),
	.w8(32'hbb11c115),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb0de7),
	.w1(32'hba90833f),
	.w2(32'hbb08a3fc),
	.w3(32'h3a2a1e0d),
	.w4(32'h3a990872),
	.w5(32'hbc838111),
	.w6(32'hbad289d3),
	.w7(32'hbb3948f8),
	.w8(32'hbc4552e1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca44803),
	.w1(32'hbc74ea19),
	.w2(32'hb9b33629),
	.w3(32'hbc8935a3),
	.w4(32'h3b21d938),
	.w5(32'hba9fce1c),
	.w6(32'hbc1cd72d),
	.w7(32'hbc7c6c5a),
	.w8(32'hbcb98f1b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938c80f),
	.w1(32'hbc2137d8),
	.w2(32'hbc5920b4),
	.w3(32'hbca1b704),
	.w4(32'hbcb70091),
	.w5(32'hbbc58291),
	.w6(32'h3bb5f83f),
	.w7(32'h3cb0857e),
	.w8(32'hbc78b941),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad3257),
	.w1(32'h3c54872f),
	.w2(32'h3b968fde),
	.w3(32'hbbc140c5),
	.w4(32'hbadb15b9),
	.w5(32'h3c00da2f),
	.w6(32'h3aaf1503),
	.w7(32'h3c89606b),
	.w8(32'h3c65a713),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89ed4e),
	.w1(32'h3c380c6c),
	.w2(32'hbbcf220b),
	.w3(32'h3bebf3d5),
	.w4(32'h3c3f8430),
	.w5(32'hbb438b3a),
	.w6(32'h3c46567e),
	.w7(32'h3c3853c6),
	.w8(32'hbbd289c7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa87acd),
	.w1(32'h3b6ebdbf),
	.w2(32'h3b0797b7),
	.w3(32'h3bacb645),
	.w4(32'h3b81fb59),
	.w5(32'hbb05c9cf),
	.w6(32'hb9c2edac),
	.w7(32'hbb902982),
	.w8(32'h3b230bc7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1738),
	.w1(32'hbb6f0899),
	.w2(32'h3ac40a4b),
	.w3(32'h3ae80852),
	.w4(32'h3bc05694),
	.w5(32'hba98c77a),
	.w6(32'h3be2e2cd),
	.w7(32'h3b138fca),
	.w8(32'hbbae6f29),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9555f),
	.w1(32'hbb69061a),
	.w2(32'hbc273c33),
	.w3(32'hbc3f9f45),
	.w4(32'h3bbacba6),
	.w5(32'h3b7649e8),
	.w6(32'h3b68fe6e),
	.w7(32'hbc662030),
	.w8(32'hbc4ce533),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24e0d1),
	.w1(32'h38fdfc7a),
	.w2(32'hbc189259),
	.w3(32'hbb9b7013),
	.w4(32'hbc0d8e64),
	.w5(32'hbc6a287e),
	.w6(32'hbc797481),
	.w7(32'hbc431c2a),
	.w8(32'hbbf43e3a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d0f5f),
	.w1(32'hbc14111e),
	.w2(32'hbca80782),
	.w3(32'hbc42d87c),
	.w4(32'hbc52f87d),
	.w5(32'hbadd46b8),
	.w6(32'h3bacf348),
	.w7(32'h3bcc06b7),
	.w8(32'hbbd69814),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3704a),
	.w1(32'hb9cf4158),
	.w2(32'hbbc3023c),
	.w3(32'hbc0a66e0),
	.w4(32'hbc47f572),
	.w5(32'hbbeee844),
	.w6(32'h3b99496a),
	.w7(32'h3c1b229a),
	.w8(32'hbc20d0b0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d5bdf),
	.w1(32'hbbf3b09b),
	.w2(32'hbc25baa0),
	.w3(32'h38dff20d),
	.w4(32'h3c03f017),
	.w5(32'hbb0d4688),
	.w6(32'h3cc3fa09),
	.w7(32'h3cc746d5),
	.w8(32'hbc074c06),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3db88),
	.w1(32'h3ab2a65d),
	.w2(32'hbc034a89),
	.w3(32'h3c09d072),
	.w4(32'hbba614cf),
	.w5(32'hbc38edc1),
	.w6(32'h3c9908b2),
	.w7(32'h3cd33b55),
	.w8(32'h3c53cea9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cba2e),
	.w1(32'hba870cb7),
	.w2(32'h3c31880f),
	.w3(32'hbca4c71a),
	.w4(32'hbb33b067),
	.w5(32'hbc585a09),
	.w6(32'hbc94806b),
	.w7(32'hbc8bb7b0),
	.w8(32'h3b59c084),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63f411),
	.w1(32'hbb62d965),
	.w2(32'hbb969e68),
	.w3(32'hbc6b3f60),
	.w4(32'hbbd24516),
	.w5(32'hbac0124d),
	.w6(32'h3ccf4830),
	.w7(32'h3bbf8044),
	.w8(32'hbca0edea),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fe82),
	.w1(32'h3b26addf),
	.w2(32'hbc23d45f),
	.w3(32'h3bfe6919),
	.w4(32'hba9fdc04),
	.w5(32'h38873254),
	.w6(32'h3ba523d5),
	.w7(32'h3b3d6301),
	.w8(32'h378838b8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae12e98),
	.w1(32'hbafc4824),
	.w2(32'hb8891e91),
	.w3(32'hbc2b00e1),
	.w4(32'hbbaef1ea),
	.w5(32'hba525e77),
	.w6(32'hbb91765a),
	.w7(32'hbafd23ba),
	.w8(32'hbc188f12),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afedeb9),
	.w1(32'h3bfca323),
	.w2(32'h3bfad4d9),
	.w3(32'h3a3f74ed),
	.w4(32'hbc66eac4),
	.w5(32'hbbcee1d4),
	.w6(32'h3c2cbf03),
	.w7(32'h3d0bdc6a),
	.w8(32'h3bd9bd2a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba056daf),
	.w1(32'h3c4c5dba),
	.w2(32'h3a31c43d),
	.w3(32'h3a4f2493),
	.w4(32'h3c344251),
	.w5(32'h3c00a201),
	.w6(32'hbbbe9b13),
	.w7(32'h3b7e5de1),
	.w8(32'h3c20deec),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20559a),
	.w1(32'hbae3a0c0),
	.w2(32'hba103fde),
	.w3(32'hbb30d9e8),
	.w4(32'hba52009b),
	.w5(32'hbb06f145),
	.w6(32'hbb02de59),
	.w7(32'h3b8da9d2),
	.w8(32'hbb8b878d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb575bc4),
	.w1(32'h3b7b00a9),
	.w2(32'hbad7aad5),
	.w3(32'hbc2e371d),
	.w4(32'h3a8844a9),
	.w5(32'h3c269fd5),
	.w6(32'hbbd56c29),
	.w7(32'hbb54566b),
	.w8(32'hbc456ddc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53b62d),
	.w1(32'h3b25911f),
	.w2(32'hba7e6ce5),
	.w3(32'h3bb5eb39),
	.w4(32'hb9a807e1),
	.w5(32'hbbf0e3b9),
	.w6(32'hbc0dc242),
	.w7(32'h3c66b66b),
	.w8(32'hbb5029dd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08685c),
	.w1(32'hbb09f99a),
	.w2(32'hbba4303e),
	.w3(32'h3b17d339),
	.w4(32'h3a72265e),
	.w5(32'h3b5d7f91),
	.w6(32'h3c359786),
	.w7(32'h3b959465),
	.w8(32'hbbaa7704),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb9635),
	.w1(32'hbb8fe703),
	.w2(32'h3b5c0761),
	.w3(32'h3bbb3fcf),
	.w4(32'hbc653736),
	.w5(32'hbb6c572b),
	.w6(32'hbc1ea4ac),
	.w7(32'hb9baee85),
	.w8(32'hbca221cd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb02946),
	.w1(32'hbc0fa3fa),
	.w2(32'hbc1595dc),
	.w3(32'hbbf06939),
	.w4(32'hbb658e8f),
	.w5(32'h3c6ef574),
	.w6(32'h3afe71fb),
	.w7(32'h3c913a09),
	.w8(32'hbc1cbdcd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4d01a),
	.w1(32'h3c388c11),
	.w2(32'h3b777e2b),
	.w3(32'h3c9e6d2e),
	.w4(32'h3c614899),
	.w5(32'h3baa0a27),
	.w6(32'h3ca2118f),
	.w7(32'h3cfddf08),
	.w8(32'h3af42a74),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b16594),
	.w1(32'h3bb4ae46),
	.w2(32'hbb27eb28),
	.w3(32'h3b389995),
	.w4(32'h3b0a1f83),
	.w5(32'hbc55ecaf),
	.w6(32'hbbcbbc95),
	.w7(32'hbb8426de),
	.w8(32'hbbdca19e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3bbb0),
	.w1(32'hbc1410bf),
	.w2(32'hbb538a9d),
	.w3(32'hbc35c22b),
	.w4(32'h3bb54890),
	.w5(32'hba91b8f1),
	.w6(32'h3bd9d8c8),
	.w7(32'h3c0d7b07),
	.w8(32'hbb547de5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca8b62),
	.w1(32'h3c5059a2),
	.w2(32'h3b857f3b),
	.w3(32'h3b4220c1),
	.w4(32'hbaf31734),
	.w5(32'hbbc398ed),
	.w6(32'hba857d68),
	.w7(32'hba79c495),
	.w8(32'hbb9d6b01),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6afae0),
	.w1(32'hbb21cdd8),
	.w2(32'h38a57078),
	.w3(32'hbbee6ba4),
	.w4(32'hba90135c),
	.w5(32'h3b5285a3),
	.w6(32'h3914db52),
	.w7(32'hba64704e),
	.w8(32'hbbd0ae61),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a59c7),
	.w1(32'h3c155d66),
	.w2(32'h3b53bb1e),
	.w3(32'hbae09359),
	.w4(32'hbbba438d),
	.w5(32'hbc61d576),
	.w6(32'hbc219881),
	.w7(32'hbc089c39),
	.w8(32'h3b157a46),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb11705),
	.w1(32'hbc3385b6),
	.w2(32'hbb62153c),
	.w3(32'hbb83938c),
	.w4(32'hbbc7433b),
	.w5(32'hbbeea884),
	.w6(32'h3bf99cef),
	.w7(32'h3bbd58bb),
	.w8(32'h3a86d866),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b716e5c),
	.w1(32'hba51747c),
	.w2(32'hbb2ea982),
	.w3(32'hbc2aa800),
	.w4(32'hbc3d41ee),
	.w5(32'h3aabe1b6),
	.w6(32'h3b211081),
	.w7(32'hbbb20f07),
	.w8(32'hbbbde020),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98ea30),
	.w1(32'h3a8446c4),
	.w2(32'hbbadd1d2),
	.w3(32'h3c366a56),
	.w4(32'h3b0a7199),
	.w5(32'hbb611a55),
	.w6(32'h3a3831d7),
	.w7(32'h3b1beebc),
	.w8(32'hbb8b955b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd512b),
	.w1(32'h3badfaef),
	.w2(32'hbaa7608e),
	.w3(32'h3bae95bc),
	.w4(32'h3c1e0118),
	.w5(32'hbaa626cc),
	.w6(32'h3bbb2591),
	.w7(32'h3bd6fe52),
	.w8(32'hb945d252),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a2f5),
	.w1(32'hb9a07511),
	.w2(32'hbbd99d8b),
	.w3(32'h395fb3d6),
	.w4(32'h3a581e3c),
	.w5(32'hbc3709c5),
	.w6(32'hbb79bc37),
	.w7(32'hbbe43829),
	.w8(32'hbc5025be),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d7545),
	.w1(32'h3b50eae1),
	.w2(32'h3af17f0f),
	.w3(32'h3c1eead2),
	.w4(32'hbb8313d3),
	.w5(32'h3bc77489),
	.w6(32'hbc2d8543),
	.w7(32'hbc5c3fde),
	.w8(32'hba734100),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3627d),
	.w1(32'h3a5f82eb),
	.w2(32'hbb08ce33),
	.w3(32'hbb53b2cd),
	.w4(32'hbc067f39),
	.w5(32'hbae27b78),
	.w6(32'hbc2b5d96),
	.w7(32'hba9d76e4),
	.w8(32'hbc252a85),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae22b0),
	.w1(32'hbb1aa6e1),
	.w2(32'h3bb0578d),
	.w3(32'hbb25d5df),
	.w4(32'hbb90f264),
	.w5(32'h3b9bff20),
	.w6(32'h3aaf730b),
	.w7(32'h3b0caafa),
	.w8(32'hbbdf15dc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be989c0),
	.w1(32'h3c6f9a6e),
	.w2(32'h3c1d2704),
	.w3(32'h3bb13876),
	.w4(32'h3b405aee),
	.w5(32'h3b978006),
	.w6(32'hbbac9ee8),
	.w7(32'h3c228b8f),
	.w8(32'hbb3157ff),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f13d),
	.w1(32'h3c08862a),
	.w2(32'h3aced411),
	.w3(32'hbc37e834),
	.w4(32'h3c229e56),
	.w5(32'hbbf5e8f4),
	.w6(32'h3bb3d701),
	.w7(32'h3b7df252),
	.w8(32'h3b7bcc89),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a0321),
	.w1(32'hbc76a158),
	.w2(32'hbbcec8f6),
	.w3(32'hbb86165a),
	.w4(32'h3c082b35),
	.w5(32'hbb1c1289),
	.w6(32'h3ca3de44),
	.w7(32'h3c60d0f3),
	.w8(32'hbc159c8f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cc51e),
	.w1(32'hbb1afe26),
	.w2(32'hbc0a6866),
	.w3(32'hbc018556),
	.w4(32'hbc0998ff),
	.w5(32'h3c2deb12),
	.w6(32'hbab48198),
	.w7(32'hbabef9b2),
	.w8(32'hbc39378c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c3711),
	.w1(32'h3b75c54d),
	.w2(32'h3b4d0c4a),
	.w3(32'h3cb8b75d),
	.w4(32'hbca6790b),
	.w5(32'h3c52b2a8),
	.w6(32'hbc7b7822),
	.w7(32'h3b173b59),
	.w8(32'h3c4f19c8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f8853),
	.w1(32'h3c857876),
	.w2(32'hbc94c292),
	.w3(32'h3c2fa3fd),
	.w4(32'h3aa68347),
	.w5(32'hbc91795c),
	.w6(32'hb81fae0a),
	.w7(32'hbb9c9f2c),
	.w8(32'hbca73204),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6eb821),
	.w1(32'hbc80050f),
	.w2(32'h3b30b608),
	.w3(32'hbb738b4f),
	.w4(32'hbc87fce9),
	.w5(32'hbbcab0de),
	.w6(32'hbd28b8a7),
	.w7(32'hbcb0d752),
	.w8(32'hbc87b48b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca774a4),
	.w1(32'hbc31b38b),
	.w2(32'hbb932f17),
	.w3(32'hbcdcb48e),
	.w4(32'hbcae9a38),
	.w5(32'hbbeaa1ba),
	.w6(32'hbc401c8e),
	.w7(32'hbc935789),
	.w8(32'hbacafdbc),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1ec43),
	.w1(32'hbb5a6cec),
	.w2(32'hbc03ead0),
	.w3(32'h3bcc7754),
	.w4(32'h3b03175d),
	.w5(32'h3ae0ea5f),
	.w6(32'h3cf278be),
	.w7(32'h3c98889e),
	.w8(32'h3a92b784),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e2871),
	.w1(32'h3beb2b70),
	.w2(32'hbb1a4c64),
	.w3(32'h3bd316b7),
	.w4(32'hba6f4de0),
	.w5(32'hbc481a2b),
	.w6(32'hbb953e1d),
	.w7(32'hbbb1b4f5),
	.w8(32'hbc45c344),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac25622),
	.w1(32'hbbbeffa5),
	.w2(32'h386037aa),
	.w3(32'hbba658ed),
	.w4(32'h3ba4e776),
	.w5(32'h3b55141c),
	.w6(32'h3bd6e9b2),
	.w7(32'h3ccdf793),
	.w8(32'h3bbb8096),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f20dd),
	.w1(32'h3c6b2656),
	.w2(32'hbb63bee7),
	.w3(32'h3c414970),
	.w4(32'h3c9529e9),
	.w5(32'hbb0f8101),
	.w6(32'h3d3996ac),
	.w7(32'h3ccb8e17),
	.w8(32'h3bd3c679),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba904ac6),
	.w1(32'h399db6f6),
	.w2(32'hb903cd41),
	.w3(32'h3ac5e90b),
	.w4(32'h3b786303),
	.w5(32'hb99465e6),
	.w6(32'h3abf3160),
	.w7(32'hbb32d505),
	.w8(32'h3ba85794),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0428a4),
	.w1(32'hba58da89),
	.w2(32'hbb87b731),
	.w3(32'hbbd7d446),
	.w4(32'hbc0ef761),
	.w5(32'hbc150adf),
	.w6(32'h3b7a3c13),
	.w7(32'h3a1f61ea),
	.w8(32'hbbb521cc),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1271),
	.w1(32'hbba28553),
	.w2(32'hbb03634c),
	.w3(32'hbbf9a29f),
	.w4(32'hbb87c993),
	.w5(32'hbc378437),
	.w6(32'hba395e75),
	.w7(32'hbb2e7d3c),
	.w8(32'hbbb0cf4d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31a8af),
	.w1(32'hbc0c6433),
	.w2(32'hbaba255d),
	.w3(32'h39b03a11),
	.w4(32'h3ba1fb13),
	.w5(32'hbcef3b14),
	.w6(32'hbbbdde22),
	.w7(32'hbba88203),
	.w8(32'h3c826600),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74a090),
	.w1(32'hbc71d944),
	.w2(32'hbb3e73c2),
	.w3(32'h3c013b84),
	.w4(32'h3d282f67),
	.w5(32'hbaca81e9),
	.w6(32'h3b7b451c),
	.w7(32'hbcbc49ce),
	.w8(32'hbc48a5ec),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4556b6),
	.w1(32'h3c0c8c9d),
	.w2(32'hbac21a54),
	.w3(32'h3afee7cc),
	.w4(32'h3b58a31f),
	.w5(32'hbb192c59),
	.w6(32'hbbbd3a53),
	.w7(32'hbbfbfabd),
	.w8(32'h3a1dd043),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77b71c),
	.w1(32'hbb651b54),
	.w2(32'hbaf96ba2),
	.w3(32'h36177ab1),
	.w4(32'h3abba1c5),
	.w5(32'hbc0fb579),
	.w6(32'h3b076d13),
	.w7(32'hba8b35a9),
	.w8(32'hbc03b778),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a4db45),
	.w1(32'hbb974135),
	.w2(32'hbbb71ccd),
	.w3(32'hbc5e5fc1),
	.w4(32'hbbb69fab),
	.w5(32'h3a7c9aba),
	.w6(32'h3a552521),
	.w7(32'h3cb54216),
	.w8(32'hbb73239e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf8d2),
	.w1(32'hbb4e4ba4),
	.w2(32'h3b4a9dc4),
	.w3(32'hbaa6d717),
	.w4(32'hbb77b5eb),
	.w5(32'h3c5ea2d1),
	.w6(32'hbc0f9c28),
	.w7(32'h3a9fc816),
	.w8(32'h3a448d66),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d193e05),
	.w1(32'h3d04276e),
	.w2(32'hbb30904b),
	.w3(32'h3ccce8b6),
	.w4(32'h3c31c509),
	.w5(32'hbb4d45c2),
	.w6(32'h3c92f9a1),
	.w7(32'h3cd1973d),
	.w8(32'hbbb8c427),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa42ad4),
	.w1(32'hbb3b1428),
	.w2(32'hbb0dc392),
	.w3(32'hbc2746b8),
	.w4(32'hbac5c7d8),
	.w5(32'h3b224933),
	.w6(32'hba040835),
	.w7(32'h3b40a22e),
	.w8(32'hba42e02d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ddd6c),
	.w1(32'hbc0f348e),
	.w2(32'hbb81d9f5),
	.w3(32'h3a8b78c5),
	.w4(32'hbc46a69f),
	.w5(32'hbb5e8b0a),
	.w6(32'hbbc24c23),
	.w7(32'h391a0897),
	.w8(32'hbb64e91d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8752f),
	.w1(32'hb9844327),
	.w2(32'hbba52015),
	.w3(32'hbb853cf4),
	.w4(32'hbb106a0f),
	.w5(32'hbc00e534),
	.w6(32'hbbdec6d5),
	.w7(32'h3ba44be0),
	.w8(32'hbb7e4874),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d93a1),
	.w1(32'h3af3e200),
	.w2(32'hbc2739e2),
	.w3(32'h3bf02139),
	.w4(32'h3c760230),
	.w5(32'hbb6f1955),
	.w6(32'h3ceba089),
	.w7(32'h3c864e5f),
	.w8(32'h3b5b37ea),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd343ff),
	.w1(32'hbb1cebd3),
	.w2(32'hbc1de1b1),
	.w3(32'h3aa30cfc),
	.w4(32'h3bd791aa),
	.w5(32'hbcb977a0),
	.w6(32'hb8853c08),
	.w7(32'hbc0623fe),
	.w8(32'hbcbc0f7e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76c6d5),
	.w1(32'hbc2b2e50),
	.w2(32'h3bee31f1),
	.w3(32'hbd21710e),
	.w4(32'hbcfd72cb),
	.w5(32'hbc101116),
	.w6(32'hbc8abbde),
	.w7(32'hbbcde7d6),
	.w8(32'h3c1ac50a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c820dd5),
	.w1(32'hbbd07e62),
	.w2(32'hba4ca878),
	.w3(32'h3b919617),
	.w4(32'h3cc3683b),
	.w5(32'h3b0ba106),
	.w6(32'h3d1f36c5),
	.w7(32'h3cb51aa2),
	.w8(32'h3b0a6358),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21a10c),
	.w1(32'hbb515154),
	.w2(32'h3b91d04f),
	.w3(32'h3bcc46e4),
	.w4(32'h3b43b35b),
	.w5(32'h3bceefaa),
	.w6(32'h3b85dd46),
	.w7(32'h39e6bb70),
	.w8(32'h3b9faec9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cedd0),
	.w1(32'hbc1ddd0b),
	.w2(32'hbb644382),
	.w3(32'hbba9c22d),
	.w4(32'hbc1a6990),
	.w5(32'hbae967b9),
	.w6(32'hbb50dc50),
	.w7(32'hbc600428),
	.w8(32'hbba88905),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af621ae),
	.w1(32'h3be20d87),
	.w2(32'h3c9f08ee),
	.w3(32'hbaaf3018),
	.w4(32'h3ba2008f),
	.w5(32'hbbf6396f),
	.w6(32'hbc155324),
	.w7(32'hbbcd40b2),
	.w8(32'hbd223637),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d97a9d2),
	.w1(32'h3d48e3d8),
	.w2(32'h3a8f3b74),
	.w3(32'h3c7f794e),
	.w4(32'h3cda8588),
	.w5(32'h3ab1f124),
	.w6(32'hbd876c9f),
	.w7(32'hbd0be14d),
	.w8(32'hb931487a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37d5ab),
	.w1(32'h39226f61),
	.w2(32'h3c4640fe),
	.w3(32'h3ba7974c),
	.w4(32'h3b40344e),
	.w5(32'h3abc494c),
	.w6(32'hbba1a661),
	.w7(32'hbb3eac3f),
	.w8(32'hbbee7751),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc457ae),
	.w1(32'h3c0826ab),
	.w2(32'h3c369dee),
	.w3(32'h3c345a1b),
	.w4(32'h3c43b289),
	.w5(32'hbccdbedc),
	.w6(32'hbc05a437),
	.w7(32'hbbc77139),
	.w8(32'hbd8e06ae),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db028b1),
	.w1(32'h3d7ff8b3),
	.w2(32'h3ade7c81),
	.w3(32'h3c13c3cb),
	.w4(32'h3cfb84b6),
	.w5(32'h3b8fdd45),
	.w6(32'hbdd5ed2d),
	.w7(32'hbd58c6b7),
	.w8(32'hbb1632be),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbdd23),
	.w1(32'h3bb31349),
	.w2(32'hbc2daa7c),
	.w3(32'h3b1a4c90),
	.w4(32'h3b989403),
	.w5(32'h3b105806),
	.w6(32'h3abcb067),
	.w7(32'hbbae71d3),
	.w8(32'h3c6cbcb8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd161321),
	.w1(32'hbc9d3b05),
	.w2(32'h3b8c441c),
	.w3(32'hbc39d21f),
	.w4(32'hbc44b280),
	.w5(32'h3bc6c66a),
	.w6(32'h3d0a2193),
	.w7(32'h3cb081ce),
	.w8(32'hbc22cc78),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c131ab7),
	.w1(32'h3bfd3c2b),
	.w2(32'h3cacfdd9),
	.w3(32'h3c1c42db),
	.w4(32'hbb4e212c),
	.w5(32'hbc8878b2),
	.w6(32'h3a70ee0e),
	.w7(32'hbbc73824),
	.w8(32'hbd5171de),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3daf3b10),
	.w1(32'h3d7b70cd),
	.w2(32'h3aa762af),
	.w3(32'h3c20ac0c),
	.w4(32'h3cf98021),
	.w5(32'h3b668c7a),
	.w6(32'hbda55691),
	.w7(32'hbd23d2ee),
	.w8(32'hbb5900f1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15bf99),
	.w1(32'hbb0c85cf),
	.w2(32'h3ae1cfe0),
	.w3(32'hbb8d819b),
	.w4(32'hbb59bb03),
	.w5(32'hbba06e50),
	.w6(32'hbbfb237f),
	.w7(32'hbb913325),
	.w8(32'hbc32d0d0),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef198d),
	.w1(32'h399da2d5),
	.w2(32'h3a99526c),
	.w3(32'hbb8eb7b9),
	.w4(32'hbc274b76),
	.w5(32'h3ba26ca1),
	.w6(32'hbc512975),
	.w7(32'hbc7bd29e),
	.w8(32'h3bae812d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaf624),
	.w1(32'h3c08e542),
	.w2(32'hbb96ab43),
	.w3(32'h3b21b899),
	.w4(32'h3c409c7b),
	.w5(32'h3b2464af),
	.w6(32'h3c357525),
	.w7(32'h3c4626ac),
	.w8(32'hbb815197),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28248b),
	.w1(32'h3c1610b7),
	.w2(32'hbb0249c8),
	.w3(32'h3bfce43e),
	.w4(32'h3beb8848),
	.w5(32'h3ae2f78d),
	.w6(32'hbc138e69),
	.w7(32'hbbb691bd),
	.w8(32'hbae481a4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbc96e),
	.w1(32'hba0ef334),
	.w2(32'hbc8141a2),
	.w3(32'hb911281b),
	.w4(32'hbb8aeb8e),
	.w5(32'h3c5ed176),
	.w6(32'hbc358cde),
	.w7(32'hbc20003b),
	.w8(32'h3d34042a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8f1f52),
	.w1(32'hbd4fc5e8),
	.w2(32'hbb1f3e70),
	.w3(32'hbbed1c07),
	.w4(32'hbd03681b),
	.w5(32'hbb8925c0),
	.w6(32'h3d908d66),
	.w7(32'h3cf52316),
	.w8(32'hbc389096),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43ddb),
	.w1(32'hbbce590d),
	.w2(32'h3b21e493),
	.w3(32'h3abb61c8),
	.w4(32'hbb8a4004),
	.w5(32'hbadd7500),
	.w6(32'h3a2618a1),
	.w7(32'hbbb2a715),
	.w8(32'hbbdc48fe),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad64128),
	.w1(32'h3c03e515),
	.w2(32'hbbd35f3e),
	.w3(32'h3b677bd0),
	.w4(32'hba090753),
	.w5(32'hbb33f0e7),
	.w6(32'hbb17fd04),
	.w7(32'h3ad42129),
	.w8(32'h39f81cee),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c064562),
	.w1(32'h3c0e742d),
	.w2(32'hbbebd369),
	.w3(32'h3c09bb3a),
	.w4(32'h3bc73d34),
	.w5(32'hbc399d25),
	.w6(32'h3c3aa8fd),
	.w7(32'hb723155a),
	.w8(32'hbc5e2af6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952e14d),
	.w1(32'hbb577c2c),
	.w2(32'hbc903a5e),
	.w3(32'hbabba1e7),
	.w4(32'hbb096992),
	.w5(32'h3c29ee0f),
	.w6(32'hbc3d5f0c),
	.w7(32'hbc454dc4),
	.w8(32'h3d417c59),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9c5808),
	.w1(32'hbd5802b8),
	.w2(32'hbc5aac5f),
	.w3(32'hbc587b8c),
	.w4(32'hbcdbbb8f),
	.w5(32'hbc8ae3b5),
	.w6(32'h3da96ac3),
	.w7(32'h3d3870e9),
	.w8(32'hbac60cfa),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135265),
	.w1(32'hb96c33fe),
	.w2(32'h3bc530f5),
	.w3(32'hbc09c19a),
	.w4(32'hbb8954dc),
	.w5(32'h3b427f49),
	.w6(32'h3a654ad9),
	.w7(32'h3b384fe7),
	.w8(32'hbba76812),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ca1de),
	.w1(32'h3ba314af),
	.w2(32'hba03576a),
	.w3(32'h3b304725),
	.w4(32'h3b9188b5),
	.w5(32'hbb5e4872),
	.w6(32'h3b8ea469),
	.w7(32'h3959150c),
	.w8(32'hbc5fc517),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62e857),
	.w1(32'h3b40187f),
	.w2(32'hbbb293a0),
	.w3(32'h3bc53e55),
	.w4(32'h3b8b8586),
	.w5(32'hbbb77c7b),
	.w6(32'h39ad2e7c),
	.w7(32'h3afb4b86),
	.w8(32'hbbbc9c39),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae84509),
	.w1(32'hba9f2213),
	.w2(32'h3be80015),
	.w3(32'hbb22c27d),
	.w4(32'h3b929fd1),
	.w5(32'hbb0e263e),
	.w6(32'hbc0c48d3),
	.w7(32'hbc12beba),
	.w8(32'hbb7b1463),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c216c),
	.w1(32'h3c3751ec),
	.w2(32'hbc13e5d4),
	.w3(32'hbb46154d),
	.w4(32'hbb0c24c9),
	.w5(32'hbb4f0702),
	.w6(32'h3a15d689),
	.w7(32'h3a98f7aa),
	.w8(32'hba8635c8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd94e5c),
	.w1(32'hbaf4f579),
	.w2(32'h3bf0c946),
	.w3(32'hbc482244),
	.w4(32'hbb9656b0),
	.w5(32'hbbff8abf),
	.w6(32'hbc22e315),
	.w7(32'hba220abd),
	.w8(32'hbc2ab329),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21db1e),
	.w1(32'h3bf4b139),
	.w2(32'hbaf4437b),
	.w3(32'hbb9b152c),
	.w4(32'hbb499021),
	.w5(32'hbaba9c7d),
	.w6(32'hbbad2f18),
	.w7(32'hbba3d561),
	.w8(32'h3bddf913),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940a03e),
	.w1(32'h3c376190),
	.w2(32'h388b53f3),
	.w3(32'h39b486fd),
	.w4(32'h3c2e2dce),
	.w5(32'h3bdc27f5),
	.w6(32'h3bb0fdec),
	.w7(32'h3c7112a0),
	.w8(32'h3b23d920),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cac2c),
	.w1(32'h3c86a8f7),
	.w2(32'hba68156a),
	.w3(32'h3bb45ca5),
	.w4(32'h3b40d597),
	.w5(32'h3aa18c2e),
	.w6(32'h3bb6cc0c),
	.w7(32'h3bd387c7),
	.w8(32'h3ccdd308),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d845c),
	.w1(32'hbb56ea97),
	.w2(32'h3bf8326f),
	.w3(32'h3a0c888d),
	.w4(32'hbba6d9be),
	.w5(32'h3bb1e54d),
	.w6(32'h3c2fc01f),
	.w7(32'h3baf8f5f),
	.w8(32'hbb293194),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3f909d),
	.w1(32'h3ce3c954),
	.w2(32'hba4a3610),
	.w3(32'h3d2f04ad),
	.w4(32'h3cfbfc04),
	.w5(32'h3baf4f11),
	.w6(32'h3d54c170),
	.w7(32'h3d046825),
	.w8(32'h3ba8dc95),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e73ca),
	.w1(32'hbbb03dd4),
	.w2(32'h3c1b22da),
	.w3(32'hbc3f053a),
	.w4(32'hbbe27f2b),
	.w5(32'hbae5d86e),
	.w6(32'hbbf0216c),
	.w7(32'hbc2563fb),
	.w8(32'hbbaea809),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c007f72),
	.w1(32'h3c455f67),
	.w2(32'hbc26b6f9),
	.w3(32'h3be751e0),
	.w4(32'h3b4d07f7),
	.w5(32'hbb97317a),
	.w6(32'hbaf1c58d),
	.w7(32'h3acfc2a0),
	.w8(32'hbab1ccba),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5018),
	.w1(32'hbb88b572),
	.w2(32'hbb19397d),
	.w3(32'hbbfb7d90),
	.w4(32'hbb9d7aeb),
	.w5(32'hbbe030c0),
	.w6(32'hbb1904ec),
	.w7(32'hbb8d5435),
	.w8(32'h3b0bee68),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac50aa8),
	.w1(32'hb9fd2da0),
	.w2(32'hbb741271),
	.w3(32'hbb3a7516),
	.w4(32'hbb9f4fd9),
	.w5(32'h39c4b9f9),
	.w6(32'h3b4b3d6f),
	.w7(32'hba0afcae),
	.w8(32'hbb5897eb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71db99),
	.w1(32'hbb61d220),
	.w2(32'h3bbe3c07),
	.w3(32'h3b50ee69),
	.w4(32'hbb3a2015),
	.w5(32'h3b34ce88),
	.w6(32'h3b3848d4),
	.w7(32'hb9cd2a1d),
	.w8(32'h3b31e26f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb2dce),
	.w1(32'h3ad97cdb),
	.w2(32'h3b2439e8),
	.w3(32'h3b4654c3),
	.w4(32'h3b37a5dd),
	.w5(32'h3c102e71),
	.w6(32'h3bd2bfe2),
	.w7(32'h3b507603),
	.w8(32'h3bdb6a6a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e2a5f),
	.w1(32'hbbecce4e),
	.w2(32'hba3290a2),
	.w3(32'h3b8dfa01),
	.w4(32'hbbbb4841),
	.w5(32'hbb41b6d4),
	.w6(32'hbc231052),
	.w7(32'hbc447847),
	.w8(32'hbc05a288),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b89b6),
	.w1(32'h3b2a2d56),
	.w2(32'h39a8c7b3),
	.w3(32'h3b8b976c),
	.w4(32'h39d3f5e3),
	.w5(32'hbb5f8c4c),
	.w6(32'hbc457a8f),
	.w7(32'hbc32748e),
	.w8(32'hbbcf8477),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb769c3f),
	.w1(32'hbb0c651e),
	.w2(32'hbb381489),
	.w3(32'hbc0f3a46),
	.w4(32'hbab9e5ce),
	.w5(32'h3b68062e),
	.w6(32'hb92df1b7),
	.w7(32'hb8a68022),
	.w8(32'h3c4bc2f1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d2360),
	.w1(32'hbbb1e3ab),
	.w2(32'h3ba0ff95),
	.w3(32'h3c02f936),
	.w4(32'h3b79ba42),
	.w5(32'hbb030c07),
	.w6(32'h3ca4d2d1),
	.w7(32'h3c73bedd),
	.w8(32'hbc1d2605),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b466a),
	.w1(32'h3a1e2f4d),
	.w2(32'h3bb45f01),
	.w3(32'h3bbd9187),
	.w4(32'h3bcef40e),
	.w5(32'hbb1deb57),
	.w6(32'h3b092edb),
	.w7(32'h3c2800df),
	.w8(32'h3b211a49),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb05edd),
	.w1(32'h3b6db87e),
	.w2(32'hb918f75e),
	.w3(32'hbbebc1b3),
	.w4(32'hbc04a988),
	.w5(32'hba792c5d),
	.w6(32'hbc195db2),
	.w7(32'hbb72e108),
	.w8(32'h39299174),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc82c8b),
	.w1(32'h3ac45a07),
	.w2(32'h3c1a550c),
	.w3(32'h3a580faa),
	.w4(32'h39f7f9e1),
	.w5(32'h3c1e570b),
	.w6(32'h3b0e9f8c),
	.w7(32'h3b9e4627),
	.w8(32'h3bafc8fd),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf94bea),
	.w1(32'hba7fb5fa),
	.w2(32'hbc34e13d),
	.w3(32'h3ba3fe4c),
	.w4(32'hbb959eb9),
	.w5(32'h3c0d999e),
	.w6(32'h3b110c8e),
	.w7(32'hbbc148d9),
	.w8(32'h3d1ac238),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd454f34),
	.w1(32'hbd04a529),
	.w2(32'h3b832811),
	.w3(32'h3acd3e38),
	.w4(32'hbc06f0fa),
	.w5(32'hbc349851),
	.w6(32'h3d8a047d),
	.w7(32'h3d2e1f03),
	.w8(32'hbbb46aa0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b32a9),
	.w1(32'h3bbc9237),
	.w2(32'hb8561ac7),
	.w3(32'hbc1eb445),
	.w4(32'hb9ac3bc5),
	.w5(32'hbb82ae45),
	.w6(32'hbca4daf5),
	.w7(32'hbc4268a2),
	.w8(32'hbc06bc41),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0415bb),
	.w1(32'hbb90b961),
	.w2(32'h3ad5ac05),
	.w3(32'hbb05264a),
	.w4(32'hbb953bfa),
	.w5(32'hbbe10ebc),
	.w6(32'hbb9975e2),
	.w7(32'hbb4c4208),
	.w8(32'hbb987116),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0bbc2),
	.w1(32'hb9d6d7ab),
	.w2(32'hbac898f2),
	.w3(32'hbb7f8ec7),
	.w4(32'hbc1bce60),
	.w5(32'hbb801a99),
	.w6(32'hbbef86dd),
	.w7(32'hbb7f59fe),
	.w8(32'h3bca2610),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb4ace),
	.w1(32'hbb558890),
	.w2(32'hbb60d4bb),
	.w3(32'hbc216534),
	.w4(32'hbae3194d),
	.w5(32'h3931467d),
	.w6(32'hbc46eb6f),
	.w7(32'hbc18a13f),
	.w8(32'hba5528dd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1abda6),
	.w1(32'hbb4d378f),
	.w2(32'hbb09e357),
	.w3(32'h3bbe5cd4),
	.w4(32'hbb2412b9),
	.w5(32'hbbd40193),
	.w6(32'h3bc3dccc),
	.w7(32'hbaf94f3c),
	.w8(32'hbbd8f142),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fd5b3),
	.w1(32'h3bfaf717),
	.w2(32'hb974fdcf),
	.w3(32'h3c5c56e3),
	.w4(32'h3c26ef0d),
	.w5(32'hba6eb33b),
	.w6(32'h3b920d4d),
	.w7(32'h3bbe2d6d),
	.w8(32'hbc945ee6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfe43c7),
	.w1(32'h3bdfc827),
	.w2(32'hbc0dc97d),
	.w3(32'h3c39b6ae),
	.w4(32'h3b36415f),
	.w5(32'hbc034bdb),
	.w6(32'hbd1e1569),
	.w7(32'hbccc1cb1),
	.w8(32'hb92b8bb1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca324dc),
	.w1(32'hbc6b0157),
	.w2(32'hbb8ab75e),
	.w3(32'hbc7048eb),
	.w4(32'hbc15a4ac),
	.w5(32'h3b3637df),
	.w6(32'hbbffdb90),
	.w7(32'hbbcfd04c),
	.w8(32'hbbbf4faf),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07457e),
	.w1(32'h3b0ade7a),
	.w2(32'h394271f3),
	.w3(32'h3b2faffc),
	.w4(32'h3a39c329),
	.w5(32'hba72a32a),
	.w6(32'hbbb471b8),
	.w7(32'hbc3a90f9),
	.w8(32'hba956548),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066618),
	.w1(32'h3c3e7d25),
	.w2(32'hbb3dfd0b),
	.w3(32'h3c2d4123),
	.w4(32'h3c84e40f),
	.w5(32'h3b9ce885),
	.w6(32'h3c951027),
	.w7(32'h3c369180),
	.w8(32'hbc3bf7ac),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3ce59),
	.w1(32'h3bf0920b),
	.w2(32'hbc1cc369),
	.w3(32'h3bc0a16b),
	.w4(32'h3c1be483),
	.w5(32'hbbb5a1ec),
	.w6(32'hbc50d368),
	.w7(32'hbb9e93bb),
	.w8(32'hbc1bd05e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07501e),
	.w1(32'h3bb1edef),
	.w2(32'h3a5e1dba),
	.w3(32'hb9064653),
	.w4(32'h3b7db961),
	.w5(32'h3ba0aeb4),
	.w6(32'h3c01fd00),
	.w7(32'h3c381639),
	.w8(32'h3bf0943f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e0d34),
	.w1(32'hbbccb94d),
	.w2(32'h3b8735f3),
	.w3(32'hba254f1b),
	.w4(32'hbb4a75a6),
	.w5(32'h3ab1e58a),
	.w6(32'h3bafd3e5),
	.w7(32'h3ade2f9a),
	.w8(32'hba544e89),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd89d4),
	.w1(32'h3be80802),
	.w2(32'h3c11a1fe),
	.w3(32'h3b4e1ea9),
	.w4(32'h3b86b735),
	.w5(32'h391587d0),
	.w6(32'hbbc6889b),
	.w7(32'h3a0480f5),
	.w8(32'hbc3accab),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c821a4d),
	.w1(32'h3c974591),
	.w2(32'h3bd70a7d),
	.w3(32'h3c251afd),
	.w4(32'h3c53fc67),
	.w5(32'hba8e2939),
	.w6(32'h3a89a2fe),
	.w7(32'h3c85f802),
	.w8(32'h3c4310a1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93de30),
	.w1(32'h3c56678b),
	.w2(32'hbbcdc354),
	.w3(32'h3c34cc49),
	.w4(32'h3c1cb1ef),
	.w5(32'hbbc6b5f0),
	.w6(32'h3cec4e16),
	.w7(32'h3ccd855d),
	.w8(32'h3bbc76da),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b80b9),
	.w1(32'hbc913be9),
	.w2(32'hbb80960a),
	.w3(32'hbc6d33df),
	.w4(32'hbc765513),
	.w5(32'hb9b8709f),
	.w6(32'h3cb30ac1),
	.w7(32'h3c4895a7),
	.w8(32'h3c15e7a4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f47076),
	.w1(32'h3c08a390),
	.w2(32'hbadbebce),
	.w3(32'hbb5654af),
	.w4(32'h3b6a3077),
	.w5(32'h3c72e931),
	.w6(32'hbb91a954),
	.w7(32'h3b864122),
	.w8(32'h3cca303b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc07d8c),
	.w1(32'hbc9fa333),
	.w2(32'hbbdf1d55),
	.w3(32'h3b731c15),
	.w4(32'hbc37a49b),
	.w5(32'hbbbce4c0),
	.w6(32'h3cdf8c01),
	.w7(32'h3bf7129c),
	.w8(32'hbb2d5036),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b0fb8),
	.w1(32'hbba7a151),
	.w2(32'h3bb18876),
	.w3(32'hbb663333),
	.w4(32'hbb89c3ab),
	.w5(32'h397b6ef8),
	.w6(32'h3b0f84df),
	.w7(32'hbbd5f0d7),
	.w8(32'h3a99f07f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3613d1),
	.w1(32'hbaa18a82),
	.w2(32'hbb4a05bc),
	.w3(32'hb8ba73f9),
	.w4(32'h3b4cfa08),
	.w5(32'hbb3039e8),
	.w6(32'h3a8412fe),
	.w7(32'h3c3843ea),
	.w8(32'h3aea0f03),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91c3b9),
	.w1(32'hbaeff601),
	.w2(32'hbc047462),
	.w3(32'hbbad2569),
	.w4(32'hb9a5a891),
	.w5(32'hbb109fa1),
	.w6(32'hbaaaf97b),
	.w7(32'hb87ee3e3),
	.w8(32'hb9993933),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab92b46),
	.w1(32'hba8447a9),
	.w2(32'h3be783d5),
	.w3(32'h3bdf7878),
	.w4(32'h3ab15443),
	.w5(32'h3b7170ca),
	.w6(32'hbb943549),
	.w7(32'hbaaf39f1),
	.w8(32'hbb9e7871),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85dbd7),
	.w1(32'h3c5ef377),
	.w2(32'hba356cb2),
	.w3(32'h3c896fc9),
	.w4(32'h3c657bd4),
	.w5(32'hbb2606d3),
	.w6(32'h3b6d71ef),
	.w7(32'h3bb14ebd),
	.w8(32'hbb66068c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62ce52),
	.w1(32'h3b766113),
	.w2(32'hbc01e50c),
	.w3(32'h39dc93ff),
	.w4(32'h3c1ff3bf),
	.w5(32'hbc789097),
	.w6(32'h3bc1699b),
	.w7(32'h3c8fd4ce),
	.w8(32'hbc94f6be),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86bc95),
	.w1(32'hba435591),
	.w2(32'hba8fe62f),
	.w3(32'hbb9d239c),
	.w4(32'hbb6d8160),
	.w5(32'hbb67ea78),
	.w6(32'hbc11fc55),
	.w7(32'hbb8df59d),
	.w8(32'hbc7074ad),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d30e3),
	.w1(32'hbb25ec3a),
	.w2(32'h3aba6505),
	.w3(32'h3a4d7d68),
	.w4(32'hbb4870c9),
	.w5(32'h3c0c9d2d),
	.w6(32'hbc3d5a0a),
	.w7(32'hbc22d8fa),
	.w8(32'h3b1eac11),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94902c),
	.w1(32'h3c79b8dd),
	.w2(32'hbc2ab2bc),
	.w3(32'h3cc9e718),
	.w4(32'h3c827ae6),
	.w5(32'h3b75226b),
	.w6(32'h3d0a3d36),
	.w7(32'h3cafbbe5),
	.w8(32'h3c1fae33),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c012354),
	.w1(32'h3bb9eb29),
	.w2(32'h39d74494),
	.w3(32'h3bb722d3),
	.w4(32'h3bbd1968),
	.w5(32'hb970abd0),
	.w6(32'h3babbb31),
	.w7(32'h3bac476d),
	.w8(32'hbc0905f1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3ae5),
	.w1(32'h3abaa34a),
	.w2(32'hbb97de45),
	.w3(32'hb9c19a27),
	.w4(32'hbb39d76f),
	.w5(32'hb8052853),
	.w6(32'hbbbf9b7d),
	.w7(32'hbba1629a),
	.w8(32'hbb28a5c3),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd4029),
	.w1(32'h36d0aa66),
	.w2(32'h3ac090d1),
	.w3(32'h3bf63368),
	.w4(32'h3b9a8b26),
	.w5(32'hbb892f19),
	.w6(32'h39d0c6a9),
	.w7(32'h3b14bb78),
	.w8(32'hbbf483f5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcbc28),
	.w1(32'hbbe2ec39),
	.w2(32'h3c3c91e0),
	.w3(32'h3b65afd4),
	.w4(32'hbb469f0d),
	.w5(32'hbaa56b9c),
	.w6(32'hbb6c01b6),
	.w7(32'hbb8bb123),
	.w8(32'h3bb17984),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87a152),
	.w1(32'h3c5e3c79),
	.w2(32'hba58d7c3),
	.w3(32'h3bf4fc6b),
	.w4(32'h3c117126),
	.w5(32'hbb40d726),
	.w6(32'hbb7f4203),
	.w7(32'h3bbab50d),
	.w8(32'hbbe6f32c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd164fd),
	.w1(32'h3c2cb115),
	.w2(32'h3c047637),
	.w3(32'hba430fd5),
	.w4(32'h3b8bc5ea),
	.w5(32'hbb46eb45),
	.w6(32'hbbc88b62),
	.w7(32'hbb2928ad),
	.w8(32'hbb8c4e1c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac34c66),
	.w1(32'h3b529e4b),
	.w2(32'hbc5994e4),
	.w3(32'hbb595357),
	.w4(32'hbbac8ccb),
	.w5(32'hbc6a2992),
	.w6(32'hbc70d364),
	.w7(32'hbbdb20de),
	.w8(32'hbb9929d6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0bbd6),
	.w1(32'hbb9fe51a),
	.w2(32'h3be217f1),
	.w3(32'hbb8e9e96),
	.w4(32'h3b219d3c),
	.w5(32'h3b51f93f),
	.w6(32'hbc5c434b),
	.w7(32'hbbcbc71f),
	.w8(32'h3c17ffdb),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08c8b8),
	.w1(32'hbad6023f),
	.w2(32'hbc61a651),
	.w3(32'h3c13702e),
	.w4(32'hb9715c5b),
	.w5(32'hbc054a0b),
	.w6(32'hbac029e7),
	.w7(32'hbbbdc20b),
	.w8(32'hbc4b92fe),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b895aa0),
	.w1(32'h3bdde9e2),
	.w2(32'hbb2eaddf),
	.w3(32'h3bac1ae3),
	.w4(32'h3be20d54),
	.w5(32'h3c17517a),
	.w6(32'h3bf4531f),
	.w7(32'h3b4671ff),
	.w8(32'hbba9ba7c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bb02d),
	.w1(32'h3c4ca2d6),
	.w2(32'h3ac5e4e3),
	.w3(32'h3c640a0b),
	.w4(32'h3c14a10b),
	.w5(32'hb992bb52),
	.w6(32'hba8bd238),
	.w7(32'hbb1e8011),
	.w8(32'hbbb3433f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76a523),
	.w1(32'h3c0067bb),
	.w2(32'h3b450983),
	.w3(32'h3bc7eb2a),
	.w4(32'h3bf238da),
	.w5(32'h3b458453),
	.w6(32'hbb7a1e9d),
	.w7(32'hbb94ab36),
	.w8(32'h3aaba257),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15f71a),
	.w1(32'h3bcd09f2),
	.w2(32'h3c3abf38),
	.w3(32'h3b9bc5ed),
	.w4(32'h3b9b4c01),
	.w5(32'h3a8bebba),
	.w6(32'h3a94bb2f),
	.w7(32'h3b218f09),
	.w8(32'h3c3788df),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea9948),
	.w1(32'h3c0e911f),
	.w2(32'h3b946e42),
	.w3(32'hbc0cf9dc),
	.w4(32'hbbd2e055),
	.w5(32'h3b376fd2),
	.w6(32'h3b10717a),
	.w7(32'h3b2034da),
	.w8(32'h3bb83e9b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c336814),
	.w1(32'h3c38d8c6),
	.w2(32'h3b87c9b4),
	.w3(32'h3bba8038),
	.w4(32'h3bb63e0e),
	.w5(32'h3a221944),
	.w6(32'h3bb66297),
	.w7(32'h3b29fd7a),
	.w8(32'hbc26bbf9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1f10c),
	.w1(32'h3b5b7605),
	.w2(32'hbb7a2d23),
	.w3(32'h3bdbed79),
	.w4(32'h3bd81fd4),
	.w5(32'hbb8dd84c),
	.w6(32'h3a58d3e1),
	.w7(32'h3b7d8a16),
	.w8(32'hbbdbf3bb),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a2b93),
	.w1(32'h3b2f40b5),
	.w2(32'hbc43fb29),
	.w3(32'hbba387ee),
	.w4(32'hbbdc2bff),
	.w5(32'hbb90e3de),
	.w6(32'hbc52e2f7),
	.w7(32'hbc3d005a),
	.w8(32'hbbd5cbf8),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e684a),
	.w1(32'hbc149364),
	.w2(32'h3c1ec327),
	.w3(32'hbb54af86),
	.w4(32'hbc02c005),
	.w5(32'hbaaab35e),
	.w6(32'hbc3c3e8d),
	.w7(32'hbc43789a),
	.w8(32'hbbedd5a7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ff76f),
	.w1(32'h3ca0d561),
	.w2(32'h3c97fcae),
	.w3(32'h3ba1051f),
	.w4(32'h3c211f24),
	.w5(32'h3b8bd563),
	.w6(32'hbc4cc20d),
	.w7(32'hba87d107),
	.w8(32'hbc3a829b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1e3ec4),
	.w1(32'h3cf31932),
	.w2(32'hbb650254),
	.w3(32'h3c3ca536),
	.w4(32'h3c8696b8),
	.w5(32'hbb106102),
	.w6(32'hbce1576a),
	.w7(32'hbc597276),
	.w8(32'h3b0b6b12),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1303e4),
	.w1(32'h3a8645f5),
	.w2(32'hba6d11af),
	.w3(32'h3c0354c7),
	.w4(32'h3bcbaf5a),
	.w5(32'h3a2ae8e4),
	.w6(32'h3bae2f69),
	.w7(32'h38b8290d),
	.w8(32'hbb01f304),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b204af2),
	.w1(32'hbaacba6a),
	.w2(32'h3c4ff38f),
	.w3(32'hba3081c0),
	.w4(32'h399f93fc),
	.w5(32'h3b447898),
	.w6(32'hbb9c7510),
	.w7(32'hbb948cd0),
	.w8(32'hb98bc1d5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f9e9),
	.w1(32'h3b8cd646),
	.w2(32'hbbdee478),
	.w3(32'h3bcf3677),
	.w4(32'h3c1c6a12),
	.w5(32'hba8b1ade),
	.w6(32'h3bc644f6),
	.w7(32'hba6be92a),
	.w8(32'hbba61a26),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a1907),
	.w1(32'h3c0bd015),
	.w2(32'h395b950d),
	.w3(32'hbb0cc07f),
	.w4(32'hbb0eee04),
	.w5(32'hbbdf186a),
	.w6(32'hbc39f523),
	.w7(32'hbb6fa633),
	.w8(32'hbc2ca808),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb5360),
	.w1(32'h3c1e6d55),
	.w2(32'h3c48d750),
	.w3(32'hbb3fdae7),
	.w4(32'h399680c1),
	.w5(32'h3c2f6a7b),
	.w6(32'hbba0447b),
	.w7(32'hbbbb08e8),
	.w8(32'hb9ac963a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule