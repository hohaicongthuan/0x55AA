module layer_10_featuremap_203(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbde2a4),
	.w1(32'h3bccc8fc),
	.w2(32'h3d0ca123),
	.w3(32'h3bb8f849),
	.w4(32'hbbef7277),
	.w5(32'h3b222a2f),
	.w6(32'h3b08e307),
	.w7(32'hbb58d428),
	.w8(32'h3b330481),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60158e),
	.w1(32'hba30e93c),
	.w2(32'hb4ffdc56),
	.w3(32'h3c48eb5f),
	.w4(32'hbba77d62),
	.w5(32'hba07fd76),
	.w6(32'h3a72a86b),
	.w7(32'h3b8b74be),
	.w8(32'h3c088a4a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf60db6),
	.w1(32'hbb0bd9b2),
	.w2(32'hbc17fc8b),
	.w3(32'h3bceff22),
	.w4(32'hbbe1dc5b),
	.w5(32'hbbea41a1),
	.w6(32'h3b04acae),
	.w7(32'hbbeefc84),
	.w8(32'hbb5edf12),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1701ec),
	.w1(32'hbc7dbe03),
	.w2(32'hba1ca5a3),
	.w3(32'h3a36c2e5),
	.w4(32'hbc5515f6),
	.w5(32'hbb455df1),
	.w6(32'hbc394e6b),
	.w7(32'hb95948d7),
	.w8(32'h3bf3708d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c3be3),
	.w1(32'hbbf55339),
	.w2(32'hbd0c9a09),
	.w3(32'h3b6ee09f),
	.w4(32'hbb28e42d),
	.w5(32'hbc1b4eb7),
	.w6(32'hbc078a64),
	.w7(32'hbc29c4ad),
	.w8(32'h3b3a4fb5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25d710),
	.w1(32'hbd2372f2),
	.w2(32'hbbd02db5),
	.w3(32'hbc04dd5f),
	.w4(32'hbccc1ce2),
	.w5(32'hbca9792a),
	.w6(32'hbc807682),
	.w7(32'h3c4d98ca),
	.w8(32'h3cd75ab2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d363217),
	.w1(32'h3bb1fb16),
	.w2(32'hbc106ee2),
	.w3(32'h3c5334c3),
	.w4(32'hbba96a63),
	.w5(32'hbad31ae8),
	.w6(32'h3a4c527f),
	.w7(32'hbb938c32),
	.w8(32'h3afb125c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05c49d),
	.w1(32'hbc21fdc9),
	.w2(32'h3b6a772d),
	.w3(32'h3ad2695e),
	.w4(32'h3b54cd81),
	.w5(32'hb9d32516),
	.w6(32'hbb079d19),
	.w7(32'h3b818443),
	.w8(32'hbad3d4cd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43b48),
	.w1(32'hbc01142b),
	.w2(32'h3c09bb35),
	.w3(32'hbb093c7d),
	.w4(32'h3b3d7cc2),
	.w5(32'hbb4e2510),
	.w6(32'h3c27499b),
	.w7(32'h3bee3e1f),
	.w8(32'hbb8d0333),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0dd6),
	.w1(32'h3ca572d9),
	.w2(32'hbc038615),
	.w3(32'hbb7f4283),
	.w4(32'hbabe4d22),
	.w5(32'hbb18b294),
	.w6(32'h3bc7cea6),
	.w7(32'hbc4040bf),
	.w8(32'hbb457aaa),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35e011),
	.w1(32'hbb0dfe6d),
	.w2(32'hbb95f82a),
	.w3(32'h3b10eed3),
	.w4(32'h3af20ae9),
	.w5(32'h3bf9d889),
	.w6(32'h3b82ea14),
	.w7(32'hba96e5e5),
	.w8(32'h3b3ff962),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10a707),
	.w1(32'hbc1500d7),
	.w2(32'hbc9f871a),
	.w3(32'h3c310f8e),
	.w4(32'hbb41460a),
	.w5(32'hbc2dfb4d),
	.w6(32'hbc1d2c9b),
	.w7(32'hbc2ce0d2),
	.w8(32'hbbfe3e9e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53d31e),
	.w1(32'hb9cbb008),
	.w2(32'hbace8e33),
	.w3(32'hbc8c939b),
	.w4(32'h3b8595c4),
	.w5(32'hbb8ac347),
	.w6(32'h3b16b70e),
	.w7(32'hbaf78ef3),
	.w8(32'hbb8f5540),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58b535),
	.w1(32'h3cc149c6),
	.w2(32'h3c6a9d09),
	.w3(32'h39db336b),
	.w4(32'h3d0aa268),
	.w5(32'h3c95ea54),
	.w6(32'h3c5add45),
	.w7(32'hbbccab69),
	.w8(32'hbce422c5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dbc3f),
	.w1(32'hbbf28cfd),
	.w2(32'hbcffb596),
	.w3(32'hbc0d54ce),
	.w4(32'h3bbb0a3f),
	.w5(32'hbb61a5dc),
	.w6(32'hbc6ecb5b),
	.w7(32'hbc18a879),
	.w8(32'hba6c4b28),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb112b71),
	.w1(32'hbc8be085),
	.w2(32'h3bf1271f),
	.w3(32'hbc07c334),
	.w4(32'hbba3b710),
	.w5(32'hbbc82c35),
	.w6(32'h3a526826),
	.w7(32'h3c444366),
	.w8(32'h3ba94fb7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3de98),
	.w1(32'hbb6a1571),
	.w2(32'h3a86b4f1),
	.w3(32'hbaed8337),
	.w4(32'h3b2b31f9),
	.w5(32'h3b6f6c8d),
	.w6(32'hb9eb8503),
	.w7(32'h3b97053c),
	.w8(32'hbab4a02b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa75dc7),
	.w1(32'h3c2f0368),
	.w2(32'hbc0605e6),
	.w3(32'hbc10c6db),
	.w4(32'hbbb01ff8),
	.w5(32'hbbc04c54),
	.w6(32'h3bc58281),
	.w7(32'hbc08d342),
	.w8(32'hbb3187b9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03de4a),
	.w1(32'hb9dc273a),
	.w2(32'h39da5b63),
	.w3(32'hb999e4a6),
	.w4(32'hbb4edaf0),
	.w5(32'h3ad45c6c),
	.w6(32'hbac7c3be),
	.w7(32'h3a7fc60b),
	.w8(32'h3bbedd78),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78b128),
	.w1(32'hbbccc2d6),
	.w2(32'h3ba56949),
	.w3(32'h3b75ac4d),
	.w4(32'hbb14846b),
	.w5(32'hbb796721),
	.w6(32'h3b251e56),
	.w7(32'h3b621fb6),
	.w8(32'hba2c2b32),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b306375),
	.w1(32'hbc59669c),
	.w2(32'h3b199ecb),
	.w3(32'hbb058f92),
	.w4(32'h3bf278f1),
	.w5(32'h3a82ac72),
	.w6(32'hbab0fc0d),
	.w7(32'h3bad5e54),
	.w8(32'h39b28052),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfea4f),
	.w1(32'hbc46fbc3),
	.w2(32'hbcc3c99d),
	.w3(32'hbb9694d6),
	.w4(32'hb9965bbf),
	.w5(32'hbb6285ab),
	.w6(32'h3ad003d1),
	.w7(32'hbc300d9f),
	.w8(32'hbbf83742),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcebea6c),
	.w1(32'hbab7d8c1),
	.w2(32'hbb8fa810),
	.w3(32'hbc141b47),
	.w4(32'h3af090fb),
	.w5(32'hbba6b856),
	.w6(32'h3b8c361f),
	.w7(32'hbbbd6718),
	.w8(32'hb9d694cc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983d726),
	.w1(32'hbc26ae99),
	.w2(32'h3bfa34d4),
	.w3(32'h388aeb36),
	.w4(32'h3bada390),
	.w5(32'hb87a4a6f),
	.w6(32'h39963e51),
	.w7(32'h3bf8ff9a),
	.w8(32'h3a1457f3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c042971),
	.w1(32'hbaf6781c),
	.w2(32'hba8c97ce),
	.w3(32'hba5dbd2c),
	.w4(32'h3aafa610),
	.w5(32'hbc07bdc2),
	.w6(32'hba9029bf),
	.w7(32'hbb837bd4),
	.w8(32'h3b267931),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c373d87),
	.w1(32'h3bc82525),
	.w2(32'h3c14f339),
	.w3(32'h3b45264c),
	.w4(32'h3bf476d5),
	.w5(32'h3bb9ecf5),
	.w6(32'hbb5a8e0f),
	.w7(32'hbb3254f9),
	.w8(32'hba94018b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e330),
	.w1(32'hbbd6cc5b),
	.w2(32'h3af7f159),
	.w3(32'h39edcefd),
	.w4(32'h3aa47dfc),
	.w5(32'hbb85ab28),
	.w6(32'h39cebb3e),
	.w7(32'h3bc254c2),
	.w8(32'h3ab59ed1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0e66e),
	.w1(32'hbb2bfc20),
	.w2(32'hbaa452b9),
	.w3(32'hbb224fde),
	.w4(32'hbbec1a9e),
	.w5(32'hbc4393a4),
	.w6(32'h399fa126),
	.w7(32'h3b0781d9),
	.w8(32'h3bfac61d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bdfc5),
	.w1(32'h3b99fa69),
	.w2(32'hbb4df00b),
	.w3(32'h3bd02970),
	.w4(32'h3b890dee),
	.w5(32'hbc18e3a3),
	.w6(32'h3bb611a6),
	.w7(32'hbbf2018a),
	.w8(32'hbc027980),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73cd591),
	.w1(32'h3b10418f),
	.w2(32'h3ad1e509),
	.w3(32'hbba1301d),
	.w4(32'h3bc55c2e),
	.w5(32'h3b7e2155),
	.w6(32'h3ad2e12b),
	.w7(32'h3aa1a7af),
	.w8(32'hbba3bb73),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a0dda),
	.w1(32'hbbf9b8d1),
	.w2(32'hb9adf21c),
	.w3(32'hbb682fe8),
	.w4(32'h3ae06ecb),
	.w5(32'hbb3ffc1f),
	.w6(32'h395cc926),
	.w7(32'h3b6be853),
	.w8(32'h3b3ad19d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc555c2),
	.w1(32'hbc08df29),
	.w2(32'hbb634252),
	.w3(32'h39a144cb),
	.w4(32'h3abee4af),
	.w5(32'hbba99942),
	.w6(32'h3a4db21e),
	.w7(32'h3b4be5f4),
	.w8(32'h3b016466),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff697),
	.w1(32'h3b85a7c3),
	.w2(32'hbc06b4f3),
	.w3(32'h3a995da4),
	.w4(32'h3ba145c1),
	.w5(32'hbc108063),
	.w6(32'h3aec1a09),
	.w7(32'hbc5476cd),
	.w8(32'hbb1c719b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4b6eb),
	.w1(32'hbba4afb7),
	.w2(32'h3b191411),
	.w3(32'hbba27808),
	.w4(32'hbb10434d),
	.w5(32'h3c2a3442),
	.w6(32'hbb930fe8),
	.w7(32'h3bcab31f),
	.w8(32'h3b98fb45),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d7dd),
	.w1(32'h3a10fd7a),
	.w2(32'hbbb9f670),
	.w3(32'hbb73d7a6),
	.w4(32'hbc01233d),
	.w5(32'hbc0578f1),
	.w6(32'h3b9bec7d),
	.w7(32'h37d25260),
	.w8(32'h3a92d6a7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10c053),
	.w1(32'hbc1b2107),
	.w2(32'hbaa2e9b2),
	.w3(32'h3b9279e2),
	.w4(32'hbae52152),
	.w5(32'hbc13b408),
	.w6(32'hbb64ddc7),
	.w7(32'h3bfd1d9b),
	.w8(32'h3bcc6eec),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71a7e1),
	.w1(32'hbc36d7c1),
	.w2(32'hbc43aa40),
	.w3(32'hbbec3c5f),
	.w4(32'hbc3e63e9),
	.w5(32'hbbd13ed2),
	.w6(32'hbc0c5dc6),
	.w7(32'h3b32c1ae),
	.w8(32'h3c45ad79),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f759e),
	.w1(32'h3be92661),
	.w2(32'hbb127ea5),
	.w3(32'h3b9aec6b),
	.w4(32'h38834e3d),
	.w5(32'h3af3ca57),
	.w6(32'h3b721c3f),
	.w7(32'hb98bce59),
	.w8(32'h3b45a19f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2666a6),
	.w1(32'hbc74b702),
	.w2(32'h3bb1fe0f),
	.w3(32'h3ae81223),
	.w4(32'hb990b14e),
	.w5(32'hbb637b53),
	.w6(32'hba2ba91d),
	.w7(32'h3c282f32),
	.w8(32'h3bbc5f8f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5dce8e),
	.w1(32'h3ac24f13),
	.w2(32'hbb343dfb),
	.w3(32'h3ab45a7e),
	.w4(32'hbb8affdb),
	.w5(32'h3b04008e),
	.w6(32'hbae88ffb),
	.w7(32'h3abc6894),
	.w8(32'h3b66a630),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a840fe6),
	.w1(32'h3bbc0cd4),
	.w2(32'h3943085e),
	.w3(32'h3b0e1684),
	.w4(32'h3c2bbb4f),
	.w5(32'h3b1b6dbc),
	.w6(32'h3a9804f9),
	.w7(32'h3a429edb),
	.w8(32'hbb8e79ea),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab84dfc),
	.w1(32'hbbb6da9a),
	.w2(32'h3b740cb0),
	.w3(32'hbb30c99f),
	.w4(32'hbc13442a),
	.w5(32'hba7df051),
	.w6(32'hbb506aa9),
	.w7(32'h3b3f34bb),
	.w8(32'h3bb71304),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3610df),
	.w1(32'hb9aa63dc),
	.w2(32'h3b5cab73),
	.w3(32'h3be1f083),
	.w4(32'h3bbc42a9),
	.w5(32'h3aa0e47e),
	.w6(32'h3b9538de),
	.w7(32'h3bb0ccee),
	.w8(32'hbb0390aa),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5e8e0),
	.w1(32'h3d0a5bf0),
	.w2(32'hbb883c9c),
	.w3(32'h3a08f73e),
	.w4(32'h3bb72b4f),
	.w5(32'h3be33dc9),
	.w6(32'h3c144703),
	.w7(32'hbc570757),
	.w8(32'hbb434285),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ff01d),
	.w1(32'h3cb66d10),
	.w2(32'h3b9f2215),
	.w3(32'h3b820eae),
	.w4(32'h3c16d364),
	.w5(32'h3a8fa4d8),
	.w6(32'h3bb4b055),
	.w7(32'hbcdd60ab),
	.w8(32'hbcd13a4c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1edaec),
	.w1(32'h3c957235),
	.w2(32'hbbb8e23e),
	.w3(32'hbc1277a2),
	.w4(32'h3be80b37),
	.w5(32'h3b956b1a),
	.w6(32'h3bb52d19),
	.w7(32'hbc3b9892),
	.w8(32'hbc6ee8a4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cde64),
	.w1(32'hbc07619f),
	.w2(32'hbcbe719c),
	.w3(32'hbbfc7403),
	.w4(32'hbbc422e1),
	.w5(32'hbbb20fa9),
	.w6(32'hbb31366a),
	.w7(32'h3b383150),
	.w8(32'hbbc158d5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8f8c),
	.w1(32'h3ba044f6),
	.w2(32'h3c09806f),
	.w3(32'hbc1537c4),
	.w4(32'h39484051),
	.w5(32'h3b21dc85),
	.w6(32'h3be07aa4),
	.w7(32'h3bfa298f),
	.w8(32'hbbb19970),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51861e),
	.w1(32'hbb4a7412),
	.w2(32'h3b50fd50),
	.w3(32'hbbe48ae5),
	.w4(32'hb6d547dc),
	.w5(32'hbb288360),
	.w6(32'h3b8526e9),
	.w7(32'h3bdc190e),
	.w8(32'h3b85e81c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cd90c),
	.w1(32'h38ecf1d5),
	.w2(32'h3bab906f),
	.w3(32'h3a8a953d),
	.w4(32'h3c237959),
	.w5(32'h3b7c8227),
	.w6(32'h3b326306),
	.w7(32'h3a9de301),
	.w8(32'hbc04f377),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4d25b),
	.w1(32'h3d3de997),
	.w2(32'hbbb16d18),
	.w3(32'hbb7bf0cd),
	.w4(32'h3c90ecd1),
	.w5(32'h3c6e4ed0),
	.w6(32'h3c2e1b0a),
	.w7(32'hbcb16f57),
	.w8(32'hbce24431),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd094828),
	.w1(32'hbb9df3ab),
	.w2(32'h3ce2ffac),
	.w3(32'hbbc1868f),
	.w4(32'hbb10405d),
	.w5(32'hbc415cb0),
	.w6(32'h3b9cc045),
	.w7(32'h3b7b96a6),
	.w8(32'h3ba359e2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86cd3e),
	.w1(32'hbd153fcb),
	.w2(32'h3c550d2c),
	.w3(32'hba27b2b7),
	.w4(32'hbcbdf16a),
	.w5(32'hbc4bd6f3),
	.w6(32'hbc79c0f0),
	.w7(32'h3c9bbcf8),
	.w8(32'h3cc9eb0e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d33506b),
	.w1(32'hbcba095d),
	.w2(32'hbcd5c64a),
	.w3(32'h3c6e09dd),
	.w4(32'hbc8a58cb),
	.w5(32'hbc732118),
	.w6(32'hbc6af6ea),
	.w7(32'hbb6f69e9),
	.w8(32'h3bb01f87),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5586d0),
	.w1(32'hbc060c79),
	.w2(32'h3ab49e3b),
	.w3(32'hb84ed383),
	.w4(32'hb9af9318),
	.w5(32'h3ab9d418),
	.w6(32'hbaadb00a),
	.w7(32'h3c08e3a5),
	.w8(32'h37ec7bf8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d0ac2),
	.w1(32'h3ba286ff),
	.w2(32'hbb162940),
	.w3(32'hbb3893bc),
	.w4(32'h3a97cbb9),
	.w5(32'hbb1cc525),
	.w6(32'h3abbe331),
	.w7(32'h3a227af4),
	.w8(32'h3bc0723f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacf155),
	.w1(32'h3c0fe309),
	.w2(32'h39c5c1fb),
	.w3(32'h3b33b6f6),
	.w4(32'h3b13e9c9),
	.w5(32'h3bf78644),
	.w6(32'h3b3822da),
	.w7(32'hbb51b330),
	.w8(32'hbc18ca77),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70ebe7),
	.w1(32'hbaa95009),
	.w2(32'hbd4d1536),
	.w3(32'hbb27b735),
	.w4(32'hbb914ef3),
	.w5(32'hbc0b7f57),
	.w6(32'hbc950f07),
	.w7(32'hbcd1fa2f),
	.w8(32'hbc56fe6d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc861038),
	.w1(32'h3bda704d),
	.w2(32'hb8bbb31c),
	.w3(32'hbc842776),
	.w4(32'h3a358f5b),
	.w5(32'hbac3c2f0),
	.w6(32'h3b7153ef),
	.w7(32'hb9cfce67),
	.w8(32'h3be880e6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70d5a4),
	.w1(32'hbc353443),
	.w2(32'h3c32ac1e),
	.w3(32'h3bf1565b),
	.w4(32'h3b0193b9),
	.w5(32'hba339321),
	.w6(32'h3b00b715),
	.w7(32'h3c20c9a4),
	.w8(32'h3b1ac5c2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4412b2),
	.w1(32'hbaeb466b),
	.w2(32'h3b352a8f),
	.w3(32'h3ad2f530),
	.w4(32'hbbe447c7),
	.w5(32'h3a62fa2b),
	.w6(32'hbad2b479),
	.w7(32'h3b10bfd4),
	.w8(32'h3b124a83),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9015a01),
	.w1(32'hb9bcd6f3),
	.w2(32'h3cad4d9c),
	.w3(32'h3babb92c),
	.w4(32'h3b417928),
	.w5(32'h3b98c6b4),
	.w6(32'h3b750f35),
	.w7(32'h3bc49596),
	.w8(32'hbbd58bbd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b08ca),
	.w1(32'hbcde7692),
	.w2(32'hbd774817),
	.w3(32'hb9b5f310),
	.w4(32'hbcb8b32f),
	.w5(32'hbd680a24),
	.w6(32'hbcb6a5b6),
	.w7(32'hbd46c50c),
	.w8(32'hbc8afb73),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d4287),
	.w1(32'h3ca750bd),
	.w2(32'hbb6d6503),
	.w3(32'hbd0550fc),
	.w4(32'h3aa6deec),
	.w5(32'h3b42a10a),
	.w6(32'h3ba5eb06),
	.w7(32'hbbf864fd),
	.w8(32'h3a85ae0e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8311b),
	.w1(32'hba1c4260),
	.w2(32'hb9b230b7),
	.w3(32'h3b740b67),
	.w4(32'hbae78a80),
	.w5(32'hbbbcd93e),
	.w6(32'h3b60f26a),
	.w7(32'h39bfcf94),
	.w8(32'h3a724294),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae305ee),
	.w1(32'h3c79de9f),
	.w2(32'hbc83e3a0),
	.w3(32'h3b78deb0),
	.w4(32'h3be40fef),
	.w5(32'h3c233c40),
	.w6(32'h3aac4719),
	.w7(32'hbb5154de),
	.w8(32'hbb57a186),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf2684),
	.w1(32'h3ab15ea2),
	.w2(32'hbb84ebd3),
	.w3(32'hbba4b0b8),
	.w4(32'h3b1121b4),
	.w5(32'h3912b310),
	.w6(32'h3a481ae0),
	.w7(32'h3b3e78a1),
	.w8(32'h3a9bd0bf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b022d08),
	.w1(32'h3b156a69),
	.w2(32'h3b30d99e),
	.w3(32'h3b1bd9f9),
	.w4(32'h3b6530bc),
	.w5(32'hbb19dd18),
	.w6(32'h3b0fd2bc),
	.w7(32'h37c2c702),
	.w8(32'hbb9e9dad),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71acef),
	.w1(32'hbc990757),
	.w2(32'h3bd9f2d6),
	.w3(32'hbbf6e5cb),
	.w4(32'h3ab9ff54),
	.w5(32'hbb567826),
	.w6(32'hbbb43cf5),
	.w7(32'h3c6f7e76),
	.w8(32'h3bdc5890),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b83f5),
	.w1(32'h3d64c299),
	.w2(32'hbcc9a8df),
	.w3(32'h39f3c6a5),
	.w4(32'h3cf754a0),
	.w5(32'h3c97bf4f),
	.w6(32'h3c197c94),
	.w7(32'hbd0109d2),
	.w8(32'hbd406bed),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd66fdbb),
	.w1(32'h3b9de57d),
	.w2(32'hba85f50e),
	.w3(32'hbcb632f8),
	.w4(32'hbb2dbd51),
	.w5(32'hbb46baa6),
	.w6(32'h3bbf2a6a),
	.w7(32'h3a5737df),
	.w8(32'h3bbb5da3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf01f2),
	.w1(32'hbc6fcc34),
	.w2(32'hbb35e63a),
	.w3(32'h3b53770b),
	.w4(32'hb92c024c),
	.w5(32'hbb943b73),
	.w6(32'hbb7719e9),
	.w7(32'h3be322bd),
	.w8(32'h3ab45af3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d2b3f),
	.w1(32'hbc5fd4bb),
	.w2(32'h3bd81e22),
	.w3(32'hba05ce5a),
	.w4(32'hba00fd4e),
	.w5(32'hbb56bd9e),
	.w6(32'hba0ccf7f),
	.w7(32'h3c2eafbe),
	.w8(32'h3b8371ec),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42cd1a),
	.w1(32'hbc104466),
	.w2(32'h386b7897),
	.w3(32'h38a85c20),
	.w4(32'h3bb3c3ab),
	.w5(32'hbb8390fe),
	.w6(32'hbb1f462c),
	.w7(32'h3bcee87c),
	.w8(32'h3b9de22e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12e58c),
	.w1(32'h3a465be2),
	.w2(32'h3ae6c14f),
	.w3(32'hbb16295f),
	.w4(32'hbb0ce105),
	.w5(32'hbb814f57),
	.w6(32'h3b34f0ca),
	.w7(32'h3b37f34a),
	.w8(32'h3b5a960c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4238e0),
	.w1(32'h3c07cece),
	.w2(32'hb9e50867),
	.w3(32'h3b8535e6),
	.w4(32'h3bb44157),
	.w5(32'h3bd3710e),
	.w6(32'h3b94ef83),
	.w7(32'hbb902eb2),
	.w8(32'hbb94b923),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8d612),
	.w1(32'hbb5f4a8b),
	.w2(32'h3b585dfe),
	.w3(32'hbc13e9c9),
	.w4(32'h3c2db552),
	.w5(32'hb9a46639),
	.w6(32'h3b606c4d),
	.w7(32'hba807566),
	.w8(32'hbc2e6d3e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a2211),
	.w1(32'hbb03c082),
	.w2(32'hbc6ada45),
	.w3(32'hbbab4dae),
	.w4(32'hbc1cce43),
	.w5(32'hbc50f615),
	.w6(32'hbb3e9c4a),
	.w7(32'hbc5553fc),
	.w8(32'h3bb005f7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab57dd8),
	.w1(32'hbc2d53fe),
	.w2(32'h3c366c94),
	.w3(32'h3b9254b4),
	.w4(32'h3afd23df),
	.w5(32'h3bfd23fc),
	.w6(32'h3b00194d),
	.w7(32'h3c64ad17),
	.w8(32'h3bac1075),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc72f0),
	.w1(32'hbc49351a),
	.w2(32'hba976fa6),
	.w3(32'hbbbabb34),
	.w4(32'h3bd8b077),
	.w5(32'hbb494f18),
	.w6(32'h3b4bbb1d),
	.w7(32'h3bc0e0fb),
	.w8(32'hbb3d58df),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c632ce),
	.w1(32'h3b704156),
	.w2(32'h3b2f08a6),
	.w3(32'hbbb997a7),
	.w4(32'h3b1c974e),
	.w5(32'hbb5e3004),
	.w6(32'h3b1fee80),
	.w7(32'h3b3e1bae),
	.w8(32'h3a8ebbb2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba88425),
	.w1(32'hbb08b904),
	.w2(32'h3bb62180),
	.w3(32'hbb6a1b93),
	.w4(32'hbc0f6d12),
	.w5(32'h3ae09dfe),
	.w6(32'hbb01e78c),
	.w7(32'h3b6b65de),
	.w8(32'h3b808263),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2a5e1),
	.w1(32'hb9fb014e),
	.w2(32'h3b48d53d),
	.w3(32'h3c0eec96),
	.w4(32'hb8e6b50c),
	.w5(32'hbb9c09ef),
	.w6(32'h3a9cb048),
	.w7(32'h3b1e5685),
	.w8(32'h3ac87bab),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7c2ee),
	.w1(32'h3a7b873a),
	.w2(32'h3bafb6be),
	.w3(32'hb9a001cc),
	.w4(32'hbbb3e15a),
	.w5(32'h3ac9b630),
	.w6(32'h3b864ab8),
	.w7(32'h3bc418cf),
	.w8(32'h3b7b5205),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac58b69),
	.w1(32'hbaa3d1b2),
	.w2(32'h3b3ce51b),
	.w3(32'h3b941746),
	.w4(32'hb87c1ad0),
	.w5(32'h3b965607),
	.w6(32'h3bf98756),
	.w7(32'h3c1b0a26),
	.w8(32'hbb5f8680),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5e982),
	.w1(32'h3ba61a86),
	.w2(32'hba8a9104),
	.w3(32'hbbba0c14),
	.w4(32'hb9477be3),
	.w5(32'h3aa409b8),
	.w6(32'h3b82b8fa),
	.w7(32'h3b133daf),
	.w8(32'h3bc2c7b0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89fb47),
	.w1(32'h3cebf86e),
	.w2(32'hbb16fab4),
	.w3(32'h3bc43531),
	.w4(32'h3c9035a6),
	.w5(32'h3c3625d2),
	.w6(32'h3c24de80),
	.w7(32'hbc32f96e),
	.w8(32'hbaba7889),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7a7a7),
	.w1(32'hbbc6eec4),
	.w2(32'h3ae0674e),
	.w3(32'h3b42883a),
	.w4(32'h3bd58af9),
	.w5(32'h3a4d348c),
	.w6(32'h3a8cc73f),
	.w7(32'h3bb3c454),
	.w8(32'h3b243cf5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9aa75),
	.w1(32'hbc407b2a),
	.w2(32'h39581162),
	.w3(32'hba249b30),
	.w4(32'hbba6e7e1),
	.w5(32'hb6d114e5),
	.w6(32'hbb78402a),
	.w7(32'h3c0b5d1c),
	.w8(32'h3b80c6a9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eeaa2),
	.w1(32'hbc2ef34c),
	.w2(32'hbb091342),
	.w3(32'h3b09e064),
	.w4(32'h3bf63454),
	.w5(32'hbb514a5d),
	.w6(32'h3b3e29c0),
	.w7(32'h3bf0c695),
	.w8(32'hba5c38de),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81f54f2),
	.w1(32'hbb9cf59c),
	.w2(32'h3b79d2eb),
	.w3(32'hbbbce490),
	.w4(32'h3b598827),
	.w5(32'h396b0858),
	.w6(32'h3883db30),
	.w7(32'h3b78d73b),
	.w8(32'h3b3d7ebc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21e16b),
	.w1(32'h3caab04e),
	.w2(32'hbbd4b34d),
	.w3(32'h3b6f009c),
	.w4(32'h3c17ea17),
	.w5(32'h3ba3fb5a),
	.w6(32'h3bf684b4),
	.w7(32'hbc2867de),
	.w8(32'hbc1c1a40),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b871e),
	.w1(32'hbc66c99d),
	.w2(32'h3b0dc2fc),
	.w3(32'hbb71b298),
	.w4(32'hbc2b0ef7),
	.w5(32'hbbce0944),
	.w6(32'h3acaef32),
	.w7(32'h3c32f58f),
	.w8(32'h3c341d04),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bb939),
	.w1(32'h3812cf1b),
	.w2(32'h3a362bce),
	.w3(32'h3bc0ae90),
	.w4(32'hba0f37b1),
	.w5(32'hbbbbbd87),
	.w6(32'hbb42e484),
	.w7(32'hbb908d70),
	.w8(32'hbb40d5cc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b889b54),
	.w1(32'hbad785ea),
	.w2(32'hbba0b22c),
	.w3(32'hbb0badc8),
	.w4(32'hbbfdfa70),
	.w5(32'hbb8d3f4c),
	.w6(32'h399c8b59),
	.w7(32'hbb5026ea),
	.w8(32'h3a88265c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14b033),
	.w1(32'hbc91fb05),
	.w2(32'h3b5c2ab2),
	.w3(32'h3a8efa14),
	.w4(32'hbcb075dc),
	.w5(32'hbc225cf9),
	.w6(32'hbab74894),
	.w7(32'hbaa86d3d),
	.w8(32'h3c2ee746),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf5106c),
	.w1(32'hbaa5a9c0),
	.w2(32'hbb6a1936),
	.w3(32'h3cb445ab),
	.w4(32'hbab3d496),
	.w5(32'hbb9aa4d6),
	.w6(32'hbab11927),
	.w7(32'hbbe530e3),
	.w8(32'hbb1ebf78),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb053888),
	.w1(32'hbb0a25ee),
	.w2(32'hbc0869ee),
	.w3(32'h3af4a8fb),
	.w4(32'hbbc2bfbb),
	.w5(32'hbcbf8c28),
	.w6(32'h3c017b1e),
	.w7(32'hbbad8dff),
	.w8(32'h3be4ee3e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c9d28),
	.w1(32'hbbaee6ca),
	.w2(32'h3b0e24d6),
	.w3(32'h398b2e8b),
	.w4(32'hbc5dcfc9),
	.w5(32'hbb16aedb),
	.w6(32'hbb4ddc31),
	.w7(32'h3be33bdd),
	.w8(32'h3bf6590c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccaca2),
	.w1(32'hbc9dbd65),
	.w2(32'h3bee1ebb),
	.w3(32'h3c078f9e),
	.w4(32'hbc572102),
	.w5(32'hbc140955),
	.w6(32'hbb2ae9e3),
	.w7(32'h3c52fcac),
	.w8(32'h3c9f884f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8456b),
	.w1(32'h3bc3dcd1),
	.w2(32'hbc522ca7),
	.w3(32'h3c1ca0c7),
	.w4(32'hbbfa45d4),
	.w5(32'h3c90f076),
	.w6(32'hbc6451fa),
	.w7(32'hb9c14675),
	.w8(32'hbc0e92f4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab49297),
	.w1(32'h3bd18f85),
	.w2(32'hbbe377ee),
	.w3(32'h3aafb91e),
	.w4(32'hbb2488f3),
	.w5(32'hba9e2764),
	.w6(32'h3bae43df),
	.w7(32'hba3b22ae),
	.w8(32'h3b81efe3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac061dd),
	.w1(32'hbb90069f),
	.w2(32'h3ba9c10f),
	.w3(32'h3bdc28ff),
	.w4(32'h3c8605c6),
	.w5(32'h39484bbb),
	.w6(32'h3bad3abc),
	.w7(32'hbaf340c9),
	.w8(32'hbc8975f9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cf65b),
	.w1(32'hbc87d222),
	.w2(32'hbc17a05b),
	.w3(32'hbc043db1),
	.w4(32'hbaf7ed51),
	.w5(32'hbc16cf83),
	.w6(32'hbb640545),
	.w7(32'h3bbc35bf),
	.w8(32'h3b69c70c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c489915),
	.w1(32'hbb8b980c),
	.w2(32'h3b25e8aa),
	.w3(32'hbab492da),
	.w4(32'h3be63552),
	.w5(32'hbab73d81),
	.w6(32'h3b0e7834),
	.w7(32'hb8129f41),
	.w8(32'hbbd9164f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd4c94),
	.w1(32'hbb8d3d6a),
	.w2(32'h3b31d74b),
	.w3(32'hbb6f0336),
	.w4(32'h3a6d0dc9),
	.w5(32'hbb3373a1),
	.w6(32'h3b35154b),
	.w7(32'h3b5e96dc),
	.w8(32'h392ccff5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8b704),
	.w1(32'hbc604688),
	.w2(32'hbc310bae),
	.w3(32'hbb7cfdb8),
	.w4(32'hbc61c835),
	.w5(32'hbc1760fe),
	.w6(32'hbb07e3ce),
	.w7(32'hbb123f39),
	.w8(32'h3a4527bd),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcaf3e),
	.w1(32'hbc0ee39c),
	.w2(32'h3bce9a60),
	.w3(32'hbb93cada),
	.w4(32'h3b96b8f0),
	.w5(32'h3b47f3d4),
	.w6(32'hbafa7b8c),
	.w7(32'h3bb83e26),
	.w8(32'h3bab99d0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33ab8c),
	.w1(32'hbafb8bf5),
	.w2(32'h3b347a26),
	.w3(32'h3b547ed5),
	.w4(32'h3c0eb177),
	.w5(32'h3a1740e3),
	.w6(32'h3b30689a),
	.w7(32'hba98e595),
	.w8(32'hbc1a7d01),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c3935),
	.w1(32'h3ca40a80),
	.w2(32'hb8e5d5d8),
	.w3(32'hbb862330),
	.w4(32'h3b0a3e24),
	.w5(32'h3a7706d4),
	.w6(32'h3be35e9c),
	.w7(32'hbc8b18bd),
	.w8(32'hbc81f232),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac4dc4),
	.w1(32'hbc6c7dce),
	.w2(32'h3c4f9b49),
	.w3(32'h39bc3e0c),
	.w4(32'hbb37f92d),
	.w5(32'hbab22f2e),
	.w6(32'hba9f2db9),
	.w7(32'h3c4eda22),
	.w8(32'h3bcba498),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58cc78),
	.w1(32'hbba0a6d1),
	.w2(32'h3c917efc),
	.w3(32'hb90439be),
	.w4(32'hbc08f423),
	.w5(32'hbc3cd70b),
	.w6(32'hbb810b60),
	.w7(32'hbccd7177),
	.w8(32'hbce6e76b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdc670a),
	.w1(32'hbcba1b8b),
	.w2(32'h3bbcb819),
	.w3(32'hbc4178b0),
	.w4(32'hbbb2a109),
	.w5(32'hbbefa474),
	.w6(32'hbbd9ddcd),
	.w7(32'h3c93b4fc),
	.w8(32'h3c81040a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5aa13),
	.w1(32'h3c4da301),
	.w2(32'hbbc02a7f),
	.w3(32'h392a78ed),
	.w4(32'hb9bdb76b),
	.w5(32'hbb0bda54),
	.w6(32'hbb2e1a92),
	.w7(32'hbc1d3da9),
	.w8(32'h3b07e02f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9588c),
	.w1(32'h3be5fd00),
	.w2(32'h3c20de00),
	.w3(32'h3bcd491f),
	.w4(32'h3c27e3f6),
	.w5(32'h3b9a48fd),
	.w6(32'h3bbb7b0a),
	.w7(32'hba3f5e68),
	.w8(32'hbc2f0724),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0d1bb),
	.w1(32'hbb75db23),
	.w2(32'h3b77b68d),
	.w3(32'hbb8ff347),
	.w4(32'h3c44fe4b),
	.w5(32'hb9ccf51a),
	.w6(32'h3b7f5d0c),
	.w7(32'hba980378),
	.w8(32'hbc47831b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56e217),
	.w1(32'hbc8072e5),
	.w2(32'h3a40ffc7),
	.w3(32'hbbc1b8af),
	.w4(32'hba80b520),
	.w5(32'hbba26777),
	.w6(32'hbb9e18df),
	.w7(32'h3b93f7c6),
	.w8(32'h3ae8ec02),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a2e1b),
	.w1(32'hbca66398),
	.w2(32'h3a1a8d8f),
	.w3(32'hb984e03b),
	.w4(32'hbb977807),
	.w5(32'hbc08d507),
	.w6(32'hbbbb6cc4),
	.w7(32'h3bbffaed),
	.w8(32'h3ba2cd22),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c790cfc),
	.w1(32'h3a34e0ca),
	.w2(32'h3b610cf2),
	.w3(32'h3a208e50),
	.w4(32'h3ac7f9a7),
	.w5(32'h3b6f8364),
	.w6(32'h3bb16ba9),
	.w7(32'hba04baa4),
	.w8(32'hbc81d994),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a966f),
	.w1(32'h3bbfd655),
	.w2(32'hbbc94bd6),
	.w3(32'h3a8cfcaa),
	.w4(32'hbb071f39),
	.w5(32'h3bad8cb2),
	.w6(32'hbc0ea1a4),
	.w7(32'hbbaf62c4),
	.w8(32'h38fbbc81),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb8b48),
	.w1(32'hbccdc23b),
	.w2(32'hbbf7aff7),
	.w3(32'h39d2553a),
	.w4(32'hbc96a429),
	.w5(32'hbc950811),
	.w6(32'hbc854f19),
	.w7(32'h3a990c7c),
	.w8(32'h3c9be6cd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc77e3c),
	.w1(32'hbc528140),
	.w2(32'h3c86d6a2),
	.w3(32'h3bf7b6bb),
	.w4(32'hbc411eec),
	.w5(32'hb9571265),
	.w6(32'hbb3d6b6c),
	.w7(32'h3c1c8570),
	.w8(32'h3c360fed),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c814306),
	.w1(32'hbc2ae30f),
	.w2(32'h3c0fc345),
	.w3(32'h3c25bf3c),
	.w4(32'h3b840acc),
	.w5(32'hb6efa8e5),
	.w6(32'h39300803),
	.w7(32'h3c00fc8f),
	.w8(32'h3a8c383b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2974b8),
	.w1(32'hbbf91e43),
	.w2(32'hbaae66de),
	.w3(32'h3a3efbd1),
	.w4(32'hbc06ea92),
	.w5(32'h3b2d222f),
	.w6(32'hbc180ae0),
	.w7(32'hb95e1a5d),
	.w8(32'hbc104eaf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56f1bd),
	.w1(32'hbd40560c),
	.w2(32'h3b6ef010),
	.w3(32'hbb971009),
	.w4(32'hbd05774b),
	.w5(32'hbcb5e690),
	.w6(32'hbc7c1782),
	.w7(32'h3c96e1be),
	.w8(32'h3d1d8e7a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d845b5d),
	.w1(32'hbc24b013),
	.w2(32'h3b693c97),
	.w3(32'h3cccd35d),
	.w4(32'h3bd1d699),
	.w5(32'hbb0615e9),
	.w6(32'h3b3748bb),
	.w7(32'h3bc41c8b),
	.w8(32'h3b849355),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8ead9),
	.w1(32'h38f9e797),
	.w2(32'hba13e60a),
	.w3(32'h38b48cd7),
	.w4(32'hb9e21600),
	.w5(32'h3b5af104),
	.w6(32'h3a2b1782),
	.w7(32'h3b6325db),
	.w8(32'h3b335283),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c03a1),
	.w1(32'h3bddf397),
	.w2(32'h3b58be84),
	.w3(32'h3b744e1d),
	.w4(32'h3b373f62),
	.w5(32'h3b8c69e7),
	.w6(32'h3b74c930),
	.w7(32'h3bca1fa6),
	.w8(32'h3aad08a1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa13bb8),
	.w1(32'hbbcabc62),
	.w2(32'hbbda77ee),
	.w3(32'h3b0be4be),
	.w4(32'hbba66de7),
	.w5(32'hbb7769b9),
	.w6(32'hbbdf72e4),
	.w7(32'hbbc26e75),
	.w8(32'hbbd50f50),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe88a2b),
	.w1(32'h39fe85da),
	.w2(32'hba2e3a80),
	.w3(32'hbbde1b85),
	.w4(32'h3a72d38c),
	.w5(32'hba865ec7),
	.w6(32'h3b1f4597),
	.w7(32'hb8af98ff),
	.w8(32'h3a0a0bf0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e8a6f),
	.w1(32'h3b14d33e),
	.w2(32'h3b1515e3),
	.w3(32'hb842011f),
	.w4(32'hba2be0ad),
	.w5(32'hba5faa2b),
	.w6(32'h3a5d7d1d),
	.w7(32'h3abd8aa1),
	.w8(32'h3ad502de),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f5552),
	.w1(32'h38a50eda),
	.w2(32'h3a9cfaca),
	.w3(32'hb9a26ed4),
	.w4(32'h3ab090a2),
	.w5(32'h3bb59382),
	.w6(32'hbb95d6e3),
	.w7(32'hbb4d5e5f),
	.w8(32'h38dfce87),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4db9e4),
	.w1(32'hbb76be13),
	.w2(32'hbb34dc0f),
	.w3(32'h3c1850b8),
	.w4(32'hbb953d9c),
	.w5(32'hbbc9cc1d),
	.w6(32'hbb95fce4),
	.w7(32'hbb824c08),
	.w8(32'hbbee8987),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb532e0c),
	.w1(32'h3b6a0699),
	.w2(32'hbb108916),
	.w3(32'hbb8cc78b),
	.w4(32'hb85cce58),
	.w5(32'hba175fb2),
	.w6(32'h3a1d87cd),
	.w7(32'h3ae8c619),
	.w8(32'hba42eaff),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb874928),
	.w1(32'hba71d8cd),
	.w2(32'h37a2fe58),
	.w3(32'hbaa2b1fc),
	.w4(32'hbac579c9),
	.w5(32'hbad6a7e6),
	.w6(32'h3a3c566e),
	.w7(32'hbb19a029),
	.w8(32'hbb1730c6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba029156),
	.w1(32'h3b93f4e0),
	.w2(32'hb953b098),
	.w3(32'hba9f0dd6),
	.w4(32'h39821055),
	.w5(32'h3a7dfcc1),
	.w6(32'h3b3ba10d),
	.w7(32'h3b9b2629),
	.w8(32'h3a31e142),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39835b30),
	.w1(32'hbaaeb2c7),
	.w2(32'hbb43bf5d),
	.w3(32'h394cdf7c),
	.w4(32'hb91cf813),
	.w5(32'h3b08f72b),
	.w6(32'hba1c40c7),
	.w7(32'h3aaf1284),
	.w8(32'h3949ae64),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d911c),
	.w1(32'hbbdf3382),
	.w2(32'h3ad7778d),
	.w3(32'h3b8e9e93),
	.w4(32'hbc12dc10),
	.w5(32'hbbf6cafc),
	.w6(32'hbb6f4cbe),
	.w7(32'hbb5db7bf),
	.w8(32'hbb306fad),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb642055),
	.w1(32'h3ab23e90),
	.w2(32'hbb82db55),
	.w3(32'hbc024c58),
	.w4(32'hbb5118ca),
	.w5(32'hbc188f75),
	.w6(32'hbb1edbfb),
	.w7(32'hbb9dacfa),
	.w8(32'hbb1caee5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd28a4),
	.w1(32'hbb9c2539),
	.w2(32'hbbaf00ff),
	.w3(32'hbc242ef9),
	.w4(32'hbbdffaaa),
	.w5(32'hbb89205b),
	.w6(32'h3a4278c4),
	.w7(32'hba17aab2),
	.w8(32'hba33d3fe),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39732c5b),
	.w1(32'h3a4e6593),
	.w2(32'hbb74b69f),
	.w3(32'hba528394),
	.w4(32'hbb149c07),
	.w5(32'hbb8c1026),
	.w6(32'h3b375fc3),
	.w7(32'h3b998c9d),
	.w8(32'h3b2ccffc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88851b),
	.w1(32'h3c10b12c),
	.w2(32'h3b718db3),
	.w3(32'hbb323e46),
	.w4(32'h3bb07499),
	.w5(32'h3b9e7bdf),
	.w6(32'h3b94d579),
	.w7(32'h3bdd54f4),
	.w8(32'h3b5d9f4e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae523e),
	.w1(32'hbbf49734),
	.w2(32'hbbebea6e),
	.w3(32'h3b517ba8),
	.w4(32'hbc147abb),
	.w5(32'hbb867131),
	.w6(32'hbb24f604),
	.w7(32'hbb9ba4d7),
	.w8(32'hbbee3280),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb99fcb),
	.w1(32'h3b0f526b),
	.w2(32'hba72677e),
	.w3(32'hbc0fb4f5),
	.w4(32'h3b59a486),
	.w5(32'h3ba43fa8),
	.w6(32'h3ae71d69),
	.w7(32'h3b669f77),
	.w8(32'h3a9c19da),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ce61),
	.w1(32'h3a249756),
	.w2(32'hbb6a5b6d),
	.w3(32'h3bb13d50),
	.w4(32'h3b1655a5),
	.w5(32'hbb8380aa),
	.w6(32'hbaf414f8),
	.w7(32'hbb8a1490),
	.w8(32'hba1ea5ac),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a070f5b),
	.w1(32'hbbc2dac1),
	.w2(32'hbb888588),
	.w3(32'hbb32c871),
	.w4(32'hbbc3a762),
	.w5(32'hbbec4ffe),
	.w6(32'hba731c62),
	.w7(32'hbb93216b),
	.w8(32'hbb4c0987),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93857f),
	.w1(32'h3a71c651),
	.w2(32'hba46b4f8),
	.w3(32'hbbd58f32),
	.w4(32'h3a3aca8f),
	.w5(32'hba08bb6b),
	.w6(32'h3a8cb2cd),
	.w7(32'hba466721),
	.w8(32'hb943edde),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be8ec8),
	.w1(32'hbaf30f77),
	.w2(32'hbbbfca87),
	.w3(32'hb6865e9e),
	.w4(32'hba619e49),
	.w5(32'hbaa02818),
	.w6(32'hba7316d8),
	.w7(32'hb9980348),
	.w8(32'hba9d32c5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c9639),
	.w1(32'h3a8a4985),
	.w2(32'h3b1b3816),
	.w3(32'h3a238b36),
	.w4(32'h3b1562fc),
	.w5(32'h3bbbf85a),
	.w6(32'h3aa46a62),
	.w7(32'h3b9df191),
	.w8(32'h3bcfa53f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9da4e),
	.w1(32'h3b948664),
	.w2(32'h3ac45b61),
	.w3(32'h3c1e8725),
	.w4(32'h3b289054),
	.w5(32'hbc19331f),
	.w6(32'h3b3f24eb),
	.w7(32'h3b8c2842),
	.w8(32'h3b388726),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d0048),
	.w1(32'hbc17e772),
	.w2(32'hbc4535b5),
	.w3(32'hbb9e45cb),
	.w4(32'hbafffb73),
	.w5(32'hbbc00fd4),
	.w6(32'hbb47ae85),
	.w7(32'hbc0f190a),
	.w8(32'hba67df6c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe3e76),
	.w1(32'h3bd2a85a),
	.w2(32'h3a57568d),
	.w3(32'h3a656c12),
	.w4(32'h3b260112),
	.w5(32'h3b31334a),
	.w6(32'h3b7f85e3),
	.w7(32'h3bb31182),
	.w8(32'h3ac4d96f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa36d41),
	.w1(32'hbae6c43c),
	.w2(32'h3a5bab4e),
	.w3(32'h3a861f66),
	.w4(32'hbabfbf84),
	.w5(32'h39bf70f0),
	.w6(32'hbb837d78),
	.w7(32'hb9a64064),
	.w8(32'hb8e9d072),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb30c4),
	.w1(32'h3a73c82f),
	.w2(32'hbc163418),
	.w3(32'h3afc23e0),
	.w4(32'h3b8d2936),
	.w5(32'h3b96a8ca),
	.w6(32'hbace2e9f),
	.w7(32'hbbf72866),
	.w8(32'hba821008),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b9dd7),
	.w1(32'hbb548b05),
	.w2(32'hbb9c9c63),
	.w3(32'h3b89b1db),
	.w4(32'hbb39a9cd),
	.w5(32'hba3329df),
	.w6(32'hbb0d2ebb),
	.w7(32'hb846fdba),
	.w8(32'hbac181ee),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2dcbc),
	.w1(32'hbb04a4db),
	.w2(32'h3a4d11cb),
	.w3(32'hba01d373),
	.w4(32'hbb12db2d),
	.w5(32'h3b260ab2),
	.w6(32'hbaf4fc6c),
	.w7(32'h3abb4ef2),
	.w8(32'h3aed1ed8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f108c),
	.w1(32'hbb9ef36c),
	.w2(32'h3aaf1742),
	.w3(32'h3bc90530),
	.w4(32'hbbcaee30),
	.w5(32'h39de1076),
	.w6(32'hbc11618e),
	.w7(32'hb908102c),
	.w8(32'hbbbd0998),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb746f4e),
	.w1(32'hbbc92758),
	.w2(32'hbbb83400),
	.w3(32'hbb86d6bd),
	.w4(32'hbba12df9),
	.w5(32'hbb961a1a),
	.w6(32'hbbc42eae),
	.w7(32'hbbaebe81),
	.w8(32'hbb922c43),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb465a5e),
	.w1(32'hba376956),
	.w2(32'h3a8e0417),
	.w3(32'hbb311601),
	.w4(32'hba0bac00),
	.w5(32'h3b3906ab),
	.w6(32'hb9d98656),
	.w7(32'h3b432b58),
	.w8(32'h3b494c34),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b809104),
	.w1(32'hbb34c01a),
	.w2(32'hbbefc016),
	.w3(32'h3b936a69),
	.w4(32'hbb909320),
	.w5(32'hbb60501a),
	.w6(32'hbb298aa4),
	.w7(32'hbb258d65),
	.w8(32'hbb308d74),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba021b3),
	.w1(32'hbbbac28b),
	.w2(32'hbbd08246),
	.w3(32'hbb4af614),
	.w4(32'hbb3fcc80),
	.w5(32'hbaee7784),
	.w6(32'hba2cf9f2),
	.w7(32'h3b14b817),
	.w8(32'h3bcdd333),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8982f1),
	.w1(32'h3bb0e1e6),
	.w2(32'hbc3ee7b6),
	.w3(32'h3baabd4f),
	.w4(32'h3b5e3028),
	.w5(32'hb9c6d72f),
	.w6(32'h3a8bcd0f),
	.w7(32'hbc0531f4),
	.w8(32'hbc503713),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc945561),
	.w1(32'hbac9e9d9),
	.w2(32'h39ac2865),
	.w3(32'hbc33f262),
	.w4(32'hbb50fb31),
	.w5(32'hbb9012ed),
	.w6(32'h3aab8c3d),
	.w7(32'hba70ec9a),
	.w8(32'h39daf36c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b6d84),
	.w1(32'hbb8683c2),
	.w2(32'hbbf9b9ea),
	.w3(32'hbb27320a),
	.w4(32'hbb8c8c71),
	.w5(32'hbac6d2cd),
	.w6(32'hbb439a3d),
	.w7(32'hbb9ff9b5),
	.w8(32'hbb8817a0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242104),
	.w1(32'hbb52af35),
	.w2(32'hbbac832a),
	.w3(32'hbb357d91),
	.w4(32'hbbb1b4e4),
	.w5(32'hbc0e9f71),
	.w6(32'h3ae16f8d),
	.w7(32'hbabf1608),
	.w8(32'hb9fbb2d8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa20f91),
	.w1(32'hb9d6ce15),
	.w2(32'hba70cdb6),
	.w3(32'hbb8ece9b),
	.w4(32'hba6bf4d2),
	.w5(32'hbb575583),
	.w6(32'h3a91f91c),
	.w7(32'hbb18ec37),
	.w8(32'hbac358a4),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359070),
	.w1(32'h3c03728b),
	.w2(32'h3b56f9c7),
	.w3(32'hbb4cb957),
	.w4(32'h3b7eb4f9),
	.w5(32'h3b9e5b97),
	.w6(32'h3b9f8408),
	.w7(32'h3bd9cfe3),
	.w8(32'h3b1c6809),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e11f6),
	.w1(32'h3a6e2745),
	.w2(32'h39aa8c0f),
	.w3(32'h3b1643f5),
	.w4(32'h3a29e0cf),
	.w5(32'hba4ea7fd),
	.w6(32'h3b2d515d),
	.w7(32'hb9253ee7),
	.w8(32'hb85e1d28),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0fd7b),
	.w1(32'hbba8bed6),
	.w2(32'hbbeae545),
	.w3(32'hb9d7eba5),
	.w4(32'hbb83ff7b),
	.w5(32'hbbc76f70),
	.w6(32'hbb98bf07),
	.w7(32'hbbfe6e58),
	.w8(32'hbba11212),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb758019),
	.w1(32'hba1c48a0),
	.w2(32'hbb0db68c),
	.w3(32'hbb7c43b8),
	.w4(32'h3ad6098d),
	.w5(32'hb9f6310d),
	.w6(32'h3b0d969f),
	.w7(32'h378479e9),
	.w8(32'h3a869ff8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56c916),
	.w1(32'hbb8684d0),
	.w2(32'hbc30a046),
	.w3(32'h3a1bd7f2),
	.w4(32'hbb917761),
	.w5(32'hbbcfd1b3),
	.w6(32'hbb023eb2),
	.w7(32'hbb14fd64),
	.w8(32'hb9fca94b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a62d5),
	.w1(32'hbc21368a),
	.w2(32'h3b5252e6),
	.w3(32'hbb26a2fc),
	.w4(32'hbc7e3b69),
	.w5(32'hbc6cb31b),
	.w6(32'hbc181b37),
	.w7(32'hbc1d364d),
	.w8(32'hbc6047c0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fb3c8),
	.w1(32'hbb104c4b),
	.w2(32'h3b950b48),
	.w3(32'hbcb5b8df),
	.w4(32'h3b5f3286),
	.w5(32'h3ba01ecb),
	.w6(32'hbbe7c901),
	.w7(32'hbba894a3),
	.w8(32'hbaef23c4),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16af9f),
	.w1(32'hbb3adc02),
	.w2(32'h39c2ca07),
	.w3(32'h3ad64d6c),
	.w4(32'hbb8c0c65),
	.w5(32'h391d35d6),
	.w6(32'hbbca0768),
	.w7(32'hbb80b391),
	.w8(32'hbb8e33a1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005416),
	.w1(32'hbb98f288),
	.w2(32'h38207d64),
	.w3(32'h3a8fa293),
	.w4(32'hbc34fced),
	.w5(32'hbb9defb6),
	.w6(32'h3a80bc11),
	.w7(32'hbb42e030),
	.w8(32'hbbade16c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac60867),
	.w1(32'hbbcc3eab),
	.w2(32'hbbd0a3c7),
	.w3(32'hbb5b49b8),
	.w4(32'hbb8e8428),
	.w5(32'hbbbe932b),
	.w6(32'hbbf8d6d0),
	.w7(32'hbbf436b5),
	.w8(32'hbbd6cb48),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd65ef4),
	.w1(32'hbb3cea92),
	.w2(32'hbc2b483b),
	.w3(32'hbbafe7ea),
	.w4(32'hbb616691),
	.w5(32'hbbb2064e),
	.w6(32'hbb2b7397),
	.w7(32'hbb7abfbb),
	.w8(32'hbb019563),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cbc6a),
	.w1(32'h3ba14825),
	.w2(32'h3aaf2c08),
	.w3(32'hbb427903),
	.w4(32'h3ad75191),
	.w5(32'h3af51910),
	.w6(32'h3b241bd1),
	.w7(32'h3b93aca0),
	.w8(32'h3acb5ca1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1c5d4),
	.w1(32'hbbe96030),
	.w2(32'h3b37e15a),
	.w3(32'h3a757b99),
	.w4(32'hbba00283),
	.w5(32'hbac0c36e),
	.w6(32'hbb8c073f),
	.w7(32'hb9aaad34),
	.w8(32'hba570846),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1a38d),
	.w1(32'hbb527c06),
	.w2(32'hbc583769),
	.w3(32'hbb47effb),
	.w4(32'hbbcbde03),
	.w5(32'hbc21c0cf),
	.w6(32'hbba72136),
	.w7(32'hbbd6925f),
	.w8(32'hbc2b61c4),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb988a8f),
	.w1(32'hbab925cf),
	.w2(32'hbbf665fd),
	.w3(32'hbb8371d9),
	.w4(32'h3a8354f9),
	.w5(32'h3a56f3bc),
	.w6(32'hba914cf9),
	.w7(32'h39aa0fa4),
	.w8(32'hb99fe9d0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb454127),
	.w1(32'h3a031de7),
	.w2(32'hbba9c680),
	.w3(32'h3b2ece60),
	.w4(32'hba264154),
	.w5(32'hbbaba127),
	.w6(32'hba02b01b),
	.w7(32'hbb827719),
	.w8(32'hbaaae57d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca7c49),
	.w1(32'hbb45b271),
	.w2(32'hbbbb76b0),
	.w3(32'h399220a0),
	.w4(32'hb9db8e0b),
	.w5(32'hbb92bd56),
	.w6(32'hbb0ca728),
	.w7(32'hbb8744e1),
	.w8(32'h3aa3cd65),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87ff528),
	.w1(32'hbb2939c6),
	.w2(32'hbbc16f28),
	.w3(32'hba07b18d),
	.w4(32'hbb46558e),
	.w5(32'hbb85ed3b),
	.w6(32'hbaefdaa2),
	.w7(32'hbb79ed39),
	.w8(32'hbb6632c4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cdb1d),
	.w1(32'hbadf0297),
	.w2(32'h3aa8013e),
	.w3(32'hbb688fbb),
	.w4(32'h3b7169f5),
	.w5(32'h3b915cb3),
	.w6(32'hba8d2a24),
	.w7(32'h39ad2e93),
	.w8(32'h3b67464a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e6708),
	.w1(32'hbaf2b2f2),
	.w2(32'h3b317d69),
	.w3(32'h3b989519),
	.w4(32'hbbc10116),
	.w5(32'h3b182b45),
	.w6(32'hbaac21e9),
	.w7(32'h3b706808),
	.w8(32'h3b6c8f76),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54fcee),
	.w1(32'h39ed50eb),
	.w2(32'h3b786165),
	.w3(32'h3b1ff800),
	.w4(32'hb9d47d0e),
	.w5(32'h3a41912d),
	.w6(32'h39d68935),
	.w7(32'h3a3dd73a),
	.w8(32'h3a5e6294),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b153da),
	.w1(32'h3bffbb2a),
	.w2(32'h3b213d2c),
	.w3(32'hba0e1f16),
	.w4(32'h3b77ad97),
	.w5(32'h3b8a8a58),
	.w6(32'h3b9e1be7),
	.w7(32'h3bcf5849),
	.w8(32'h3b023ffb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13016f),
	.w1(32'h3abff62b),
	.w2(32'hba76b2d6),
	.w3(32'h3b075759),
	.w4(32'h3a8b724b),
	.w5(32'hbaba604d),
	.w6(32'h3b4828e5),
	.w7(32'hba86dc15),
	.w8(32'hba0c037e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d5524),
	.w1(32'h3b954886),
	.w2(32'h3aec73d0),
	.w3(32'h38659a7a),
	.w4(32'h3b0ea9a7),
	.w5(32'hb945165b),
	.w6(32'h3b28d3c7),
	.w7(32'h3b6cc321),
	.w8(32'h39b158de),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a28dc),
	.w1(32'hbb81c0cd),
	.w2(32'hbc31213a),
	.w3(32'h3a9278b4),
	.w4(32'hb8be5a76),
	.w5(32'hba8f678c),
	.w6(32'h3ad24b8c),
	.w7(32'hb9c0c681),
	.w8(32'h3bc50be3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc190d7),
	.w1(32'hbbd06ee9),
	.w2(32'h3b1191f8),
	.w3(32'h3bc5c557),
	.w4(32'hbc20b190),
	.w5(32'hbc159f92),
	.w6(32'hbbc03590),
	.w7(32'hbbc79f48),
	.w8(32'hbc0b64a2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf24f2e),
	.w1(32'h3acd6c07),
	.w2(32'h3af67103),
	.w3(32'hbc644ac6),
	.w4(32'hba5ddf76),
	.w5(32'h3a67bdd0),
	.w6(32'h3947c5a4),
	.w7(32'h3aa05815),
	.w8(32'h3a2d2a41),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d63db),
	.w1(32'hba01effb),
	.w2(32'h3ba069d3),
	.w3(32'h3a8529b3),
	.w4(32'hbbb39233),
	.w5(32'h3b13d7ac),
	.w6(32'hbb943635),
	.w7(32'h3bb4ebd4),
	.w8(32'h3ae8859b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fba9a),
	.w1(32'hbabe8c65),
	.w2(32'hbb9632bd),
	.w3(32'h3ab7ac9f),
	.w4(32'hb9adc68b),
	.w5(32'hbb6bcf1a),
	.w6(32'h3a8fd17b),
	.w7(32'hbae9ff57),
	.w8(32'hba162332),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf03c60),
	.w1(32'hbc160081),
	.w2(32'hbc30d23e),
	.w3(32'hbb220173),
	.w4(32'hbb75c5ad),
	.w5(32'hbbfc7b79),
	.w6(32'hbbb62e22),
	.w7(32'hbc2d2942),
	.w8(32'hbb90bdfb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde60aa),
	.w1(32'h3ba603c1),
	.w2(32'h3a633411),
	.w3(32'hbb1ff3ac),
	.w4(32'h3b51d047),
	.w5(32'h3bc71536),
	.w6(32'h3b8257d3),
	.w7(32'h3ba8dbdd),
	.w8(32'h3b120fd7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56834c),
	.w1(32'hbb9d3903),
	.w2(32'h3bd717b7),
	.w3(32'h3bbac4fa),
	.w4(32'hbc24bda9),
	.w5(32'hbb01e24f),
	.w6(32'hbbec9e94),
	.w7(32'hba0efbde),
	.w8(32'h39fe5a5f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a677e),
	.w1(32'hbb28f947),
	.w2(32'hbb091e35),
	.w3(32'h39d2dce1),
	.w4(32'hbb055d8b),
	.w5(32'hbb2c7aae),
	.w6(32'hba85a1f7),
	.w7(32'hbb648e0c),
	.w8(32'hbb0b5b2a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cc139),
	.w1(32'h3bd05141),
	.w2(32'h3b279bdd),
	.w3(32'hbb7e5264),
	.w4(32'h3b4c1d99),
	.w5(32'h3b75e847),
	.w6(32'h3b886843),
	.w7(32'h3bc4b2ff),
	.w8(32'h3a4ed00e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a2014),
	.w1(32'h3beb57c6),
	.w2(32'h3b1d05cd),
	.w3(32'h3ae466a5),
	.w4(32'h3b6d821d),
	.w5(32'h3b8c1a94),
	.w6(32'h3b98da0e),
	.w7(32'h3bbed09e),
	.w8(32'h3b0dc9e5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f93b4),
	.w1(32'hbba381d8),
	.w2(32'hbc1d838d),
	.w3(32'h3b0dda62),
	.w4(32'hbbcdf78c),
	.w5(32'hbb9c2717),
	.w6(32'hbb72dabe),
	.w7(32'hbb7a6661),
	.w8(32'hbb3ae59d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9545b3),
	.w1(32'h3988477e),
	.w2(32'h3b4a52dd),
	.w3(32'hbb88f832),
	.w4(32'hb9022399),
	.w5(32'h3a88f689),
	.w6(32'hb912ba64),
	.w7(32'h3a9ab516),
	.w8(32'h3aa7fc40),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abee2d5),
	.w1(32'hbb37e533),
	.w2(32'hbc1b567d),
	.w3(32'h3a2b901c),
	.w4(32'h389dd0f6),
	.w5(32'h3af73eb4),
	.w6(32'h3b9a1cab),
	.w7(32'hba8e2ed9),
	.w8(32'hba68b879),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba50be8),
	.w1(32'h3aa34bfb),
	.w2(32'hbacba408),
	.w3(32'h3b854151),
	.w4(32'hbb9c572c),
	.w5(32'hbb4277e7),
	.w6(32'hbb2887a8),
	.w7(32'h3aef4921),
	.w8(32'hbb5655ee),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e8ce0),
	.w1(32'hb8655cad),
	.w2(32'hb9943d0f),
	.w3(32'hbb9c2d21),
	.w4(32'h3ab595fe),
	.w5(32'hb9eea434),
	.w6(32'h3a5261a8),
	.w7(32'hba91c96e),
	.w8(32'hbaf10ae1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ac9a3),
	.w1(32'hbc2424cb),
	.w2(32'hbc98ec4e),
	.w3(32'hbb176c9e),
	.w4(32'hbb2a1cf5),
	.w5(32'hbc0d41b4),
	.w6(32'hbbdc41b2),
	.w7(32'hbc1dee87),
	.w8(32'h39916108),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40b26a),
	.w1(32'hbb12930d),
	.w2(32'h3a8c45aa),
	.w3(32'hb74479f0),
	.w4(32'hbafb5ee5),
	.w5(32'h3bb19981),
	.w6(32'hbaf9611a),
	.w7(32'h3b961d31),
	.w8(32'h3bb83cb3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe76e6),
	.w1(32'hbb82eeed),
	.w2(32'hbb943a9a),
	.w3(32'h3c04eaf6),
	.w4(32'hbb19631d),
	.w5(32'hbb8ec363),
	.w6(32'hbb845b33),
	.w7(32'hbbea707c),
	.w8(32'hbb8e637b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f6bfb),
	.w1(32'h3b1a8c61),
	.w2(32'h3b27aefe),
	.w3(32'hbb0c297a),
	.w4(32'h3b32ceb8),
	.w5(32'h3a6eae9c),
	.w6(32'h3b292d36),
	.w7(32'h3ac16f72),
	.w8(32'h39d0fb21),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6e909),
	.w1(32'hbb69ea7e),
	.w2(32'hbb6d845c),
	.w3(32'h3aa715e3),
	.w4(32'hbaf27967),
	.w5(32'hba9baf6b),
	.w6(32'hbba7738d),
	.w7(32'hbb8b68d9),
	.w8(32'hbb687dd0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae6f9b),
	.w1(32'h39a8d624),
	.w2(32'h3a82a304),
	.w3(32'hbaa6b83b),
	.w4(32'h392315d5),
	.w5(32'h397a3c20),
	.w6(32'h3a9f3eb1),
	.w7(32'hba1e5082),
	.w8(32'hba152e45),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6abff1),
	.w1(32'hbb6616fc),
	.w2(32'hbc1d3408),
	.w3(32'hb94a2833),
	.w4(32'hb973e52d),
	.w5(32'hbbff6baf),
	.w6(32'hbb001658),
	.w7(32'hbbfca79f),
	.w8(32'hbad20efc),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8d070),
	.w1(32'h3b7c73ca),
	.w2(32'h3b3ae8a9),
	.w3(32'hbb273d76),
	.w4(32'h3b8b4026),
	.w5(32'h3b104236),
	.w6(32'h3b3156b4),
	.w7(32'h3a9f38d0),
	.w8(32'hb9cce2ab),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a419a01),
	.w1(32'hbbc1204a),
	.w2(32'hbbc7ac6e),
	.w3(32'h397e20b9),
	.w4(32'hbba528cb),
	.w5(32'hbb9b6c34),
	.w6(32'hbb862dea),
	.w7(32'hbbfdcc24),
	.w8(32'hbbfa6046),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10528e),
	.w1(32'h3a02d460),
	.w2(32'h3a8315df),
	.w3(32'hbbf3349e),
	.w4(32'h38798c3b),
	.w5(32'h3b292666),
	.w6(32'h39fa2c71),
	.w7(32'h3b46c50c),
	.w8(32'h3b253562),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4be865),
	.w1(32'hb8415216),
	.w2(32'hbb42d907),
	.w3(32'h3b811c1e),
	.w4(32'h3a7ff217),
	.w5(32'hbaff27fe),
	.w6(32'h37c657c7),
	.w7(32'hbb101879),
	.w8(32'h3ac35dd9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15f36f),
	.w1(32'h3a99969b),
	.w2(32'h3af1978e),
	.w3(32'h389bcb38),
	.w4(32'h3a9a9815),
	.w5(32'h3bc7f1a2),
	.w6(32'h3aee4473),
	.w7(32'h3ba4dbe1),
	.w8(32'h3bc50f47),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb330e),
	.w1(32'hba2ce825),
	.w2(32'hbb43cf01),
	.w3(32'h3bfde0fb),
	.w4(32'hbaf3074e),
	.w5(32'hbaf89bbb),
	.w6(32'hbb090659),
	.w7(32'hbaeeee7c),
	.w8(32'hbb260fe9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65c394),
	.w1(32'hbc0372cb),
	.w2(32'hbbb4028f),
	.w3(32'hba10535b),
	.w4(32'hbba84ae9),
	.w5(32'hbbeb2424),
	.w6(32'hbb94a798),
	.w7(32'hbbf2da21),
	.w8(32'hbb8ba9d8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe7b2b),
	.w1(32'hbb5333c5),
	.w2(32'hbbbe20a7),
	.w3(32'hbbd204c8),
	.w4(32'hbae01c5b),
	.w5(32'hbb51bcf3),
	.w6(32'hbac04eb4),
	.w7(32'hbb71b27b),
	.w8(32'hba5cbe2a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb831551),
	.w1(32'hbb1435d1),
	.w2(32'h38f700bb),
	.w3(32'hbac46639),
	.w4(32'hbb02e2eb),
	.w5(32'h39a2d5ea),
	.w6(32'hbb74ca65),
	.w7(32'hbaaec876),
	.w8(32'hbb8a2b30),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567808),
	.w1(32'h3a454a14),
	.w2(32'hba3eb83f),
	.w3(32'hbb4e0414),
	.w4(32'hba30abd6),
	.w5(32'hbaea0702),
	.w6(32'h3b047b9e),
	.w7(32'h3a027c97),
	.w8(32'h3a5a45de),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa4666),
	.w1(32'hba84fd94),
	.w2(32'hbb7ee50b),
	.w3(32'hba4617be),
	.w4(32'hbb8aa2b9),
	.w5(32'hbb4994b4),
	.w6(32'hbb62c36d),
	.w7(32'hbbae9370),
	.w8(32'hbba10583),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb748dbd),
	.w1(32'hbb97571f),
	.w2(32'hbc845c8d),
	.w3(32'hbb2ba677),
	.w4(32'h3b036bb5),
	.w5(32'hbc232aa9),
	.w6(32'h3b60b1fa),
	.w7(32'hbc360546),
	.w8(32'h3aced435),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c9b3),
	.w1(32'hbb5fc2b3),
	.w2(32'hba47f2bd),
	.w3(32'h3b756c89),
	.w4(32'hbbada4c0),
	.w5(32'h3ac2451f),
	.w6(32'hbb9dac7d),
	.w7(32'h3ab67216),
	.w8(32'h3bd90e2b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3f19f),
	.w1(32'h3b43f081),
	.w2(32'h3a42ecaf),
	.w3(32'h3bf5d4ae),
	.w4(32'h3b67dfeb),
	.w5(32'h3a3ded36),
	.w6(32'h3b90ea99),
	.w7(32'h3ab11779),
	.w8(32'h3b2a90ec),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af80a66),
	.w1(32'hbbdc9449),
	.w2(32'hbc09407b),
	.w3(32'h3ab16e0e),
	.w4(32'hbbce1ec0),
	.w5(32'hbbcc50c3),
	.w6(32'hbc06951a),
	.w7(32'hbbb96ecc),
	.w8(32'hbb8496aa),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8105c2),
	.w1(32'hba296050),
	.w2(32'hbba717f1),
	.w3(32'hbaca518c),
	.w4(32'h3b60c8c5),
	.w5(32'h3b98c1aa),
	.w6(32'h3a867ac4),
	.w7(32'h399ca4a6),
	.w8(32'h3996f470),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fe5b6),
	.w1(32'h3bc68291),
	.w2(32'h3be5d1c6),
	.w3(32'h39d10902),
	.w4(32'h3b66931c),
	.w5(32'h3a44c79e),
	.w6(32'h3a39dbbe),
	.w7(32'h3b353f47),
	.w8(32'h398487b7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfeb96f),
	.w1(32'h3afc43a4),
	.w2(32'hbb0c6729),
	.w3(32'h3b543404),
	.w4(32'hbbee106a),
	.w5(32'hbb934883),
	.w6(32'hbb761c3e),
	.w7(32'h3b37f0ed),
	.w8(32'hbba17a8e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b5d64),
	.w1(32'h3ba8e0d4),
	.w2(32'h3abd2afe),
	.w3(32'hbbebcdc9),
	.w4(32'h3af24257),
	.w5(32'h3b81b6a5),
	.w6(32'h3b3b8c6d),
	.w7(32'h3b97e6cb),
	.w8(32'hb89836d5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d1beb),
	.w1(32'h3a852600),
	.w2(32'hba9f0695),
	.w3(32'h3ac8b9ae),
	.w4(32'hbb61d1d0),
	.w5(32'hbb04fdf9),
	.w6(32'hbafbf9bf),
	.w7(32'h3ac2d15b),
	.w8(32'hbb24dacf),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6b286),
	.w1(32'hbb4c88e6),
	.w2(32'hbbcf58cc),
	.w3(32'hbb6758d0),
	.w4(32'hbb0361c9),
	.w5(32'hbac49237),
	.w6(32'hbaaeca33),
	.w7(32'hba8972a6),
	.w8(32'hb9bdf004),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393db439),
	.w1(32'h3aafbf13),
	.w2(32'h3b0ac25d),
	.w3(32'h3a824d33),
	.w4(32'hba272a0d),
	.w5(32'hbacde587),
	.w6(32'h3a6a7105),
	.w7(32'h3ae7501a),
	.w8(32'h3b2a7f37),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5fa64),
	.w1(32'h3b0b8ced),
	.w2(32'h3b13f726),
	.w3(32'hba60be24),
	.w4(32'h3b373c55),
	.w5(32'h3b87b4ff),
	.w6(32'h3accf2b7),
	.w7(32'h3b6e81f0),
	.w8(32'h3b7671a6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba55316),
	.w1(32'h3a90d6fb),
	.w2(32'hba8c336a),
	.w3(32'h3bbea583),
	.w4(32'hbb6f0d86),
	.w5(32'hbb1209f9),
	.w6(32'hbb0010e8),
	.w7(32'h3ac78b14),
	.w8(32'hbb220050),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae08d8d),
	.w1(32'h3962e449),
	.w2(32'h3a8b65fb),
	.w3(32'hbb697e6a),
	.w4(32'h3a25440c),
	.w5(32'hb9f0ecdb),
	.w6(32'hbab1fb05),
	.w7(32'hbb22dbc0),
	.w8(32'hbba27864),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb416b),
	.w1(32'h3b6266e2),
	.w2(32'hbac76c24),
	.w3(32'hbb937b74),
	.w4(32'h3aab8524),
	.w5(32'h3b42d056),
	.w6(32'h3aeb992a),
	.w7(32'h3b2cbe48),
	.w8(32'h38e19419),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39437dd9),
	.w1(32'h3b3436a2),
	.w2(32'hbc82fd11),
	.w3(32'h3acfcfbf),
	.w4(32'h3bf86817),
	.w5(32'hbbbfb2a8),
	.w6(32'hbb467e8c),
	.w7(32'hbc2a23e5),
	.w8(32'hbc4a745f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc05a7),
	.w1(32'h3b4c1004),
	.w2(32'hb9d39177),
	.w3(32'hbbee281b),
	.w4(32'h3ac5d666),
	.w5(32'h3b85415a),
	.w6(32'h3a93c538),
	.w7(32'h3b20256a),
	.w8(32'h38ad8d35),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a291be6),
	.w1(32'hb95e974e),
	.w2(32'h3a1ac0a2),
	.w3(32'h3b290112),
	.w4(32'h3aac0725),
	.w5(32'hba876db0),
	.w6(32'h3a9cde23),
	.w7(32'hb999d55e),
	.w8(32'h39cbc0d7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad56b33),
	.w1(32'h3b52859b),
	.w2(32'hbbbb10d9),
	.w3(32'hbb5af264),
	.w4(32'h3bdc9df1),
	.w5(32'h3b1140c9),
	.w6(32'h3ba0f165),
	.w7(32'h3ba7d450),
	.w8(32'h3c0d6e00),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea17aa),
	.w1(32'h3ab8da0a),
	.w2(32'hbae46f49),
	.w3(32'h3c2404a0),
	.w4(32'hbbb17ab3),
	.w5(32'hbb5bebfd),
	.w6(32'hbb3f9c9c),
	.w7(32'h3b072432),
	.w8(32'hbb734d34),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34c7be),
	.w1(32'h3b7bd374),
	.w2(32'hb961eb34),
	.w3(32'hbbb1557a),
	.w4(32'h3ac41bd7),
	.w5(32'h3aa64bd4),
	.w6(32'h3ae4a7ff),
	.w7(32'h3b7b1d80),
	.w8(32'h3ab2ba52),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76d432),
	.w1(32'h3b69d0d5),
	.w2(32'h3991a51f),
	.w3(32'h3a362dcd),
	.w4(32'h3a6ca838),
	.w5(32'h3a8dc48d),
	.w6(32'h3a9df8c4),
	.w7(32'h3b9053a2),
	.w8(32'h3a7c8218),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f30cd9),
	.w1(32'h3aaad38b),
	.w2(32'h3a7b7756),
	.w3(32'h38b6f38e),
	.w4(32'h38a65900),
	.w5(32'hbb9180f5),
	.w6(32'h3ae7719a),
	.w7(32'h3b72f3ac),
	.w8(32'h3b9e2862),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce7903),
	.w1(32'hbb10a9e2),
	.w2(32'hbaad71dd),
	.w3(32'hba18e8ed),
	.w4(32'hbb4f3986),
	.w5(32'hba8e99d6),
	.w6(32'hbb0378e8),
	.w7(32'hbad85b6a),
	.w8(32'hbad4eb01),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9df6d),
	.w1(32'hbb70dacb),
	.w2(32'hbb9ef474),
	.w3(32'hba0da859),
	.w4(32'hbb5aa809),
	.w5(32'hbaaa5320),
	.w6(32'hbb4cc0d0),
	.w7(32'hbaa3070d),
	.w8(32'hbb48d335),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bfda2),
	.w1(32'h3a8b2e1c),
	.w2(32'hba4aabed),
	.w3(32'hbb208875),
	.w4(32'h3b157b1e),
	.w5(32'h3a5bac6e),
	.w6(32'h3a9dfd0c),
	.w7(32'h3b9c66fd),
	.w8(32'h3a330e50),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefb071),
	.w1(32'h3be9c1e3),
	.w2(32'h3acf9653),
	.w3(32'h3b27e6ac),
	.w4(32'h3b4665d0),
	.w5(32'h3b40c0f4),
	.w6(32'h3b8e5f03),
	.w7(32'h3bc22fe7),
	.w8(32'h3ad6d5cc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb7cfd),
	.w1(32'hbbc977de),
	.w2(32'hbb3d10ac),
	.w3(32'h3ab53169),
	.w4(32'hbab16586),
	.w5(32'hbb2eb2c3),
	.w6(32'hbc36546a),
	.w7(32'hbc2d9051),
	.w8(32'hbb65a881),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af68f41),
	.w1(32'hbb91a04f),
	.w2(32'hbc2bdd91),
	.w3(32'hb9b2de31),
	.w4(32'hbbd00104),
	.w5(32'hbbf60f18),
	.w6(32'hbbcd9f05),
	.w7(32'hbb4a0a50),
	.w8(32'hbbb93f38),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e74d9),
	.w1(32'hbba9e60d),
	.w2(32'hbb80a9b0),
	.w3(32'hbbbb888b),
	.w4(32'hbb926223),
	.w5(32'hba03d47c),
	.w6(32'hbbaf204c),
	.w7(32'hba2424a7),
	.w8(32'hbae8c976),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f23e0b),
	.w1(32'hb96d7502),
	.w2(32'hba6fa054),
	.w3(32'h3a82cdfe),
	.w4(32'hba23dba1),
	.w5(32'hba77f774),
	.w6(32'hb879e726),
	.w7(32'hba0a4cc6),
	.w8(32'hb8df2d72),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a93ea5),
	.w1(32'h3a86705a),
	.w2(32'h39c4d9c7),
	.w3(32'hb9841b96),
	.w4(32'h3a873541),
	.w5(32'h3a216fdc),
	.w6(32'h3a9e1eff),
	.w7(32'h3a6584e0),
	.w8(32'h3a5eb18b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule