module layer_10_featuremap_251(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb332),
	.w1(32'hbc0ce1d8),
	.w2(32'hbb00d70a),
	.w3(32'hbbc372b3),
	.w4(32'hba827ad5),
	.w5(32'hbbbca4bf),
	.w6(32'hbc6b8dfd),
	.w7(32'hbb1e9079),
	.w8(32'hbb5083ff),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93e167),
	.w1(32'h389a98c8),
	.w2(32'h3b20976a),
	.w3(32'hbbc0c26e),
	.w4(32'hbb212020),
	.w5(32'hbab68742),
	.w6(32'h3c052388),
	.w7(32'hbb1f450e),
	.w8(32'hba109479),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a50f8f),
	.w1(32'h3c93a6cd),
	.w2(32'h3c0275e6),
	.w3(32'h3c157473),
	.w4(32'hbb079535),
	.w5(32'hbb75e9c3),
	.w6(32'hbc2244f1),
	.w7(32'hbba7f414),
	.w8(32'hba779961),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0b8f1),
	.w1(32'h3b05d924),
	.w2(32'h397e5aef),
	.w3(32'hbba2faf7),
	.w4(32'hbba44422),
	.w5(32'h3b01e1b7),
	.w6(32'h3bcb1666),
	.w7(32'h39d4ac82),
	.w8(32'h3a6f6e6e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d05628),
	.w1(32'hbc8a33c4),
	.w2(32'hbb1c2f16),
	.w3(32'hbb5379fe),
	.w4(32'h3b0e7040),
	.w5(32'hbb3bd530),
	.w6(32'hbc1eb8a1),
	.w7(32'hbacba278),
	.w8(32'hbbaccffe),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91346a),
	.w1(32'h3a795cec),
	.w2(32'hba3f8f2a),
	.w3(32'hbb859234),
	.w4(32'hbb932eab),
	.w5(32'hbc0c9b10),
	.w6(32'h3b06f1e1),
	.w7(32'h3a99b5ce),
	.w8(32'hbbecc7bc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf02ba3),
	.w1(32'hbbb8cb2b),
	.w2(32'hbbfba536),
	.w3(32'hbc1d3aa2),
	.w4(32'hbbde79d0),
	.w5(32'hbb075cbc),
	.w6(32'h3b9fb20a),
	.w7(32'hbb732555),
	.w8(32'hbb315081),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb671a54),
	.w1(32'hbb8d0215),
	.w2(32'hbae0b3a7),
	.w3(32'hbbecd306),
	.w4(32'hbb57d2f3),
	.w5(32'hbae94b5c),
	.w6(32'hbb847439),
	.w7(32'hb9fc6146),
	.w8(32'hbb8bc7c1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25ce18),
	.w1(32'hbaaa1339),
	.w2(32'hba413e02),
	.w3(32'hbb38118c),
	.w4(32'hb993eab9),
	.w5(32'hbaf13be8),
	.w6(32'hbba19890),
	.w7(32'hbb95c911),
	.w8(32'hbb22f753),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0520e),
	.w1(32'hbad228b7),
	.w2(32'hba0edd3a),
	.w3(32'hbbc56d81),
	.w4(32'hbba3da8c),
	.w5(32'hbb3a2039),
	.w6(32'h3a9e085c),
	.w7(32'hbab56997),
	.w8(32'hbb2e38eb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d47803),
	.w1(32'h3b133e2a),
	.w2(32'hbac20483),
	.w3(32'hbb27c1c2),
	.w4(32'hbb42d3ce),
	.w5(32'hbae3fefd),
	.w6(32'h3c1f6e51),
	.w7(32'h3a74e91e),
	.w8(32'hbbb259ce),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e8ec5),
	.w1(32'h3cd45edd),
	.w2(32'h3cb3977c),
	.w3(32'h3baebe07),
	.w4(32'h390487ac),
	.w5(32'hbbf5c8ff),
	.w6(32'hbc387012),
	.w7(32'h3ba6450f),
	.w8(32'hba95fda9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39f927),
	.w1(32'hbc5ca25a),
	.w2(32'hbc32b927),
	.w3(32'hbc56f32d),
	.w4(32'hbbc2fc0e),
	.w5(32'hbb9a7056),
	.w6(32'hba92a978),
	.w7(32'hbbaa9bd3),
	.w8(32'hbb8b3302),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfa066),
	.w1(32'hb9658226),
	.w2(32'hbb5f4207),
	.w3(32'hba8c8e58),
	.w4(32'hbac4db79),
	.w5(32'hbb01bb31),
	.w6(32'h37e07ebe),
	.w7(32'hbbaf2477),
	.w8(32'h3a94c83a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d80cd),
	.w1(32'hbb27ae5f),
	.w2(32'hb99d01cc),
	.w3(32'hbadd3333),
	.w4(32'hb9265c22),
	.w5(32'hbba4fb7b),
	.w6(32'h3c4d8ea0),
	.w7(32'h39e76407),
	.w8(32'hbc38288d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e46b8),
	.w1(32'hbc53b215),
	.w2(32'hbb3549a6),
	.w3(32'hbc1e505c),
	.w4(32'h3746d66f),
	.w5(32'hbb863ce7),
	.w6(32'hbbc0f1ce),
	.w7(32'hb9ee4a81),
	.w8(32'hbbf754bf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba147e7),
	.w1(32'h3ba61981),
	.w2(32'h3b74b18f),
	.w3(32'hbbbdcc12),
	.w4(32'hbae4a9e0),
	.w5(32'hbba7cfdf),
	.w6(32'hb8b87dff),
	.w7(32'h3a414eb2),
	.w8(32'h3a51fe3a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb867334),
	.w1(32'hbbdb8a9a),
	.w2(32'hbc12febe),
	.w3(32'hbb04934f),
	.w4(32'hbb24bdaa),
	.w5(32'hba09f5b4),
	.w6(32'hba7ef1f9),
	.w7(32'hbb59acc9),
	.w8(32'h3c9ae3af),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cb210),
	.w1(32'h39706afa),
	.w2(32'h3b374c08),
	.w3(32'hbb19d2c3),
	.w4(32'h3bb7d948),
	.w5(32'hba482d6e),
	.w6(32'h3cfad8fd),
	.w7(32'h3caed476),
	.w8(32'hbc0137b2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9f414),
	.w1(32'hba45ed3b),
	.w2(32'hbbc6d7e1),
	.w3(32'hba5583c5),
	.w4(32'h3adcd4e0),
	.w5(32'hbb99e45b),
	.w6(32'h3b7d0ec3),
	.w7(32'hbb10cefe),
	.w8(32'hbbbb16f5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc518c4),
	.w1(32'hbc0718ff),
	.w2(32'hbae9ce3d),
	.w3(32'hbb828244),
	.w4(32'hbbac2aac),
	.w5(32'h39911321),
	.w6(32'hbc2ede00),
	.w7(32'hbab9503d),
	.w8(32'hbb6e6418),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07e500),
	.w1(32'hbb9bd198),
	.w2(32'hba037997),
	.w3(32'h3ba4e0e6),
	.w4(32'h3b16e9f3),
	.w5(32'hba983917),
	.w6(32'hbba93f38),
	.w7(32'hba3c8df3),
	.w8(32'h39b8c088),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89277e),
	.w1(32'h3a357ae1),
	.w2(32'h3ab387cc),
	.w3(32'h3b31723e),
	.w4(32'hbb4994e3),
	.w5(32'hbb8afc7b),
	.w6(32'hbb020f7f),
	.w7(32'hbadefa5f),
	.w8(32'hbbe43bed),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1cb6),
	.w1(32'hbc6b8a3c),
	.w2(32'hbbed6720),
	.w3(32'hbbba80ce),
	.w4(32'h3ba0b916),
	.w5(32'h3a79f69c),
	.w6(32'h3b3ddac8),
	.w7(32'hbbb64e0c),
	.w8(32'h3b0b4d02),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2024e7),
	.w1(32'h3c0965c8),
	.w2(32'h3b66f8ad),
	.w3(32'h3bb88883),
	.w4(32'hbb53bfc3),
	.w5(32'hbb1a47a6),
	.w6(32'h38adbe41),
	.w7(32'hbada4fba),
	.w8(32'hbb2e1288),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89566e),
	.w1(32'hbab77466),
	.w2(32'h382a59a6),
	.w3(32'hbbd1ebbe),
	.w4(32'h3a4a370a),
	.w5(32'hbb34d958),
	.w6(32'h3c0f0e32),
	.w7(32'h39ab1cd2),
	.w8(32'h3baee452),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aea3c),
	.w1(32'hb7aa8449),
	.w2(32'h3b005886),
	.w3(32'hba9882b3),
	.w4(32'hbb8b2ed4),
	.w5(32'h3ac2bb04),
	.w6(32'h3c7d6869),
	.w7(32'h3b85d76a),
	.w8(32'h39259df4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fddfe),
	.w1(32'hbbd21460),
	.w2(32'hbaed4fbd),
	.w3(32'hbb2859b6),
	.w4(32'hbab6103b),
	.w5(32'hbc06a568),
	.w6(32'hbc10dd5c),
	.w7(32'hbac9c131),
	.w8(32'hbb0a8c74),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b250ff0),
	.w1(32'hbb0d5a17),
	.w2(32'hbc32e06c),
	.w3(32'hbb898b5b),
	.w4(32'hbb22215c),
	.w5(32'h3b2fc0d4),
	.w6(32'hbb02a014),
	.w7(32'hbac95e70),
	.w8(32'hbb70d321),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07b9a8),
	.w1(32'hbc0210ab),
	.w2(32'h39959944),
	.w3(32'hbb886d1e),
	.w4(32'hbb13ca0e),
	.w5(32'h3b7904f9),
	.w6(32'hbbda8b35),
	.w7(32'hbb3c0f10),
	.w8(32'hbc021ebb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ab57d),
	.w1(32'h39f7430c),
	.w2(32'h3a10219d),
	.w3(32'hbc16b36f),
	.w4(32'h3b295606),
	.w5(32'hbb56bdf5),
	.w6(32'h3c5b13c4),
	.w7(32'hbc070a1e),
	.w8(32'hbb54c097),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac19c),
	.w1(32'h3c6f67bf),
	.w2(32'hbc2d24cc),
	.w3(32'h3a1ce4d6),
	.w4(32'h3c040e57),
	.w5(32'hbbbb96ad),
	.w6(32'hbca4b8d4),
	.w7(32'hbb81888e),
	.w8(32'hbae33050),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe59e2),
	.w1(32'hbb04232c),
	.w2(32'h3b81959b),
	.w3(32'hbc91974e),
	.w4(32'h3bfb0e59),
	.w5(32'hbae5be96),
	.w6(32'h3bccd789),
	.w7(32'hbb872a90),
	.w8(32'hbbb4e320),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb219f),
	.w1(32'h3b824f08),
	.w2(32'hbc0d4274),
	.w3(32'h39a4985b),
	.w4(32'hb89ddf8a),
	.w5(32'h3ad50ece),
	.w6(32'h3a324541),
	.w7(32'hbbd9f283),
	.w8(32'hbb1d64d1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32e9df),
	.w1(32'h3b63945a),
	.w2(32'hbb5ebac4),
	.w3(32'h3b3c0d1e),
	.w4(32'hbac49744),
	.w5(32'h3bfcb33e),
	.w6(32'hba0664ba),
	.w7(32'hbb92ab9d),
	.w8(32'h3c003965),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a17c7),
	.w1(32'h3c925b46),
	.w2(32'h3b8ecde2),
	.w3(32'h3bef4b98),
	.w4(32'hbb2cccf2),
	.w5(32'h3b5876bf),
	.w6(32'h3ab97f68),
	.w7(32'h39f1bf6f),
	.w8(32'hbabae6d9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a8a35),
	.w1(32'h3a9eb5bf),
	.w2(32'h3ba83399),
	.w3(32'hbbae55b4),
	.w4(32'h3abf2c71),
	.w5(32'h3a3bc1c4),
	.w6(32'hbbe73035),
	.w7(32'hbb5c0bef),
	.w8(32'h398c66a5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18df20),
	.w1(32'h3b822658),
	.w2(32'h3c0e836e),
	.w3(32'hbb3035bd),
	.w4(32'hbbc38cbf),
	.w5(32'h3a1772c4),
	.w6(32'h3c160a6a),
	.w7(32'h3c2f56b2),
	.w8(32'hbac12293),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4343c9),
	.w1(32'hbc2d14f0),
	.w2(32'hbadac033),
	.w3(32'hbb6dacb5),
	.w4(32'hbb6cce99),
	.w5(32'hbba30058),
	.w6(32'h3c041ad5),
	.w7(32'h3c166c59),
	.w8(32'hbbfd0a9d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b7a7c),
	.w1(32'hbc8d4511),
	.w2(32'hbb40b320),
	.w3(32'hba80e66d),
	.w4(32'hbc7926ab),
	.w5(32'hbb460ccf),
	.w6(32'hbc970f0d),
	.w7(32'hbc180bee),
	.w8(32'h3b2cc340),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba85eef),
	.w1(32'hba9bb576),
	.w2(32'hbb208385),
	.w3(32'hbb1bc46d),
	.w4(32'hbafdfbd4),
	.w5(32'hba9ec8a4),
	.w6(32'h39f205c6),
	.w7(32'hbb87f594),
	.w8(32'hbc010442),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb683da7),
	.w1(32'hb9f3c4f3),
	.w2(32'h3b564168),
	.w3(32'hbb3e2ca5),
	.w4(32'hbb30c139),
	.w5(32'hbb8d50cc),
	.w6(32'h3adf9e15),
	.w7(32'hbbd68df8),
	.w8(32'h3c2dee42),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61d551),
	.w1(32'hbb8cf777),
	.w2(32'h3c24c62b),
	.w3(32'h3a8a6560),
	.w4(32'hba0f166a),
	.w5(32'hbab0da8c),
	.w6(32'h3c0e2291),
	.w7(32'h3c427bf7),
	.w8(32'hbb1a2f22),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6dcc3),
	.w1(32'h3ca089e5),
	.w2(32'h3b250176),
	.w3(32'hbc23c215),
	.w4(32'h3b6b2864),
	.w5(32'hbb8c5b4f),
	.w6(32'h3d10fc52),
	.w7(32'h3abb68e1),
	.w8(32'h3b4c58f2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2f18d),
	.w1(32'hbaa144e2),
	.w2(32'h3b5b1b25),
	.w3(32'hbb58f6b0),
	.w4(32'hbb51f989),
	.w5(32'h3accc47d),
	.w6(32'hb9b47884),
	.w7(32'h3ba2b95d),
	.w8(32'hbc38e3ea),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd78806),
	.w1(32'hbbeeadde),
	.w2(32'hbc476c16),
	.w3(32'hbbe07c99),
	.w4(32'hbb3a62e2),
	.w5(32'hb9946630),
	.w6(32'hbbe3d89b),
	.w7(32'hbc6dd80a),
	.w8(32'hbb08ed45),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb921592),
	.w1(32'hba712030),
	.w2(32'hbb4d5cc2),
	.w3(32'hbad39f61),
	.w4(32'hbbb78ffd),
	.w5(32'h3b9d321e),
	.w6(32'hbae09d9a),
	.w7(32'hbbd7dbe0),
	.w8(32'h3b15b7fe),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d3e66),
	.w1(32'h3b60d562),
	.w2(32'h3baf7725),
	.w3(32'h3be6aa63),
	.w4(32'h3c381a91),
	.w5(32'h3b8ec388),
	.w6(32'h3a3ee745),
	.w7(32'h3b7fc991),
	.w8(32'h3c19c249),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb9fcd),
	.w1(32'h3c266280),
	.w2(32'h3bc97079),
	.w3(32'h3ae0decf),
	.w4(32'h3bd59576),
	.w5(32'h3a10cca6),
	.w6(32'h3c6b39eb),
	.w7(32'h3c17d21b),
	.w8(32'hbbf69657),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f7be4),
	.w1(32'hbb39a477),
	.w2(32'hbae7c8f3),
	.w3(32'h3b0e5b7e),
	.w4(32'hb95c4058),
	.w5(32'h3c082376),
	.w6(32'hbb837aad),
	.w7(32'hbb81f510),
	.w8(32'h3b1db204),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c091e6e),
	.w1(32'h3cb57749),
	.w2(32'hbb45ca44),
	.w3(32'h39d838b1),
	.w4(32'hbbd411ce),
	.w5(32'hbbb34446),
	.w6(32'h3c7372fe),
	.w7(32'h3ba5d225),
	.w8(32'h3c68491b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb7746),
	.w1(32'h3c167f3a),
	.w2(32'hbb8979e8),
	.w3(32'hbb9b4504),
	.w4(32'h3b8380b0),
	.w5(32'h3b18ccdb),
	.w6(32'h3cb357e8),
	.w7(32'h3b9d3d5f),
	.w8(32'h3bc4671f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2049d9),
	.w1(32'hbb2d29df),
	.w2(32'hbb54070e),
	.w3(32'h3c0ee07e),
	.w4(32'h3b9af89a),
	.w5(32'h3bdcc7d9),
	.w6(32'h3b6d2275),
	.w7(32'hbb39c74b),
	.w8(32'h3aa43181),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f78f2),
	.w1(32'hbbeac47e),
	.w2(32'h3acc4fd2),
	.w3(32'hbb2d4362),
	.w4(32'hba739622),
	.w5(32'hba41cc13),
	.w6(32'hbbdab44c),
	.w7(32'hbc5bd6a8),
	.w8(32'hbc1f0c94),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb588220),
	.w1(32'hbb47d277),
	.w2(32'hbb880c9e),
	.w3(32'h3b0b5fa8),
	.w4(32'h3b1a02a0),
	.w5(32'hbbf8026d),
	.w6(32'hbb2267fa),
	.w7(32'hbaf4d3e0),
	.w8(32'hbbad9f66),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9326e0),
	.w1(32'hbb14170d),
	.w2(32'hbc05e3f9),
	.w3(32'h3b3e0986),
	.w4(32'h3bd6b0b0),
	.w5(32'hbb6fa10b),
	.w6(32'h3b2900a0),
	.w7(32'hba8cf496),
	.w8(32'hbbd2ce5f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd461b0),
	.w1(32'hba31db2b),
	.w2(32'h3af1cf16),
	.w3(32'hba874cdb),
	.w4(32'h3b249701),
	.w5(32'h3b504cbe),
	.w6(32'hbbe11f15),
	.w7(32'hbae1d157),
	.w8(32'hb94cfd6d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b030691),
	.w1(32'hbbaede6d),
	.w2(32'h3b2d41b6),
	.w3(32'hbbc34e16),
	.w4(32'h3be359d2),
	.w5(32'hbb11022d),
	.w6(32'hbc275565),
	.w7(32'h3a53fc55),
	.w8(32'hbc1c794f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb201e3e),
	.w1(32'hbacc73dd),
	.w2(32'hba3e0d29),
	.w3(32'h3b3a857e),
	.w4(32'h3a5fd5ae),
	.w5(32'h3b6dd919),
	.w6(32'hbbcae097),
	.w7(32'hbbef2b7b),
	.w8(32'h3bee4638),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be56e0e),
	.w1(32'h3b21aec5),
	.w2(32'h3c4d39cd),
	.w3(32'h3c8389c1),
	.w4(32'h3c522198),
	.w5(32'hbae25ac7),
	.w6(32'hbbfe6842),
	.w7(32'h3c26f489),
	.w8(32'h3b382aa0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe548e3),
	.w1(32'hbc024a0c),
	.w2(32'hbc12f1ee),
	.w3(32'hbbd4ee40),
	.w4(32'hbb7bad21),
	.w5(32'hbc229a01),
	.w6(32'h3c48f968),
	.w7(32'h3afc3490),
	.w8(32'hbb8aa08d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd341a),
	.w1(32'hb9225499),
	.w2(32'hbbfa8b85),
	.w3(32'hbc8adb22),
	.w4(32'hbc09bc2f),
	.w5(32'h3b4a7f74),
	.w6(32'h3bf5067e),
	.w7(32'hbbc09d94),
	.w8(32'h3bd2c8dc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c98ad),
	.w1(32'hbb9433de),
	.w2(32'hba7a96aa),
	.w3(32'h3aaae06e),
	.w4(32'h3aae01e2),
	.w5(32'hba837199),
	.w6(32'h3c0760da),
	.w7(32'h3b734efa),
	.w8(32'hb9cf20f2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79b7e9),
	.w1(32'h3bbac660),
	.w2(32'hbac89994),
	.w3(32'hb92a7e4a),
	.w4(32'hbb08a8e0),
	.w5(32'hb9fcb4be),
	.w6(32'h3b255a88),
	.w7(32'hbb9049f7),
	.w8(32'hbbaecb36),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e2a06),
	.w1(32'hbaa9da63),
	.w2(32'hbc303762),
	.w3(32'hbb33698c),
	.w4(32'h3aa8074e),
	.w5(32'h3a4ae45d),
	.w6(32'h3bda3baa),
	.w7(32'hbbf7d70d),
	.w8(32'h3abdf2ed),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0183e4),
	.w1(32'hbc06e13d),
	.w2(32'hbc0a9ab9),
	.w3(32'h3bdfb142),
	.w4(32'hbb086836),
	.w5(32'hbb478583),
	.w6(32'h3ab333d1),
	.w7(32'h3b1c1647),
	.w8(32'h3b769af9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23e2cb),
	.w1(32'h3a84bdc4),
	.w2(32'hbb4b4aa5),
	.w3(32'hbbc10549),
	.w4(32'hbbef7e4a),
	.w5(32'hbb956136),
	.w6(32'h3bc20f75),
	.w7(32'hba643998),
	.w8(32'hbba42daa),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9451fa),
	.w1(32'h3c843ed2),
	.w2(32'h3b3de94e),
	.w3(32'hbbbceaba),
	.w4(32'hbb814187),
	.w5(32'h3a530b96),
	.w6(32'h3ca5a1b0),
	.w7(32'hbb0bb3af),
	.w8(32'h3b1a5451),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb967061),
	.w1(32'hbb9c4e2f),
	.w2(32'h3a229061),
	.w3(32'hbb4f62d2),
	.w4(32'h3ae4017b),
	.w5(32'h3c68f92e),
	.w6(32'h3b16be13),
	.w7(32'h3ba99e34),
	.w8(32'h3b997985),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5876e1),
	.w1(32'h3c5bb863),
	.w2(32'h3bbb127b),
	.w3(32'h3bede9f5),
	.w4(32'h3bf49fab),
	.w5(32'hbb68e5bf),
	.w6(32'h3c98b1d3),
	.w7(32'h3baf1884),
	.w8(32'h3c3f32c1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf061c6),
	.w1(32'h3b8b616e),
	.w2(32'h3c446dbd),
	.w3(32'h3ab356fc),
	.w4(32'hb903685f),
	.w5(32'hbb68588a),
	.w6(32'h3ca34302),
	.w7(32'h3c787448),
	.w8(32'hbc1b29e1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb261142),
	.w1(32'hbb0d54b6),
	.w2(32'hbba8dddc),
	.w3(32'hbad61c7d),
	.w4(32'hbbb2fd19),
	.w5(32'hb80926d5),
	.w6(32'hbbcb64a9),
	.w7(32'h3c194e00),
	.w8(32'h3b92ac8e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a80a2),
	.w1(32'h3c209365),
	.w2(32'h3b1c67f9),
	.w3(32'hbb261752),
	.w4(32'h3b4b0c37),
	.w5(32'hbb2c5085),
	.w6(32'h3be426ca),
	.w7(32'h3c84ab58),
	.w8(32'hbac546e1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b68d8a),
	.w1(32'h3a11e83e),
	.w2(32'hbb31a12d),
	.w3(32'hbbde21e5),
	.w4(32'hbb1aba30),
	.w5(32'hba9bc386),
	.w6(32'hbb3a883b),
	.w7(32'hbb8f73a7),
	.w8(32'hbaf743da),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b12b6),
	.w1(32'h3c1527d3),
	.w2(32'h3b9f4de6),
	.w3(32'hbbfc8bee),
	.w4(32'hbb821651),
	.w5(32'hbbf48f3b),
	.w6(32'h3a0a55fa),
	.w7(32'hbb28e30b),
	.w8(32'h3b0b533a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba224d97),
	.w1(32'hb98b94a5),
	.w2(32'h3b922fee),
	.w3(32'hbaf4fca3),
	.w4(32'h3b90cc4a),
	.w5(32'hbb27c2fe),
	.w6(32'hbb666192),
	.w7(32'h3ba87f4d),
	.w8(32'h3ba5983d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51bfd4),
	.w1(32'hbb3f29b9),
	.w2(32'hba4a06ce),
	.w3(32'h3b381c4d),
	.w4(32'hbb570395),
	.w5(32'hbb32e1dd),
	.w6(32'h3b9f10b0),
	.w7(32'h3af68f15),
	.w8(32'hbb10dfe3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2af68),
	.w1(32'h3c0b950b),
	.w2(32'h3a92c086),
	.w3(32'hbb506541),
	.w4(32'hba1fd8d8),
	.w5(32'hbc3f8deb),
	.w6(32'h3b811417),
	.w7(32'hbb292946),
	.w8(32'h3afe5a56),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f2cb),
	.w1(32'hbaf488f0),
	.w2(32'hbb865688),
	.w3(32'hbbcb6f96),
	.w4(32'hbbb55e0a),
	.w5(32'hbc0da165),
	.w6(32'h3b545eaf),
	.w7(32'h3b9b0aa0),
	.w8(32'hbc0a65d8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb01b57),
	.w1(32'hb974b7f8),
	.w2(32'hbb7f3093),
	.w3(32'hbc4a0889),
	.w4(32'hbc0d8518),
	.w5(32'hbb8235bd),
	.w6(32'h3b4dd177),
	.w7(32'hbbe8dbcf),
	.w8(32'h3a5ce69a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb873ef12),
	.w1(32'hbb7921a1),
	.w2(32'h3c1c9f29),
	.w3(32'h3b6dc60a),
	.w4(32'hb9ea143f),
	.w5(32'h3a8a517b),
	.w6(32'hbc0b6aa4),
	.w7(32'h39a0a2c1),
	.w8(32'h3be69c06),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62b210),
	.w1(32'h3a9ef7fb),
	.w2(32'h3b1c4d44),
	.w3(32'h3b5ff71c),
	.w4(32'h3b9f6b85),
	.w5(32'hbb6fd21d),
	.w6(32'hbbd3027a),
	.w7(32'h3bc07fe3),
	.w8(32'h3b04a39b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1f385),
	.w1(32'hbbfdcb74),
	.w2(32'hbb883800),
	.w3(32'h3b08e969),
	.w4(32'hbbca90cc),
	.w5(32'hbab0306e),
	.w6(32'h3b2e80fa),
	.w7(32'h3a9b78c2),
	.w8(32'h3b7be41c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cfeaa),
	.w1(32'h3c061470),
	.w2(32'h3b39d321),
	.w3(32'h3b1e74ba),
	.w4(32'hbb84c4e5),
	.w5(32'hbb5a9b11),
	.w6(32'h3c905864),
	.w7(32'h3bb9a3ed),
	.w8(32'h3b61d418),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe97f4e),
	.w1(32'hbbb5bc84),
	.w2(32'hba92c597),
	.w3(32'h3b0c0295),
	.w4(32'h3aeb994f),
	.w5(32'hbb909311),
	.w6(32'h3b867650),
	.w7(32'h3a623196),
	.w8(32'hbb6117ee),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d8936),
	.w1(32'h3bc5b7c2),
	.w2(32'hbb9e228b),
	.w3(32'hbbed85c8),
	.w4(32'hbc03fc5a),
	.w5(32'hba519154),
	.w6(32'h3c535202),
	.w7(32'h3be586cc),
	.w8(32'hbbaf9d12),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb471a4e),
	.w1(32'h3aafe833),
	.w2(32'h3bb2f3bf),
	.w3(32'hba4a9262),
	.w4(32'hbbbfb5fc),
	.w5(32'hb9962aa2),
	.w6(32'hbbe762f9),
	.w7(32'hbb2229c6),
	.w8(32'hb97a2474),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a494f2e),
	.w1(32'h3b490e13),
	.w2(32'h3baa8e54),
	.w3(32'hba533e50),
	.w4(32'h3b6b86e0),
	.w5(32'hbb9ea2f1),
	.w6(32'hbaa91fd3),
	.w7(32'h3b7d819e),
	.w8(32'hbc0f118a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc130594),
	.w1(32'hbb976516),
	.w2(32'hbb9d31ed),
	.w3(32'hbc0d9537),
	.w4(32'hbbe9b27c),
	.w5(32'hbab71f9d),
	.w6(32'hbace398f),
	.w7(32'hbc131ec2),
	.w8(32'hbbe0367c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec7179),
	.w1(32'hbc02e733),
	.w2(32'hbbe2020b),
	.w3(32'hbaccf187),
	.w4(32'hbb3f690a),
	.w5(32'h3a0cff55),
	.w6(32'hbbd57f9c),
	.w7(32'hbbafba7c),
	.w8(32'hbc1d17f1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae1065),
	.w1(32'hbb54d89f),
	.w2(32'hbbcf62e2),
	.w3(32'h3a88067a),
	.w4(32'h3ad60f44),
	.w5(32'hbba52292),
	.w6(32'hbbc8f8dc),
	.w7(32'hbbc9f158),
	.w8(32'hba89deba),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22d68a),
	.w1(32'hbbc8a39e),
	.w2(32'hbb496315),
	.w3(32'hbbb9f9ac),
	.w4(32'hbaf5972a),
	.w5(32'hbbb6cf90),
	.w6(32'hbb2fe9b3),
	.w7(32'hba493a3a),
	.w8(32'hbaf7e8f0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7216a),
	.w1(32'h3bb10b51),
	.w2(32'hbb7ae281),
	.w3(32'hbb9a08c2),
	.w4(32'h3bf9a731),
	.w5(32'hbb4ffaa6),
	.w6(32'h3b6ca3e4),
	.w7(32'h3bd66906),
	.w8(32'h3ca43f63),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aca89),
	.w1(32'h3b4a5da7),
	.w2(32'h3b0f0e85),
	.w3(32'hbb8b71cd),
	.w4(32'hbb8943f0),
	.w5(32'hbba810e8),
	.w6(32'h3c73b1a8),
	.w7(32'h3c63842f),
	.w8(32'hbbd71363),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ee46e),
	.w1(32'hba9602d7),
	.w2(32'h3ac0c704),
	.w3(32'hbc24d4cf),
	.w4(32'hbb8a40f1),
	.w5(32'h3b7c4fe4),
	.w6(32'hbc0cdba2),
	.w7(32'hba4391ae),
	.w8(32'h3bbb4a28),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f8252),
	.w1(32'h3ca9282a),
	.w2(32'h3c68857f),
	.w3(32'h3bab7c5b),
	.w4(32'h3b5fa7bc),
	.w5(32'hbc1cad06),
	.w6(32'hbbe69ca9),
	.w7(32'h3c0f7d64),
	.w8(32'hba9d1421),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01963a),
	.w1(32'hbbedad5b),
	.w2(32'hbb0ad32e),
	.w3(32'hbb196a7f),
	.w4(32'hbc092ad1),
	.w5(32'hbbc92c8d),
	.w6(32'hbafb9c3b),
	.w7(32'h3ba7d7b6),
	.w8(32'h3af6f0de),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ca571),
	.w1(32'h3ab3b441),
	.w2(32'h3b671a22),
	.w3(32'hbbeb2d79),
	.w4(32'h3bcc24f1),
	.w5(32'h3b20b5ca),
	.w6(32'h3bf54ea0),
	.w7(32'h3b59c31f),
	.w8(32'hb9dbbdd6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e69ff),
	.w1(32'h3a17503d),
	.w2(32'hba785f47),
	.w3(32'hbb109e09),
	.w4(32'hb71ab8f5),
	.w5(32'hbb5be548),
	.w6(32'hbad50624),
	.w7(32'h3b58ff03),
	.w8(32'hbb825ded),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2dbcb),
	.w1(32'h3b269d66),
	.w2(32'h3b281def),
	.w3(32'hbc227344),
	.w4(32'hbbb4c2e6),
	.w5(32'hbad139fc),
	.w6(32'h3b59baac),
	.w7(32'hbab75092),
	.w8(32'hbb85d729),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e0310),
	.w1(32'hbb915d8a),
	.w2(32'hbb6daa12),
	.w3(32'h3b70d79e),
	.w4(32'h3bf4608f),
	.w5(32'h3b588c52),
	.w6(32'hbbe3e6f8),
	.w7(32'h3b2cf9bf),
	.w8(32'hbb6bf152),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98f34f),
	.w1(32'hb99be042),
	.w2(32'hb99b1ef6),
	.w3(32'hbbecda2f),
	.w4(32'hba51d671),
	.w5(32'h3c0226fa),
	.w6(32'h3c5eeb3a),
	.w7(32'hbb289f62),
	.w8(32'hbc1d85db),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3bb38),
	.w1(32'h3b7d2fe7),
	.w2(32'h3bf8e6d6),
	.w3(32'hbba79bf7),
	.w4(32'hbc437ce4),
	.w5(32'hbb612171),
	.w6(32'hbbb25509),
	.w7(32'hbc1f447f),
	.w8(32'hbb5b69dc),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb656858),
	.w1(32'hbaf2e64d),
	.w2(32'hbb5b469e),
	.w3(32'hba9b9a53),
	.w4(32'hbb1526cf),
	.w5(32'h3b53e7c1),
	.w6(32'hb9eb400b),
	.w7(32'hbb418218),
	.w8(32'h3a64bfe2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb091fd7),
	.w1(32'hbb06d896),
	.w2(32'hba86a582),
	.w3(32'hbb2bd31f),
	.w4(32'hb911e253),
	.w5(32'h3b4546e6),
	.w6(32'h3adaf6cf),
	.w7(32'h3bcf4016),
	.w8(32'hba9b0698),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4453f9),
	.w1(32'hba89aecb),
	.w2(32'hbad0925b),
	.w3(32'h3a956251),
	.w4(32'h3a81c630),
	.w5(32'h3b924377),
	.w6(32'hbb98c3f9),
	.w7(32'hbace7c43),
	.w8(32'hbc2bc448),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33e421),
	.w1(32'hbb1b5a92),
	.w2(32'hbb9583ab),
	.w3(32'hbaefdac4),
	.w4(32'hbb3bb5b4),
	.w5(32'h3af4fdcd),
	.w6(32'h3bb3b086),
	.w7(32'hbb9f3b9d),
	.w8(32'h3abd69d8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1434b8),
	.w1(32'h3ad405da),
	.w2(32'h3b839cba),
	.w3(32'h3965fa5b),
	.w4(32'hbb3c6807),
	.w5(32'h3b0b611b),
	.w6(32'h3a69e339),
	.w7(32'hbaa9a389),
	.w8(32'h3a95b547),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a39e3),
	.w1(32'h3b88c35b),
	.w2(32'h3b6cbbf3),
	.w3(32'hbad13655),
	.w4(32'h3b8d58ea),
	.w5(32'hb99aa05e),
	.w6(32'hba899e3a),
	.w7(32'h3c1b75e1),
	.w8(32'hbb29daca),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e41cda),
	.w1(32'hbb73c7a9),
	.w2(32'hbad23269),
	.w3(32'hbb7e35b5),
	.w4(32'h3ac07272),
	.w5(32'hb8e60d72),
	.w6(32'hbbe7a1aa),
	.w7(32'hbb2085f1),
	.w8(32'hb8d53192),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb836d7c),
	.w1(32'h3a345516),
	.w2(32'h3ba46371),
	.w3(32'hbb9aeb22),
	.w4(32'hbba4c170),
	.w5(32'hbc3c8c2e),
	.w6(32'hbb9dbdac),
	.w7(32'h3b8670cf),
	.w8(32'h3c08f0db),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96044a),
	.w1(32'h392b0330),
	.w2(32'hbb9547f2),
	.w3(32'hbc1ee160),
	.w4(32'h3c602485),
	.w5(32'h39cab38b),
	.w6(32'h3c218cec),
	.w7(32'h3c36d9a1),
	.w8(32'h3b42569e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cadf0),
	.w1(32'hba503b72),
	.w2(32'hbb20dc65),
	.w3(32'hb8ca65ea),
	.w4(32'hbaad680a),
	.w5(32'h3c4e91c3),
	.w6(32'hbac237b1),
	.w7(32'hbac37c75),
	.w8(32'hbb9f1bdb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8708e5),
	.w1(32'hbbbaabd8),
	.w2(32'h39e2e37e),
	.w3(32'h3c140d09),
	.w4(32'h3cb1ed4e),
	.w5(32'hbb1286a6),
	.w6(32'h363e9ecc),
	.w7(32'hbb3303a3),
	.w8(32'hbb9af7c8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389933ab),
	.w1(32'hb9e099f5),
	.w2(32'h3b1c57f6),
	.w3(32'hb9925bd7),
	.w4(32'h3b617e06),
	.w5(32'hbc1758cd),
	.w6(32'hbb268978),
	.w7(32'hbaac4916),
	.w8(32'h3bc49ec6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68731e),
	.w1(32'h3c26f468),
	.w2(32'hbbd5bbf8),
	.w3(32'hbc826eed),
	.w4(32'h3aaac235),
	.w5(32'h3ad4308d),
	.w6(32'h3c7559a0),
	.w7(32'h3bac09be),
	.w8(32'hb884270c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9afab),
	.w1(32'h3b334fa6),
	.w2(32'h3b3bceee),
	.w3(32'h3aa78b12),
	.w4(32'h392bb0ea),
	.w5(32'h3ba6219a),
	.w6(32'hba72a549),
	.w7(32'hb772fc12),
	.w8(32'h39c3c3eb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48e3f0),
	.w1(32'hbb7083cc),
	.w2(32'h38ca0b29),
	.w3(32'h3b1498a8),
	.w4(32'hbb0e0ed8),
	.w5(32'hbabf8ba2),
	.w6(32'h3af300c4),
	.w7(32'h3b306e90),
	.w8(32'hba7e357b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a531467),
	.w1(32'h3b6262cd),
	.w2(32'h3b53ffc3),
	.w3(32'hbb5d9799),
	.w4(32'hbbb8111c),
	.w5(32'h3a9079f8),
	.w6(32'h3a991900),
	.w7(32'h3a9bcdc7),
	.w8(32'h3b2056f2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b87bc),
	.w1(32'h3a59d207),
	.w2(32'hba144e0d),
	.w3(32'h3aeb9b51),
	.w4(32'hbb8c8c46),
	.w5(32'hbbf16cfe),
	.w6(32'h3bf9211b),
	.w7(32'h3bb68c9e),
	.w8(32'h3c75e983),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf15852),
	.w1(32'h3c981fbe),
	.w2(32'h3b4ae22d),
	.w3(32'hbc879695),
	.w4(32'h3c46571e),
	.w5(32'hbb9b1ee6),
	.w6(32'h3bb0d2d6),
	.w7(32'h3c922109),
	.w8(32'hbb799705),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24c529),
	.w1(32'hbab94fdf),
	.w2(32'hba1b0f85),
	.w3(32'hbbcdaba8),
	.w4(32'hbbed6b94),
	.w5(32'h3b602c88),
	.w6(32'hbb4e0e5d),
	.w7(32'h3a194f68),
	.w8(32'h3b00d106),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf80e27),
	.w1(32'h3c5375fc),
	.w2(32'h3c27ff60),
	.w3(32'h3bbc8ff6),
	.w4(32'h3be9cf3d),
	.w5(32'hbba59659),
	.w6(32'h3c291a38),
	.w7(32'h3b855f63),
	.w8(32'hb9db99bc),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec1c4d),
	.w1(32'h3ab849f6),
	.w2(32'h3b00f819),
	.w3(32'h38104ddf),
	.w4(32'h3adcc04b),
	.w5(32'hba91234e),
	.w6(32'h3ada2e95),
	.w7(32'h3b02900f),
	.w8(32'hb8d2acb5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6e9bd),
	.w1(32'h3c54ccc2),
	.w2(32'h3b2664b2),
	.w3(32'hbbf61a89),
	.w4(32'hbb2c5ff6),
	.w5(32'hba9bfe80),
	.w6(32'h3bf30ac7),
	.w7(32'h3bd5ce12),
	.w8(32'hbc0fcab9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c041b2b),
	.w1(32'hbc1449cf),
	.w2(32'hbb38e6bf),
	.w3(32'hbb8febfe),
	.w4(32'h3c7eaf75),
	.w5(32'hba5488df),
	.w6(32'h3a4971f2),
	.w7(32'hbb32b459),
	.w8(32'hba351d90),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98beccd),
	.w1(32'h3b8b4fcd),
	.w2(32'h3af61de1),
	.w3(32'h387e96d4),
	.w4(32'h3aa49b2d),
	.w5(32'h3b7e2fc1),
	.w6(32'hbab98078),
	.w7(32'hbb03738d),
	.w8(32'hbb06c9ab),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb538e8d),
	.w1(32'hbc29a6fd),
	.w2(32'hbc0f0795),
	.w3(32'h3a7068b8),
	.w4(32'h3b8cdae1),
	.w5(32'hbab2c266),
	.w6(32'hbbb0cf10),
	.w7(32'hbc0a50b5),
	.w8(32'hbbd07e78),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14ea64),
	.w1(32'hbb255d52),
	.w2(32'hba8cde43),
	.w3(32'hbbc3f9cf),
	.w4(32'hbbbdad8d),
	.w5(32'hbb36fb7a),
	.w6(32'hbb8fa2ad),
	.w7(32'hbbc5746b),
	.w8(32'hbb619e67),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16f676),
	.w1(32'hb8e45ff6),
	.w2(32'hbaa7c911),
	.w3(32'hbb0b7c57),
	.w4(32'hb9bccd14),
	.w5(32'hbc00e719),
	.w6(32'hbb4682ca),
	.w7(32'hbb8926ce),
	.w8(32'h3abc0417),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d517f),
	.w1(32'h3bfdb00e),
	.w2(32'h3984dc35),
	.w3(32'hbc26e9af),
	.w4(32'hbc025bd6),
	.w5(32'hba9a6e06),
	.w6(32'h3bf0e483),
	.w7(32'h3bb7a1db),
	.w8(32'h3a188f70),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5abad),
	.w1(32'h3b286553),
	.w2(32'h3af9a3d6),
	.w3(32'hba283afb),
	.w4(32'hba0bc34b),
	.w5(32'hbba21cba),
	.w6(32'h3b3174b4),
	.w7(32'h3a76583a),
	.w8(32'hbbbf46f0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049e35),
	.w1(32'hbaf23bdb),
	.w2(32'hbc114012),
	.w3(32'hbbccba59),
	.w4(32'hbb832cda),
	.w5(32'hb8d4d40c),
	.w6(32'h3b9a623f),
	.w7(32'hbbe9c0f5),
	.w8(32'hbaf9041a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee8710),
	.w1(32'hba98deeb),
	.w2(32'hbad8a525),
	.w3(32'hbb3bf3b9),
	.w4(32'hbaf51992),
	.w5(32'hbb19c995),
	.w6(32'hbb18129e),
	.w7(32'hbb4b1de1),
	.w8(32'hba435e58),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38896b15),
	.w1(32'h3b609e2b),
	.w2(32'h3ad3f742),
	.w3(32'h389a2c01),
	.w4(32'h3b03726b),
	.w5(32'h3b1e3c29),
	.w6(32'h3ac1c520),
	.w7(32'h3ad169e7),
	.w8(32'h3adf463a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b47ba),
	.w1(32'h3ab4dfa0),
	.w2(32'h3bb245a5),
	.w3(32'h389ed0ee),
	.w4(32'hbb9dad27),
	.w5(32'h393ac805),
	.w6(32'h3b00beca),
	.w7(32'h39bc0834),
	.w8(32'h3942516c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f50cae),
	.w1(32'hbb1af000),
	.w2(32'hbae0fcce),
	.w3(32'hbad3dad2),
	.w4(32'hba4baa56),
	.w5(32'hbb10c143),
	.w6(32'hbb941d62),
	.w7(32'hbaadd9a9),
	.w8(32'hbb18c7f3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50cbbe),
	.w1(32'h398c8f94),
	.w2(32'h3aa589bd),
	.w3(32'hbaeaae63),
	.w4(32'h396c2f67),
	.w5(32'hba28269d),
	.w6(32'hbb413387),
	.w7(32'hbb55d09f),
	.w8(32'hbb9601d2),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12aab8),
	.w1(32'hbb0ee618),
	.w2(32'hbb3b3449),
	.w3(32'hbb8e1a29),
	.w4(32'hbb92f6d2),
	.w5(32'h3b069a6a),
	.w6(32'hba538bcb),
	.w7(32'hbbb92696),
	.w8(32'hbb1661d5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb322bd5),
	.w1(32'hbb141a74),
	.w2(32'hbb74fe47),
	.w3(32'h3bbeb297),
	.w4(32'h3b2795cd),
	.w5(32'h3b5d5e79),
	.w6(32'hbb8e7bf7),
	.w7(32'h3a8a4bfb),
	.w8(32'hbaac4403),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec6453),
	.w1(32'hbb7cc918),
	.w2(32'hbbdf2f29),
	.w3(32'h3ac273a1),
	.w4(32'h3b56ab35),
	.w5(32'hbc6dc807),
	.w6(32'h3a402c9e),
	.w7(32'h3b28ba9b),
	.w8(32'hbc0019a6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81da7e),
	.w1(32'hbc8850ec),
	.w2(32'hbc8b2190),
	.w3(32'hbc2b8cda),
	.w4(32'h3c3dd783),
	.w5(32'h3b02013c),
	.w6(32'hbbb2f72a),
	.w7(32'hbc0cd4d6),
	.w8(32'h3b6b5bbe),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18e8f7),
	.w1(32'h3b3c1184),
	.w2(32'h3b64a95b),
	.w3(32'h3902bbdf),
	.w4(32'h3a66a0c9),
	.w5(32'hba16fbcd),
	.w6(32'h3ad05481),
	.w7(32'h3b807052),
	.w8(32'h3b427279),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad188dd),
	.w1(32'h3b008fa5),
	.w2(32'hba9f995b),
	.w3(32'h39cf769a),
	.w4(32'hbafad9e6),
	.w5(32'h3a93e1a6),
	.w6(32'h3bbf52e5),
	.w7(32'hbb5ece44),
	.w8(32'h3a0eacaa),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afedbe1),
	.w1(32'h3a02cc02),
	.w2(32'h3a2cdd9e),
	.w3(32'hba8d577c),
	.w4(32'h3b1b0486),
	.w5(32'hbb8f6b0b),
	.w6(32'hbb0330d6),
	.w7(32'h3a984957),
	.w8(32'hba1da4c2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4a241),
	.w1(32'h3b0a20dc),
	.w2(32'h3b56593b),
	.w3(32'hbbd22244),
	.w4(32'hbbafb5e1),
	.w5(32'hbb10293b),
	.w6(32'h3ac8e931),
	.w7(32'h3addd394),
	.w8(32'h3b932d11),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772ad1c),
	.w1(32'h3a9366ec),
	.w2(32'hbabfdab7),
	.w3(32'hbb87269d),
	.w4(32'hbbbcdbc7),
	.w5(32'hbc0e4c0e),
	.w6(32'h3bc23979),
	.w7(32'h3a9b4ed5),
	.w8(32'hbc3205d9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c959),
	.w1(32'hbb93546b),
	.w2(32'hbb9dcc2e),
	.w3(32'hbbf319b7),
	.w4(32'h3b51afc7),
	.w5(32'h3aa50e44),
	.w6(32'hb70499f1),
	.w7(32'hbc1068fd),
	.w8(32'hb9e3b69e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbf8a6),
	.w1(32'hb9fbce0a),
	.w2(32'h38e7c873),
	.w3(32'hba9c1557),
	.w4(32'hbaf9762c),
	.w5(32'h3b708a02),
	.w6(32'hb9c0d44d),
	.w7(32'hbb8d2169),
	.w8(32'h3a6e4fbc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b8d7e),
	.w1(32'hba769cbf),
	.w2(32'h3b305170),
	.w3(32'h3b3bc770),
	.w4(32'h3b88d814),
	.w5(32'h3c12dd24),
	.w6(32'hbb8a02c3),
	.w7(32'h3a247fa5),
	.w8(32'hbbdc5c9b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6cb2c),
	.w1(32'hbbfa77e5),
	.w2(32'h3bc0f7ab),
	.w3(32'h3b963a8b),
	.w4(32'h3b5bc654),
	.w5(32'hbb213a6f),
	.w6(32'hbbfb8721),
	.w7(32'hbb6f3f91),
	.w8(32'hbb1205af),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98881ff),
	.w1(32'hba8ba8ea),
	.w2(32'h3a25a2d9),
	.w3(32'hbbb9c244),
	.w4(32'hbb490541),
	.w5(32'h3bf16cb1),
	.w6(32'h3b42d94a),
	.w7(32'hbb581320),
	.w8(32'h3c88e185),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba319d6),
	.w1(32'h3bc9c715),
	.w2(32'h3b9cb9c4),
	.w3(32'hbb194a6d),
	.w4(32'hba7defcb),
	.w5(32'h3885dbc4),
	.w6(32'h3d2a1fe7),
	.w7(32'h3c7ce6b0),
	.w8(32'h3b673d04),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17b1c1),
	.w1(32'hba33f56c),
	.w2(32'h3aac1721),
	.w3(32'hbb1ad1ca),
	.w4(32'hbaad0b6f),
	.w5(32'h39d8e034),
	.w6(32'hba824e5c),
	.w7(32'hba19271c),
	.w8(32'h397ad27e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e406),
	.w1(32'hbb81de5f),
	.w2(32'hbaf798e2),
	.w3(32'h3b0dec6d),
	.w4(32'h3b1f1667),
	.w5(32'hb9a9141a),
	.w6(32'hbb59f941),
	.w7(32'h3b98b1e1),
	.w8(32'hbb256737),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a5f76),
	.w1(32'hbadabcca),
	.w2(32'hbaedb6d5),
	.w3(32'hbb8afcbd),
	.w4(32'h393e1edb),
	.w5(32'hbc4db919),
	.w6(32'hbbe40463),
	.w7(32'hbb7e3988),
	.w8(32'hbc71f798),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0dba3),
	.w1(32'hbc2f1cd0),
	.w2(32'hbb91d462),
	.w3(32'hbc32c568),
	.w4(32'hbb32000b),
	.w5(32'hbb53f54a),
	.w6(32'hbaf65d5c),
	.w7(32'hbc1977cb),
	.w8(32'hbb2fe02f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9960f),
	.w1(32'h395b1a45),
	.w2(32'hbb6d6de7),
	.w3(32'hbc114c2f),
	.w4(32'hbc1351ed),
	.w5(32'hbb516b43),
	.w6(32'hbac7e739),
	.w7(32'hbb8dbd5a),
	.w8(32'hbb73daf0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc074e9),
	.w1(32'hbba838b4),
	.w2(32'hbbdfe1d4),
	.w3(32'hbb399d23),
	.w4(32'h3bc01d18),
	.w5(32'hb9bd142b),
	.w6(32'h3bb89920),
	.w7(32'hbbc56584),
	.w8(32'h3c088a5a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85be4d),
	.w1(32'h3be79e6f),
	.w2(32'h3b8f1b64),
	.w3(32'h3b49e09f),
	.w4(32'hbb70a10d),
	.w5(32'hbbb37d6b),
	.w6(32'h3c49a7b8),
	.w7(32'h3b43f0b5),
	.w8(32'hba05363f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2d22),
	.w1(32'hbc05f1fb),
	.w2(32'hbc00bc0c),
	.w3(32'hbbafb15d),
	.w4(32'hba98be9f),
	.w5(32'hbb98c278),
	.w6(32'hbb8a226f),
	.w7(32'hbbee8333),
	.w8(32'h3b2e65b3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b853e72),
	.w1(32'h3a57c9fb),
	.w2(32'h3b1c69ea),
	.w3(32'hbc0cc3f6),
	.w4(32'hbb9d066d),
	.w5(32'h3cd1b359),
	.w6(32'h3b900506),
	.w7(32'h3ad1d725),
	.w8(32'h3c991538),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9603e3),
	.w1(32'h3c49b80d),
	.w2(32'h3cc3ad5b),
	.w3(32'h3ccbbe9c),
	.w4(32'hba3ac496),
	.w5(32'hbaf07575),
	.w6(32'h3d415f1d),
	.w7(32'h3cc0d23f),
	.w8(32'hbadc8f2c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01c3d2),
	.w1(32'h3b91dd07),
	.w2(32'h3b9a5021),
	.w3(32'hbc0dd646),
	.w4(32'hbc0924fb),
	.w5(32'hbb51a806),
	.w6(32'h3ae51015),
	.w7(32'hba9cd445),
	.w8(32'hbac8e02d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa3c46),
	.w1(32'hba063a8f),
	.w2(32'hb8fbef23),
	.w3(32'h3bc83fc1),
	.w4(32'hba80c86b),
	.w5(32'hba07177f),
	.w6(32'h3aefd287),
	.w7(32'h3b06bd12),
	.w8(32'h3afaa351),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade81e8),
	.w1(32'h3ac5ab6a),
	.w2(32'h3b11df1e),
	.w3(32'hbb14b82a),
	.w4(32'hba87f745),
	.w5(32'hbb33ca07),
	.w6(32'h3a65a9d7),
	.w7(32'hba832cf6),
	.w8(32'hbbaf0ce1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab60fae),
	.w1(32'hbb111324),
	.w2(32'h3aecf257),
	.w3(32'hba44400f),
	.w4(32'h3b1173cf),
	.w5(32'hba9f7a8c),
	.w6(32'h3b2858e9),
	.w7(32'hbbaa46da),
	.w8(32'hbbcb6d9d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bc9a2),
	.w1(32'hba753002),
	.w2(32'h3aa754b3),
	.w3(32'hbafcda33),
	.w4(32'h3b7909ea),
	.w5(32'hbc23b584),
	.w6(32'hbc0cb7b5),
	.w7(32'hbb72b7b7),
	.w8(32'hbc2e3e3c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0109b),
	.w1(32'hbac589a2),
	.w2(32'h3b6b175e),
	.w3(32'hbc0dee1d),
	.w4(32'hbb2739c0),
	.w5(32'hba2b2255),
	.w6(32'hbc3dada7),
	.w7(32'hbc0d1a99),
	.w8(32'h3b61b953),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923ad54),
	.w1(32'h3abc84fd),
	.w2(32'h382859b7),
	.w3(32'h38f19ac2),
	.w4(32'hb9f88f81),
	.w5(32'hbaea6472),
	.w6(32'h3b15d289),
	.w7(32'h3b69a920),
	.w8(32'h3b497881),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a948c41),
	.w1(32'h3a5862cb),
	.w2(32'h3b32c30a),
	.w3(32'hbba16460),
	.w4(32'hbbde78ca),
	.w5(32'h3ad057f5),
	.w6(32'h3b567996),
	.w7(32'h3ad9e372),
	.w8(32'hbaf6448c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb63e18),
	.w1(32'hbc0ba988),
	.w2(32'h3a97773b),
	.w3(32'hb9faf06f),
	.w4(32'h3b990cff),
	.w5(32'hbb6927e7),
	.w6(32'h3bcb2c4b),
	.w7(32'h3bc53c25),
	.w8(32'hbb887add),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab96a83),
	.w1(32'h3b6ce947),
	.w2(32'h3bc1bea1),
	.w3(32'h3b40492b),
	.w4(32'hba61eae8),
	.w5(32'h3a15570b),
	.w6(32'hbb14bc7a),
	.w7(32'h3b416e40),
	.w8(32'hbabf316c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63854a),
	.w1(32'hbbe55172),
	.w2(32'hb8304f77),
	.w3(32'h3a9547d5),
	.w4(32'h3b79bf3a),
	.w5(32'h38a5112c),
	.w6(32'hbb6778c4),
	.w7(32'h3b043381),
	.w8(32'h3afc4b10),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0566a),
	.w1(32'hbbd563f2),
	.w2(32'hbb370e63),
	.w3(32'hbac97b49),
	.w4(32'h3abf9242),
	.w5(32'h3b87080f),
	.w6(32'hbac64f99),
	.w7(32'h3bc0efc0),
	.w8(32'hb99c47de),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6646e8),
	.w1(32'hb7258a9c),
	.w2(32'hb933a5fe),
	.w3(32'h3b1c6208),
	.w4(32'h3b8f9fae),
	.w5(32'h3b3b9130),
	.w6(32'hbaedd4a2),
	.w7(32'h397650ae),
	.w8(32'h3a8c149e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0a1c8),
	.w1(32'h3ae742c7),
	.w2(32'h3aedb8fb),
	.w3(32'h3ae34ef1),
	.w4(32'h399e0baa),
	.w5(32'h3a479556),
	.w6(32'h39591e0a),
	.w7(32'h376d2e70),
	.w8(32'h3a7f5e36),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e8fda),
	.w1(32'hba9993f7),
	.w2(32'hba869168),
	.w3(32'hba9d7413),
	.w4(32'hb8a3fa35),
	.w5(32'h3a836913),
	.w6(32'hb80606f0),
	.w7(32'h3900a78e),
	.w8(32'h3c08aad8),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cc2ae),
	.w1(32'h3bef04fd),
	.w2(32'hbc178f30),
	.w3(32'hbc6166ef),
	.w4(32'h3bf2d978),
	.w5(32'hbb085f0d),
	.w6(32'h3b7509b0),
	.w7(32'h3c24a895),
	.w8(32'hbb124cb2),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b2fa3),
	.w1(32'hbbdd6a68),
	.w2(32'hbb1d9c57),
	.w3(32'hbb44ff7b),
	.w4(32'h3b2bb654),
	.w5(32'hbca74f86),
	.w6(32'h3a976600),
	.w7(32'h3a4f46fe),
	.w8(32'h3aadbadb),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5b563),
	.w1(32'h3b9c32c6),
	.w2(32'hbc5322b6),
	.w3(32'hbc9efc92),
	.w4(32'hbb90b9fc),
	.w5(32'hbbcc0d5d),
	.w6(32'h3c18c179),
	.w7(32'h3afc326b),
	.w8(32'hbb050ade),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba51d00),
	.w1(32'h39765ff6),
	.w2(32'hbb6fe864),
	.w3(32'h3b190238),
	.w4(32'hbbb855e6),
	.w5(32'hbbad934a),
	.w6(32'hbaa6a4b8),
	.w7(32'hbb28eb2e),
	.w8(32'hbbc93563),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce1aa2),
	.w1(32'hbb9bebc1),
	.w2(32'hbb857a4e),
	.w3(32'hbb87d70a),
	.w4(32'hbbf121d6),
	.w5(32'h3c1ddae3),
	.w6(32'h3c2be272),
	.w7(32'hbbed17db),
	.w8(32'h3c0734f0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c97df),
	.w1(32'h3c3c48af),
	.w2(32'h3c7e7ca7),
	.w3(32'h3b8ff737),
	.w4(32'hbc8be2ae),
	.w5(32'h3b6d1da2),
	.w6(32'h3d13f5e2),
	.w7(32'h3be2e64f),
	.w8(32'h3bf15bee),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b934d4e),
	.w1(32'h3bda59e6),
	.w2(32'h3c63dcf2),
	.w3(32'h3b9ceacc),
	.w4(32'hbb32e8f5),
	.w5(32'hbbf08327),
	.w6(32'h3c08a842),
	.w7(32'h3bec4dc6),
	.w8(32'hbbfa7035),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58fc16),
	.w1(32'h3a6b6622),
	.w2(32'hbb78f8ac),
	.w3(32'hbc0fd72b),
	.w4(32'hbc0cdffa),
	.w5(32'hbb3234e9),
	.w6(32'h3b801f7d),
	.w7(32'hbc2bae78),
	.w8(32'h3a002136),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5a4a7),
	.w1(32'hb9b558bc),
	.w2(32'hbafa1e74),
	.w3(32'hbb251f52),
	.w4(32'hbb0ccb61),
	.w5(32'h3b2f3707),
	.w6(32'h3aad854e),
	.w7(32'h3897fdde),
	.w8(32'hb8fd5c08),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aef65),
	.w1(32'hbb849911),
	.w2(32'hbb6cc91c),
	.w3(32'hba84de23),
	.w4(32'hb9bb4237),
	.w5(32'h3a599afa),
	.w6(32'h3ac2c7ae),
	.w7(32'h3a31053f),
	.w8(32'hbb435d53),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d1f5a),
	.w1(32'hbb169e72),
	.w2(32'h3ad9fe4c),
	.w3(32'h3a760fc2),
	.w4(32'h3b7e294a),
	.w5(32'hbb2e1309),
	.w6(32'h3a004570),
	.w7(32'hba9f05db),
	.w8(32'hba717b94),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab14709),
	.w1(32'h385ee63c),
	.w2(32'hbad45c8c),
	.w3(32'h3a053f9b),
	.w4(32'h3b170d8d),
	.w5(32'h3c5347e6),
	.w6(32'h3abe932e),
	.w7(32'hba971355),
	.w8(32'h3c768ab0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b476),
	.w1(32'h3c11ff2a),
	.w2(32'h3ad21746),
	.w3(32'h3c73133e),
	.w4(32'h3c425a94),
	.w5(32'h3c08b888),
	.w6(32'h3d3ba185),
	.w7(32'h3c868b32),
	.w8(32'h3b58b2d2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bbfa2),
	.w1(32'h3c00664e),
	.w2(32'h3c8747c9),
	.w3(32'h3baab5d6),
	.w4(32'hbc37d98d),
	.w5(32'h3cc42032),
	.w6(32'h3c5e9610),
	.w7(32'h3bd65720),
	.w8(32'h3c1b932c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bfa9f),
	.w1(32'h3c9f40ed),
	.w2(32'h3c95059e),
	.w3(32'h3bfbde19),
	.w4(32'hbca1f4e5),
	.w5(32'hbc047a98),
	.w6(32'h3d0153cd),
	.w7(32'h3aa642a0),
	.w8(32'h3b8a52c0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a68bc),
	.w1(32'h369d3ace),
	.w2(32'hbb059300),
	.w3(32'hbbce76c9),
	.w4(32'hbbb761da),
	.w5(32'h39e95a9d),
	.w6(32'h3ce6923b),
	.w7(32'hba96bc9c),
	.w8(32'h3b108ced),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf745df),
	.w1(32'h3b1fda42),
	.w2(32'h3acb6550),
	.w3(32'hbab7176f),
	.w4(32'h39e2c41e),
	.w5(32'hbb7eea3a),
	.w6(32'h3b9b7969),
	.w7(32'h3b8b1cb2),
	.w8(32'hb9393153),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccc033),
	.w1(32'hbb536b41),
	.w2(32'hbba21d09),
	.w3(32'h3b3f82a8),
	.w4(32'h3bd14532),
	.w5(32'hbb9d5094),
	.w6(32'hbb3df8e8),
	.w7(32'hb99256e2),
	.w8(32'hbbf3858d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0906f7),
	.w1(32'h399b4a05),
	.w2(32'hba903035),
	.w3(32'hbc67e9c0),
	.w4(32'hbc95c392),
	.w5(32'h3b357965),
	.w6(32'hbb39cccb),
	.w7(32'hbc38ddef),
	.w8(32'hbac5f47e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40ee17),
	.w1(32'hbb481f77),
	.w2(32'h3b750eb9),
	.w3(32'hbaae9a33),
	.w4(32'h399399b5),
	.w5(32'h3aa63f7a),
	.w6(32'hbc5ae62e),
	.w7(32'h3b0899bf),
	.w8(32'h3adfd97c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e30aed),
	.w1(32'h3b42d20b),
	.w2(32'h3af3fd24),
	.w3(32'h3bb057e3),
	.w4(32'h3b214bee),
	.w5(32'hbadb716e),
	.w6(32'hba5bafbb),
	.w7(32'h3bbe3321),
	.w8(32'hbb98b6ab),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb354108),
	.w1(32'hbb920d17),
	.w2(32'hbb2c4d38),
	.w3(32'hbaa1c2a7),
	.w4(32'hbb520714),
	.w5(32'hbb399c39),
	.w6(32'h3aac6518),
	.w7(32'hbb14a316),
	.w8(32'hbb8c932d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8b6a1),
	.w1(32'hbbd61bec),
	.w2(32'hbb3c2ba0),
	.w3(32'hbbc4d3f8),
	.w4(32'hbbf69208),
	.w5(32'h3ab07da7),
	.w6(32'h3b453586),
	.w7(32'hba6de7f9),
	.w8(32'h381c4c43),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccea2b),
	.w1(32'hba8c6276),
	.w2(32'hbad92e59),
	.w3(32'hbb0a699a),
	.w4(32'hbb145b44),
	.w5(32'hbb0e5f83),
	.w6(32'hbaf3b4bc),
	.w7(32'hbb0c1197),
	.w8(32'h3a0e6709),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d90b94),
	.w1(32'hbb5d7b26),
	.w2(32'hbb73938e),
	.w3(32'hbb2c82f8),
	.w4(32'hbb71843c),
	.w5(32'h3ad600d7),
	.w6(32'hbaab3b75),
	.w7(32'hbb8bdb8f),
	.w8(32'hba8fa667),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb574a42),
	.w1(32'hbbc15095),
	.w2(32'hbb1a3464),
	.w3(32'h39b18f06),
	.w4(32'hb969a9f8),
	.w5(32'h3b0ca8a3),
	.w6(32'h3a06ceb7),
	.w7(32'hba90968c),
	.w8(32'hbb69d05f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2287f),
	.w1(32'h3b1de0cc),
	.w2(32'h3b9df6ae),
	.w3(32'hbb9fa3d7),
	.w4(32'hbb87327f),
	.w5(32'hb9a7b094),
	.w6(32'h39fb278c),
	.w7(32'hbbed30f4),
	.w8(32'hbbb7d018),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39cc43),
	.w1(32'hbaf924d0),
	.w2(32'h3b9f1db1),
	.w3(32'h3a2610dc),
	.w4(32'h3abb0a7f),
	.w5(32'hbb0567d2),
	.w6(32'h3b32fba4),
	.w7(32'h3b3b8c07),
	.w8(32'h3b506518),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7522d2),
	.w1(32'h37069913),
	.w2(32'h3b10f89e),
	.w3(32'h3a3ab7cd),
	.w4(32'h3911e218),
	.w5(32'h3b94da97),
	.w6(32'hb9e26cbe),
	.w7(32'h3ab85b20),
	.w8(32'h3b0aeca5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b69d23),
	.w1(32'h3b5e3253),
	.w2(32'h3b76efea),
	.w3(32'h3b7aa258),
	.w4(32'h3bb339a9),
	.w5(32'h3ba838b3),
	.w6(32'hbac1827d),
	.w7(32'hb9c4007b),
	.w8(32'h3a51b14a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0558c5),
	.w1(32'h3a9ec874),
	.w2(32'h3a013085),
	.w3(32'h3bdaf367),
	.w4(32'hba23b575),
	.w5(32'hba4e926a),
	.w6(32'h3b27059b),
	.w7(32'hbb074d99),
	.w8(32'hba16f703),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b027ded),
	.w1(32'h3b929f45),
	.w2(32'hba1d864d),
	.w3(32'hbba39539),
	.w4(32'hbbd5ccb3),
	.w5(32'h3bcbe35d),
	.w6(32'hbad02e71),
	.w7(32'hbbaba66a),
	.w8(32'hbc3f1cd2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a698c),
	.w1(32'hbb4473c1),
	.w2(32'h3b60087c),
	.w3(32'hbc324815),
	.w4(32'hbc9c6475),
	.w5(32'hbb4be5e2),
	.w6(32'hbc13c9bd),
	.w7(32'hbc64bfeb),
	.w8(32'hbb9f3a0b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2faf25),
	.w1(32'h3a85e872),
	.w2(32'h3a8cbf12),
	.w3(32'hbac23ead),
	.w4(32'h3b4fa5b0),
	.w5(32'h3baf00be),
	.w6(32'hbb2253fa),
	.w7(32'h3ac91e25),
	.w8(32'hbbd05507),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bc82a),
	.w1(32'hbc1931c1),
	.w2(32'h3a056d3f),
	.w3(32'hbb72d6fc),
	.w4(32'h3b309bbc),
	.w5(32'hbab2e122),
	.w6(32'hbc0a0362),
	.w7(32'hbbb61b68),
	.w8(32'hbc04342b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1db3d9),
	.w1(32'hb9feb056),
	.w2(32'hb9933008),
	.w3(32'hba745cd2),
	.w4(32'hba487e5e),
	.w5(32'hbb71a169),
	.w6(32'h3b335b17),
	.w7(32'hbbf89134),
	.w8(32'hbab80193),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac6a1),
	.w1(32'h3bad5068),
	.w2(32'hbb7e018c),
	.w3(32'hbafe7e8f),
	.w4(32'hbbcce1a1),
	.w5(32'hbbea833e),
	.w6(32'hbb014435),
	.w7(32'h3b363f1d),
	.w8(32'h3aa81522),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0edaf4),
	.w1(32'hbbba7aff),
	.w2(32'hbaebc7e7),
	.w3(32'hbc2cc423),
	.w4(32'hbb1058f6),
	.w5(32'hba229841),
	.w6(32'h3c397ebb),
	.w7(32'h3afec479),
	.w8(32'h3b6afdc4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b50e9),
	.w1(32'hba4678ba),
	.w2(32'hb947a7e1),
	.w3(32'h38950072),
	.w4(32'h3b4697bf),
	.w5(32'hbb810986),
	.w6(32'hbadb0727),
	.w7(32'h3b51475f),
	.w8(32'hbadd3ff0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc77183),
	.w1(32'h3b60eb23),
	.w2(32'h3b49c77f),
	.w3(32'hbb8a81a9),
	.w4(32'hb97bd2bd),
	.w5(32'h3a88d401),
	.w6(32'hbb5dce03),
	.w7(32'hbad95ba8),
	.w8(32'hbb7a38cb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68e9a1),
	.w1(32'h3b50c702),
	.w2(32'h3b5b92d2),
	.w3(32'h3b249d47),
	.w4(32'h3bb4be9e),
	.w5(32'hbb892341),
	.w6(32'hbb4b0212),
	.w7(32'h3a3737e6),
	.w8(32'hbaa7bb11),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e9272),
	.w1(32'h398486cb),
	.w2(32'hbac64e87),
	.w3(32'hbb85b29e),
	.w4(32'hbbb23636),
	.w5(32'hbb298ad5),
	.w6(32'h3c1d6b61),
	.w7(32'hbb86f863),
	.w8(32'h3ab30c32),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc031635),
	.w1(32'h3b97caa4),
	.w2(32'h3c01b58d),
	.w3(32'h3a241d2b),
	.w4(32'hbb4bd7ec),
	.w5(32'hbb86f849),
	.w6(32'h3c2747d5),
	.w7(32'h3b7e69ee),
	.w8(32'h3abaaace),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8335e),
	.w1(32'hbbf83b8c),
	.w2(32'hbaef296b),
	.w3(32'hbba26d14),
	.w4(32'hbb12068e),
	.w5(32'hbb66431e),
	.w6(32'h3bc26eb3),
	.w7(32'h3b10a9b9),
	.w8(32'hbaf832fc),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51892c),
	.w1(32'hba2b225a),
	.w2(32'hbac004ef),
	.w3(32'hbb882e8f),
	.w4(32'hba845e3d),
	.w5(32'hb9e63112),
	.w6(32'hbab4da4e),
	.w7(32'hbbbaf77b),
	.w8(32'h3a6c75a2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bef6af),
	.w1(32'hbbf1ab23),
	.w2(32'hbb938c54),
	.w3(32'h3a9a3413),
	.w4(32'h3a09a4c1),
	.w5(32'hba247560),
	.w6(32'h3b19c573),
	.w7(32'hb9b1e03a),
	.w8(32'h39d50af6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86dd33),
	.w1(32'hbb11fe62),
	.w2(32'hb8d7bb63),
	.w3(32'hbaad0dac),
	.w4(32'h3b062ae8),
	.w5(32'h3b5b72b9),
	.w6(32'hbbbfaadd),
	.w7(32'hbb0f837f),
	.w8(32'h3b9cc950),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb542f3b),
	.w1(32'h3a9df39e),
	.w2(32'hbac382c3),
	.w3(32'hbabc2eab),
	.w4(32'h398f2c0e),
	.w5(32'hb9d4c0a7),
	.w6(32'h3be92474),
	.w7(32'hbb587ad1),
	.w8(32'hb980baff),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb639c82a),
	.w1(32'h3997ec2e),
	.w2(32'h39ce847b),
	.w3(32'h39736d1b),
	.w4(32'h392641a1),
	.w5(32'hba96e40d),
	.w6(32'hb8d2a18b),
	.w7(32'h39765a3b),
	.w8(32'h39fe957c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba400a7c),
	.w1(32'hbb5b7fc3),
	.w2(32'hbb024906),
	.w3(32'hba788663),
	.w4(32'hbaaa3750),
	.w5(32'h35ed39d2),
	.w6(32'hbb4478f3),
	.w7(32'hbb4c985f),
	.w8(32'hbb5ea65a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fc443),
	.w1(32'h392a2ef5),
	.w2(32'hba1cf24c),
	.w3(32'h3a016e9b),
	.w4(32'hb8f1d834),
	.w5(32'h37682ed7),
	.w6(32'hb94f46d6),
	.w7(32'hb93e8406),
	.w8(32'hbac232c6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39338ee7),
	.w1(32'h3a434b2b),
	.w2(32'hba43c850),
	.w3(32'h3988f6b4),
	.w4(32'h394dcb13),
	.w5(32'h39935c33),
	.w6(32'h398d0453),
	.w7(32'h3a28fb70),
	.w8(32'h3946fa54),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba441cef),
	.w1(32'hba17ca70),
	.w2(32'hb9c69f88),
	.w3(32'h389a486f),
	.w4(32'hb808be14),
	.w5(32'hbaa631d1),
	.w6(32'h38d83a74),
	.w7(32'hb9a1a1a6),
	.w8(32'hba2d75e7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad57592),
	.w1(32'hbaa3f75a),
	.w2(32'hbabe286c),
	.w3(32'hbb0ab1b4),
	.w4(32'hbb112547),
	.w5(32'h396ccc10),
	.w6(32'hba96cc67),
	.w7(32'hbac00253),
	.w8(32'hbb3a2854),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fef2b),
	.w1(32'hbad238bf),
	.w2(32'hb9d63b22),
	.w3(32'hba40d7f2),
	.w4(32'h3895555f),
	.w5(32'hb984ea54),
	.w6(32'hbac41403),
	.w7(32'hba5859b1),
	.w8(32'hb9bd66ef),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9f86a),
	.w1(32'hbb14a8c1),
	.w2(32'hbae35ec2),
	.w3(32'hbad47c06),
	.w4(32'hba0f19fc),
	.w5(32'hba174f4e),
	.w6(32'hbb19b146),
	.w7(32'hbaba1339),
	.w8(32'hb83a8936),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52b37e),
	.w1(32'hbae4e627),
	.w2(32'hb963b021),
	.w3(32'hba934d88),
	.w4(32'h39998642),
	.w5(32'h39af2898),
	.w6(32'h3a19ef06),
	.w7(32'h3ad3853b),
	.w8(32'h3a0cc40d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d211de),
	.w1(32'h3ab2d7be),
	.w2(32'h3a8d6456),
	.w3(32'h3aa52e5f),
	.w4(32'h3abc773b),
	.w5(32'hbab03820),
	.w6(32'h3adf8613),
	.w7(32'h3a7cee83),
	.w8(32'hbb01a942),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0b014),
	.w1(32'hbac959c9),
	.w2(32'hba855ddf),
	.w3(32'hba841453),
	.w4(32'hbaacea43),
	.w5(32'h37ec2eac),
	.w6(32'hbaff1a99),
	.w7(32'hbaa02a7f),
	.w8(32'hb8ee5a63),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3951d4b8),
	.w1(32'h3ab8b568),
	.w2(32'h3a328f21),
	.w3(32'h3ad30115),
	.w4(32'h3a5c0f42),
	.w5(32'hbb189de9),
	.w6(32'h3ad6a6d9),
	.w7(32'h3a8c0b68),
	.w8(32'hba8ecf0b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37580cf4),
	.w1(32'h3966cad0),
	.w2(32'hbade1239),
	.w3(32'hbaf21602),
	.w4(32'hba55243d),
	.w5(32'hb9692b0c),
	.w6(32'hba6626d5),
	.w7(32'hbafbc9d5),
	.w8(32'h3a384134),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e61bf),
	.w1(32'h39f9053a),
	.w2(32'h398c2357),
	.w3(32'hbaa70850),
	.w4(32'hba5d6508),
	.w5(32'h38d10c7d),
	.w6(32'h3a7802cf),
	.w7(32'hb9253df5),
	.w8(32'hba6d450e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70f6dc),
	.w1(32'h39cbdc97),
	.w2(32'h3a13f965),
	.w3(32'h382acd22),
	.w4(32'h399dd4a7),
	.w5(32'h3a6bc97d),
	.w6(32'h3a80d368),
	.w7(32'h38a115d2),
	.w8(32'hba909425),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a75b43),
	.w1(32'h3a972055),
	.w2(32'h3a955ab0),
	.w3(32'h39316e02),
	.w4(32'h39bd68e9),
	.w5(32'h3983c958),
	.w6(32'hba5b0c17),
	.w7(32'hba18d72b),
	.w8(32'h395bda50),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67eba2),
	.w1(32'h39160455),
	.w2(32'h397d0572),
	.w3(32'h3a1424d1),
	.w4(32'h3b193ca4),
	.w5(32'hb9bb9f60),
	.w6(32'hba9f89c4),
	.w7(32'hb77aa95b),
	.w8(32'h3a0eb417),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a750726),
	.w1(32'h3a88f8b2),
	.w2(32'hb9110fd9),
	.w3(32'hbaa2234c),
	.w4(32'hba83c8f2),
	.w5(32'h3b02f4fd),
	.w6(32'h3a8a02e9),
	.w7(32'h3a3dbb63),
	.w8(32'h3b16c715),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13fbac),
	.w1(32'h3ac57159),
	.w2(32'h3ade9324),
	.w3(32'h3ab386f4),
	.w4(32'h3aaf69ca),
	.w5(32'h3b44cfb0),
	.w6(32'h3a73e867),
	.w7(32'h3aca177a),
	.w8(32'h3a4aab6a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae647ed),
	.w1(32'hbb107114),
	.w2(32'hb9be16c6),
	.w3(32'h3a9c568b),
	.w4(32'h3a04e234),
	.w5(32'h3940587a),
	.w6(32'h3a8b6a6b),
	.w7(32'h3a01c121),
	.w8(32'hba373143),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab8255),
	.w1(32'hb9fc6aeb),
	.w2(32'hba89b20e),
	.w3(32'h3a61d840),
	.w4(32'h3a1b911d),
	.w5(32'hba49c651),
	.w6(32'hb9df6562),
	.w7(32'hb9564863),
	.w8(32'hba5996fc),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36af23),
	.w1(32'h3a3bed4c),
	.w2(32'h3a142b5e),
	.w3(32'hb9b124e7),
	.w4(32'hb75bb0d7),
	.w5(32'hbaa9732d),
	.w6(32'hba1af87c),
	.w7(32'h3ad90b37),
	.w8(32'hbb042cef),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3697e048),
	.w1(32'h3b017f2f),
	.w2(32'h3a7cf0bc),
	.w3(32'hba8ab2e7),
	.w4(32'hba853e90),
	.w5(32'hb961c26a),
	.w6(32'hba776a58),
	.w7(32'h39c8d41d),
	.w8(32'hba977077),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50c233),
	.w1(32'hba913065),
	.w2(32'hb92d958a),
	.w3(32'hb98ce389),
	.w4(32'hba1b9638),
	.w5(32'hbb05fdba),
	.w6(32'hb8864a64),
	.w7(32'h39b21835),
	.w8(32'hbaa7dd7b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad45b47),
	.w1(32'hba1c6ffb),
	.w2(32'hba06eb9d),
	.w3(32'hbaeeafd1),
	.w4(32'hb9b2c20f),
	.w5(32'hb9ce824b),
	.w6(32'hba2c561c),
	.w7(32'hba237942),
	.w8(32'hba3055c5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993afe2),
	.w1(32'hbaafd155),
	.w2(32'hba602653),
	.w3(32'hb98a570a),
	.w4(32'hb93a9b99),
	.w5(32'hba82d37c),
	.w6(32'h39e40db0),
	.w7(32'hb8cea2ee),
	.w8(32'hba7a0134),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d0c96),
	.w1(32'h3a54df1c),
	.w2(32'hba1f8ef1),
	.w3(32'h3907aca6),
	.w4(32'h396c5d80),
	.w5(32'hb9d3ac3e),
	.w6(32'h3a673bf1),
	.w7(32'h3928de27),
	.w8(32'hbaeec6d7),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba341654),
	.w1(32'hba83f5ab),
	.w2(32'hba954d12),
	.w3(32'h38925dca),
	.w4(32'hb90bed56),
	.w5(32'h3acc750c),
	.w6(32'hb9a89b06),
	.w7(32'h39c490e4),
	.w8(32'h3aa5be9b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab14e4b),
	.w1(32'h3a13b793),
	.w2(32'hb8ad4047),
	.w3(32'h3b1c4ec2),
	.w4(32'h3ad3261a),
	.w5(32'hba01b7bb),
	.w6(32'h3ae73bbe),
	.w7(32'h3ac8645f),
	.w8(32'hb905bf36),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3872ac),
	.w1(32'hb9f42038),
	.w2(32'hba40be36),
	.w3(32'hba037955),
	.w4(32'hb8e99a6d),
	.w5(32'hba1ac316),
	.w6(32'hb97cff32),
	.w7(32'h398b0100),
	.w8(32'hb9b26e9a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule