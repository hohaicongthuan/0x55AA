module layer_10_featuremap_100(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64e4d9b),
	.w1(32'h35c37afa),
	.w2(32'hb5a454ab),
	.w3(32'hb5f21276),
	.w4(32'h357a6244),
	.w5(32'hb64f609b),
	.w6(32'h3576917c),
	.w7(32'hb50991ce),
	.w8(32'hb6be1a41),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7e50b),
	.w1(32'h38d049e1),
	.w2(32'h38feae6b),
	.w3(32'h38ecbc06),
	.w4(32'h38d7df92),
	.w5(32'h38a046ea),
	.w6(32'h390ed453),
	.w7(32'h3844b875),
	.w8(32'hb8149d6e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e5ed31),
	.w1(32'hb647a30e),
	.w2(32'hb5b8aab0),
	.w3(32'h36c0eca2),
	.w4(32'hb67015ae),
	.w5(32'h35ea9909),
	.w6(32'hb667551b),
	.w7(32'hb6e56393),
	.w8(32'hb6a9d7c6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371e78f5),
	.w1(32'hb710fa16),
	.w2(32'h386a1b19),
	.w3(32'h37196560),
	.w4(32'h384df045),
	.w5(32'h38b771bc),
	.w6(32'h3792fab7),
	.w7(32'h376e5011),
	.w8(32'h38894646),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3715fbf8),
	.w1(32'hb6b720a4),
	.w2(32'h3708cbf6),
	.w3(32'h374a6900),
	.w4(32'hb6c6140d),
	.w5(32'h36ea913c),
	.w6(32'hb462901c),
	.w7(32'hb6854781),
	.w8(32'hb5b64af6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3688f44b),
	.w1(32'hb7059d86),
	.w2(32'hb758ab86),
	.w3(32'h36b83585),
	.w4(32'hb7022784),
	.w5(32'hb75fd5be),
	.w6(32'h36f6271e),
	.w7(32'hb63300fc),
	.w8(32'hb69b537c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384f4580),
	.w1(32'h39840508),
	.w2(32'hb82831dc),
	.w3(32'h3991e900),
	.w4(32'h39c46969),
	.w5(32'h38aef876),
	.w6(32'h398f0977),
	.w7(32'h3990bd13),
	.w8(32'hb7e5f4bf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb802d792),
	.w1(32'hb9ff1037),
	.w2(32'hba4d2e72),
	.w3(32'hb8ec29bd),
	.w4(32'hb999e2d1),
	.w5(32'hba1fc451),
	.w6(32'h3982de21),
	.w7(32'hba4161fd),
	.w8(32'hb9b8504a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba039e6a),
	.w1(32'hb9522d80),
	.w2(32'hb849669c),
	.w3(32'hb9ff4990),
	.w4(32'h3887ee42),
	.w5(32'h39053a0c),
	.w6(32'hb9f9e5a6),
	.w7(32'h38c87975),
	.w8(32'h39569e5b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba971614),
	.w1(32'hba8a83b6),
	.w2(32'hba727568),
	.w3(32'hba4eab74),
	.w4(32'hb9cb40bc),
	.w5(32'hba197c4d),
	.w6(32'hb953803b),
	.w7(32'h39214100),
	.w8(32'hb97e0baf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dbe5a0),
	.w1(32'hb98e07aa),
	.w2(32'hb99db9dc),
	.w3(32'h3815f1a6),
	.w4(32'hb8574f16),
	.w5(32'hb99a8637),
	.w6(32'h391fb85e),
	.w7(32'h3908579b),
	.w8(32'h38a66ecb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f173a0),
	.w1(32'hb75ff0ad),
	.w2(32'hb9b35ad6),
	.w3(32'h398e5622),
	.w4(32'h399c8f9d),
	.w5(32'h387bf121),
	.w6(32'h39d34f48),
	.w7(32'h39ccad89),
	.w8(32'h398586b1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993b15c),
	.w1(32'h397c3269),
	.w2(32'hb908357d),
	.w3(32'h39a4209d),
	.w4(32'h3822edbb),
	.w5(32'hb95e07e9),
	.w6(32'h39bc01c3),
	.w7(32'h39934870),
	.w8(32'hb91b1c26),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ac2f7a),
	.w1(32'hb82ff60c),
	.w2(32'hb956758a),
	.w3(32'hb89b2a3f),
	.w4(32'hb6ddde15),
	.w5(32'hb91d9bf7),
	.w6(32'h38a22c95),
	.w7(32'h383512dc),
	.w8(32'hb91b6b8c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c9d05),
	.w1(32'h392e743a),
	.w2(32'h38ac895f),
	.w3(32'hba220a19),
	.w4(32'hb98ea937),
	.w5(32'hb90cc4e8),
	.w6(32'hba0a0169),
	.w7(32'hb85122d8),
	.w8(32'hb933bd0e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387825ba),
	.w1(32'hb90a58f6),
	.w2(32'hba230b8d),
	.w3(32'hb982b041),
	.w4(32'hb99457f1),
	.w5(32'hba453955),
	.w6(32'hb9b5f874),
	.w7(32'hb93e2048),
	.w8(32'hb9eb000d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9929e0a),
	.w1(32'hb9445cd3),
	.w2(32'hb945514d),
	.w3(32'hb9c69aeb),
	.w4(32'hb881a626),
	.w5(32'hb8b56f38),
	.w6(32'hba101232),
	.w7(32'hb9820056),
	.w8(32'hb79e1795),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994d277),
	.w1(32'hba19567c),
	.w2(32'hba930a1d),
	.w3(32'h37a6a281),
	.w4(32'hb9dd6838),
	.w5(32'hba4cce10),
	.w6(32'h3996b54a),
	.w7(32'h375db2d3),
	.w8(32'hb9967a3e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3893760d),
	.w1(32'hb8ea8dab),
	.w2(32'hb9bfa2d7),
	.w3(32'hb75616e6),
	.w4(32'hb8b6b055),
	.w5(32'hb9b19924),
	.w6(32'h38eba3a4),
	.w7(32'h37848921),
	.w8(32'hb96a3311),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3624082c),
	.w1(32'hb5826511),
	.w2(32'h372d9259),
	.w3(32'h36eb7250),
	.w4(32'h370b1e28),
	.w5(32'h37662b33),
	.w6(32'h36f97dc1),
	.w7(32'h368e86c1),
	.w8(32'h370ff257),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374b7168),
	.w1(32'h35d16f56),
	.w2(32'h362d39df),
	.w3(32'h3745c852),
	.w4(32'hb5d31eff),
	.w5(32'hb689b0ca),
	.w6(32'h372a56bc),
	.w7(32'h363069a7),
	.w8(32'hb5bbeb73),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895486d),
	.w1(32'h382b10c3),
	.w2(32'h38a5aea8),
	.w3(32'h37259846),
	.w4(32'hb86b49a3),
	.w5(32'hb638f597),
	.w6(32'hb53e2d78),
	.w7(32'hb85bf74a),
	.w8(32'hb7ab6b46),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2c225),
	.w1(32'h3a026cf3),
	.w2(32'h39c702bc),
	.w3(32'h3a0fc836),
	.w4(32'h39aaea5c),
	.w5(32'h390beaa3),
	.w6(32'hb88ffd24),
	.w7(32'h3980fe0f),
	.w8(32'h3797a7e6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f8866),
	.w1(32'hb9940075),
	.w2(32'hb921b0c0),
	.w3(32'hba0aa777),
	.w4(32'h385b73db),
	.w5(32'h389a086f),
	.w6(32'hb8a9026f),
	.w7(32'h3a115bf2),
	.w8(32'h3a12282c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f2aa0),
	.w1(32'h3acdcddc),
	.w2(32'h3ab8673a),
	.w3(32'h3a185213),
	.w4(32'h3a681494),
	.w5(32'h3a51b194),
	.w6(32'h39bfc711),
	.w7(32'h3a1e7e81),
	.w8(32'h39cedec9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810d0a8),
	.w1(32'h37d39298),
	.w2(32'h37016618),
	.w3(32'hb6a1e7e6),
	.w4(32'hb62113dc),
	.w5(32'hb81e32b8),
	.w6(32'hb862a85a),
	.w7(32'hb7a0ae73),
	.w8(32'h37163197),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385d28b3),
	.w1(32'h362b58d2),
	.w2(32'hb7b3bd5b),
	.w3(32'h37e8eb3b),
	.w4(32'hb7e2056c),
	.w5(32'hb82a671f),
	.w6(32'h380e7b57),
	.w7(32'hb6b58108),
	.w8(32'hb7c360e0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1566e),
	.w1(32'h386824ca),
	.w2(32'hb7ffee7d),
	.w3(32'hb7dfe4f8),
	.w4(32'hb9443621),
	.w5(32'hb9b4a671),
	.w6(32'hb9e961a1),
	.w7(32'hb980ca4b),
	.w8(32'hb9b0a32c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994b823),
	.w1(32'hb8f42f11),
	.w2(32'hb9c29380),
	.w3(32'h39ccb899),
	.w4(32'hb92a206b),
	.w5(32'hba500897),
	.w6(32'h3a6b14dd),
	.w7(32'h3a52e78d),
	.w8(32'h39c4545b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba067ae1),
	.w1(32'hb93bb564),
	.w2(32'h39b9831f),
	.w3(32'hba1e21a6),
	.w4(32'hb918c40e),
	.w5(32'hb8bf7d49),
	.w6(32'hba07a889),
	.w7(32'h38c8b793),
	.w8(32'h3742e35d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37548309),
	.w1(32'hb5f0ae10),
	.w2(32'hb72ff24d),
	.w3(32'h37314bcf),
	.w4(32'hb47711fa),
	.w5(32'hb66dcc1e),
	.w6(32'hb5347e02),
	.w7(32'h3725757c),
	.w8(32'h370d35ff),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a9fe5d),
	.w1(32'hb7f5d03f),
	.w2(32'hb8656d3b),
	.w3(32'hb81c5172),
	.w4(32'h37365ad4),
	.w5(32'h3785e619),
	.w6(32'hb8182f46),
	.w7(32'h38acff63),
	.w8(32'h3820e5cd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49d351),
	.w1(32'hb9a4bbb2),
	.w2(32'hb92a9004),
	.w3(32'hba02bbfe),
	.w4(32'h37f7ff6c),
	.w5(32'hb7d6953a),
	.w6(32'hb97b7087),
	.w7(32'h39bcc100),
	.w8(32'h39bce334),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37275024),
	.w1(32'h3953e385),
	.w2(32'h39abc048),
	.w3(32'hb863bc8f),
	.w4(32'h38302cc6),
	.w5(32'h3953a66d),
	.w6(32'hb959ecde),
	.w7(32'hb832d7c6),
	.w8(32'h36d92aaf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb832ce57),
	.w1(32'hb82b3abc),
	.w2(32'hb875b191),
	.w3(32'h3835c903),
	.w4(32'h3801ed58),
	.w5(32'h3546fa23),
	.w6(32'hb786cd42),
	.w7(32'hb85f8442),
	.w8(32'hb815dac7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37863471),
	.w1(32'h3836bd25),
	.w2(32'hb7548100),
	.w3(32'h38d1c916),
	.w4(32'hb7aa8819),
	.w5(32'hb828ed5a),
	.w6(32'h3931e974),
	.w7(32'h38f82721),
	.w8(32'hb59d03c0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbafca),
	.w1(32'hb9ea960a),
	.w2(32'hb8fad1b9),
	.w3(32'h38ef3d4d),
	.w4(32'hba53e504),
	.w5(32'h3979db6c),
	.w6(32'h3a46b1fc),
	.w7(32'h394958d4),
	.w8(32'h3a0350b5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f0cfb),
	.w1(32'hba5d45f6),
	.w2(32'hb9706697),
	.w3(32'hb9cd6903),
	.w4(32'hba2443d6),
	.w5(32'hba549524),
	.w6(32'h399e93f5),
	.w7(32'h39daac5a),
	.w8(32'h3a0cfbdb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaab16),
	.w1(32'h3a871b3a),
	.w2(32'h399bda1d),
	.w3(32'h3a930da7),
	.w4(32'hb91231b6),
	.w5(32'hba8dc399),
	.w6(32'h3a189678),
	.w7(32'hba09f433),
	.w8(32'hba9b65b8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ccaab),
	.w1(32'h386b53bd),
	.w2(32'h38c6a5c9),
	.w3(32'h37d68573),
	.w4(32'h376be50e),
	.w5(32'h38a0b1cc),
	.w6(32'h3887c62c),
	.w7(32'h37e6b0e1),
	.w8(32'h38b0335f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885fc5d),
	.w1(32'hb5e1cc5b),
	.w2(32'hb7253964),
	.w3(32'hb8a56251),
	.w4(32'hb6a0c267),
	.w5(32'h3465bd8a),
	.w6(32'hb33b2818),
	.w7(32'hb63b6fd4),
	.w8(32'h38343697),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384cb5ee),
	.w1(32'h383f594b),
	.w2(32'h388c3bf0),
	.w3(32'hb884ebde),
	.w4(32'hb5b7b177),
	.w5(32'h388360fc),
	.w6(32'hb9288588),
	.w7(32'hb76ef6d9),
	.w8(32'h3851ec8c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914a711),
	.w1(32'hb770519b),
	.w2(32'hb7e69402),
	.w3(32'h37d557f1),
	.w4(32'hb8816dcd),
	.w5(32'hb6ca8fab),
	.w6(32'h37e3557d),
	.w7(32'hb6ddedb0),
	.w8(32'h3849e5ae),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa54f03),
	.w1(32'h38869edd),
	.w2(32'hb9a71f33),
	.w3(32'hba672757),
	.w4(32'h38f33a67),
	.w5(32'h381d9287),
	.w6(32'h39a24b17),
	.w7(32'h3a9e5e43),
	.w8(32'h3a7d2077),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba319109),
	.w1(32'hb978d027),
	.w2(32'h396f35e7),
	.w3(32'hba5493e7),
	.w4(32'hb942fd20),
	.w5(32'h398ac809),
	.w6(32'hba2ede97),
	.w7(32'h38b90729),
	.w8(32'h39eafff7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3863a90e),
	.w1(32'h3a0f3fce),
	.w2(32'h3a56997d),
	.w3(32'hb827899a),
	.w4(32'h39c70fc9),
	.w5(32'h3a0f5518),
	.w6(32'h38957f85),
	.w7(32'h39d6ea88),
	.w8(32'h3a050c34),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf2e80),
	.w1(32'hb9d59bca),
	.w2(32'h39378bf2),
	.w3(32'hbaaddbdb),
	.w4(32'hb9ccbe50),
	.w5(32'h3992fa88),
	.w6(32'hba84333c),
	.w7(32'hb996be6c),
	.w8(32'h39f0c946),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9c34d),
	.w1(32'hb89c466b),
	.w2(32'hba440859),
	.w3(32'h3a251be0),
	.w4(32'hb928ca6f),
	.w5(32'hba6a9271),
	.w6(32'h3a819d7b),
	.w7(32'h38d803f9),
	.w8(32'hb9f44123),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39898360),
	.w1(32'h3a02af74),
	.w2(32'h39eadd67),
	.w3(32'h39a722da),
	.w4(32'h3a035273),
	.w5(32'h39fb82f9),
	.w6(32'h39aca363),
	.w7(32'h39e2ee8d),
	.w8(32'h399e8592),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a547b2b),
	.w1(32'h3a89874a),
	.w2(32'h3a60172b),
	.w3(32'h3a480cb6),
	.w4(32'h3a51b15e),
	.w5(32'h3a765726),
	.w6(32'h3975a62a),
	.w7(32'h396d1945),
	.w8(32'h39b70ee0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ccc32),
	.w1(32'h3a102d0c),
	.w2(32'h39bb5346),
	.w3(32'h3a2cd13b),
	.w4(32'h39e70326),
	.w5(32'h39649523),
	.w6(32'h3a3c686c),
	.w7(32'h3a311d5f),
	.w8(32'h39b9595e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb872acf0),
	.w1(32'hb93a73fb),
	.w2(32'hb950c2e4),
	.w3(32'h35482e84),
	.w4(32'hb8eb1275),
	.w5(32'hb908f18c),
	.w6(32'h36cf41c5),
	.w7(32'h38e414b0),
	.w8(32'h3777c610),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391aaa0c),
	.w1(32'h38a555fa),
	.w2(32'hb7c7b488),
	.w3(32'h38fbf280),
	.w4(32'h372837d8),
	.w5(32'hb78bd620),
	.w6(32'hb82facfd),
	.w7(32'hb8e62218),
	.w8(32'hb902b3dc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e49f7c),
	.w1(32'hb9fce25a),
	.w2(32'hba850ac8),
	.w3(32'h396cc0eb),
	.w4(32'hb90acd01),
	.w5(32'hba341ce7),
	.w6(32'h39c6680f),
	.w7(32'h38b6565d),
	.w8(32'hb9a21f99),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f66659),
	.w1(32'hb895b4f8),
	.w2(32'hb91ec905),
	.w3(32'hb8dbf07a),
	.w4(32'hb884e6dc),
	.w5(32'hb9188193),
	.w6(32'h38a200d7),
	.w7(32'h38ec589e),
	.w8(32'h378712e7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372558c0),
	.w1(32'h37a659eb),
	.w2(32'h370aca65),
	.w3(32'h362a6251),
	.w4(32'h36d86eef),
	.w5(32'hb6ff1831),
	.w6(32'h37849d1c),
	.w7(32'h36d3ae84),
	.w8(32'h3663a9a0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360fc1f1),
	.w1(32'h36e2abc9),
	.w2(32'h350d951b),
	.w3(32'h36175c81),
	.w4(32'hb4e655cc),
	.w5(32'h350df51e),
	.w6(32'h37226105),
	.w7(32'h361b0ab2),
	.w8(32'h3624f24e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f715a4),
	.w1(32'h38678718),
	.w2(32'h38852578),
	.w3(32'h3723b9d9),
	.w4(32'hb604b095),
	.w5(32'hb53da0b8),
	.w6(32'h38203b92),
	.w7(32'hb60b18a7),
	.w8(32'hb79a0e6d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9506d45),
	.w1(32'hb953dde5),
	.w2(32'hb90e49c5),
	.w3(32'hb90020dd),
	.w4(32'hb8f2ee77),
	.w5(32'hb8f73923),
	.w6(32'hb9a074a2),
	.w7(32'hb9903449),
	.w8(32'hb9483a31),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d5ce9),
	.w1(32'hb88b7ad8),
	.w2(32'hb873888c),
	.w3(32'hb90fe6d6),
	.w4(32'hb7df1b60),
	.w5(32'h3616ebe8),
	.w6(32'hb78ed8c3),
	.w7(32'hb7d1c80c),
	.w8(32'h386cbac5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c7822),
	.w1(32'hb8c01fed),
	.w2(32'hb9844b3f),
	.w3(32'hb7f5b073),
	.w4(32'hb8798e0a),
	.w5(32'hb96e494f),
	.w6(32'h38dd1928),
	.w7(32'h38a8f7e1),
	.w8(32'hb93e3d14),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9865b69),
	.w1(32'hb987a143),
	.w2(32'hb9ad9f59),
	.w3(32'hb9bd8146),
	.w4(32'hb96d77e2),
	.w5(32'hb98857be),
	.w6(32'hb9c26e7b),
	.w7(32'hb9278848),
	.w8(32'hb983e010),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381d5f9c),
	.w1(32'h38021e63),
	.w2(32'h37b5f57b),
	.w3(32'h38045240),
	.w4(32'h380352cb),
	.w5(32'h37e02a0b),
	.w6(32'h38144d77),
	.w7(32'h379c2ec0),
	.w8(32'h3799ca1b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b693f2),
	.w1(32'hb6904d96),
	.w2(32'h359b8e6a),
	.w3(32'hb66f6767),
	.w4(32'hb5d6b895),
	.w5(32'h367ffd0d),
	.w6(32'hb6c43b79),
	.w7(32'hb6ad35f6),
	.w8(32'hb70718cf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926f4ba),
	.w1(32'h3919481d),
	.w2(32'h38fe4c4e),
	.w3(32'h3902112b),
	.w4(32'h38b0eb7d),
	.w5(32'h37ec7302),
	.w6(32'h381286bb),
	.w7(32'h37f7ded8),
	.w8(32'hb80308e5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7948caa),
	.w1(32'hb6bdad81),
	.w2(32'hb661bdd3),
	.w3(32'hb72fea49),
	.w4(32'hb5383e1a),
	.w5(32'hb60fc0c2),
	.w6(32'hb64127ae),
	.w7(32'hb56a1ff7),
	.w8(32'hb6bbe042),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a5d39),
	.w1(32'hb98b0523),
	.w2(32'hba9dd99f),
	.w3(32'h39b25908),
	.w4(32'hb8a3c42b),
	.w5(32'hba5747dc),
	.w6(32'hb793df6c),
	.w7(32'hb9a895f0),
	.w8(32'hba486487),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d2e44),
	.w1(32'h3908305d),
	.w2(32'hb95042d5),
	.w3(32'h39734288),
	.w4(32'h38399462),
	.w5(32'hb9a2c2fe),
	.w6(32'h39eb4479),
	.w7(32'h39a8d015),
	.w8(32'hb600b9da),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990485a),
	.w1(32'h39d3ebcb),
	.w2(32'h39497363),
	.w3(32'h38a39f6c),
	.w4(32'h3949a975),
	.w5(32'h38e09d2d),
	.w6(32'h389f1ff5),
	.w7(32'h39b51b1c),
	.w8(32'h383a48c9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379908e3),
	.w1(32'h39bf43a4),
	.w2(32'h3a4b7812),
	.w3(32'hb91f538b),
	.w4(32'h39820fd8),
	.w5(32'h3a0f14a5),
	.w6(32'h37e97ecd),
	.w7(32'h39e54110),
	.w8(32'h39e4d19c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37566831),
	.w1(32'h36dd9aaf),
	.w2(32'h36abb60d),
	.w3(32'h372f35ce),
	.w4(32'h36acf1f2),
	.w5(32'h36f67878),
	.w6(32'h37015520),
	.w7(32'hb20a30cc),
	.w8(32'hb5d40448),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c14afe),
	.w1(32'h370f3cd8),
	.w2(32'h36aaaf8c),
	.w3(32'h379f35c0),
	.w4(32'h3690c46f),
	.w5(32'h36731698),
	.w6(32'h37122123),
	.w7(32'hb63229ff),
	.w8(32'hb655d0b3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b5857),
	.w1(32'h366bacaa),
	.w2(32'h379ce78f),
	.w3(32'h36ea3dde),
	.w4(32'h36116d92),
	.w5(32'hb69ed696),
	.w6(32'h371f4781),
	.w7(32'hb78bedfc),
	.w8(32'hb7736a8d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe9805),
	.w1(32'hb96639fa),
	.w2(32'hb9b3862d),
	.w3(32'hb940d97b),
	.w4(32'hb91971ac),
	.w5(32'hb96ce62b),
	.w6(32'hb7e6792b),
	.w7(32'hb867a528),
	.w8(32'hb92436b0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b59dd2),
	.w1(32'h385a7305),
	.w2(32'h387ba9ab),
	.w3(32'hb5eba51c),
	.w4(32'h380a6ddb),
	.w5(32'h384022a6),
	.w6(32'hb8452592),
	.w7(32'h377b8cc8),
	.w8(32'h381e15c6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a986f),
	.w1(32'hb981725d),
	.w2(32'hb9d352e6),
	.w3(32'h38cb7ce5),
	.w4(32'hb8500c9e),
	.w5(32'hb9556aa9),
	.w6(32'h3955e7bd),
	.w7(32'hb88df96e),
	.w8(32'hb8998879),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37948316),
	.w1(32'hb955e004),
	.w2(32'hba024291),
	.w3(32'h3946c5c7),
	.w4(32'hb8b04e85),
	.w5(32'hb98e656e),
	.w6(32'h39fe993f),
	.w7(32'h38dadd32),
	.w8(32'hb908118c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f22c75),
	.w1(32'h391f0c23),
	.w2(32'h390ad149),
	.w3(32'h3824bdb3),
	.w4(32'h38a5dc60),
	.w5(32'hb885bda0),
	.w6(32'h391a6060),
	.w7(32'h3912d6d7),
	.w8(32'h376d0eac),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902c2d1),
	.w1(32'hb8866203),
	.w2(32'hb99f4616),
	.w3(32'h37f4f1fd),
	.w4(32'hb857da63),
	.w5(32'hb976df24),
	.w6(32'h39426d67),
	.w7(32'h393a86b5),
	.w8(32'hb6f9ca15),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378de5e8),
	.w1(32'hb894e0f6),
	.w2(32'hb9ca3a6c),
	.w3(32'h395e449a),
	.w4(32'h38edac49),
	.w5(32'hb8f84803),
	.w6(32'h390ae527),
	.w7(32'hb89dc67d),
	.w8(32'hb8fb72c0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2532f5),
	.w1(32'hb9d8d8a6),
	.w2(32'hb9a3add0),
	.w3(32'hba2f5ab4),
	.w4(32'hb9c0bab1),
	.w5(32'hb998aa77),
	.w6(32'hb9dd354a),
	.w7(32'h381766bb),
	.w8(32'h3840f6a0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e3b1c),
	.w1(32'hb964cfdf),
	.w2(32'hb9da8994),
	.w3(32'hb7a38172),
	.w4(32'hb88600ca),
	.w5(32'hb998cfb8),
	.w6(32'h38b6d912),
	.w7(32'h379ac471),
	.w8(32'hb91c033c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3584eec),
	.w1(32'h3663e18a),
	.w2(32'h36985a7e),
	.w3(32'h34b7db84),
	.w4(32'h3675aae0),
	.w5(32'h369f3953),
	.w6(32'h36ab3acb),
	.w7(32'h36869f02),
	.w8(32'h36e06965),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37349c2a),
	.w1(32'hb6a0beb8),
	.w2(32'hb70eebcf),
	.w3(32'h3728aff8),
	.w4(32'hb67833c6),
	.w5(32'hb7365dfd),
	.w6(32'h362d8581),
	.w7(32'hb632164c),
	.w8(32'hb7067ed9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb684da40),
	.w1(32'h373887e3),
	.w2(32'h36878d8d),
	.w3(32'hb6846ee0),
	.w4(32'h370cc88f),
	.w5(32'hb5646a4d),
	.w6(32'h3764ec25),
	.w7(32'h36c0fc1a),
	.w8(32'hb68fa021),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373b3b94),
	.w1(32'h37f6abb7),
	.w2(32'h3822d218),
	.w3(32'h376488ca),
	.w4(32'h37ba4eef),
	.w5(32'h37d7e78d),
	.w6(32'h37aa9d39),
	.w7(32'h3575baa9),
	.w8(32'h37795143),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a037af),
	.w1(32'hb814a3a1),
	.w2(32'h39890664),
	.w3(32'hb99988e7),
	.w4(32'hb6f57c88),
	.w5(32'h39795725),
	.w6(32'hb8d3e452),
	.w7(32'h38a49226),
	.w8(32'h39530f39),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d7a266),
	.w1(32'h358b0bb5),
	.w2(32'h382d346e),
	.w3(32'h36d3e5f0),
	.w4(32'hb8043a50),
	.w5(32'hb7631fcd),
	.w6(32'hb739989d),
	.w7(32'hb8903884),
	.w8(32'hb8458637),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6aca1),
	.w1(32'hb4e2e303),
	.w2(32'h38d2ba58),
	.w3(32'h38810877),
	.w4(32'h37b1187d),
	.w5(32'h37973a6e),
	.w6(32'h39870865),
	.w7(32'h3947afbc),
	.w8(32'h396211b4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db8bcc),
	.w1(32'h38f46ebd),
	.w2(32'hb90942a2),
	.w3(32'h398ac76c),
	.w4(32'hb7c8789a),
	.w5(32'hb974af9f),
	.w6(32'h39658f70),
	.w7(32'hb8b9f993),
	.w8(32'hb96fb510),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a65483),
	.w1(32'h39c3676f),
	.w2(32'h39cd52f3),
	.w3(32'h398b1a60),
	.w4(32'h39431d7a),
	.w5(32'h397ced20),
	.w6(32'h364d97c5),
	.w7(32'hb871e0b3),
	.w8(32'h38867152),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8daa44b),
	.w1(32'hb9c6b3a0),
	.w2(32'hba1167e0),
	.w3(32'h3814ad4a),
	.w4(32'hb8ae25a8),
	.w5(32'hb8ed0453),
	.w6(32'h39785f08),
	.w7(32'h3986d558),
	.w8(32'h36bb2006),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cb48d),
	.w1(32'hb915bcd3),
	.w2(32'hb8df4656),
	.w3(32'hb933cc44),
	.w4(32'hb8cab17c),
	.w5(32'hb93c2c14),
	.w6(32'hb9827688),
	.w7(32'h378d5dc7),
	.w8(32'h3903d340),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a149410),
	.w1(32'h3a14ec3d),
	.w2(32'hb8087723),
	.w3(32'h39be088a),
	.w4(32'h399d7ad3),
	.w5(32'hb8bfb828),
	.w6(32'h39c6c7fc),
	.w7(32'h3907e107),
	.w8(32'hb919dbfe),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf1f7c),
	.w1(32'h399de0e2),
	.w2(32'h388261a0),
	.w3(32'h397dcba1),
	.w4(32'h398be38a),
	.w5(32'h388f0623),
	.w6(32'h398f141d),
	.w7(32'h398b9a13),
	.w8(32'h38983102),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84ebc19),
	.w1(32'h383deb83),
	.w2(32'h395a7092),
	.w3(32'hb91d2ddb),
	.w4(32'h38e20895),
	.w5(32'h39a7928c),
	.w6(32'hb99b2da7),
	.w7(32'hb8d9b2c9),
	.w8(32'h39004d14),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a406082),
	.w1(32'h3a87a436),
	.w2(32'h3a434af6),
	.w3(32'h3a5f85d9),
	.w4(32'h3a94ad3c),
	.w5(32'h3a8a8a88),
	.w6(32'h3a3a6746),
	.w7(32'h3a6db615),
	.w8(32'h3a2020ad),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea91b5),
	.w1(32'h3b061f83),
	.w2(32'h3ab85fa1),
	.w3(32'h3acb88d6),
	.w4(32'h3aab67cb),
	.w5(32'h3add2999),
	.w6(32'h3a014c78),
	.w7(32'h3a099fbf),
	.w8(32'h3a6b96c0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2405e9),
	.w1(32'h3a6c565d),
	.w2(32'h3a6f28b5),
	.w3(32'h3a40d680),
	.w4(32'h3a3a7345),
	.w5(32'h3a6194a0),
	.w6(32'hba2983f5),
	.w7(32'hba46007e),
	.w8(32'hba334bd0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b10c3a),
	.w1(32'h38c83d61),
	.w2(32'h398cd236),
	.w3(32'h395a1306),
	.w4(32'hb9105eaf),
	.w5(32'h39583ee9),
	.w6(32'h39c16124),
	.w7(32'h39c2ac4b),
	.w8(32'h39a5b06b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a94d2),
	.w1(32'h392fcc5f),
	.w2(32'h3a94dee8),
	.w3(32'hb8d40ae6),
	.w4(32'h39d21cef),
	.w5(32'h3a85cd71),
	.w6(32'hbad51e09),
	.w7(32'hbab37128),
	.w8(32'hba197473),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2e79d),
	.w1(32'h3ac307c5),
	.w2(32'h3acb8e30),
	.w3(32'h3a71b3df),
	.w4(32'h3a0d32c1),
	.w5(32'h3a72c75f),
	.w6(32'h399a562d),
	.w7(32'h3a246940),
	.w8(32'h3a60dff2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bbb3b),
	.w1(32'hb8ee60cd),
	.w2(32'hb8ec200a),
	.w3(32'h38443ae5),
	.w4(32'h39de72af),
	.w5(32'h39942cbc),
	.w6(32'h39f1529f),
	.w7(32'h39efc355),
	.w8(32'h39d16431),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391cf032),
	.w1(32'h3a14b974),
	.w2(32'h3a1651e0),
	.w3(32'h39099283),
	.w4(32'h3a478268),
	.w5(32'h3a1da3aa),
	.w6(32'h3983211a),
	.w7(32'h358184e0),
	.w8(32'hb979c7cf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbfb4a),
	.w1(32'h39386297),
	.w2(32'h36e9415e),
	.w3(32'h39d2d6a3),
	.w4(32'h390dffcf),
	.w5(32'h39af65b5),
	.w6(32'h3a469ba0),
	.w7(32'h39dd07d8),
	.w8(32'h3990a576),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9510ae0),
	.w1(32'h38b03f87),
	.w2(32'h39c95b52),
	.w3(32'hb8ddf36c),
	.w4(32'h398895ce),
	.w5(32'h39ee2663),
	.w6(32'h38de7970),
	.w7(32'h39fe8b69),
	.w8(32'h39f3bc66),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901999f),
	.w1(32'hb8db4800),
	.w2(32'hb8c76ecc),
	.w3(32'hb8ab4ea5),
	.w4(32'hb8997dcb),
	.w5(32'hb8607bfc),
	.w6(32'hb904437b),
	.w7(32'hb89300c9),
	.w8(32'hb82eef7d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d5ed3),
	.w1(32'h394c08f4),
	.w2(32'h38c9fb4c),
	.w3(32'h3962b00b),
	.w4(32'h391e2c97),
	.w5(32'h382b8649),
	.w6(32'h38877e7a),
	.w7(32'hb8d18e10),
	.w8(32'hb9188134),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8521e5),
	.w1(32'h3a8aa86a),
	.w2(32'h3a8bcbe0),
	.w3(32'h3a993d13),
	.w4(32'h3a01076d),
	.w5(32'h3a158d6c),
	.w6(32'h3a6dc710),
	.w7(32'h39b560ab),
	.w8(32'h399610e4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06db7c),
	.w1(32'h3b137ba5),
	.w2(32'h3afc51cf),
	.w3(32'h3ad60469),
	.w4(32'h3a9f44cd),
	.w5(32'h3a9a6481),
	.w6(32'h3a7e622c),
	.w7(32'h3a2381a3),
	.w8(32'h3a0038a9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80d3bd5),
	.w1(32'hb78b6a26),
	.w2(32'h376cb807),
	.w3(32'h381383f0),
	.w4(32'h38018138),
	.w5(32'h380db8ed),
	.w6(32'hb8e6cb58),
	.w7(32'hb9146865),
	.w8(32'hb9574ad9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f0f365),
	.w1(32'h39c1530d),
	.w2(32'h39f2d797),
	.w3(32'h38ceff19),
	.w4(32'h39c9ab0c),
	.w5(32'h39ce02d9),
	.w6(32'h398d3c92),
	.w7(32'h398a4788),
	.w8(32'h3965f58c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c7265),
	.w1(32'hb88c9563),
	.w2(32'hb906b9bc),
	.w3(32'hb7e5f1e6),
	.w4(32'hb85bd0eb),
	.w5(32'hb90ae84b),
	.w6(32'h39cee0fa),
	.w7(32'h39c2362d),
	.w8(32'h394bbaaa),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba099263),
	.w1(32'hba2c90a3),
	.w2(32'hba95fdb3),
	.w3(32'hb9b1a6c3),
	.w4(32'hb9c60469),
	.w5(32'hba6dd151),
	.w6(32'hb78ab851),
	.w7(32'hb9e967a4),
	.w8(32'hba1032b0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87f75c1),
	.w1(32'h395864fb),
	.w2(32'h39859dc9),
	.w3(32'hb88e58cc),
	.w4(32'h39442731),
	.w5(32'h39528a25),
	.w6(32'hb85fe948),
	.w7(32'h39320e62),
	.w8(32'h395955d4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d22285),
	.w1(32'hb8377eab),
	.w2(32'hb8175d0e),
	.w3(32'hb8609d94),
	.w4(32'hb8073aad),
	.w5(32'hb670abb1),
	.w6(32'hb7c36828),
	.w7(32'h37596502),
	.w8(32'h3799d59a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380645fd),
	.w1(32'hb77625f8),
	.w2(32'hb82bab15),
	.w3(32'h370c1041),
	.w4(32'hb7b9be9f),
	.w5(32'hb864b340),
	.w6(32'h37326783),
	.w7(32'hb7a580a1),
	.w8(32'hb8a7835b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b0478b),
	.w1(32'hb610e8c4),
	.w2(32'hb6dde57c),
	.w3(32'h357245eb),
	.w4(32'h36a6ec94),
	.w5(32'h35faac59),
	.w6(32'h35f0ccc2),
	.w7(32'h363b286b),
	.w8(32'h34ac4156),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60f7433),
	.w1(32'h372bfdce),
	.w2(32'hb735eff5),
	.w3(32'hb7b06a67),
	.w4(32'hb70d4bc1),
	.w5(32'hb6f1f0ce),
	.w6(32'h3782be53),
	.w7(32'h370fff51),
	.w8(32'h38152a63),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b64b6f),
	.w1(32'hb93b311f),
	.w2(32'hb9012fbe),
	.w3(32'hb9c14ae6),
	.w4(32'hb8945c6d),
	.w5(32'hb8d0e2b1),
	.w6(32'hb96590fe),
	.w7(32'h395e3234),
	.w8(32'h394cac4c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9532775),
	.w1(32'hb923517b),
	.w2(32'hb7493323),
	.w3(32'hb95032f1),
	.w4(32'hb8466cca),
	.w5(32'h37bcebbc),
	.w6(32'hb91b4edc),
	.w7(32'h377e9d67),
	.w8(32'h388a766f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378aaad1),
	.w1(32'hb6195826),
	.w2(32'hb91138ff),
	.w3(32'h39280e9e),
	.w4(32'h38c2054c),
	.w5(32'hb8479d40),
	.w6(32'h39806228),
	.w7(32'h38e4c4de),
	.w8(32'h38225821),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3774fce4),
	.w1(32'h394ec905),
	.w2(32'h39a93d7a),
	.w3(32'h3874a39b),
	.w4(32'h393f3bd2),
	.w5(32'h38efb5c7),
	.w6(32'h38ebddf4),
	.w7(32'h3811b6c7),
	.w8(32'hb8c445b4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33bac3f8),
	.w1(32'hb5692845),
	.w2(32'hb6930957),
	.w3(32'hb4fee127),
	.w4(32'hb7118c39),
	.w5(32'hb730ff2a),
	.w6(32'h36d4b812),
	.w7(32'hb5369583),
	.w8(32'hb693fc81),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fba48d),
	.w1(32'h37ebd334),
	.w2(32'h386301b1),
	.w3(32'h35aaeadc),
	.w4(32'h37e28280),
	.w5(32'h38815f78),
	.w6(32'h37098347),
	.w7(32'h37092ba2),
	.w8(32'h38347c02),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377b3fa1),
	.w1(32'hb725376e),
	.w2(32'hb708d27b),
	.w3(32'h37aa08f9),
	.w4(32'h366b7bf6),
	.w5(32'hb79900fa),
	.w6(32'hb842299d),
	.w7(32'hb7981be4),
	.w8(32'hb674cfea),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f4b649),
	.w1(32'hb7be2bd5),
	.w2(32'h375e605e),
	.w3(32'h389680ad),
	.w4(32'h3780abb8),
	.w5(32'h37ea6585),
	.w6(32'h389b2fdf),
	.w7(32'h36fae9bc),
	.w8(32'h38705a70),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f0580),
	.w1(32'h38f95fb5),
	.w2(32'hb90bc628),
	.w3(32'h39b3fd4b),
	.w4(32'h38644ab9),
	.w5(32'hb9445880),
	.w6(32'h3a21fd84),
	.w7(32'h398dfbd9),
	.w8(32'hb8b6fcea),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81bd69b),
	.w1(32'hb9b22710),
	.w2(32'hba51443e),
	.w3(32'hb7907eaa),
	.w4(32'hb8b49c91),
	.w5(32'hba004e05),
	.w6(32'hb8c1abf1),
	.w7(32'hb954b703),
	.w8(32'hb9fc7c0f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37954f13),
	.w1(32'hb7961b92),
	.w2(32'hb840600c),
	.w3(32'h380ff9a5),
	.w4(32'h36ace7df),
	.w5(32'hb7aa0d30),
	.w6(32'h3828902c),
	.w7(32'h3766991c),
	.w8(32'hb7edebbd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937e555),
	.w1(32'hb9834a48),
	.w2(32'hb9b6fefb),
	.w3(32'hb9885f53),
	.w4(32'hb8363dc9),
	.w5(32'hb9451e10),
	.w6(32'h38717c40),
	.w7(32'h37c60322),
	.w8(32'hb8325437),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372428f8),
	.w1(32'h38519919),
	.w2(32'h3865b3f9),
	.w3(32'h36250ce5),
	.w4(32'h37ed797f),
	.w5(32'h38471d90),
	.w6(32'hb6d10b5c),
	.w7(32'h38126845),
	.w8(32'h3814fb64),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39671e05),
	.w1(32'h38ed8a21),
	.w2(32'hb748dbc2),
	.w3(32'hb7187f80),
	.w4(32'hb74ebdac),
	.w5(32'hb8440828),
	.w6(32'h38a78ee1),
	.w7(32'h38223fb3),
	.w8(32'hb863adb1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ebba6f),
	.w1(32'hb85fede2),
	.w2(32'hb8dd7246),
	.w3(32'h37ea8f43),
	.w4(32'h37ba740f),
	.w5(32'hb8c43428),
	.w6(32'h37e06c84),
	.w7(32'h38df85e9),
	.w8(32'hb7884697),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987255e),
	.w1(32'hb9d1d6cb),
	.w2(32'hba5e46c2),
	.w3(32'h3921b8db),
	.w4(32'hb881de33),
	.w5(32'hb9f76481),
	.w6(32'h395d25a6),
	.w7(32'hb666f296),
	.w8(32'hb95bae40),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82dfc14),
	.w1(32'h38875ca2),
	.w2(32'h395758e1),
	.w3(32'hb82372bb),
	.w4(32'h37f9e8cb),
	.w5(32'h38d5023a),
	.w6(32'hb78992bf),
	.w7(32'h38751410),
	.w8(32'h3926c1df),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397983f2),
	.w1(32'h398b1f3f),
	.w2(32'h3987ab81),
	.w3(32'h39ba7c2e),
	.w4(32'h3912983c),
	.w5(32'h38999d20),
	.w6(32'h398d7cac),
	.w7(32'h392f0aa8),
	.w8(32'h36d4f89c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d85024),
	.w1(32'hb934bb14),
	.w2(32'hb9c682eb),
	.w3(32'h3907d18a),
	.w4(32'h3941ccc9),
	.w5(32'hb92676a5),
	.w6(32'h39889b27),
	.w7(32'h398745e0),
	.w8(32'hb7eaf57f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8772c80),
	.w1(32'h35d711db),
	.w2(32'h3908af95),
	.w3(32'hb6eb0ae9),
	.w4(32'h3820337d),
	.w5(32'h3945794a),
	.w6(32'h3748cce3),
	.w7(32'h38a3f1ba),
	.w8(32'h397905ff),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a552a3),
	.w1(32'hb95e7bc1),
	.w2(32'hb9b1c04c),
	.w3(32'hb945247b),
	.w4(32'hb66e7fcc),
	.w5(32'hb925fd00),
	.w6(32'hb7686db3),
	.w7(32'hb760a2a6),
	.w8(32'hb9392568),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5d522),
	.w1(32'h37f79034),
	.w2(32'h38c785c7),
	.w3(32'hb72e62f6),
	.w4(32'h38905ed3),
	.w5(32'h38ba465d),
	.w6(32'h33385534),
	.w7(32'h38b9a074),
	.w8(32'h38d3f330),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b90345),
	.w1(32'h39a85eb3),
	.w2(32'h39dd52b4),
	.w3(32'h3939b34e),
	.w4(32'h388f6df8),
	.w5(32'hb9180ed2),
	.w6(32'h37b8f7e3),
	.w7(32'hb91cd41c),
	.w8(32'hb95d37e2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38045036),
	.w1(32'h37eacbbe),
	.w2(32'h386099c7),
	.w3(32'h38d3d67c),
	.w4(32'h38b12426),
	.w5(32'h38bed5df),
	.w6(32'h39224c5d),
	.w7(32'h39048ee1),
	.w8(32'h38cd1dff),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e8d95a),
	.w1(32'hb6d8fc76),
	.w2(32'hb7249ad4),
	.w3(32'h371ce798),
	.w4(32'hb6369fd9),
	.w5(32'hb6ee2c8e),
	.w6(32'h373a8491),
	.w7(32'h366ea895),
	.w8(32'hb70be5f6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374387f2),
	.w1(32'h373edda0),
	.w2(32'h375347b0),
	.w3(32'h373d60ec),
	.w4(32'h36ff7320),
	.w5(32'h371c467d),
	.w6(32'h3793b80e),
	.w7(32'h37423b71),
	.w8(32'hb5ee36d4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76a005c),
	.w1(32'hb7a37340),
	.w2(32'hb7738ba8),
	.w3(32'h38044fc3),
	.w4(32'h35b47514),
	.w5(32'h3758ca25),
	.w6(32'h38563ee4),
	.w7(32'h3759a21d),
	.w8(32'h37c247bf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916c2ad),
	.w1(32'h396d56a0),
	.w2(32'h39929de0),
	.w3(32'h3920e414),
	.w4(32'h3905b37f),
	.w5(32'h39789553),
	.w6(32'h39b32989),
	.w7(32'h393bc0ab),
	.w8(32'h3983d48d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0517c),
	.w1(32'hb8eebfb3),
	.w2(32'hb99ee9a2),
	.w3(32'h374f720b),
	.w4(32'hb885a4e6),
	.w5(32'hb9ade2d9),
	.w6(32'h39583b52),
	.w7(32'h3928d848),
	.w8(32'hb930ea67),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb613499a),
	.w1(32'h36b658e3),
	.w2(32'h36f5c18c),
	.w3(32'hb6d8aef1),
	.w4(32'hb4ce2d89),
	.w5(32'h35de112a),
	.w6(32'hb6a9b594),
	.w7(32'h35f3b65b),
	.w8(32'hb688d15f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943510b),
	.w1(32'hb629aedc),
	.w2(32'hb983fd43),
	.w3(32'hb9536437),
	.w4(32'hb8dbbacc),
	.w5(32'hb968b373),
	.w6(32'hb916835d),
	.w7(32'hb738dca9),
	.w8(32'hb8ae04d7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89e1e9),
	.w1(32'h3a8e0a4d),
	.w2(32'h3a40b6af),
	.w3(32'h3a1b295e),
	.w4(32'h39b00b26),
	.w5(32'h386ff744),
	.w6(32'h3a1531ce),
	.w7(32'h399af738),
	.w8(32'h37bcfae4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17205e),
	.w1(32'hba1552c0),
	.w2(32'hba1c1aa6),
	.w3(32'hb91e0b43),
	.w4(32'hb8aa3ca2),
	.w5(32'hb9fccbec),
	.w6(32'h380bac55),
	.w7(32'hb8da8a94),
	.w8(32'hb9bc342e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c5769),
	.w1(32'h3992375c),
	.w2(32'h39f03bfa),
	.w3(32'hb9425ef4),
	.w4(32'h384287de),
	.w5(32'h37985abd),
	.w6(32'hb89b2c19),
	.w7(32'h3819e836),
	.w8(32'hb8c34c9e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1affe2),
	.w1(32'h3a30b225),
	.w2(32'h3a17de11),
	.w3(32'h3a183536),
	.w4(32'h3a128ea5),
	.w5(32'h3a021cd0),
	.w6(32'h398a6afc),
	.w7(32'h387c630d),
	.w8(32'hb8fa9054),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a012c),
	.w1(32'h3a185b3a),
	.w2(32'h39ea2c8a),
	.w3(32'h3ac6fb9e),
	.w4(32'h3ab3938e),
	.w5(32'h3a888e0c),
	.w6(32'h3add2651),
	.w7(32'h3a366b41),
	.w8(32'h39a12de7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab39fa),
	.w1(32'hba005dc4),
	.w2(32'h396203e8),
	.w3(32'hbaa79ce3),
	.w4(32'hb9c9b827),
	.w5(32'h38950123),
	.w6(32'hba4bf996),
	.w7(32'hb83c3fac),
	.w8(32'h3986768c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bd119c),
	.w1(32'h38d34484),
	.w2(32'h39bedbb0),
	.w3(32'h389927fb),
	.w4(32'h38d4ca30),
	.w5(32'h39b29d35),
	.w6(32'h380c17b0),
	.w7(32'h3903e2a3),
	.w8(32'h3973d67c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940369e),
	.w1(32'h3935c531),
	.w2(32'h3933d524),
	.w3(32'h38b06820),
	.w4(32'h36c9f6f5),
	.w5(32'h384809aa),
	.w6(32'hb6c5288b),
	.w7(32'hb750f0b7),
	.w8(32'h38578328),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e48f67),
	.w1(32'hb81041b6),
	.w2(32'hb8c54874),
	.w3(32'hb635a406),
	.w4(32'h35c8940a),
	.w5(32'hb8249d60),
	.w6(32'h3831909b),
	.w7(32'h38200bdc),
	.w8(32'hb7861b7a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3685074c),
	.w1(32'h378df486),
	.w2(32'h374ce4b5),
	.w3(32'h3764e20f),
	.w4(32'h378301db),
	.w5(32'h35cf470b),
	.w6(32'h36d911c1),
	.w7(32'h36a93518),
	.w8(32'hb6c1b856),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3839868b),
	.w1(32'h36f87b03),
	.w2(32'hb91bdb38),
	.w3(32'h3913c4a6),
	.w4(32'h3956eae6),
	.w5(32'h38091d2a),
	.w6(32'h3900b61b),
	.w7(32'h394f4516),
	.w8(32'h38ff5f90),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38381ae2),
	.w1(32'h38686042),
	.w2(32'h378dafd7),
	.w3(32'h3810d1d5),
	.w4(32'h3885562c),
	.w5(32'h37f60311),
	.w6(32'h38778ab0),
	.w7(32'h385800d5),
	.w8(32'h38581679),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9671986),
	.w1(32'hb865e71e),
	.w2(32'h3902ee27),
	.w3(32'hb9a857f6),
	.w4(32'hb7ad3c8b),
	.w5(32'h38cee3b3),
	.w6(32'hb91168c6),
	.w7(32'h39632b9c),
	.w8(32'h39509578),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84c3e81),
	.w1(32'hb95c69d4),
	.w2(32'hb9b17ee2),
	.w3(32'hb88a00a2),
	.w4(32'hb92c5074),
	.w5(32'hb93bc211),
	.w6(32'hb6cb602b),
	.w7(32'hb8258e95),
	.w8(32'hb8f92e95),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9b6da),
	.w1(32'h39c30cce),
	.w2(32'hb8085a80),
	.w3(32'h3a03ebc4),
	.w4(32'h39882a79),
	.w5(32'hb911cf17),
	.w6(32'h39e8d92c),
	.w7(32'h396e6baa),
	.w8(32'hb95d944f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb879b83a),
	.w1(32'hb515c0a2),
	.w2(32'h38127902),
	.w3(32'h3785ae9c),
	.w4(32'h3819f9c7),
	.w5(32'h382c12a1),
	.w6(32'h38c812fc),
	.w7(32'h394184f6),
	.w8(32'h3916654e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3ad19),
	.w1(32'hb984f0a7),
	.w2(32'hb99af79f),
	.w3(32'hb7e18877),
	.w4(32'hb9007b77),
	.w5(32'hb984d9b3),
	.w6(32'hb8a6f46a),
	.w7(32'hb8b6d1ba),
	.w8(32'hb9559e99),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e6ea7),
	.w1(32'h3950fe2e),
	.w2(32'h39c95d25),
	.w3(32'hb96df9ea),
	.w4(32'h39867bfa),
	.w5(32'h39ca08d9),
	.w6(32'h392eddcf),
	.w7(32'h39d007a4),
	.w8(32'h39be6bb0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba757755),
	.w1(32'hba268b2c),
	.w2(32'hb91bf69f),
	.w3(32'hba0cfe63),
	.w4(32'hb9a4afb8),
	.w5(32'hb92ef6f3),
	.w6(32'hb9aab39b),
	.w7(32'h39020b05),
	.w8(32'h3996eac3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00a9d6),
	.w1(32'h38fcf643),
	.w2(32'hba064546),
	.w3(32'h39b83d1f),
	.w4(32'hb70733da),
	.w5(32'hba2f9e44),
	.w6(32'h39f21b1c),
	.w7(32'h3994abfc),
	.w8(32'h380e721d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ecffe),
	.w1(32'h39a2fd69),
	.w2(32'h38f47492),
	.w3(32'h3999736c),
	.w4(32'h3a092a5b),
	.w5(32'h3913bc86),
	.w6(32'hb9257b2d),
	.w7(32'h361e21e1),
	.w8(32'h37957bff),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aaade7),
	.w1(32'h3800076a),
	.w2(32'hb899bc8a),
	.w3(32'h37a5494f),
	.w4(32'hb7b85c2f),
	.w5(32'hb923fe8d),
	.w6(32'hb9017b54),
	.w7(32'hb8977985),
	.w8(32'hb901a9c0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00fad3),
	.w1(32'hba028f16),
	.w2(32'hba0cd837),
	.w3(32'hb9b82a12),
	.w4(32'hb9b0d2e6),
	.w5(32'hb99d5d43),
	.w6(32'hb9cdacb4),
	.w7(32'hb8071cf4),
	.w8(32'hb9404dba),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384b648b),
	.w1(32'h38d2080c),
	.w2(32'hb879734f),
	.w3(32'hb8cfa621),
	.w4(32'h383a72c9),
	.w5(32'h385a8cb4),
	.w6(32'hb8f4646b),
	.w7(32'h38aaf378),
	.w8(32'hb898b513),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d714e),
	.w1(32'h390f461f),
	.w2(32'h382877e8),
	.w3(32'h392997b5),
	.w4(32'h3a08f777),
	.w5(32'h39850535),
	.w6(32'h38e5fccc),
	.w7(32'h380a0f43),
	.w8(32'h3803fdd7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e0a75),
	.w1(32'h3956a7e7),
	.w2(32'h39797845),
	.w3(32'hb9156787),
	.w4(32'h3941b32e),
	.w5(32'h3983e8a7),
	.w6(32'h390d2e92),
	.w7(32'h39b5ee23),
	.w8(32'h39a729c6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecece9),
	.w1(32'hb96c948b),
	.w2(32'hb98ecbcf),
	.w3(32'hb9b116bc),
	.w4(32'hb8c61482),
	.w5(32'hb98d96f1),
	.w6(32'hb93fa9ed),
	.w7(32'h36b169fe),
	.w8(32'hb882d6b1),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3752371e),
	.w1(32'h36420326),
	.w2(32'hb5e15561),
	.w3(32'h3764de3b),
	.w4(32'h35da7bef),
	.w5(32'hb68c107e),
	.w6(32'h3750c9fe),
	.w7(32'h36085fb7),
	.w8(32'hb69f6ed2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a9d432),
	.w1(32'h389453db),
	.w2(32'h378daecb),
	.w3(32'h388316a3),
	.w4(32'h383f50ae),
	.w5(32'h37cb97f4),
	.w6(32'h386656dc),
	.w7(32'h38065f87),
	.w8(32'hb771128e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f49bb1),
	.w1(32'h381ec92e),
	.w2(32'hb82ad717),
	.w3(32'hb7de50f2),
	.w4(32'h370c2861),
	.w5(32'hb833366d),
	.w6(32'h378f0126),
	.w7(32'h375ffefc),
	.w8(32'hb7e42966),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac3df6),
	.w1(32'hb81b768f),
	.w2(32'hb99ef631),
	.w3(32'h3899d06a),
	.w4(32'hb87e9a80),
	.w5(32'hb9aa3972),
	.w6(32'hb8b06ebf),
	.w7(32'hb90bbc75),
	.w8(32'hb9a4633f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66f2208),
	.w1(32'h359e9322),
	.w2(32'h359f3219),
	.w3(32'hb64fa4aa),
	.w4(32'hb6a0d32d),
	.w5(32'h34f185e0),
	.w6(32'h352b6752),
	.w7(32'hb5a41ca9),
	.w8(32'hb62e0a9e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b7962),
	.w1(32'h396a0410),
	.w2(32'h395cd2cc),
	.w3(32'h394e1c54),
	.w4(32'h3951055c),
	.w5(32'h394bfbbc),
	.w6(32'h38ab6bb8),
	.w7(32'h38d143b4),
	.w8(32'h38074b86),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78e19ce),
	.w1(32'hb7cddad5),
	.w2(32'h3715416d),
	.w3(32'hb89c92b2),
	.w4(32'h370db51e),
	.w5(32'h38495c02),
	.w6(32'h37c2c44a),
	.w7(32'h38bd692a),
	.w8(32'h38183cca),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398935cf),
	.w1(32'h391cc89b),
	.w2(32'h38386c14),
	.w3(32'h39e0c437),
	.w4(32'h3951ed7c),
	.w5(32'h3865bddb),
	.w6(32'h394a43ea),
	.w7(32'h39118681),
	.w8(32'hb8b792c0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c3c6a),
	.w1(32'h3893caaa),
	.w2(32'h395dc1a4),
	.w3(32'h3845bc4d),
	.w4(32'hb73ea274),
	.w5(32'h39a349d3),
	.w6(32'h392df333),
	.w7(32'h38377067),
	.w8(32'h392ea0a4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f04379),
	.w1(32'hb8a65acc),
	.w2(32'hb89ed7d8),
	.w3(32'h3644d7a2),
	.w4(32'hb8b5d852),
	.w5(32'hb89b56fa),
	.w6(32'h3706fc27),
	.w7(32'h37dfb2c8),
	.w8(32'h380680e0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78836e),
	.w1(32'h3a80d313),
	.w2(32'h36d6816e),
	.w3(32'h3a823af4),
	.w4(32'h3a5b9dff),
	.w5(32'h37f95200),
	.w6(32'h3a14add4),
	.w7(32'h39e9b7f2),
	.w8(32'hb98df36d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba459de1),
	.w1(32'hb88cfa58),
	.w2(32'h39b1b53e),
	.w3(32'hb99d8046),
	.w4(32'hb8b321b9),
	.w5(32'h39870861),
	.w6(32'hb88eabd0),
	.w7(32'h3853ef57),
	.w8(32'h399cab14),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382439d0),
	.w1(32'hb78318ca),
	.w2(32'hb834792c),
	.w3(32'h38c6ff44),
	.w4(32'h38e172ec),
	.w5(32'h38df3644),
	.w6(32'h3956bd09),
	.w7(32'h3985d4bc),
	.w8(32'h38e2030c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33c11d2c),
	.w1(32'hb7855c44),
	.w2(32'hb658d925),
	.w3(32'h361be67d),
	.w4(32'hb55ab110),
	.w5(32'h36d0270c),
	.w6(32'hb76860d6),
	.w7(32'hb7a510dd),
	.w8(32'hb775b466),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03e318),
	.w1(32'h39b5658a),
	.w2(32'h3982dc04),
	.w3(32'h39f0badc),
	.w4(32'h399d058b),
	.w5(32'h399322bd),
	.w6(32'h3914371f),
	.w7(32'hb9000586),
	.w8(32'hb8c506e2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3805ffc4),
	.w1(32'h37198fe9),
	.w2(32'h36b73041),
	.w3(32'h379fbe32),
	.w4(32'hb5b46dd0),
	.w5(32'hb690b98c),
	.w6(32'hb8a45570),
	.w7(32'hb83003ad),
	.w8(32'hb744d850),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390cf055),
	.w1(32'h3957826f),
	.w2(32'h39091989),
	.w3(32'h398bab93),
	.w4(32'h39649294),
	.w5(32'h394eaa64),
	.w6(32'h397179f0),
	.w7(32'h392d8d72),
	.w8(32'h38df3d42),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9891df4),
	.w1(32'hb9c5e2b1),
	.w2(32'hb99b2ecd),
	.w3(32'h391933d1),
	.w4(32'h3987c3c8),
	.w5(32'hb8d421bc),
	.w6(32'h397024f8),
	.w7(32'h39e6d0bd),
	.w8(32'h39287576),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d88f4),
	.w1(32'h3976226c),
	.w2(32'h393e2026),
	.w3(32'h394357b6),
	.w4(32'h390d104f),
	.w5(32'h38f85b94),
	.w6(32'h39205767),
	.w7(32'h38dc6e10),
	.w8(32'h388c9915),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9048a74),
	.w1(32'hb84691a2),
	.w2(32'h388cb18e),
	.w3(32'h364d1b8e),
	.w4(32'h379ae8a4),
	.w5(32'h38db873f),
	.w6(32'h3826a2eb),
	.w7(32'h3876d3ce),
	.w8(32'h38dad37b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11de74),
	.w1(32'h39e89ffc),
	.w2(32'h39de44d3),
	.w3(32'h3990a1d2),
	.w4(32'hb79e69c8),
	.w5(32'hb8ec1e3e),
	.w6(32'h39fc2798),
	.w7(32'h39631888),
	.w8(32'hb896c0c9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c173a),
	.w1(32'hb9b3551e),
	.w2(32'hb9429ce1),
	.w3(32'hb8618a72),
	.w4(32'hb9bd6ba1),
	.w5(32'hb907e05c),
	.w6(32'h3930e504),
	.w7(32'h3904d445),
	.w8(32'h390aaff4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6693774),
	.w1(32'hb69095ad),
	.w2(32'hb4bc0132),
	.w3(32'hb6aa8f1b),
	.w4(32'hb66e62dc),
	.w5(32'hb506dad3),
	.w6(32'h362b507d),
	.w7(32'hb52db183),
	.w8(32'hb52271c5),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39315110),
	.w1(32'hb91ea757),
	.w2(32'hb99fdbba),
	.w3(32'h393085ca),
	.w4(32'hb8a478bb),
	.w5(32'hb97801e4),
	.w6(32'h388c1978),
	.w7(32'hb8e999aa),
	.w8(32'hb9a1ac82),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3779e398),
	.w1(32'hb5e44025),
	.w2(32'hb6ac5e19),
	.w3(32'h375a2948),
	.w4(32'hb613bc85),
	.w5(32'hb7220e9d),
	.w6(32'h37124e28),
	.w7(32'hb6e5525e),
	.w8(32'hb7456f00),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38701813),
	.w1(32'hb8484e33),
	.w2(32'hb8fa37a4),
	.w3(32'h387110ad),
	.w4(32'h38219c73),
	.w5(32'h36e18198),
	.w6(32'h39039436),
	.w7(32'h3977bbbb),
	.w8(32'h38cd6bff),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e1ab11),
	.w1(32'h37d40d90),
	.w2(32'h397e263b),
	.w3(32'hb941cbae),
	.w4(32'hb8ea8364),
	.w5(32'h38f02010),
	.w6(32'hb9725c15),
	.w7(32'hb8c845a9),
	.w8(32'hb7e2b88d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb862eee5),
	.w1(32'h38cde363),
	.w2(32'h38f54f15),
	.w3(32'hb8990786),
	.w4(32'h386353eb),
	.w5(32'h358e60c5),
	.w6(32'h3854bd58),
	.w7(32'h398bd63f),
	.w8(32'h398419d7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8250fe1),
	.w1(32'h3708bf78),
	.w2(32'h383ef5fa),
	.w3(32'hb7ff8928),
	.w4(32'h34f26908),
	.w5(32'h3875df43),
	.w6(32'hb7132c36),
	.w7(32'h3584cb21),
	.w8(32'h381094d5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898a8ec),
	.w1(32'h37682a34),
	.w2(32'h395ed7f7),
	.w3(32'hb9044d39),
	.w4(32'hb740fc24),
	.w5(32'h38604d5d),
	.w6(32'h3880cdb9),
	.w7(32'h39221e57),
	.w8(32'h3970c868),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbf562),
	.w1(32'h3a09e409),
	.w2(32'h398851bf),
	.w3(32'h39e801fe),
	.w4(32'h39c37594),
	.w5(32'h39a4cdd3),
	.w6(32'h3999ea46),
	.w7(32'h38c99e0f),
	.w8(32'h38fb7830),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36121f),
	.w1(32'hb9b499ac),
	.w2(32'hb9b83ecc),
	.w3(32'hba2cb446),
	.w4(32'hb9a0eb79),
	.w5(32'hba043aba),
	.w6(32'hb92c2465),
	.w7(32'h38b2f06f),
	.w8(32'hb953f2c1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382df17d),
	.w1(32'h36c5bb31),
	.w2(32'hb7314d45),
	.w3(32'h37b9e421),
	.w4(32'h37ec0db6),
	.w5(32'h36df9995),
	.w6(32'h37a56e1e),
	.w7(32'h37f1b360),
	.w8(32'h34af04ce),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370689e0),
	.w1(32'hb68349c0),
	.w2(32'hb6838b5a),
	.w3(32'hb60722ba),
	.w4(32'hb5ebe84f),
	.w5(32'hb6854b4a),
	.w6(32'hb68d0a49),
	.w7(32'hb6a449f8),
	.w8(32'hb73cb7f5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f81ea),
	.w1(32'h3884a450),
	.w2(32'h38b27a04),
	.w3(32'hb914b073),
	.w4(32'hb87521df),
	.w5(32'h38c91109),
	.w6(32'h3931a559),
	.w7(32'h39708dc2),
	.w8(32'h39545293),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b69acf),
	.w1(32'hb99f13fb),
	.w2(32'hb9c9db51),
	.w3(32'hb997d048),
	.w4(32'hb9a221a9),
	.w5(32'hb9afa159),
	.w6(32'hb8881b1f),
	.w7(32'h396d5f7e),
	.w8(32'h39130dfd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82edd63),
	.w1(32'h3867c95b),
	.w2(32'hb8c12311),
	.w3(32'hb9d1818a),
	.w4(32'hb8f88993),
	.w5(32'hb9495bae),
	.w6(32'h384f8a67),
	.w7(32'h3947ee1a),
	.w8(32'hb57d3c0c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372da404),
	.w1(32'h3880351a),
	.w2(32'hb9d1007f),
	.w3(32'h39ac13b9),
	.w4(32'h399f61e4),
	.w5(32'hb759e97d),
	.w6(32'h3930df97),
	.w7(32'h3820bca5),
	.w8(32'hb8b71077),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3818cc6e),
	.w1(32'hb726c73c),
	.w2(32'hb869fe04),
	.w3(32'h37fa35cd),
	.w4(32'hb790608c),
	.w5(32'hb85dee07),
	.w6(32'h380aeb99),
	.w7(32'hb7790f00),
	.w8(32'hb897f633),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386e969a),
	.w1(32'hb718d98b),
	.w2(32'hb9033526),
	.w3(32'h36bae714),
	.w4(32'hb8357e1d),
	.w5(32'hb8f79669),
	.w6(32'hb8b3b469),
	.w7(32'hb7ca73dc),
	.w8(32'hb8c32808),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88e3c0d),
	.w1(32'h39c2c5b2),
	.w2(32'h39feb545),
	.w3(32'h38fceaaa),
	.w4(32'h3940c6c0),
	.w5(32'h39a80789),
	.w6(32'h394fb88f),
	.w7(32'h39bc6cc4),
	.w8(32'h3930b24c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9857528),
	.w1(32'hba10194a),
	.w2(32'hba635e0e),
	.w3(32'hb9638d28),
	.w4(32'hb9d2c364),
	.w5(32'hba3aab4a),
	.w6(32'h394a2235),
	.w7(32'h39863dac),
	.w8(32'hb98487ad),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392bcb47),
	.w1(32'hb83fc7a9),
	.w2(32'hb915413a),
	.w3(32'h39a808b2),
	.w4(32'h389cad6e),
	.w5(32'hb851fe46),
	.w6(32'h3a0ef376),
	.w7(32'h3984c0e8),
	.w8(32'h38e10f53),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89709d9),
	.w1(32'h382c7578),
	.w2(32'h39a677db),
	.w3(32'hb9068baa),
	.w4(32'h37bea399),
	.w5(32'h396d5649),
	.w6(32'hb79a5b72),
	.w7(32'hb6eacb22),
	.w8(32'h390f5ea4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e0e07),
	.w1(32'h39843ef0),
	.w2(32'h39f77470),
	.w3(32'hb9134d00),
	.w4(32'h3888911c),
	.w5(32'h39820fd9),
	.w6(32'hb93f5740),
	.w7(32'hb87fd129),
	.w8(32'h37be4b34),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e4db7c),
	.w1(32'hb664b2a7),
	.w2(32'hb6c964a2),
	.w3(32'h34fa6b0e),
	.w4(32'hb6ac2f94),
	.w5(32'hb738113f),
	.w6(32'h360ba188),
	.w7(32'hb5907108),
	.w8(32'hb65e5fa4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35158d54),
	.w1(32'hb4a023e1),
	.w2(32'hb53c6987),
	.w3(32'hb627ee43),
	.w4(32'hb63038cd),
	.w5(32'hb5cd35ba),
	.w6(32'hb41c2816),
	.w7(32'hb5ab50a5),
	.w8(32'h34ade17d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dd3a9e),
	.w1(32'h37004f37),
	.w2(32'h36cedbc5),
	.w3(32'h3837f969),
	.w4(32'h38880f21),
	.w5(32'h38487b4e),
	.w6(32'h378bda7f),
	.w7(32'h36c94578),
	.w8(32'h36bd5c01),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3592ddca),
	.w1(32'hb736d2ce),
	.w2(32'h3600175d),
	.w3(32'h371b7c9a),
	.w4(32'hb68fd797),
	.w5(32'hb52eeec5),
	.w6(32'h36a4a43a),
	.w7(32'h35dc0b21),
	.w8(32'hb6a9f14a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a0ee8),
	.w1(32'h38be214a),
	.w2(32'h37c146ad),
	.w3(32'h38877dad),
	.w4(32'h38948ce3),
	.w5(32'h3833869f),
	.w6(32'h38c66f49),
	.w7(32'h381138d2),
	.w8(32'hb6a6b371),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ceab9),
	.w1(32'hb9a36555),
	.w2(32'hba165572),
	.w3(32'hb98a9e70),
	.w4(32'hb9c028e7),
	.w5(32'hba04be62),
	.w6(32'hb9554e08),
	.w7(32'hb8eb9f1d),
	.w8(32'hb99c5fef),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972ccd9),
	.w1(32'hb8cfbbc3),
	.w2(32'hb6e2be7e),
	.w3(32'hb980aae6),
	.w4(32'hb90933e0),
	.w5(32'h36df8e7a),
	.w6(32'hb90b6bea),
	.w7(32'h38800133),
	.w8(32'h3911bb5c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69d6672),
	.w1(32'h35a5dbb2),
	.w2(32'h36d0944e),
	.w3(32'hb6a4ed7d),
	.w4(32'h35858f1e),
	.w5(32'h3709b0f0),
	.w6(32'h372a5ce4),
	.w7(32'h370e7558),
	.w8(32'h3721d6c3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf0484),
	.w1(32'hb99897d2),
	.w2(32'hb9d2d7ab),
	.w3(32'h37832e69),
	.w4(32'hb920222b),
	.w5(32'hb9199fff),
	.w6(32'h39140de4),
	.w7(32'h3821f9e6),
	.w8(32'h39258d82),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37baf2b0),
	.w1(32'h38d4ee00),
	.w2(32'hb8446d74),
	.w3(32'h38aac2ae),
	.w4(32'h3909206a),
	.w5(32'h371d40a8),
	.w6(32'h38f2b8b5),
	.w7(32'h3922b82a),
	.w8(32'hb6ef7ed4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f2c697),
	.w1(32'h37958f54),
	.w2(32'h37168d66),
	.w3(32'h3704fbe7),
	.w4(32'h375fd82e),
	.w5(32'h36e8a58f),
	.w6(32'h3714358b),
	.w7(32'h3748d0cd),
	.w8(32'h3709bc05),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1a0b3),
	.w1(32'hb98c7608),
	.w2(32'hb98bb371),
	.w3(32'hb8debb37),
	.w4(32'hb88b2d58),
	.w5(32'hb90ae145),
	.w6(32'h3909fe61),
	.w7(32'h3962c9ca),
	.w8(32'h38e975cd),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee6b33),
	.w1(32'h3890cb04),
	.w2(32'h378b8891),
	.w3(32'h3899a175),
	.w4(32'h386d4bf0),
	.w5(32'h375f3c50),
	.w6(32'hb826c31f),
	.w7(32'hb86ab691),
	.w8(32'hb883149e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981df3d),
	.w1(32'hb90a39cf),
	.w2(32'hb80b3fd1),
	.w3(32'hb90dab89),
	.w4(32'hb7fdb9b0),
	.w5(32'hb6b1d5fb),
	.w6(32'hb7ea1d04),
	.w7(32'h380eb293),
	.w8(32'h387afb29),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c0c0f1),
	.w1(32'h370a4409),
	.w2(32'h3702ae4b),
	.w3(32'hb63146fe),
	.w4(32'h366c48df),
	.w5(32'h370ae470),
	.w6(32'h36a6f4a7),
	.w7(32'h36aa84e2),
	.w8(32'h35bc24de),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66ffd12),
	.w1(32'hb683e227),
	.w2(32'hb6b967a7),
	.w3(32'h34413545),
	.w4(32'hb700a6a0),
	.w5(32'hb76899ee),
	.w6(32'h362745a7),
	.w7(32'hb6145b6e),
	.w8(32'hb52ac26a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d6a9f),
	.w1(32'h3928af8f),
	.w2(32'h393fd8e2),
	.w3(32'hb7a34b49),
	.w4(32'h379cbc5b),
	.w5(32'h38fbc277),
	.w6(32'h368f95ac),
	.w7(32'hb7c084c5),
	.w8(32'h3832ed94),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6c64d),
	.w1(32'hb9aeafed),
	.w2(32'hba3886d9),
	.w3(32'hb99c893a),
	.w4(32'hb8f7d2fd),
	.w5(32'hba14c580),
	.w6(32'hb9844956),
	.w7(32'h37aa9725),
	.w8(32'hb9a4ab38),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8274f),
	.w1(32'hb948a943),
	.w2(32'hb9b10074),
	.w3(32'hb8ecf6dc),
	.w4(32'h384ecfaf),
	.w5(32'hb8b46476),
	.w6(32'h3946dd4e),
	.w7(32'h39c32228),
	.w8(32'h394566d4),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a6efa),
	.w1(32'hba45addb),
	.w2(32'hba60abb6),
	.w3(32'hb9e2d798),
	.w4(32'hb9d66b3b),
	.w5(32'hba03a528),
	.w6(32'hb69e123a),
	.w7(32'h38ccf2d0),
	.w8(32'hb92bc56a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb649cd7f),
	.w1(32'hb7607437),
	.w2(32'hb68e01bc),
	.w3(32'hb732128a),
	.w4(32'hb789f2d8),
	.w5(32'hb46ab5a5),
	.w6(32'h3616761c),
	.w7(32'hb6e30c4e),
	.w8(32'h3755343e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809c1e8),
	.w1(32'hb6fe7e6c),
	.w2(32'hb855f010),
	.w3(32'h37e9952c),
	.w4(32'hb7830d4d),
	.w5(32'hb845141e),
	.w6(32'h37614428),
	.w7(32'hb7d66210),
	.w8(32'hb86a89c7),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a5177b),
	.w1(32'hb5992d2f),
	.w2(32'hb5f54b0d),
	.w3(32'h37063f08),
	.w4(32'h36b48633),
	.w5(32'h37ba5eab),
	.w6(32'h375b8a21),
	.w7(32'h3597647e),
	.w8(32'h364b30df),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb44a2202),
	.w1(32'h354b21b6),
	.w2(32'h35d96c3b),
	.w3(32'h36368f5e),
	.w4(32'h36ae037e),
	.w5(32'h36f3133c),
	.w6(32'h3696468c),
	.w7(32'h36969b38),
	.w8(32'h36972040),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c47fb4),
	.w1(32'hb8afb214),
	.w2(32'hba0020f9),
	.w3(32'h38b2653e),
	.w4(32'hb7e90633),
	.w5(32'hb9a29b41),
	.w6(32'h3934c5a0),
	.w7(32'hb83ef0c9),
	.w8(32'hb9585620),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39045782),
	.w1(32'h393f3fa4),
	.w2(32'h39341ec6),
	.w3(32'h3968e7c4),
	.w4(32'h393c94a4),
	.w5(32'h395400b3),
	.w6(32'hb73e9883),
	.w7(32'hb93257d3),
	.w8(32'hb81f4f04),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f79798),
	.w1(32'hb748cf2f),
	.w2(32'hb91d4a97),
	.w3(32'h391e88f8),
	.w4(32'h3841e2cf),
	.w5(32'hb8811f49),
	.w6(32'h391ea17f),
	.w7(32'h38a193fc),
	.w8(32'hb7ead58e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922c9cb),
	.w1(32'hb7fba1cd),
	.w2(32'hb9092697),
	.w3(32'h38395223),
	.w4(32'hb897cb8d),
	.w5(32'hb91d625c),
	.w6(32'hb91211c0),
	.w7(32'hb92305dd),
	.w8(32'hb9532803),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a60fd3),
	.w1(32'h3837bf1b),
	.w2(32'h368c7b83),
	.w3(32'h38e0360f),
	.w4(32'h37c97cca),
	.w5(32'hb75c4e25),
	.w6(32'h3827e631),
	.w7(32'hb8602a3b),
	.w8(32'hb8369cf2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a7f854),
	.w1(32'hb739c1cf),
	.w2(32'hb9009b31),
	.w3(32'h38805b4d),
	.w4(32'h370c7044),
	.w5(32'hb90f8034),
	.w6(32'h390da08b),
	.w7(32'h38a11650),
	.w8(32'hb89e1954),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b90152),
	.w1(32'h371b4e18),
	.w2(32'hb7b0d20c),
	.w3(32'h36c38398),
	.w4(32'hb73cb651),
	.w5(32'hb802ac4e),
	.w6(32'h35971e49),
	.w7(32'hb7efa16b),
	.w8(32'hb8367278),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968b16e),
	.w1(32'hb9f09884),
	.w2(32'hba637f2b),
	.w3(32'hb95a4ffd),
	.w4(32'hb98e5789),
	.w5(32'hba573333),
	.w6(32'hb9a6cb05),
	.w7(32'hb977ec63),
	.w8(32'hba1a4879),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3736b9dc),
	.w1(32'hbb20c09a),
	.w2(32'hbaf9cc20),
	.w3(32'h37273949),
	.w4(32'hbafa5f6d),
	.w5(32'hba70bb75),
	.w6(32'hbb42bfae),
	.w7(32'hbaca14c1),
	.w8(32'hba4b119b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c4a3),
	.w1(32'h3a488070),
	.w2(32'hb9780eaf),
	.w3(32'hbb1485af),
	.w4(32'h3948a5a9),
	.w5(32'h39e9db39),
	.w6(32'h39dfbc5c),
	.w7(32'hb9862897),
	.w8(32'hb9350988),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule