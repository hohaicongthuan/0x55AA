module layer_10_featuremap_366(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29d8dc),
	.w1(32'h3a11f89c),
	.w2(32'hbbdf4668),
	.w3(32'h393c35a1),
	.w4(32'hbb090d68),
	.w5(32'hbb2145eb),
	.w6(32'hbb589abd),
	.w7(32'h3998089a),
	.w8(32'hbb6ce751),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfa786),
	.w1(32'hb8e54f5b),
	.w2(32'h3b08effd),
	.w3(32'hb9e332b1),
	.w4(32'h3ae36d72),
	.w5(32'h3b6ff894),
	.w6(32'hbc9618ce),
	.w7(32'hbc3972be),
	.w8(32'hbc283659),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f4a9f),
	.w1(32'hb9dc3dae),
	.w2(32'hba77bbb0),
	.w3(32'h3bd9f5ef),
	.w4(32'h3c6ed7bb),
	.w5(32'hb9936374),
	.w6(32'hbcf785d0),
	.w7(32'hbc8812c9),
	.w8(32'hbbd0b599),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0de062),
	.w1(32'h3cae67e4),
	.w2(32'h3ad001a9),
	.w3(32'hbcc271ae),
	.w4(32'hbcf6fd26),
	.w5(32'h3c4c8047),
	.w6(32'h3af28f75),
	.w7(32'hbbb15ca0),
	.w8(32'hbba37f28),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b78a0),
	.w1(32'h3cb2de7f),
	.w2(32'hbb937882),
	.w3(32'hbcddae2e),
	.w4(32'hbb4627ec),
	.w5(32'hba8b54b5),
	.w6(32'h3c50d929),
	.w7(32'hbc3dd178),
	.w8(32'hbd49e782),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07f3ce),
	.w1(32'h3c5c00ce),
	.w2(32'hbb1146a5),
	.w3(32'h3be28631),
	.w4(32'h3bd95079),
	.w5(32'h3c193749),
	.w6(32'hbb809e31),
	.w7(32'hbb87240b),
	.w8(32'h3b1a9465),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad05fa7),
	.w1(32'hbb59893f),
	.w2(32'hba881130),
	.w3(32'hbcbaaf7f),
	.w4(32'h3cdf4296),
	.w5(32'hbb3cfa0f),
	.w6(32'hbb86338d),
	.w7(32'h3bd7a9ad),
	.w8(32'hbb1cfb9f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb62a27),
	.w1(32'h3a912e53),
	.w2(32'h3aa1a1f2),
	.w3(32'h3c07c007),
	.w4(32'hba1f8e81),
	.w5(32'hbbb5070f),
	.w6(32'hba43a3ba),
	.w7(32'hbb25c748),
	.w8(32'hbb9077da),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7180c0),
	.w1(32'h3a70dfca),
	.w2(32'hbb188c16),
	.w3(32'hbb25bd77),
	.w4(32'h3c238fa8),
	.w5(32'h3c2264dd),
	.w6(32'hbb042d83),
	.w7(32'hbc190430),
	.w8(32'h3a0d33cd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01583e),
	.w1(32'hba095b97),
	.w2(32'h3c7790d8),
	.w3(32'h3a4eed53),
	.w4(32'h3b9087cb),
	.w5(32'h3b30c003),
	.w6(32'h3bbf072c),
	.w7(32'h3c0cd3f6),
	.w8(32'hbbdf2af6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b8edb),
	.w1(32'hbc803488),
	.w2(32'h3bbfc5a6),
	.w3(32'h3b8763a0),
	.w4(32'hbc07e862),
	.w5(32'h3c4df10f),
	.w6(32'hbc366aaf),
	.w7(32'h3b43f6c5),
	.w8(32'hbb85f556),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9c04e),
	.w1(32'hbb892432),
	.w2(32'h3cd7b619),
	.w3(32'hbbb6909f),
	.w4(32'h3d03c656),
	.w5(32'h3b695ae2),
	.w6(32'h3a7afb0c),
	.w7(32'h3912607a),
	.w8(32'h3b1336c9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62ce8d),
	.w1(32'h3bd4d23f),
	.w2(32'h3c118af0),
	.w3(32'hbb9f8cf4),
	.w4(32'h3b0f68d8),
	.w5(32'h3c16fa23),
	.w6(32'h3bd20ff5),
	.w7(32'h3be6aa85),
	.w8(32'hbc9f7d92),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a36c8),
	.w1(32'h3c249e6b),
	.w2(32'hbaf8351f),
	.w3(32'h3ba3fb0c),
	.w4(32'hbd459045),
	.w5(32'hba9b3d83),
	.w6(32'h3ce8c990),
	.w7(32'h3c25f0cd),
	.w8(32'h3ab6c7d8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e43ab),
	.w1(32'hbb4d476f),
	.w2(32'h3bdaf6a3),
	.w3(32'hbae23f7e),
	.w4(32'hb96d2bad),
	.w5(32'hbb6cdd69),
	.w6(32'hbae0469a),
	.w7(32'h3bc092d7),
	.w8(32'h3ad9da7c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b348a09),
	.w1(32'h3b56aa53),
	.w2(32'h3a0e201d),
	.w3(32'h3c0058b3),
	.w4(32'hbc01735e),
	.w5(32'hba3c9525),
	.w6(32'hba217c33),
	.w7(32'hbc27fe60),
	.w8(32'hbc62b305),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdee58),
	.w1(32'h3bbc5ded),
	.w2(32'h3c1607f4),
	.w3(32'hbc2e79a6),
	.w4(32'hb8b87e4c),
	.w5(32'hbc07d58a),
	.w6(32'hbc0e3ee3),
	.w7(32'h3b140e3b),
	.w8(32'hba2cec21),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d72da),
	.w1(32'h3bbd4bb6),
	.w2(32'hbbfdf461),
	.w3(32'h3a023832),
	.w4(32'h3c09b77f),
	.w5(32'hbb4df197),
	.w6(32'h3bc8c7d8),
	.w7(32'hbd3a607a),
	.w8(32'hba373336),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8446d9),
	.w1(32'h3c1255c6),
	.w2(32'hba37c115),
	.w3(32'hbbd705ad),
	.w4(32'hbb8b9ef0),
	.w5(32'h3c91b9a5),
	.w6(32'hbc001e3b),
	.w7(32'h3c02c2bd),
	.w8(32'hbb94b3b9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41eac4),
	.w1(32'hbc8da39e),
	.w2(32'hbc1cf1dc),
	.w3(32'hbb9af40a),
	.w4(32'h3d0299e1),
	.w5(32'hbc357d7d),
	.w6(32'hbca1b4f1),
	.w7(32'hbb587b0a),
	.w8(32'hb9671089),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeb77f),
	.w1(32'h3b58dc47),
	.w2(32'h3c73a323),
	.w3(32'hbbd7091f),
	.w4(32'h3bf06a73),
	.w5(32'hbbed6654),
	.w6(32'h3a9484f2),
	.w7(32'hb84db450),
	.w8(32'h3c89cebf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bfd8a),
	.w1(32'hbd21e036),
	.w2(32'hbb72b571),
	.w3(32'hbb625ee8),
	.w4(32'hbb2d4ac8),
	.w5(32'hbc7175d8),
	.w6(32'hbd032339),
	.w7(32'hba9a45bb),
	.w8(32'hba414d91),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc563e3),
	.w1(32'h39b0d1d6),
	.w2(32'hbd792afc),
	.w3(32'h3b452230),
	.w4(32'h3995d21c),
	.w5(32'h3b96e2b8),
	.w6(32'hba8744a1),
	.w7(32'hbaec7c86),
	.w8(32'h3b69d4eb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc382542),
	.w1(32'hbbf93632),
	.w2(32'hbbb119e3),
	.w3(32'hbab471d1),
	.w4(32'hb9ed6de0),
	.w5(32'h3941ad09),
	.w6(32'h3c3df80f),
	.w7(32'hbb8e8f3c),
	.w8(32'hbc0dad0f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2658d),
	.w1(32'h3c574a88),
	.w2(32'hba45bd31),
	.w3(32'h3c09e11a),
	.w4(32'h3cb6835f),
	.w5(32'h3b659166),
	.w6(32'h3ac012fb),
	.w7(32'h39820ec5),
	.w8(32'hbc8767c0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8c24c),
	.w1(32'h3af15386),
	.w2(32'h3c42c035),
	.w3(32'hbc39421f),
	.w4(32'hbb6b5006),
	.w5(32'h3b10475e),
	.w6(32'hbb1f2fc9),
	.w7(32'hbb6c450a),
	.w8(32'h3a3803bc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ace0e3),
	.w1(32'hbab7799d),
	.w2(32'h3bcf4e70),
	.w3(32'hbb52f3e0),
	.w4(32'hbb866a82),
	.w5(32'h3b327cbd),
	.w6(32'hbc3ca39e),
	.w7(32'h3a541f17),
	.w8(32'hbbf39b82),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b20793),
	.w1(32'hba91508b),
	.w2(32'h3b75fb4b),
	.w3(32'hbbcb19d6),
	.w4(32'h3a894866),
	.w5(32'h3b977a75),
	.w6(32'h3a1b1bb4),
	.w7(32'h3b9c658f),
	.w8(32'h3b69e2d8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b91f),
	.w1(32'h39e07cff),
	.w2(32'h3bf8016d),
	.w3(32'hbb81e6e5),
	.w4(32'h3a90c521),
	.w5(32'h3ba0fe0c),
	.w6(32'h3b0a8181),
	.w7(32'hbb407fc3),
	.w8(32'hbbb13c43),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89ad05),
	.w1(32'h3bce3118),
	.w2(32'h39aac94b),
	.w3(32'h3bed71b6),
	.w4(32'hbc467158),
	.w5(32'hbb22ceeb),
	.w6(32'h3c4242ed),
	.w7(32'h3911287f),
	.w8(32'h3be8daa1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf3f70),
	.w1(32'hbb0f8692),
	.w2(32'hbd21626c),
	.w3(32'h3b6d7545),
	.w4(32'h3c1c7e1d),
	.w5(32'hbbb50c5a),
	.w6(32'h3a25e386),
	.w7(32'hbab564fd),
	.w8(32'h3c7c2648),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70d4ee),
	.w1(32'h3b0a5911),
	.w2(32'hbb8ce2ec),
	.w3(32'h3cc0c590),
	.w4(32'hbb830cec),
	.w5(32'hbb209bcf),
	.w6(32'h3c46b471),
	.w7(32'hbd60d671),
	.w8(32'hbc9eadaf),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0322b9),
	.w1(32'hbb19b3c5),
	.w2(32'h3c5239a5),
	.w3(32'h3b767992),
	.w4(32'h3bb210e0),
	.w5(32'h3b8f0963),
	.w6(32'hbc0ca152),
	.w7(32'h38096d37),
	.w8(32'hbacf5bd0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea4f83),
	.w1(32'h3c8f7b48),
	.w2(32'hba970c09),
	.w3(32'hbc2163bd),
	.w4(32'h3c64eafa),
	.w5(32'hbad6677e),
	.w6(32'h39af6d77),
	.w7(32'hbb90f0c4),
	.w8(32'h3bf61289),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e0f68),
	.w1(32'hbb922941),
	.w2(32'h3b2b43d8),
	.w3(32'hba4488fc),
	.w4(32'hbc724e13),
	.w5(32'hbc122e86),
	.w6(32'h3ae6f513),
	.w7(32'hba6808e2),
	.w8(32'hbc6ee4c2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf3062),
	.w1(32'h3bcb419d),
	.w2(32'h3af0c7aa),
	.w3(32'h3c2cac3b),
	.w4(32'h3c0f4108),
	.w5(32'hbc645601),
	.w6(32'h3ba03394),
	.w7(32'hbc918498),
	.w8(32'h3c14e6ae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39887144),
	.w1(32'hbc7b019e),
	.w2(32'h3a397972),
	.w3(32'hbc23ce30),
	.w4(32'hbc3c3189),
	.w5(32'hbbebb68a),
	.w6(32'hbb6b7520),
	.w7(32'hbbf5a989),
	.w8(32'hbb7bfbb7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac51f2b),
	.w1(32'h3a8b46da),
	.w2(32'h3c1ae2fa),
	.w3(32'h3b10f60b),
	.w4(32'h3d74c2dc),
	.w5(32'hba986565),
	.w6(32'h3bb5441c),
	.w7(32'h3b9d20f7),
	.w8(32'hb90c7db6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe7116),
	.w1(32'h3b83da58),
	.w2(32'h3b80e66f),
	.w3(32'hba2149b0),
	.w4(32'h3b063664),
	.w5(32'hbc0baa9d),
	.w6(32'hbbbe190e),
	.w7(32'hbc1710c0),
	.w8(32'hb8e497c6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2feb56),
	.w1(32'hbc2df54c),
	.w2(32'hba9aad47),
	.w3(32'h3a495d06),
	.w4(32'h3ab276c4),
	.w5(32'h3b211d91),
	.w6(32'hbb2919d0),
	.w7(32'h3b4b1634),
	.w8(32'h3d331141),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bf936),
	.w1(32'h3b07e654),
	.w2(32'h3c638ebe),
	.w3(32'h3d8513d8),
	.w4(32'h3b4d6a6f),
	.w5(32'hbb0adb56),
	.w6(32'h3a3e6d85),
	.w7(32'hbb590856),
	.w8(32'hbc026d74),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed64af),
	.w1(32'hbcb15e2f),
	.w2(32'hbc21be7c),
	.w3(32'hbab93cf0),
	.w4(32'h3ca40347),
	.w5(32'h3cec0005),
	.w6(32'hba7254c8),
	.w7(32'hbcc4c1f4),
	.w8(32'hbda59c18),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca189a6),
	.w1(32'hbba677db),
	.w2(32'h3c26aa01),
	.w3(32'h3c0384a4),
	.w4(32'hbc69699e),
	.w5(32'hbb64bd00),
	.w6(32'h3b8ab4ec),
	.w7(32'hbbb34df4),
	.w8(32'hbb29516a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc35f36),
	.w1(32'h3bb539f0),
	.w2(32'hba27f359),
	.w3(32'h3bd258f3),
	.w4(32'hbbadef23),
	.w5(32'hb8ff59de),
	.w6(32'h3bc11eff),
	.w7(32'h3c1536aa),
	.w8(32'hb9d20b89),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a5932),
	.w1(32'h3c0dabce),
	.w2(32'h3b0476d9),
	.w3(32'hbb9eff90),
	.w4(32'hbb58cede),
	.w5(32'h3c14f241),
	.w6(32'hba2e62c8),
	.w7(32'hbbac6681),
	.w8(32'h3a563dd7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12effc),
	.w1(32'h3a1ddb9f),
	.w2(32'h3b4fd980),
	.w3(32'h3bd8eed0),
	.w4(32'hbb312aa8),
	.w5(32'hbc2aae7e),
	.w6(32'hbc6885b0),
	.w7(32'h3a90f34f),
	.w8(32'hbc1d1573),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d8fc9),
	.w1(32'h3aa91693),
	.w2(32'hbbe29073),
	.w3(32'hbaf4f3e6),
	.w4(32'h3b8a2889),
	.w5(32'h3c42b92b),
	.w6(32'hbb1ae22d),
	.w7(32'hbae0e1e6),
	.w8(32'hb8d5564b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b3f0d),
	.w1(32'hbb9d6992),
	.w2(32'hbb638c00),
	.w3(32'h3c02804c),
	.w4(32'h3c73f3b6),
	.w5(32'hbcc97b10),
	.w6(32'hbcc43855),
	.w7(32'hbbac38c6),
	.w8(32'h3c18fb4b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5142e3),
	.w1(32'hbb021bbb),
	.w2(32'h3bfd6bf1),
	.w3(32'hbb3b14d3),
	.w4(32'h3acb3915),
	.w5(32'h3c3f8abc),
	.w6(32'h3c26ca90),
	.w7(32'hbb32065b),
	.w8(32'hbb2d0c00),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc564ee8),
	.w1(32'h3c4e579e),
	.w2(32'h3c398ef1),
	.w3(32'hbbf2799b),
	.w4(32'hbd2c7e74),
	.w5(32'hbc33c216),
	.w6(32'h3ad8aca0),
	.w7(32'hbb5b7f0b),
	.w8(32'hb9b95181),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10c053),
	.w1(32'h3b7fea68),
	.w2(32'hb956757f),
	.w3(32'h3abb9369),
	.w4(32'hbb89f8d3),
	.w5(32'h3a033ded),
	.w6(32'hbbd0a8b9),
	.w7(32'h3ba255ca),
	.w8(32'h3a62edb7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd5c45),
	.w1(32'hbce3b441),
	.w2(32'h3c51cdbd),
	.w3(32'hbd124e00),
	.w4(32'hbb1032d8),
	.w5(32'h3b0f10ad),
	.w6(32'h3c1f240b),
	.w7(32'hba8d5fb3),
	.w8(32'h3bd746ec),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bd21b),
	.w1(32'h3bbf7afd),
	.w2(32'h3bea0b9b),
	.w3(32'hbb6338d5),
	.w4(32'h3ba15874),
	.w5(32'hbc8b90a8),
	.w6(32'hba4394c0),
	.w7(32'h3bce1451),
	.w8(32'h3bbe5eca),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8268ed),
	.w1(32'h3aa162bb),
	.w2(32'hbb1309e6),
	.w3(32'hbaacecd7),
	.w4(32'hbbf40d88),
	.w5(32'hbb71174a),
	.w6(32'hbb31c6ab),
	.w7(32'hbd0466a7),
	.w8(32'h3c44888b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ee44),
	.w1(32'h3b8fd080),
	.w2(32'hba51496a),
	.w3(32'h3c580fa8),
	.w4(32'hbb8dea68),
	.w5(32'hbcd4a1f7),
	.w6(32'h39ed13fe),
	.w7(32'hbb9bd662),
	.w8(32'hbbb78a5e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b3561),
	.w1(32'h3c8a5f2c),
	.w2(32'h3c770bce),
	.w3(32'h3c56e622),
	.w4(32'hbc41089c),
	.w5(32'hbba28554),
	.w6(32'h3aac883f),
	.w7(32'hbadd0d2f),
	.w8(32'hbb408205),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39faf2a4),
	.w1(32'hbb97eeb5),
	.w2(32'h3c9e188e),
	.w3(32'h3ba745ab),
	.w4(32'h3bdb0027),
	.w5(32'h3c7f2f53),
	.w6(32'h3b8c2b9c),
	.w7(32'h3bf26a2c),
	.w8(32'hba5fd3a1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb82303),
	.w1(32'hbae0e9ee),
	.w2(32'hbc024adc),
	.w3(32'hbb038ffe),
	.w4(32'h3cd8628b),
	.w5(32'h3bd5193d),
	.w6(32'h3bbdc3fd),
	.w7(32'hbc004b5b),
	.w8(32'hbb7cdc16),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c685080),
	.w1(32'hbbc901f3),
	.w2(32'hbb20ad49),
	.w3(32'hbc4fac05),
	.w4(32'h3ca6073d),
	.w5(32'h3b8bed65),
	.w6(32'hbc2168a7),
	.w7(32'hbc327308),
	.w8(32'hbb3d1def),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf8af5),
	.w1(32'hbbeebef9),
	.w2(32'hb954598d),
	.w3(32'hbc506bb1),
	.w4(32'hbae6f2e5),
	.w5(32'hbc299d95),
	.w6(32'hbc753716),
	.w7(32'hbc4d2284),
	.w8(32'h3c30c447),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c116097),
	.w1(32'h3ade0be7),
	.w2(32'hbc804027),
	.w3(32'hbbb19465),
	.w4(32'hbc1de6e7),
	.w5(32'h3a97af80),
	.w6(32'hbac87219),
	.w7(32'hbc004a1a),
	.w8(32'h3a868042),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddad4d),
	.w1(32'hbbd9d27d),
	.w2(32'hb8949bed),
	.w3(32'hbbd9e298),
	.w4(32'h3ade5c70),
	.w5(32'h3c16e404),
	.w6(32'h3c8aedc3),
	.w7(32'hbbdc1d39),
	.w8(32'h3c49a4a1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b7ed3),
	.w1(32'h3bd63610),
	.w2(32'hba104eb2),
	.w3(32'h3b05b1f4),
	.w4(32'hbc49496e),
	.w5(32'h3bbe50ac),
	.w6(32'hba570a1e),
	.w7(32'h3b307b74),
	.w8(32'hbbbc68f3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbff842),
	.w1(32'hbc81f22a),
	.w2(32'h3bebde99),
	.w3(32'hbc84bf40),
	.w4(32'h3bcdc7a7),
	.w5(32'h3cc2220b),
	.w6(32'hbb8e72f9),
	.w7(32'hb9ba64f0),
	.w8(32'h36a1d1f1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc510637),
	.w1(32'h3b356481),
	.w2(32'hb78a5c02),
	.w3(32'h3c0adc57),
	.w4(32'hbb8ed582),
	.w5(32'h3c8c55df),
	.w6(32'h3b7bf3b9),
	.w7(32'hbb5255d6),
	.w8(32'hbac1a8ad),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38d2b3),
	.w1(32'h3c4fc57d),
	.w2(32'h3c463c38),
	.w3(32'hbc6dd37a),
	.w4(32'h3abf7a90),
	.w5(32'h3b8e0f09),
	.w6(32'h3c04b18b),
	.w7(32'hbc16d408),
	.w8(32'h3b5d21bc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4fbdc),
	.w1(32'h3cf7a9bd),
	.w2(32'hbc1086e8),
	.w3(32'hbba4c435),
	.w4(32'hbc27c468),
	.w5(32'h3be1845d),
	.w6(32'h3ad6325b),
	.w7(32'h3bdf2c65),
	.w8(32'hbbfffe7b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f7688),
	.w1(32'h3c5584d6),
	.w2(32'hbc7a81a4),
	.w3(32'hbc23f31e),
	.w4(32'hb9db2737),
	.w5(32'hbc4fbe1b),
	.w6(32'h3ae985ee),
	.w7(32'h3a041971),
	.w8(32'h3c41251e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad324c),
	.w1(32'h3be11901),
	.w2(32'h3aafdeaf),
	.w3(32'h3b070bc5),
	.w4(32'h3933c4a5),
	.w5(32'h3a722f3a),
	.w6(32'h3bb34ae2),
	.w7(32'hbc83c3e1),
	.w8(32'h3c9b71c2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be875),
	.w1(32'hba81cb58),
	.w2(32'hbcc08782),
	.w3(32'hbbbbf09a),
	.w4(32'hbb9960cc),
	.w5(32'h3bd35f1a),
	.w6(32'h3bceb7d9),
	.w7(32'h3a33364f),
	.w8(32'h3c6d796d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b624),
	.w1(32'hbb936ba7),
	.w2(32'h3bae9ac0),
	.w3(32'hbc7c25af),
	.w4(32'h3cc9ec69),
	.w5(32'hbc828078),
	.w6(32'h3c19ec60),
	.w7(32'h3d06d857),
	.w8(32'hbbbc27ef),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2791a),
	.w1(32'hbc01f78a),
	.w2(32'h3bb7dc5a),
	.w3(32'h3b999dfe),
	.w4(32'h3c140f7c),
	.w5(32'h3b1bb721),
	.w6(32'h3c1f50b7),
	.w7(32'hbbd92965),
	.w8(32'hbc4c35ec),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75e37a),
	.w1(32'hb9b8c788),
	.w2(32'hbb65775a),
	.w3(32'h3c0cb3f2),
	.w4(32'h3b334364),
	.w5(32'hba9725bc),
	.w6(32'h3bed527a),
	.w7(32'h3921ae67),
	.w8(32'h3b9c9fc5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf533fd),
	.w1(32'h382ea34d),
	.w2(32'hbbaf40c5),
	.w3(32'h3ac4a489),
	.w4(32'hbbab25b9),
	.w5(32'hbb390ddc),
	.w6(32'h3b2ad4ad),
	.w7(32'hbb79eda2),
	.w8(32'hbaa5e936),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1848b),
	.w1(32'hbc00cca6),
	.w2(32'h3b5c2da2),
	.w3(32'hbc019c6a),
	.w4(32'h3be90db2),
	.w5(32'h3a6b2c46),
	.w6(32'hbbe8eb62),
	.w7(32'h3bc995fe),
	.w8(32'h3924468e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5db9a1),
	.w1(32'hbbd7ac36),
	.w2(32'h3c42e3c9),
	.w3(32'hbbdf92a9),
	.w4(32'hbc9d1bd3),
	.w5(32'hbb002a5c),
	.w6(32'h3c3e6018),
	.w7(32'hbc654ae1),
	.w8(32'h3c08e501),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5526c1),
	.w1(32'hbb5ff392),
	.w2(32'hbbb6ada0),
	.w3(32'hbc3a125e),
	.w4(32'h3b2464a7),
	.w5(32'hbc88c206),
	.w6(32'h3c4d304c),
	.w7(32'hbbbda152),
	.w8(32'h3ae8d9cb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12d78f),
	.w1(32'h39cb49c4),
	.w2(32'hbc2292dc),
	.w3(32'hbb1ffe5b),
	.w4(32'hbb36cb7f),
	.w5(32'hbc3bfc7c),
	.w6(32'h3c15a8a5),
	.w7(32'hbc2dcec8),
	.w8(32'hbc14a83e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0817f5),
	.w1(32'h38e99d9c),
	.w2(32'hba100d17),
	.w3(32'h391c35be),
	.w4(32'hbab0b4e5),
	.w5(32'hbbd1dea9),
	.w6(32'hbc5d893b),
	.w7(32'hbb8a26be),
	.w8(32'h3d330cf4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a167466),
	.w1(32'hbb3d9176),
	.w2(32'h3c15c5ba),
	.w3(32'h3b422788),
	.w4(32'h3aa4f1b0),
	.w5(32'hbc0c7d55),
	.w6(32'h3a7dd029),
	.w7(32'hbc5aefbd),
	.w8(32'hbbd7e556),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ca645),
	.w1(32'hbb52a100),
	.w2(32'h3be3f52c),
	.w3(32'h3b031a34),
	.w4(32'hbbae98ab),
	.w5(32'h3bff5993),
	.w6(32'hbca63570),
	.w7(32'h3a1a088f),
	.w8(32'hbbb1bf07),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f6b5a),
	.w1(32'h3bb2c114),
	.w2(32'hbbf688d7),
	.w3(32'hbb63d94f),
	.w4(32'hbacc1bd8),
	.w5(32'hbbec07ee),
	.w6(32'h3b9f459c),
	.w7(32'hb98282cd),
	.w8(32'hbca25782),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56e02e),
	.w1(32'h3bd0ed01),
	.w2(32'hbba6dbf9),
	.w3(32'h3961e757),
	.w4(32'hbc62cb33),
	.w5(32'hb9f69ae7),
	.w6(32'h3c5a61fc),
	.w7(32'h3c875062),
	.w8(32'h3bcde9a4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc282196),
	.w1(32'h3b71e9de),
	.w2(32'hbb8f7f69),
	.w3(32'h39fffc01),
	.w4(32'h3c3bcc98),
	.w5(32'h3b08565a),
	.w6(32'hbb4ba47b),
	.w7(32'h3b0b8b30),
	.w8(32'hbc086d6b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf74607),
	.w1(32'h3ad349cb),
	.w2(32'h3c494c55),
	.w3(32'hbb9c9084),
	.w4(32'hbb8442dc),
	.w5(32'h3985a39a),
	.w6(32'hbb4fd4a5),
	.w7(32'h3c1db09e),
	.w8(32'hbba05fcf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc00e02),
	.w1(32'hbbc133bb),
	.w2(32'h3b67731f),
	.w3(32'hbb1b8391),
	.w4(32'h38eb0cf4),
	.w5(32'hbc0da890),
	.w6(32'h3bd1cc40),
	.w7(32'h3c393bd3),
	.w8(32'hbc61c074),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5cb4),
	.w1(32'h3c421213),
	.w2(32'hbc51f829),
	.w3(32'h3bb3f6d7),
	.w4(32'h3b3e6399),
	.w5(32'hbada77ed),
	.w6(32'hbb69bac0),
	.w7(32'hbc3eb93b),
	.w8(32'h3bbd960c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfa73b),
	.w1(32'hbc194464),
	.w2(32'h39857603),
	.w3(32'h3c039e64),
	.w4(32'hbc34d9f5),
	.w5(32'h3b87fb76),
	.w6(32'h39fe76f1),
	.w7(32'hbce152aa),
	.w8(32'hbbac5c4c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c519b),
	.w1(32'hbb885408),
	.w2(32'hbcf0921d),
	.w3(32'hbba730f6),
	.w4(32'hbbd663ee),
	.w5(32'hbbe9cbe8),
	.w6(32'h3b3bcbd8),
	.w7(32'hba9d7389),
	.w8(32'h3bb124e1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46c9dd),
	.w1(32'hbbcd3d26),
	.w2(32'hba221011),
	.w3(32'hb8e49aeb),
	.w4(32'hbc9f0b1b),
	.w5(32'h3b653026),
	.w6(32'hb9fb7179),
	.w7(32'hbc5ad2ae),
	.w8(32'h3b8f9199),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb461a2),
	.w1(32'hbb66567f),
	.w2(32'hbb133efc),
	.w3(32'h3b8900eb),
	.w4(32'hbbbb560b),
	.w5(32'h3bd9cd07),
	.w6(32'hbccfd9c9),
	.w7(32'hbbe8d582),
	.w8(32'hbbb97a22),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca97a4),
	.w1(32'h3c40586a),
	.w2(32'hbb8c2d8f),
	.w3(32'h3c05540d),
	.w4(32'hbbb1d60c),
	.w5(32'h3c66e6b8),
	.w6(32'hbc29e67c),
	.w7(32'hbbe9a889),
	.w8(32'hbad5bf60),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaafab2),
	.w1(32'h3b954b75),
	.w2(32'h3b290348),
	.w3(32'h3b7e1965),
	.w4(32'h3b1bd8bb),
	.w5(32'h3c20fd4c),
	.w6(32'h3c7bc845),
	.w7(32'h3c339aff),
	.w8(32'h3c2c0f43),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08e3ce),
	.w1(32'h3ab7bfb9),
	.w2(32'h3d17d7fe),
	.w3(32'h3ab184fd),
	.w4(32'h3c3b549e),
	.w5(32'h3bd6cc7d),
	.w6(32'h3ba0b880),
	.w7(32'hbc39b519),
	.w8(32'hbb877a46),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc309b33),
	.w1(32'h3b8c8f6f),
	.w2(32'h3b89ac6d),
	.w3(32'h3b1d69bb),
	.w4(32'h3beff5fa),
	.w5(32'hbc8e8da9),
	.w6(32'h3bdbf927),
	.w7(32'hbcdfefc0),
	.w8(32'hbba6e168),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2953de),
	.w1(32'hbc04de23),
	.w2(32'h390a304e),
	.w3(32'hbbb2de1f),
	.w4(32'h3b66570e),
	.w5(32'hbbed35fd),
	.w6(32'hbc2b937f),
	.w7(32'hba1a1fe7),
	.w8(32'h3c2a7cc0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba562c0),
	.w1(32'h3c184e7b),
	.w2(32'h3ac3f011),
	.w3(32'hbb450b39),
	.w4(32'h3b614519),
	.w5(32'h3c802f83),
	.w6(32'hbbbed718),
	.w7(32'h3b6fba2e),
	.w8(32'h35219576),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b825957),
	.w1(32'hbc1ea2d2),
	.w2(32'hbb0cf753),
	.w3(32'h3a892c04),
	.w4(32'h3a85cdf2),
	.w5(32'h3a0eccae),
	.w6(32'h3a95f930),
	.w7(32'hbaaa8b05),
	.w8(32'hbaca5fb0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128ece),
	.w1(32'h3c1a2266),
	.w2(32'hbc6ec444),
	.w3(32'h3c904e4c),
	.w4(32'hbbfca178),
	.w5(32'hbc31f164),
	.w6(32'h3be8e881),
	.w7(32'hbb722376),
	.w8(32'h3c9544e8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4c40d),
	.w1(32'hbc6ba591),
	.w2(32'h39c35bad),
	.w3(32'hbab09c72),
	.w4(32'h3b819327),
	.w5(32'h3c004820),
	.w6(32'h3c00d384),
	.w7(32'hbbb1f7b2),
	.w8(32'hbafff9bd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff57a7),
	.w1(32'h3ba09225),
	.w2(32'h3b6481b5),
	.w3(32'hba4e0d75),
	.w4(32'hbc443806),
	.w5(32'hb85b39c4),
	.w6(32'h3b1825e8),
	.w7(32'h3b00ca4d),
	.w8(32'hbbd0861a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e8f0f),
	.w1(32'h3a03f694),
	.w2(32'h3c6bdae7),
	.w3(32'hbb997eb5),
	.w4(32'hbc18ddda),
	.w5(32'h3a1eeda8),
	.w6(32'h3c355494),
	.w7(32'hbb2c0ec0),
	.w8(32'hb9264723),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1380c8),
	.w1(32'h3ba63cc4),
	.w2(32'h3c09e621),
	.w3(32'hbc4a0995),
	.w4(32'h3b4ff388),
	.w5(32'hbc60b963),
	.w6(32'hbb317abb),
	.w7(32'h3c56d990),
	.w8(32'hbc20510e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dce51),
	.w1(32'h3b8a76e8),
	.w2(32'h3c859907),
	.w3(32'h3c082aad),
	.w4(32'hbb85ccb3),
	.w5(32'hbc0731a6),
	.w6(32'hbc245138),
	.w7(32'hbc20cfaa),
	.w8(32'h3b2206d3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd71fbc),
	.w1(32'h3ccd6cab),
	.w2(32'hbb13a0fe),
	.w3(32'hbc6730f9),
	.w4(32'hbca333c2),
	.w5(32'h3c09d7b5),
	.w6(32'h3c071147),
	.w7(32'hba1fc26d),
	.w8(32'hbba2ad56),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cb1e0),
	.w1(32'hbb399a56),
	.w2(32'h3b101b2c),
	.w3(32'hbb55e97c),
	.w4(32'hbbb62406),
	.w5(32'h3be6311a),
	.w6(32'h3a398295),
	.w7(32'hbbeebe2b),
	.w8(32'hbb904827),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce2a705),
	.w1(32'h3c9cbb2d),
	.w2(32'hbc21d016),
	.w3(32'h3afd50f8),
	.w4(32'h3b0f88ab),
	.w5(32'hb91a83c1),
	.w6(32'h3a35e5ab),
	.w7(32'h3cd5a19a),
	.w8(32'h3b843b56),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a358d),
	.w1(32'h3abe5ae0),
	.w2(32'h395bb31b),
	.w3(32'hbc11f3ed),
	.w4(32'hbaf041f2),
	.w5(32'hbbdcaea0),
	.w6(32'h3b04518e),
	.w7(32'h3b6fd2b1),
	.w8(32'h3b307150),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2efb9),
	.w1(32'h3c8848ee),
	.w2(32'h3c2909d8),
	.w3(32'h3b4d0cc8),
	.w4(32'h3ba6ecd2),
	.w5(32'hbb622d91),
	.w6(32'hbc04399e),
	.w7(32'hb782502f),
	.w8(32'hbbf14ee9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b3a38),
	.w1(32'h3b5032a9),
	.w2(32'hbbd09513),
	.w3(32'hb9851f9a),
	.w4(32'h38c8d1c1),
	.w5(32'hbba3d86f),
	.w6(32'hbc61f0ca),
	.w7(32'hbc3db595),
	.w8(32'h3bad05cc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2562f8),
	.w1(32'hbc12a2ef),
	.w2(32'hbb79d521),
	.w3(32'h3c55f28c),
	.w4(32'hbb1f5322),
	.w5(32'hbb1eee1f),
	.w6(32'hbc068924),
	.w7(32'hbb655a6d),
	.w8(32'hbc4aa1d9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02c67f),
	.w1(32'h3c53f00b),
	.w2(32'h3aeabb9e),
	.w3(32'hbb64e9cf),
	.w4(32'h3c3c2a26),
	.w5(32'hbbca7416),
	.w6(32'hb7bfc7b3),
	.w7(32'h3b844055),
	.w8(32'hb9c20308),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80db91),
	.w1(32'hbc2d96db),
	.w2(32'h3c0718cf),
	.w3(32'hba9d1936),
	.w4(32'hbc82f2d7),
	.w5(32'hbc67a895),
	.w6(32'hbc2230c5),
	.w7(32'hba4e320f),
	.w8(32'h3b183403),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd6275),
	.w1(32'h39cd5fa8),
	.w2(32'hbc24ead5),
	.w3(32'hbc716ff8),
	.w4(32'h3bc987d2),
	.w5(32'hbb1266ad),
	.w6(32'hbb41c4e6),
	.w7(32'hba67d3ec),
	.w8(32'h3b41b53b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58fc34),
	.w1(32'hbb272220),
	.w2(32'hb98e903c),
	.w3(32'h39e99d2a),
	.w4(32'hbc8e488f),
	.w5(32'h3a99b9e6),
	.w6(32'h3a1eb4bf),
	.w7(32'h3a1de792),
	.w8(32'h3b9ad85d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b3630),
	.w1(32'h3bb358fa),
	.w2(32'hbb31ec9d),
	.w3(32'hbbbd85c4),
	.w4(32'hb9a76180),
	.w5(32'hbba69091),
	.w6(32'h3c0deb73),
	.w7(32'h3b6646b5),
	.w8(32'hbc97953d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12fea3),
	.w1(32'hbbbd3cd9),
	.w2(32'h3c33658c),
	.w3(32'hbbca7288),
	.w4(32'h3c7129e4),
	.w5(32'h3c1845bf),
	.w6(32'hba4c7544),
	.w7(32'h3ba83fd2),
	.w8(32'h3bcd6602),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f26a4),
	.w1(32'hbcb05a4e),
	.w2(32'hbb9d1b37),
	.w3(32'h3c38bf61),
	.w4(32'h3aa8d06b),
	.w5(32'hbbfac5d8),
	.w6(32'hbc3b87f7),
	.w7(32'hbc316f45),
	.w8(32'hba165e6e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca80d4),
	.w1(32'h3c12b068),
	.w2(32'h3b8d0410),
	.w3(32'h3c479329),
	.w4(32'h3c1aecf0),
	.w5(32'hbbea8409),
	.w6(32'hbc5ce946),
	.w7(32'h3b08ac30),
	.w8(32'hbb770d8a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54e299),
	.w1(32'hbb1101e4),
	.w2(32'hbc31deb3),
	.w3(32'hbaada192),
	.w4(32'hbc0bd238),
	.w5(32'h3ceea7ec),
	.w6(32'h3b90e8e0),
	.w7(32'hb9d2d17a),
	.w8(32'h3c44dc7d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8140c5),
	.w1(32'hb9a09c48),
	.w2(32'hbc75fe6a),
	.w3(32'h3a8d998b),
	.w4(32'hbc34bae3),
	.w5(32'hbc04a467),
	.w6(32'hbc92c518),
	.w7(32'hbc08ffa9),
	.w8(32'hbb3522e9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d65f4),
	.w1(32'hbb22814f),
	.w2(32'h3bb13119),
	.w3(32'hba0ffbcf),
	.w4(32'h3cc7ec8f),
	.w5(32'hbbaf778b),
	.w6(32'hbc27af3b),
	.w7(32'h3709b41d),
	.w8(32'h3b996c17),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc831c14),
	.w1(32'hbc12cd20),
	.w2(32'hbaa01cb1),
	.w3(32'h3c98f529),
	.w4(32'hbc7534c8),
	.w5(32'hbb9221c0),
	.w6(32'h3a13c08c),
	.w7(32'h3a25f736),
	.w8(32'h3c1cee4a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84c3b3),
	.w1(32'hbc291d11),
	.w2(32'h3ada713a),
	.w3(32'h3ba4658d),
	.w4(32'hbc5f9392),
	.w5(32'h3b37530f),
	.w6(32'h3bbee292),
	.w7(32'hbbaaab68),
	.w8(32'h3b0fecf0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aa7f6),
	.w1(32'hbbfde351),
	.w2(32'hbccd4c1b),
	.w3(32'hbaf90685),
	.w4(32'hbae5d936),
	.w5(32'h3bda59a3),
	.w6(32'hbb11ce3f),
	.w7(32'hb9cb81ba),
	.w8(32'h37d91a34),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd029c4),
	.w1(32'h39b9a2cb),
	.w2(32'hbbfc1e6e),
	.w3(32'h39958c5f),
	.w4(32'hbb82c68b),
	.w5(32'h3ca13671),
	.w6(32'hba1e41ed),
	.w7(32'hbb195f45),
	.w8(32'hbb9825db),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff2f41),
	.w1(32'hbb9357f0),
	.w2(32'h3b705e22),
	.w3(32'hbc2782c4),
	.w4(32'h3c797a25),
	.w5(32'hbbf26dba),
	.w6(32'hbb5556ee),
	.w7(32'hbcfd7040),
	.w8(32'hbafe1aa5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2460ee),
	.w1(32'hbc5c5498),
	.w2(32'h3a76e5b4),
	.w3(32'hbbe15925),
	.w4(32'h3d1faafe),
	.w5(32'hbc54d2b8),
	.w6(32'hbacce3c4),
	.w7(32'h3c034fad),
	.w8(32'hbb833eb1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd5202c),
	.w1(32'hba7468b9),
	.w2(32'h3a775e12),
	.w3(32'h3b3f9061),
	.w4(32'h3bc70ed8),
	.w5(32'h3c23555a),
	.w6(32'hbc21f185),
	.w7(32'hbb94e836),
	.w8(32'hbc07dd0b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6a52a),
	.w1(32'hbbed3df9),
	.w2(32'h3c072eda),
	.w3(32'hbafb26a6),
	.w4(32'h3bf84a4d),
	.w5(32'h3b59bcc7),
	.w6(32'hbad85cdf),
	.w7(32'hbc5ca775),
	.w8(32'hbb8fffc1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e32f9),
	.w1(32'hba96df25),
	.w2(32'hbb4dd343),
	.w3(32'hbc5c09b1),
	.w4(32'hbc8d4414),
	.w5(32'hbb38a9ee),
	.w6(32'h387e3426),
	.w7(32'h3b851b26),
	.w8(32'hbbf162d2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87f983),
	.w1(32'h3c1084ae),
	.w2(32'h3b07ab51),
	.w3(32'hbc6a0c37),
	.w4(32'h3c566110),
	.w5(32'h3bc2f128),
	.w6(32'h3d68f36a),
	.w7(32'h3b570504),
	.w8(32'hbc1233a0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba40752),
	.w1(32'h3c3ee104),
	.w2(32'h3a6e82a7),
	.w3(32'hbb6e555d),
	.w4(32'hbbfabe34),
	.w5(32'h3b59200d),
	.w6(32'hbc53c4f3),
	.w7(32'hba88e8a8),
	.w8(32'h3c214e1d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9486c3),
	.w1(32'hba5400a6),
	.w2(32'hbb565f36),
	.w3(32'hbbc5004f),
	.w4(32'hbc8e0b73),
	.w5(32'h3bdeebc2),
	.w6(32'hbc3584dc),
	.w7(32'h3aea7291),
	.w8(32'hbc4a0179),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba04964),
	.w1(32'hbc1d6f34),
	.w2(32'hbc4400b9),
	.w3(32'hbc0dec78),
	.w4(32'h389ab9db),
	.w5(32'h3bc191be),
	.w6(32'hba34fb7b),
	.w7(32'hbaecd33e),
	.w8(32'h3aed8a5f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c41ff),
	.w1(32'h3b61cd30),
	.w2(32'h3c0f580a),
	.w3(32'h3bfb72e2),
	.w4(32'hbb8ec183),
	.w5(32'h3bbf5c38),
	.w6(32'h39a4e9b1),
	.w7(32'hbba9611d),
	.w8(32'hbc1ea552),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386fcf56),
	.w1(32'hbbd50098),
	.w2(32'hbc6f606d),
	.w3(32'h39a4d232),
	.w4(32'h3bc907f6),
	.w5(32'h3a07245a),
	.w6(32'hbbbad365),
	.w7(32'hbca7ec32),
	.w8(32'h3a416561),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7d88f),
	.w1(32'h39ca7bd6),
	.w2(32'hbb62d578),
	.w3(32'h3bdf4e2a),
	.w4(32'h3b4bf2ac),
	.w5(32'hbbc04148),
	.w6(32'h3b58773a),
	.w7(32'h3a62a9e6),
	.w8(32'h39a53d13),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b804f08),
	.w1(32'hbc309234),
	.w2(32'h3c5b5c7f),
	.w3(32'h3cacfea1),
	.w4(32'h3b73c37a),
	.w5(32'h3b49f570),
	.w6(32'hbb8a833e),
	.w7(32'hbb07698b),
	.w8(32'hba2d7a6f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6356f),
	.w1(32'h3c1dcff1),
	.w2(32'hbc27f5f5),
	.w3(32'hb7993cf3),
	.w4(32'h3cd675de),
	.w5(32'h3aebb6fa),
	.w6(32'h3bfb5d24),
	.w7(32'hbbfcc941),
	.w8(32'hbaeaff39),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0467d5),
	.w1(32'h3c0ef966),
	.w2(32'hb9f264eb),
	.w3(32'hbc186d15),
	.w4(32'hba9b0690),
	.w5(32'hba36a677),
	.w6(32'hbb85e5a9),
	.w7(32'h3b16b4d5),
	.w8(32'h3ba536f5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ba22b),
	.w1(32'hbbede630),
	.w2(32'h3afcf537),
	.w3(32'h3a14c0ef),
	.w4(32'hbaeffbe8),
	.w5(32'hbbf9d488),
	.w6(32'h3c07a62f),
	.w7(32'hbbbcfef6),
	.w8(32'h3bb9fe06),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc215ea6),
	.w1(32'hbb829aab),
	.w2(32'hbbb9f159),
	.w3(32'h3c13b5f2),
	.w4(32'hbc391c17),
	.w5(32'hbcb0d900),
	.w6(32'hbbb1e7d2),
	.w7(32'hbbd535db),
	.w8(32'h3b4593d3),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30e7f6),
	.w1(32'hbb6ded91),
	.w2(32'h3b87e968),
	.w3(32'h3c1128fe),
	.w4(32'h3c4425af),
	.w5(32'hbd267952),
	.w6(32'hbb5cdf5f),
	.w7(32'hbb9679bf),
	.w8(32'h3c108dc9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10fe5a),
	.w1(32'hbb81326c),
	.w2(32'hbc7af5fa),
	.w3(32'hba9dfed7),
	.w4(32'h3bea2b4a),
	.w5(32'h3c058731),
	.w6(32'h3c2d1185),
	.w7(32'hbbef666e),
	.w8(32'h3c918be2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84029f),
	.w1(32'hbd047165),
	.w2(32'hbc8173e4),
	.w3(32'h3b2bf132),
	.w4(32'hbc187744),
	.w5(32'h3c946670),
	.w6(32'hbc773e20),
	.w7(32'h3b9c0dcc),
	.w8(32'hbbcbeb2f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2a3a8),
	.w1(32'h3b0135c0),
	.w2(32'hbb154c19),
	.w3(32'hbae445a6),
	.w4(32'hbb831a5d),
	.w5(32'hbb2d36c2),
	.w6(32'h3b7e543a),
	.w7(32'hba9181fd),
	.w8(32'hbc3c6b89),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0ee4),
	.w1(32'hbba0ebd3),
	.w2(32'hba491133),
	.w3(32'h3bb713a4),
	.w4(32'h3b5d4a74),
	.w5(32'h3bd12e23),
	.w6(32'hbc7e9584),
	.w7(32'hbb83898d),
	.w8(32'h3c012363),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb24a2),
	.w1(32'h3c399561),
	.w2(32'h3c2dda7e),
	.w3(32'h3d1f4a0c),
	.w4(32'hbb650707),
	.w5(32'hbba9eca1),
	.w6(32'hbb8d135b),
	.w7(32'hbc074f53),
	.w8(32'hbbd94310),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71423c),
	.w1(32'hbd072a9a),
	.w2(32'hbb34a582),
	.w3(32'hbad88e72),
	.w4(32'hbbacb60f),
	.w5(32'hbb69c64d),
	.w6(32'hbb1583bd),
	.w7(32'hbb93b4a1),
	.w8(32'hbae62c73),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc318606),
	.w1(32'h3c600ee3),
	.w2(32'hbccf7184),
	.w3(32'hbb825ea7),
	.w4(32'hbc38b0c0),
	.w5(32'hba88e53c),
	.w6(32'h3c47d2ad),
	.w7(32'h3ca0cc14),
	.w8(32'h3a98f86c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4db598),
	.w1(32'h3cd9a2e0),
	.w2(32'hba77e18d),
	.w3(32'hbb549738),
	.w4(32'hb86e1d79),
	.w5(32'hbc4952e4),
	.w6(32'h3cb20662),
	.w7(32'h3a834e28),
	.w8(32'hbbe0c9fd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04e909),
	.w1(32'h3c8c2433),
	.w2(32'h3bba002e),
	.w3(32'hbb910898),
	.w4(32'hbc90c019),
	.w5(32'h3b3252d9),
	.w6(32'hbca818cd),
	.w7(32'hbb14f8c5),
	.w8(32'hbb551692),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89d46),
	.w1(32'h3be5d042),
	.w2(32'h3bb9c102),
	.w3(32'hbc97762c),
	.w4(32'h3c38eb7b),
	.w5(32'h39880d0d),
	.w6(32'hbae9bb98),
	.w7(32'h3c3193e7),
	.w8(32'h3be23ca8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f33a5),
	.w1(32'h3c296c70),
	.w2(32'hbb99b757),
	.w3(32'hbbb5b70f),
	.w4(32'h3c896d8a),
	.w5(32'h3cc39584),
	.w6(32'h3bbfde7a),
	.w7(32'h3c22710f),
	.w8(32'hbb8bc14d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf2707),
	.w1(32'h3a281d71),
	.w2(32'hbb4ba03b),
	.w3(32'h3c720298),
	.w4(32'hbc78b0e8),
	.w5(32'hba306b79),
	.w6(32'hba1295f4),
	.w7(32'h3c375450),
	.w8(32'hbc87c8df),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbba81),
	.w1(32'hbc1184c3),
	.w2(32'h3cff9e85),
	.w3(32'h3b7501ed),
	.w4(32'h3b6b60ab),
	.w5(32'hbc80a7bf),
	.w6(32'hbcb9ed16),
	.w7(32'h3b7bb23a),
	.w8(32'h3c6d128c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f7e0c),
	.w1(32'hbb109d14),
	.w2(32'h3a77367e),
	.w3(32'h3b64d277),
	.w4(32'h3babdb9a),
	.w5(32'hbba3f8b9),
	.w6(32'h3c4e08d6),
	.w7(32'h3c0041c1),
	.w8(32'h3a897388),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd41fb8),
	.w1(32'h3c7b1738),
	.w2(32'h3a591a3f),
	.w3(32'hbab5520f),
	.w4(32'hbc4a59a0),
	.w5(32'h3aebff0a),
	.w6(32'hbb4b5b84),
	.w7(32'h3b5676cd),
	.w8(32'hbc02ee94),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d81c4),
	.w1(32'h3cb46231),
	.w2(32'hbc709020),
	.w3(32'hbb444e33),
	.w4(32'h3bd2d24a),
	.w5(32'h3baf4e66),
	.w6(32'h3c45c42a),
	.w7(32'hbb5b28d0),
	.w8(32'hb903ad69),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b235114),
	.w1(32'hbc9fcb73),
	.w2(32'h3b937a4d),
	.w3(32'hbbc81095),
	.w4(32'hbab58ffe),
	.w5(32'hbaeee7f8),
	.w6(32'h3c06eec8),
	.w7(32'hbb686e2b),
	.w8(32'h3c81ec39),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb928766),
	.w1(32'hb8538e60),
	.w2(32'hbbd1b382),
	.w3(32'h3c381af9),
	.w4(32'h3cebbec0),
	.w5(32'hbc44117b),
	.w6(32'h3acc2abf),
	.w7(32'hbac75a17),
	.w8(32'hbb030e4a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca850fb),
	.w1(32'h3bdf5cc5),
	.w2(32'h3c54fd94),
	.w3(32'hbb24ac90),
	.w4(32'hba8188d8),
	.w5(32'h3c25375f),
	.w6(32'h3b3d5bb6),
	.w7(32'hb8e90e3f),
	.w8(32'h3a9cc58c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23748c),
	.w1(32'h3b072d67),
	.w2(32'h39668eb4),
	.w3(32'h3cf4f014),
	.w4(32'h3c1aba9a),
	.w5(32'h3b40f7c9),
	.w6(32'hbc0c413a),
	.w7(32'hbce370dc),
	.w8(32'hbb5e7092),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce81610),
	.w1(32'hbb46460c),
	.w2(32'h3a7c7b72),
	.w3(32'hbc13e0d3),
	.w4(32'h3b89813c),
	.w5(32'h3b307727),
	.w6(32'hbae2595c),
	.w7(32'h3989c36e),
	.w8(32'hbbbdf0f8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6569d0),
	.w1(32'hba84643e),
	.w2(32'h3bf459ae),
	.w3(32'hbc375139),
	.w4(32'hbb88238c),
	.w5(32'h3c004ef0),
	.w6(32'h39f8edbc),
	.w7(32'hbb24247d),
	.w8(32'hbb699423),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c802f),
	.w1(32'hbc1c1ae3),
	.w2(32'h3b460709),
	.w3(32'hbb26b17e),
	.w4(32'h3a4251d8),
	.w5(32'h3be8d236),
	.w6(32'hbb3f5bf3),
	.w7(32'hbcc4779c),
	.w8(32'h3ad1a3e5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84661c),
	.w1(32'hbb8ddcc5),
	.w2(32'hbc04bd28),
	.w3(32'hbb5df1bf),
	.w4(32'hba307a9d),
	.w5(32'hbbed6a62),
	.w6(32'hba93f58f),
	.w7(32'hbbe84f4d),
	.w8(32'h3a9f5eda),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6cee9),
	.w1(32'hbcdafe07),
	.w2(32'hbc5b38e0),
	.w3(32'hbba777cc),
	.w4(32'hbc301443),
	.w5(32'hbb0f9436),
	.w6(32'h3b2e415d),
	.w7(32'h3c537ddf),
	.w8(32'hbbdcf88b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf06818),
	.w1(32'hbbade56f),
	.w2(32'hbb953b72),
	.w3(32'hbaf3e180),
	.w4(32'h3ba8d559),
	.w5(32'hbbd21666),
	.w6(32'h3b5d026b),
	.w7(32'hbbdf5e54),
	.w8(32'h399c1945),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcee03a),
	.w1(32'hbc98353f),
	.w2(32'hbb6c979b),
	.w3(32'hbb98de65),
	.w4(32'hbba75483),
	.w5(32'hbc41f8ce),
	.w6(32'hbc038e93),
	.w7(32'h3a3f96dd),
	.w8(32'hbb64c520),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829cdc),
	.w1(32'hba9c4245),
	.w2(32'hbcc01978),
	.w3(32'hbb3a3479),
	.w4(32'h3b378829),
	.w5(32'h3b5d84c4),
	.w6(32'hbbfc0c96),
	.w7(32'hb9b9fa0c),
	.w8(32'h3ba8abf2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf31951),
	.w1(32'hbcff46b8),
	.w2(32'hbb3b1135),
	.w3(32'h3c0a7835),
	.w4(32'h3a502c03),
	.w5(32'hbbeff7d2),
	.w6(32'hb9b15c39),
	.w7(32'h3b62d34c),
	.w8(32'h3d42c35a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b106b56),
	.w1(32'hbb2226e7),
	.w2(32'hbb8c452a),
	.w3(32'h3cdc45ce),
	.w4(32'hbb1f6e4d),
	.w5(32'hbcd6dd25),
	.w6(32'hbc0b37a6),
	.w7(32'h3be9e6d3),
	.w8(32'h3aa5f5ab),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae01daf),
	.w1(32'hbb55ecc8),
	.w2(32'hbb3e3c6f),
	.w3(32'hbbbb7627),
	.w4(32'h3c1ab6dc),
	.w5(32'hbb8687a3),
	.w6(32'hbc16efc9),
	.w7(32'h3c24e096),
	.w8(32'hbbec597f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f25a),
	.w1(32'h3ab11fbd),
	.w2(32'hbbb92cfb),
	.w3(32'hbc4b5b0a),
	.w4(32'hba5f3553),
	.w5(32'h3b68fffb),
	.w6(32'hba1bc4d1),
	.w7(32'h3a740593),
	.w8(32'h3c003af4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc694513),
	.w1(32'hbbdf0212),
	.w2(32'hbc85faad),
	.w3(32'hba8436b6),
	.w4(32'h3bfbec85),
	.w5(32'h3b0902ae),
	.w6(32'h3aa9bc02),
	.w7(32'h3bffed5f),
	.w8(32'h3c1dce72),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2abbb4),
	.w1(32'h3bf98f91),
	.w2(32'h3ba58a96),
	.w3(32'h3be6a9ca),
	.w4(32'hb9ee3fa0),
	.w5(32'hbb8363fc),
	.w6(32'hbb85daf3),
	.w7(32'h39ed7a2a),
	.w8(32'h3a6f9a3d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ee2cb),
	.w1(32'hb9f00ee9),
	.w2(32'hbc658fa3),
	.w3(32'hbbadf8f2),
	.w4(32'h3af5b449),
	.w5(32'hbb95efae),
	.w6(32'hbb5c29ff),
	.w7(32'hbc0cb941),
	.w8(32'h3a7cc60d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47cb1e),
	.w1(32'hba411abc),
	.w2(32'hbd4e136b),
	.w3(32'h3b5c0621),
	.w4(32'h3ba0dc35),
	.w5(32'h3c7a3efb),
	.w6(32'h3a59ad0f),
	.w7(32'h3b77f312),
	.w8(32'hbc63b465),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7f6c4),
	.w1(32'hbc413369),
	.w2(32'hbc36083e),
	.w3(32'hbb9d374f),
	.w4(32'h3b859ffa),
	.w5(32'hbaf81ec6),
	.w6(32'hbb82fc62),
	.w7(32'h3bc32a1c),
	.w8(32'hbb2bde9e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb27e53),
	.w1(32'hb8942e0f),
	.w2(32'h39b16533),
	.w3(32'hbc695f75),
	.w4(32'hbceb7f80),
	.w5(32'h3bab26aa),
	.w6(32'h3c36bad4),
	.w7(32'hbbe90fa6),
	.w8(32'h3a6e3975),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36a280),
	.w1(32'hbd0742d5),
	.w2(32'hbc30c844),
	.w3(32'hbd1f41d3),
	.w4(32'hbabecd48),
	.w5(32'h3abbec2c),
	.w6(32'hb974b28e),
	.w7(32'h3b8c49b4),
	.w8(32'h3b9bad3e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97bb16),
	.w1(32'h3c2bf074),
	.w2(32'h3c6e4bff),
	.w3(32'hbb5494a1),
	.w4(32'h3c1144a8),
	.w5(32'hbc885c49),
	.w6(32'h3b3e9138),
	.w7(32'hbb616c89),
	.w8(32'h3b5f7df8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9696a),
	.w1(32'hba0acd80),
	.w2(32'hbd4911ad),
	.w3(32'h3d31f703),
	.w4(32'h3be2af73),
	.w5(32'h3bd1beb9),
	.w6(32'h3b441ff5),
	.w7(32'hbcae085e),
	.w8(32'h3c2ff4d6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9c5e7),
	.w1(32'h3bc31751),
	.w2(32'h3a8fc835),
	.w3(32'h3b13e6f9),
	.w4(32'h3a474cd4),
	.w5(32'h3ba1113d),
	.w6(32'hb96cf267),
	.w7(32'hbaf3dd98),
	.w8(32'h3b68a520),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ac03),
	.w1(32'h3c2c452f),
	.w2(32'h3a3b77af),
	.w3(32'h3b8c64ba),
	.w4(32'hba88766a),
	.w5(32'h3ade4d4b),
	.w6(32'hbb740ddb),
	.w7(32'h3c5ce800),
	.w8(32'h3b94f0a8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b4116),
	.w1(32'hbc0e1835),
	.w2(32'h3be05f9a),
	.w3(32'h3865d3a6),
	.w4(32'hbc2cb59e),
	.w5(32'h3a420417),
	.w6(32'hbc179a77),
	.w7(32'hbb2db1f7),
	.w8(32'hbc860819),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84c905),
	.w1(32'hbce73b9d),
	.w2(32'h3a838af5),
	.w3(32'hbbfe0eac),
	.w4(32'hbc6660b2),
	.w5(32'h3b39ace4),
	.w6(32'h3b533c42),
	.w7(32'hbad1ba74),
	.w8(32'h3a0ae069),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26b97e),
	.w1(32'h3acdea4f),
	.w2(32'h3c786030),
	.w3(32'h3bcb4ddb),
	.w4(32'hbd141c6f),
	.w5(32'hbb42f24f),
	.w6(32'hbbf2ec2b),
	.w7(32'hba62fc8c),
	.w8(32'hbb41cc96),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d3019),
	.w1(32'hbc156359),
	.w2(32'hbad77c27),
	.w3(32'h3bc426bd),
	.w4(32'h3c308437),
	.w5(32'h3b49e188),
	.w6(32'h3bb34e45),
	.w7(32'hbabb7eb1),
	.w8(32'hbbc258d7),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d9572),
	.w1(32'hbcdff348),
	.w2(32'hbc4ec322),
	.w3(32'h3bf37390),
	.w4(32'h3c05949e),
	.w5(32'hbc40dbe0),
	.w6(32'hbcadacb8),
	.w7(32'hbbef828f),
	.w8(32'hbd2b91c9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1ea71),
	.w1(32'hba33176c),
	.w2(32'hbbe5efab),
	.w3(32'hbbef057c),
	.w4(32'h3bd4f164),
	.w5(32'hba972981),
	.w6(32'hbb03b177),
	.w7(32'h3b2570d0),
	.w8(32'hba839699),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07d1af),
	.w1(32'h3c89ebd9),
	.w2(32'hbc11c135),
	.w3(32'hbb9daa48),
	.w4(32'h3ca3be97),
	.w5(32'h3c366905),
	.w6(32'h3c3bc696),
	.w7(32'hbcc54dd5),
	.w8(32'h3ba000bf),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995b12c),
	.w1(32'hbc33558f),
	.w2(32'h3bba80a7),
	.w3(32'h3cb7a584),
	.w4(32'h3b7208a0),
	.w5(32'h3c2dcf48),
	.w6(32'hbcd74420),
	.w7(32'hbb181919),
	.w8(32'h3b4399cd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab466b4),
	.w1(32'h3b2b4961),
	.w2(32'hbb58c485),
	.w3(32'hbc6af264),
	.w4(32'h3a76029f),
	.w5(32'hbc4a1dd2),
	.w6(32'hbbb6071e),
	.w7(32'hbcf65859),
	.w8(32'hbbb7f1fc),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34f2d6),
	.w1(32'h3bba9738),
	.w2(32'h3c4acd4d),
	.w3(32'h3c98a658),
	.w4(32'hbb1db984),
	.w5(32'h3b9c2dbc),
	.w6(32'hbc4878fd),
	.w7(32'h3ab29745),
	.w8(32'hbc0eadab),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcef5a81),
	.w1(32'h3aa5b6c9),
	.w2(32'h3b0696a1),
	.w3(32'hbb033f1c),
	.w4(32'hba348ab1),
	.w5(32'hbb808716),
	.w6(32'h3b847c49),
	.w7(32'h3bbfb8ad),
	.w8(32'h39e05928),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2a08f),
	.w1(32'h3b074bec),
	.w2(32'h3b3a6104),
	.w3(32'hbc119834),
	.w4(32'hbb9534bf),
	.w5(32'hbca9ea2b),
	.w6(32'h399b6e2f),
	.w7(32'h3b912615),
	.w8(32'h3b227b0c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b155d51),
	.w1(32'hbbb6b91b),
	.w2(32'h3bb0c9ce),
	.w3(32'hbc3fa863),
	.w4(32'hb9cdb3ea),
	.w5(32'h3b819cc7),
	.w6(32'hbb968f80),
	.w7(32'hbb1989b1),
	.w8(32'h3a087eab),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909679),
	.w1(32'h3b6ea099),
	.w2(32'hbaaa3df1),
	.w3(32'h3d4be3c1),
	.w4(32'hbc1bb84d),
	.w5(32'hbdb2b181),
	.w6(32'hb9aa9ea7),
	.w7(32'h3bb836f3),
	.w8(32'h3a98499a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be58eea),
	.w1(32'h3b7bd550),
	.w2(32'h3c1b201d),
	.w3(32'h3beadf1c),
	.w4(32'hbb38cc31),
	.w5(32'h3a243e07),
	.w6(32'h3bb0cbd9),
	.w7(32'h3bd2e0f2),
	.w8(32'hba859438),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b78a0),
	.w1(32'hb9bc2077),
	.w2(32'h3ac79710),
	.w3(32'hbbbe3f81),
	.w4(32'h3b3bcb04),
	.w5(32'hbb0762fd),
	.w6(32'hbd1dd804),
	.w7(32'hbc383e4e),
	.w8(32'hbb8761b6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcff0ab),
	.w1(32'h3c219536),
	.w2(32'h3b6ac0cb),
	.w3(32'h3a530084),
	.w4(32'hb96929c2),
	.w5(32'h3b353055),
	.w6(32'hba51883e),
	.w7(32'h3a8b45bc),
	.w8(32'h3aca8dd4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c652491),
	.w1(32'h3af380f4),
	.w2(32'h3b8e58a1),
	.w3(32'h3ad1d230),
	.w4(32'h3bca31db),
	.w5(32'h3c2914b4),
	.w6(32'h3ae3c22e),
	.w7(32'h3a1149db),
	.w8(32'h3c1fb88f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85ccd6),
	.w1(32'h3b1e3ccf),
	.w2(32'hb8a2fdbd),
	.w3(32'hbc4878bb),
	.w4(32'hbb689c22),
	.w5(32'h3b415a03),
	.w6(32'h3b7ba1d9),
	.w7(32'h3c56a76f),
	.w8(32'h3c35546a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e6f14),
	.w1(32'hbb990c82),
	.w2(32'h3bbe1b58),
	.w3(32'hbaf30acf),
	.w4(32'hbc02782d),
	.w5(32'h3c274591),
	.w6(32'h3b1f58e2),
	.w7(32'h3c24027c),
	.w8(32'hbaf125d7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe346eb),
	.w1(32'h3b543eb8),
	.w2(32'hbbd6fd55),
	.w3(32'hbbce77d3),
	.w4(32'h3a4fd954),
	.w5(32'h3acaa345),
	.w6(32'hbc2001d8),
	.w7(32'hbc59b097),
	.w8(32'h3b64c22e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7eb323),
	.w1(32'h3ab68c11),
	.w2(32'h3b81aa7a),
	.w3(32'hbc4b5ab4),
	.w4(32'hb97ebc85),
	.w5(32'hbc1e58a4),
	.w6(32'h3bdbde82),
	.w7(32'hbba02835),
	.w8(32'h3be850d2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28eeda),
	.w1(32'hbbb13a48),
	.w2(32'h3bb0eeaa),
	.w3(32'hb996cd1d),
	.w4(32'hbbe55b59),
	.w5(32'h3b53c975),
	.w6(32'hba94c390),
	.w7(32'hbb06b6cb),
	.w8(32'hbda9b8f9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60f977),
	.w1(32'h3b79ab00),
	.w2(32'h38f65d66),
	.w3(32'h3be996cd),
	.w4(32'h3b3e309a),
	.w5(32'hbb8e5bbe),
	.w6(32'h3a0f0165),
	.w7(32'hbcf8a2d0),
	.w8(32'h3b00cb90),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15f0c1),
	.w1(32'h3b159776),
	.w2(32'h3c00745c),
	.w3(32'h3b6a0bc1),
	.w4(32'h3b94a411),
	.w5(32'hbbcde096),
	.w6(32'h3a02204c),
	.w7(32'h3a73b3be),
	.w8(32'hbb1e7277),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4890cf),
	.w1(32'h3be90db2),
	.w2(32'h3c616746),
	.w3(32'hbd381d58),
	.w4(32'hbb783da9),
	.w5(32'hbbf94c4b),
	.w6(32'hbb980795),
	.w7(32'hbc8b2dc8),
	.w8(32'hbb7902f7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0877ae),
	.w1(32'h3b2dea11),
	.w2(32'hbc41a5a6),
	.w3(32'hbda3b12a),
	.w4(32'h3c290384),
	.w5(32'h3b8a2099),
	.w6(32'h3afc8f81),
	.w7(32'hbab63ca9),
	.w8(32'h3a3f57b5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb133f9),
	.w1(32'h3b4a2772),
	.w2(32'hbba3645e),
	.w3(32'hbaedbb82),
	.w4(32'h3aa3deab),
	.w5(32'hbac84572),
	.w6(32'hbc121298),
	.w7(32'h3bc41b59),
	.w8(32'hbbfa3910),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a5d0c),
	.w1(32'hbada0fa8),
	.w2(32'hb91a1fd1),
	.w3(32'hbaf227d1),
	.w4(32'h3c248796),
	.w5(32'hbbeb1c1e),
	.w6(32'h3bd16fe3),
	.w7(32'hba12520e),
	.w8(32'h3aff1096),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aba5b),
	.w1(32'hbc159e87),
	.w2(32'h3bc20533),
	.w3(32'h3c130c74),
	.w4(32'hbc915630),
	.w5(32'hbc351a8a),
	.w6(32'h3bac244f),
	.w7(32'hbc66ec7d),
	.w8(32'hbb581124),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39200fab),
	.w1(32'hbba107a8),
	.w2(32'hbbf734aa),
	.w3(32'h3a93d683),
	.w4(32'h3ba25c5f),
	.w5(32'hbb4da1f6),
	.w6(32'h3b341ac8),
	.w7(32'hbad533a7),
	.w8(32'hbcbf15bf),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ff89),
	.w1(32'h3ba845f4),
	.w2(32'h3931046a),
	.w3(32'hbd7601dc),
	.w4(32'h3a93e87e),
	.w5(32'hbc6ed66d),
	.w6(32'h3b8a94af),
	.w7(32'hbb3363b9),
	.w8(32'h3b9d9964),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a757a46),
	.w1(32'hbaf59094),
	.w2(32'hbadc2ffb),
	.w3(32'h38d66637),
	.w4(32'hb9ad14ce),
	.w5(32'hba8a0ffc),
	.w6(32'h3b545e33),
	.w7(32'hb9f78787),
	.w8(32'h3c21cf4f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0907),
	.w1(32'hbc0c3996),
	.w2(32'hba287724),
	.w3(32'hbaac0adc),
	.w4(32'hb9f26d6c),
	.w5(32'h3bbfba41),
	.w6(32'hbb0358ac),
	.w7(32'h3b88418a),
	.w8(32'h3b91929f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c556e6c),
	.w1(32'h3badbd1e),
	.w2(32'h3c086056),
	.w3(32'h3a972460),
	.w4(32'hb8b975e4),
	.w5(32'h3ca8818d),
	.w6(32'hbac45ed3),
	.w7(32'h3af91d94),
	.w8(32'h3ca20775),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf87fd3),
	.w1(32'h3b93c978),
	.w2(32'hbd50ec62),
	.w3(32'hbc5ad725),
	.w4(32'hbbc98bfe),
	.w5(32'hb912cff6),
	.w6(32'h3b57c55d),
	.w7(32'h3b678e4a),
	.w8(32'h3a385fe3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf4892),
	.w1(32'h3b4612f3),
	.w2(32'hbac3113d),
	.w3(32'hbb0c469d),
	.w4(32'h3a8c2e9c),
	.w5(32'h3bb49634),
	.w6(32'h39258e3b),
	.w7(32'h39f928cc),
	.w8(32'h3b6b3294),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec84f3),
	.w1(32'hbb4809e0),
	.w2(32'hbc04cdbf),
	.w3(32'h3c4b2664),
	.w4(32'hbb735558),
	.w5(32'h3a140a01),
	.w6(32'h3bb9bd4b),
	.w7(32'hbb134361),
	.w8(32'h3a1ccaec),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b210db5),
	.w1(32'hbbb73da9),
	.w2(32'hbc17f029),
	.w3(32'h3a9b0927),
	.w4(32'h3c3f83ec),
	.w5(32'hbcde18a9),
	.w6(32'h3c8a44dd),
	.w7(32'h3b659609),
	.w8(32'h3b22e434),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25a486),
	.w1(32'h3be8cfc2),
	.w2(32'hbb8a34c0),
	.w3(32'hbc24db6c),
	.w4(32'h3a1fb77e),
	.w5(32'h3b01afca),
	.w6(32'h3b042a7b),
	.w7(32'h3bb70b5a),
	.w8(32'hbb9e19fb),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b78ea7),
	.w1(32'h3b890206),
	.w2(32'h3bd4ddb0),
	.w3(32'h3bc9d347),
	.w4(32'hbb07fff9),
	.w5(32'h3b15bdd1),
	.w6(32'h3bc68436),
	.w7(32'hbbd982cb),
	.w8(32'h3b8832f2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2096e2),
	.w1(32'hbb02d179),
	.w2(32'hbb8eb01d),
	.w3(32'h3d5b49db),
	.w4(32'h3b6d09c1),
	.w5(32'h3bda0591),
	.w6(32'h3a9ad385),
	.w7(32'hbc110d1e),
	.w8(32'hbc430ace),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eb12d),
	.w1(32'hbb2caed5),
	.w2(32'h3bc2fda0),
	.w3(32'h3c088868),
	.w4(32'h3ba06ef8),
	.w5(32'hbae685c5),
	.w6(32'hbb04c9ce),
	.w7(32'h3bd1d407),
	.w8(32'h3c04bfac),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad1b77),
	.w1(32'h3ab86d6c),
	.w2(32'hbd0a5fb2),
	.w3(32'hbabe7a7b),
	.w4(32'h3af09f3d),
	.w5(32'h3b863afc),
	.w6(32'hbc5d0d9d),
	.w7(32'hbb6a6039),
	.w8(32'h3b99400a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05cad1),
	.w1(32'h3a83f1bd),
	.w2(32'hbbaa4f5f),
	.w3(32'h3c336b9f),
	.w4(32'hbc0951a2),
	.w5(32'h3c1e908b),
	.w6(32'h3ae5dcea),
	.w7(32'hbc46f341),
	.w8(32'h38d86bfa),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5c92e),
	.w1(32'hb9cf7cd4),
	.w2(32'hbc0bb586),
	.w3(32'hbc32f25b),
	.w4(32'h3bfe7da6),
	.w5(32'h3c5a5a11),
	.w6(32'hbc1a45f4),
	.w7(32'hbcbcf8b5),
	.w8(32'hbbee890f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1ded8),
	.w1(32'h3cc95013),
	.w2(32'h3be6ae3e),
	.w3(32'hbcf4be07),
	.w4(32'h3c29efd4),
	.w5(32'hbbb0bfb0),
	.w6(32'h3bad1b60),
	.w7(32'h3c1d3b9c),
	.w8(32'h3b231f87),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e080),
	.w1(32'hbacd976d),
	.w2(32'hbc97c710),
	.w3(32'hba8a9ccc),
	.w4(32'hbbc69a7b),
	.w5(32'h3bf23a7b),
	.w6(32'h3bb62057),
	.w7(32'h3bc407e5),
	.w8(32'hbc20e13c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb014bda),
	.w1(32'hbb9e9c83),
	.w2(32'h3ad24612),
	.w3(32'hbb722fc5),
	.w4(32'h3c5e28f4),
	.w5(32'hbbb37435),
	.w6(32'h3c2316d4),
	.w7(32'h39fa3ff6),
	.w8(32'hbae1d362),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d264c),
	.w1(32'h3ca0f9ca),
	.w2(32'h3d2cb3ee),
	.w3(32'h3bbe88ee),
	.w4(32'hbbbc8069),
	.w5(32'hba52bd93),
	.w6(32'h3c99fdf4),
	.w7(32'h3b6cc40a),
	.w8(32'hb9abd01b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94e099),
	.w1(32'hbadc243f),
	.w2(32'h3c0e47f4),
	.w3(32'hbbd10cf1),
	.w4(32'h3b19113a),
	.w5(32'hbbdd107b),
	.w6(32'hbc19450c),
	.w7(32'hbca277fb),
	.w8(32'h3c7a499a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e28bb),
	.w1(32'h3a211ddd),
	.w2(32'hbc3e8364),
	.w3(32'hbc031162),
	.w4(32'hbc4683a4),
	.w5(32'hbbc26f87),
	.w6(32'h3b95a986),
	.w7(32'h3aeede4c),
	.w8(32'hba9d9a3a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbfac1c),
	.w1(32'h3bb71799),
	.w2(32'h3ba9cd7f),
	.w3(32'hb932241a),
	.w4(32'h3c4d709c),
	.w5(32'h3bfe1fa7),
	.w6(32'hbc87dae3),
	.w7(32'hbc1264e6),
	.w8(32'h3bd8a357),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b438b0b),
	.w1(32'h3cbba50c),
	.w2(32'hbc07d3d7),
	.w3(32'h3a55f55a),
	.w4(32'hbc148c7e),
	.w5(32'hbcca6f05),
	.w6(32'hbbccc091),
	.w7(32'h3bfc1dbc),
	.w8(32'h3c4d3f2c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb522b0),
	.w1(32'hbb3e4208),
	.w2(32'hbbb2a5f1),
	.w3(32'h3ba68a1c),
	.w4(32'hbc582e0a),
	.w5(32'hbc0c8b08),
	.w6(32'hbbdcf147),
	.w7(32'h3b2d5ec9),
	.w8(32'h3c5e7c2c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f772f),
	.w1(32'h3bfb7fe9),
	.w2(32'h3bdb1bd7),
	.w3(32'hbbf08ce8),
	.w4(32'h3ae63b21),
	.w5(32'hb99b0497),
	.w6(32'h3cb20b5f),
	.w7(32'h3a4af93f),
	.w8(32'h3c48c3b8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd8926),
	.w1(32'h3a7a340a),
	.w2(32'hbc0f22c3),
	.w3(32'hbc00a3f0),
	.w4(32'hbb0454d1),
	.w5(32'hbc03aea1),
	.w6(32'hbb43c79c),
	.w7(32'h39e13f5c),
	.w8(32'hbb1b323d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399273a2),
	.w1(32'h3aefe68e),
	.w2(32'h3ce71dfd),
	.w3(32'hb99be836),
	.w4(32'hbb8eb6e3),
	.w5(32'hbc0bb863),
	.w6(32'hbca66b47),
	.w7(32'h3c5b2650),
	.w8(32'hbbfb3143),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3583eb),
	.w1(32'h3bdb4ebb),
	.w2(32'hbbf4a263),
	.w3(32'h3c0daadd),
	.w4(32'hbc00e116),
	.w5(32'hbbbaecb0),
	.w6(32'hbb57878a),
	.w7(32'h3bdc1acd),
	.w8(32'hbb3a3856),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cedda5),
	.w1(32'h3d411b3a),
	.w2(32'hbbce4970),
	.w3(32'hbb3f34ef),
	.w4(32'h3c3d6db8),
	.w5(32'hbbc69057),
	.w6(32'h3b7920d9),
	.w7(32'hbc12c5b8),
	.w8(32'h3caf6f79),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95bc28),
	.w1(32'hbba4cf03),
	.w2(32'h3bb0f014),
	.w3(32'h398d1f64),
	.w4(32'h3aad6874),
	.w5(32'h3c076e64),
	.w6(32'h3bd25a40),
	.w7(32'hbc99058e),
	.w8(32'h3a4f8104),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b906805),
	.w1(32'hbb942be7),
	.w2(32'h3b1ee55f),
	.w3(32'h3bb8b8f6),
	.w4(32'h3c2e5873),
	.w5(32'hbc239c18),
	.w6(32'h3bd9a309),
	.w7(32'hbc79f60b),
	.w8(32'hbd23549f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b702df4),
	.w1(32'hbc3e1ad7),
	.w2(32'hbaa50d9e),
	.w3(32'h35682a7a),
	.w4(32'hbc9fde40),
	.w5(32'h3b9679de),
	.w6(32'h3ba2b2ea),
	.w7(32'h3c903bb3),
	.w8(32'hba011e15),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b500f48),
	.w1(32'h3c6933d0),
	.w2(32'hbb2f91d6),
	.w3(32'hba37d264),
	.w4(32'hbb841a78),
	.w5(32'h3ba53caa),
	.w6(32'hbbe6789e),
	.w7(32'h3b0eab60),
	.w8(32'hbb7a76e9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a332f),
	.w1(32'h3a226322),
	.w2(32'hbb45d7d4),
	.w3(32'h3c0105b1),
	.w4(32'hbbf56d94),
	.w5(32'h3b88231d),
	.w6(32'h3c27ce93),
	.w7(32'h3939ad71),
	.w8(32'h3c7c82b0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba51416),
	.w1(32'h3b9b16b1),
	.w2(32'h3b172d72),
	.w3(32'h3bb48534),
	.w4(32'hbbcfd209),
	.w5(32'h3ab04237),
	.w6(32'h3cd73683),
	.w7(32'hbbc5d2b7),
	.w8(32'h3b02397c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c83a9),
	.w1(32'hba632ad7),
	.w2(32'hbd176b08),
	.w3(32'hbbeb93fb),
	.w4(32'hbb18bc00),
	.w5(32'hbba0c5be),
	.w6(32'h3bc0f380),
	.w7(32'hbc0379a6),
	.w8(32'hbb47d872),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77931e),
	.w1(32'h3b862529),
	.w2(32'h3bbc0cb8),
	.w3(32'hbbfa836f),
	.w4(32'h3aeacd38),
	.w5(32'h3b81fd7b),
	.w6(32'hbbb1dd2e),
	.w7(32'hbc05d5f3),
	.w8(32'hbc917ce4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcfaed),
	.w1(32'h3c13a65c),
	.w2(32'hbb87bd43),
	.w3(32'h3b4558e8),
	.w4(32'hbafaef14),
	.w5(32'h3aab03c0),
	.w6(32'hbcc25481),
	.w7(32'hbb34e228),
	.w8(32'hbb038c12),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule