module layer_8_featuremap_37(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e36f5),
	.w1(32'hbb62bee6),
	.w2(32'hba9ffb04),
	.w3(32'hbbf06ae5),
	.w4(32'hbc343bb6),
	.w5(32'hbbcd30fa),
	.w6(32'hbc07f302),
	.w7(32'hbb8c4a4d),
	.w8(32'h3b2b4acc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ecb1c),
	.w1(32'h391ab808),
	.w2(32'hb9e8e92d),
	.w3(32'hbbc5f5e8),
	.w4(32'hbb02b226),
	.w5(32'hbb2d49fe),
	.w6(32'hbb320b45),
	.w7(32'h398a5f00),
	.w8(32'hbbd38450),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f3a6),
	.w1(32'h3b6fb3e3),
	.w2(32'h3a977645),
	.w3(32'hbbaa1b41),
	.w4(32'h3bb5ab56),
	.w5(32'h3a2adf87),
	.w6(32'hbba74ac0),
	.w7(32'h3b5aa8e5),
	.w8(32'hbb474bfd),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81b706),
	.w1(32'h3a86572d),
	.w2(32'hbcaa0329),
	.w3(32'hbb6b093e),
	.w4(32'h3bd38c3d),
	.w5(32'hbc629b29),
	.w6(32'hbc32544c),
	.w7(32'hbbe80338),
	.w8(32'hbc517f02),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71660),
	.w1(32'hba67c5c3),
	.w2(32'hbc0f3a6b),
	.w3(32'hbc4ccad7),
	.w4(32'hbb9fef17),
	.w5(32'hbc51e8d3),
	.w6(32'hbb6accd2),
	.w7(32'hbba0f3e0),
	.w8(32'hbb880b8e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7d23b),
	.w1(32'hbc2a0bcc),
	.w2(32'hbd26b53f),
	.w3(32'hbd204c79),
	.w4(32'hbcf0b681),
	.w5(32'hbcff45aa),
	.w6(32'hbc976807),
	.w7(32'hbca07137),
	.w8(32'hbc19c7a7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dacdae),
	.w1(32'hbad210dd),
	.w2(32'h3ad780b1),
	.w3(32'hbb0540ab),
	.w4(32'hbb232a94),
	.w5(32'hbb2793c1),
	.w6(32'h3a972e1d),
	.w7(32'hba4fed55),
	.w8(32'hba105a9b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc466e35),
	.w1(32'h3b452ff4),
	.w2(32'hbc1220d1),
	.w3(32'hbcb948a4),
	.w4(32'hbc340ae4),
	.w5(32'hbc9aa018),
	.w6(32'hbc45e738),
	.w7(32'hbb85b99a),
	.w8(32'hbc01cb38),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf57abf),
	.w1(32'hbc265e05),
	.w2(32'hba23cc4b),
	.w3(32'hbc3d5b09),
	.w4(32'hbc2ff76d),
	.w5(32'hbc1649c3),
	.w6(32'hbc0caa4a),
	.w7(32'hbc11165c),
	.w8(32'hbb9c155f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1181b3),
	.w1(32'h3ca17957),
	.w2(32'hbc15d44c),
	.w3(32'h3b46678d),
	.w4(32'h3b6b7ca7),
	.w5(32'hbc0c4daf),
	.w6(32'h3b467425),
	.w7(32'hba16e7d8),
	.w8(32'hbb9af5d1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92c3f7),
	.w1(32'h3be7059b),
	.w2(32'h3aae2f9e),
	.w3(32'hbbed2697),
	.w4(32'hbb45dc09),
	.w5(32'hbc4a18bf),
	.w6(32'hbb972e1d),
	.w7(32'hbb5df9fa),
	.w8(32'hba8d7adb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9b0f),
	.w1(32'hbc0e2fa3),
	.w2(32'hbc46d7e8),
	.w3(32'hbc13f5e1),
	.w4(32'hbbbb4ce2),
	.w5(32'hbc411bd4),
	.w6(32'hbbf1f088),
	.w7(32'hbba9b2f1),
	.w8(32'hbc49750d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ed210),
	.w1(32'h3b3c821e),
	.w2(32'hbb51379a),
	.w3(32'hbc484cfd),
	.w4(32'h3b0de50f),
	.w5(32'hbc05a628),
	.w6(32'hbc28f281),
	.w7(32'hbacd4e57),
	.w8(32'hbba7c9a0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d053),
	.w1(32'hbbe96d21),
	.w2(32'hbd2e00b4),
	.w3(32'hbcd29e53),
	.w4(32'hbd2926e8),
	.w5(32'hbd086865),
	.w6(32'hba681602),
	.w7(32'hbce30d22),
	.w8(32'hb9bca678),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362b55b9),
	.w1(32'hbba1575f),
	.w2(32'hbc3a3ff8),
	.w3(32'hbbed8259),
	.w4(32'hbc296dee),
	.w5(32'hbc0a811c),
	.w6(32'hbad3c2bb),
	.w7(32'hbc0b2883),
	.w8(32'h3b8e334c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27b072),
	.w1(32'h3b19886f),
	.w2(32'h3b660fa5),
	.w3(32'h3a0187e4),
	.w4(32'hbbc564c2),
	.w5(32'hbac4b3bd),
	.w6(32'h3a01508b),
	.w7(32'hbae1b8a1),
	.w8(32'h3c2f3228),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88e83f),
	.w1(32'h3c31d855),
	.w2(32'hbcad021f),
	.w3(32'hbbf62c61),
	.w4(32'hbb8d10b2),
	.w5(32'hbbabd658),
	.w6(32'h3c9b2477),
	.w7(32'hbc883fd8),
	.w8(32'h3a8895b9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0f89),
	.w1(32'h3bcb4706),
	.w2(32'hbbf21f89),
	.w3(32'hbc2577c3),
	.w4(32'h3b12dd51),
	.w5(32'hbc17c8d5),
	.w6(32'hbc098682),
	.w7(32'h3b0cdd5c),
	.w8(32'hbb84dde2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee4be3),
	.w1(32'h3c4178ab),
	.w2(32'hbbb1d796),
	.w3(32'hbd06068f),
	.w4(32'hbc184f80),
	.w5(32'hbce926d9),
	.w6(32'hbd1ae892),
	.w7(32'hbb544a9b),
	.w8(32'h3c82ffa3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f013e),
	.w1(32'h3c57c87c),
	.w2(32'hbccd5221),
	.w3(32'hbd1349fb),
	.w4(32'hbbf5caf8),
	.w5(32'hbcaa56e3),
	.w6(32'hbc8a17bf),
	.w7(32'hbb9b8f7b),
	.w8(32'hbca11a96),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05e298),
	.w1(32'h3803c804),
	.w2(32'hba980c9b),
	.w3(32'hbc45ff01),
	.w4(32'hbc75c98b),
	.w5(32'hbc54a301),
	.w6(32'hbc08cf3d),
	.w7(32'hbad8172a),
	.w8(32'hbb687974),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22717c),
	.w1(32'h3c3f9e6c),
	.w2(32'hb94ae7ed),
	.w3(32'h39625548),
	.w4(32'h3c06da37),
	.w5(32'hbb7d80aa),
	.w6(32'h3b5ad563),
	.w7(32'h3b4c0810),
	.w8(32'hbb96b182),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd1e7b),
	.w1(32'hba7d3805),
	.w2(32'hbd16cf6f),
	.w3(32'hbcf8d568),
	.w4(32'hbd6b044e),
	.w5(32'hbd2632e2),
	.w6(32'hbc4e1d5f),
	.w7(32'hbcb36d6a),
	.w8(32'h3c903685),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa563fb),
	.w1(32'h3ba2fd04),
	.w2(32'h3b15cfc3),
	.w3(32'hbc1be222),
	.w4(32'hbc08a332),
	.w5(32'hbc05e1ca),
	.w6(32'hbbbc772a),
	.w7(32'hbbb81258),
	.w8(32'h3b878957),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3341d6),
	.w1(32'h3c60c217),
	.w2(32'hbb022706),
	.w3(32'hbb8b12a6),
	.w4(32'hbc3f8b04),
	.w5(32'hbb8e2c99),
	.w6(32'h3af27f6c),
	.w7(32'hbb198799),
	.w8(32'hbb5a4047),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d723c),
	.w1(32'hbc1bed86),
	.w2(32'hbd5b97c1),
	.w3(32'hbd1277bb),
	.w4(32'hbd595bf0),
	.w5(32'hbd4d8265),
	.w6(32'hbc8a8dc6),
	.w7(32'hbcea61f1),
	.w8(32'hbc2a4588),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5fd45),
	.w1(32'hbaad95c4),
	.w2(32'hbd11e439),
	.w3(32'hbc900680),
	.w4(32'hbd08d33f),
	.w5(32'hbcdc7c98),
	.w6(32'hbbbfbe52),
	.w7(32'hbc914f88),
	.w8(32'h3bf35734),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3c24fa),
	.w1(32'h3c998fc2),
	.w2(32'h3b789060),
	.w3(32'hbd95ff99),
	.w4(32'hbca6e709),
	.w5(32'hbd996adf),
	.w6(32'hbda3195d),
	.w7(32'hbd68982c),
	.w8(32'hbd6ddfce),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58bb4e),
	.w1(32'h3b3b42ea),
	.w2(32'h3b576089),
	.w3(32'hbc708ac0),
	.w4(32'hbcf4a635),
	.w5(32'hbca1f294),
	.w6(32'hbc670270),
	.w7(32'hbbeb309d),
	.w8(32'hbb476772),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706411),
	.w1(32'hbaaffdec),
	.w2(32'h39716875),
	.w3(32'hbaf4c57d),
	.w4(32'h3acf6334),
	.w5(32'hbaeb4b5e),
	.w6(32'hbb44924b),
	.w7(32'hba78af50),
	.w8(32'h3c14a796),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b142f),
	.w1(32'h3c5ad86b),
	.w2(32'hbca6f105),
	.w3(32'h3acaec04),
	.w4(32'h3b647f19),
	.w5(32'hbc103cc0),
	.w6(32'h3cc11c9c),
	.w7(32'hbc33c53f),
	.w8(32'hbb8863cd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29cc17),
	.w1(32'h3bf2eae0),
	.w2(32'hbbe12205),
	.w3(32'hbc147cd6),
	.w4(32'hbc198411),
	.w5(32'hbc32ed97),
	.w6(32'hbc6c63b7),
	.w7(32'h3a334878),
	.w8(32'hbb034f15),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f276),
	.w1(32'hbb18dc74),
	.w2(32'hbc5e2360),
	.w3(32'hbadb6679),
	.w4(32'h3b9faa17),
	.w5(32'hbc1b3493),
	.w6(32'h3c387717),
	.w7(32'hbbd83f6f),
	.w8(32'hbb9ea8d3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb65116),
	.w1(32'h3b0f6456),
	.w2(32'hbb1a117a),
	.w3(32'hbaf2572f),
	.w4(32'h3b8d38b4),
	.w5(32'h3b9d6acd),
	.w6(32'hbbb8072f),
	.w7(32'hbbe0b55d),
	.w8(32'h3b4289be),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf91eb4),
	.w1(32'h3be8c544),
	.w2(32'hbd22421e),
	.w3(32'hbd0da9c3),
	.w4(32'hbcc3cf28),
	.w5(32'hbd06c1fe),
	.w6(32'hbc6617b0),
	.w7(32'hbc7839d4),
	.w8(32'hbbbd4b86),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86bb98),
	.w1(32'h3b702100),
	.w2(32'h3b8da643),
	.w3(32'hbc3f0c98),
	.w4(32'hbbfc01c1),
	.w5(32'hbbf3383d),
	.w6(32'hbc00a15f),
	.w7(32'hbb013921),
	.w8(32'h3c4a1c5d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9158f),
	.w1(32'h3c42feac),
	.w2(32'hbb9716fc),
	.w3(32'hbbe677d2),
	.w4(32'hbc10f36f),
	.w5(32'hbbcd9430),
	.w6(32'h3b35c3d2),
	.w7(32'hbba9b0c4),
	.w8(32'hbb091412),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1633fb),
	.w1(32'h3a1ac2df),
	.w2(32'h3b086e9a),
	.w3(32'h3af78519),
	.w4(32'h3accfdb3),
	.w5(32'hbb0e07a4),
	.w6(32'h3b48b553),
	.w7(32'h3b16c56e),
	.w8(32'hba13035b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57009e),
	.w1(32'hbbe20e06),
	.w2(32'hbc93ec91),
	.w3(32'hbc3dbe59),
	.w4(32'hbc712454),
	.w5(32'hbc6b104b),
	.w6(32'hbb3ade86),
	.w7(32'hbc6de9fb),
	.w8(32'h3c3b8cc7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ae2fe),
	.w1(32'h3c3a2d79),
	.w2(32'hb976bede),
	.w3(32'h3af122ff),
	.w4(32'hbb913596),
	.w5(32'hbb160169),
	.w6(32'h3badd3b1),
	.w7(32'hb9f1ad2f),
	.w8(32'hba83cede),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7e3d00),
	.w1(32'hbca37e34),
	.w2(32'hbd60eee6),
	.w3(32'hbda643e9),
	.w4(32'hbd06ede4),
	.w5(32'hbd5b3165),
	.w6(32'hbdab9120),
	.w7(32'hbcf2a678),
	.w8(32'hbd29a5bd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5700e),
	.w1(32'h3b8a9c63),
	.w2(32'hbb2bc9de),
	.w3(32'hbc937dca),
	.w4(32'hbc89f73a),
	.w5(32'hbbfbe24f),
	.w6(32'hbab6ea73),
	.w7(32'h3bbf5b1d),
	.w8(32'h3af20ffa),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7fe65),
	.w1(32'hbbb2328f),
	.w2(32'h3a9c3b04),
	.w3(32'h3be36b72),
	.w4(32'h3cd00f4b),
	.w5(32'hbc8e6d58),
	.w6(32'hbc6cbfa1),
	.w7(32'h3cd93131),
	.w8(32'h3bd14e03),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ba27f),
	.w1(32'hbb82c425),
	.w2(32'hbb2f390f),
	.w3(32'hbcb92bf7),
	.w4(32'hbcdbb82f),
	.w5(32'hbc65225c),
	.w6(32'h3b85ab64),
	.w7(32'h37c39260),
	.w8(32'h3c7f92b3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fc281),
	.w1(32'h3b531c52),
	.w2(32'hbbe9f741),
	.w3(32'hbc93fb7a),
	.w4(32'hbcea96af),
	.w5(32'hbcf818ba),
	.w6(32'h3ca25f58),
	.w7(32'h3c969448),
	.w8(32'hb9fdd941),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7652c4),
	.w1(32'hbbca1f7c),
	.w2(32'hbbb1aa49),
	.w3(32'hbcd0ee06),
	.w4(32'hbc9081ea),
	.w5(32'hbc6bddcc),
	.w6(32'h3a6f7310),
	.w7(32'h3c1cf03f),
	.w8(32'hbc09f341),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e6e6f),
	.w1(32'hbc0a7fe9),
	.w2(32'h3c14320d),
	.w3(32'hbc467e59),
	.w4(32'hbb344850),
	.w5(32'h3a4ccba4),
	.w6(32'h3a2996c1),
	.w7(32'h3c95a3ed),
	.w8(32'h3bfcb4eb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b480e5e),
	.w1(32'hbbd96c5b),
	.w2(32'hbcb9e532),
	.w3(32'hbc572574),
	.w4(32'hbd0fb33a),
	.w5(32'hbcc0015e),
	.w6(32'h3b836e43),
	.w7(32'hbc425d29),
	.w8(32'hbc6f8bea),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c45a5),
	.w1(32'h3b5572e7),
	.w2(32'hbc040694),
	.w3(32'h3c122f1a),
	.w4(32'h3d41266b),
	.w5(32'h3c883885),
	.w6(32'hbd53900d),
	.w7(32'hbc936e65),
	.w8(32'h3c75125a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d44c9),
	.w1(32'h3ba44183),
	.w2(32'hbbe0ff99),
	.w3(32'hbc855971),
	.w4(32'hbce23121),
	.w5(32'hbcd8aa6d),
	.w6(32'h3c689fca),
	.w7(32'h3c0cf33c),
	.w8(32'h3b578444),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40dc0d),
	.w1(32'hb9af9180),
	.w2(32'hbc53dead),
	.w3(32'hbc2e85e4),
	.w4(32'hbc98ff2f),
	.w5(32'hbcefaefc),
	.w6(32'h3c6e6ea8),
	.w7(32'h3af80059),
	.w8(32'hbc20251a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd26863f),
	.w1(32'hbb240897),
	.w2(32'hbc26005e),
	.w3(32'hbd924814),
	.w4(32'hbd4a2434),
	.w5(32'hbd2c49fc),
	.w6(32'hbc7e4b94),
	.w7(32'h3c3f48c8),
	.w8(32'hbc0e5944),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bb0d5),
	.w1(32'hbc960777),
	.w2(32'hbc0e7295),
	.w3(32'hbcce197e),
	.w4(32'hbcfa9d12),
	.w5(32'hbc0da60a),
	.w6(32'hbc1edfaf),
	.w7(32'hbb97a104),
	.w8(32'h3b1613eb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b3239),
	.w1(32'h3c073550),
	.w2(32'h3b0b836d),
	.w3(32'hbc866092),
	.w4(32'hbae62e4c),
	.w5(32'hbc23e35a),
	.w6(32'h3a994b7a),
	.w7(32'h3c6a924e),
	.w8(32'hbbae7c63),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c490e4a),
	.w1(32'hbb19d8c4),
	.w2(32'h3bdb1481),
	.w3(32'h3c93cc4d),
	.w4(32'hbc9b3d34),
	.w5(32'hbc2dcf8e),
	.w6(32'h3bff4cd5),
	.w7(32'h3c91a88f),
	.w8(32'hbc02231c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fefb5),
	.w1(32'hbc686ede),
	.w2(32'hbca71541),
	.w3(32'hbbafbd70),
	.w4(32'hbc7f3de8),
	.w5(32'hbc2b2577),
	.w6(32'hbc478e72),
	.w7(32'hbccde6d3),
	.w8(32'hbbddd2e8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb442f0),
	.w1(32'h3c031061),
	.w2(32'h3be07f1e),
	.w3(32'hbc9b4592),
	.w4(32'hbc1a4335),
	.w5(32'h3bb3e050),
	.w6(32'h3a2fa139),
	.w7(32'hbb93249a),
	.w8(32'hbc903d57),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab5bf6),
	.w1(32'h3c6f6970),
	.w2(32'hbc02c50c),
	.w3(32'hbc775c96),
	.w4(32'h3ac0c0be),
	.w5(32'hbc37aa6a),
	.w6(32'hbbfdc155),
	.w7(32'h3c397bdd),
	.w8(32'h3b174dc0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8a185),
	.w1(32'hba00b000),
	.w2(32'hbb241ef8),
	.w3(32'h3b93b353),
	.w4(32'h3c3b00c3),
	.w5(32'h3c0d4110),
	.w6(32'h3c653965),
	.w7(32'h3b139a70),
	.w8(32'h3ca56115),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb773220),
	.w1(32'hbbe80949),
	.w2(32'hbbbe83e0),
	.w3(32'hbc8b72bd),
	.w4(32'hbc86118f),
	.w5(32'hbc9a0a1c),
	.w6(32'hbc40b653),
	.w7(32'h3c17ae58),
	.w8(32'hbc17dee7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcacb4),
	.w1(32'hbcac008d),
	.w2(32'hbbe53a85),
	.w3(32'hbc82d712),
	.w4(32'hbc814b6b),
	.w5(32'hbae22a03),
	.w6(32'hbc987e86),
	.w7(32'hbaa78268),
	.w8(32'hbb8c936c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48d208),
	.w1(32'hbbb540a7),
	.w2(32'hbc5d84e8),
	.w3(32'hbc7ce190),
	.w4(32'hbcaa9f6a),
	.w5(32'hbc642721),
	.w6(32'h3bad6243),
	.w7(32'hbb975de3),
	.w8(32'h3cf8efb7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78960e),
	.w1(32'h3b221c6a),
	.w2(32'hbc4368a1),
	.w3(32'hbd3189f4),
	.w4(32'hbcad041f),
	.w5(32'hbcd9f800),
	.w6(32'h3bec634e),
	.w7(32'h3cfa1de8),
	.w8(32'hbca72da5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d45d5),
	.w1(32'h3c43491f),
	.w2(32'h3bf2715c),
	.w3(32'hbc46d52b),
	.w4(32'hbb3de002),
	.w5(32'h3c0c8d71),
	.w6(32'hb9a95072),
	.w7(32'h3be8058f),
	.w8(32'h3c62f10b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c7ba),
	.w1(32'h39d18534),
	.w2(32'h39b1de3f),
	.w3(32'hbbc2fe85),
	.w4(32'hbc9535cb),
	.w5(32'hbc1ed913),
	.w6(32'h3c96f5cb),
	.w7(32'h3b9951f8),
	.w8(32'h37c3d85e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc110228),
	.w1(32'hbb09daab),
	.w2(32'hba90af7d),
	.w3(32'hbc77b9ba),
	.w4(32'hbc740b82),
	.w5(32'hbbe6cf6f),
	.w6(32'hba7ae179),
	.w7(32'h3b0f7a27),
	.w8(32'h3b75a3eb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc96c66),
	.w1(32'hba7c82e6),
	.w2(32'hbc0c7fd9),
	.w3(32'hbc7125b7),
	.w4(32'hbc102698),
	.w5(32'hbc51be9e),
	.w6(32'h39872b40),
	.w7(32'h3b793ab7),
	.w8(32'hbc81c7d0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdeb43c),
	.w1(32'hbc8d1632),
	.w2(32'hbccd7403),
	.w3(32'hbbd973c3),
	.w4(32'h3ba3555e),
	.w5(32'h3c278a35),
	.w6(32'hbc15e733),
	.w7(32'hbc3ab307),
	.w8(32'h3c0c8ee7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbffa96),
	.w1(32'h3b9448ad),
	.w2(32'h392d309c),
	.w3(32'hbc06d203),
	.w4(32'hbca21fa1),
	.w5(32'hbc70daba),
	.w6(32'h3cc00d8c),
	.w7(32'h3c3a7ae9),
	.w8(32'h3cf36d7a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbebbe),
	.w1(32'hbb5bfb87),
	.w2(32'hbc25ffea),
	.w3(32'hbd151635),
	.w4(32'hbd216445),
	.w5(32'hbcf8b7ab),
	.w6(32'h3d283a43),
	.w7(32'h3c537803),
	.w8(32'h3b1ce51c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba01a10),
	.w1(32'h3b584261),
	.w2(32'h3a3bfc31),
	.w3(32'hbb894a4f),
	.w4(32'hbc5c5a70),
	.w5(32'hbbb67624),
	.w6(32'h3c485794),
	.w7(32'h3ba2311e),
	.w8(32'h3c869ace),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da39e),
	.w1(32'h3bb510cb),
	.w2(32'hbc112fdf),
	.w3(32'hbcca1b4e),
	.w4(32'hbcc625c6),
	.w5(32'hbcd72d8d),
	.w6(32'h3c44775f),
	.w7(32'h3c0ec7ac),
	.w8(32'hbb546576),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba89156),
	.w1(32'h3ae63207),
	.w2(32'hb9e7d086),
	.w3(32'hbc0f56c5),
	.w4(32'hbcaaff1d),
	.w5(32'hbc34d93e),
	.w6(32'h3c7dd09f),
	.w7(32'h3bf13e23),
	.w8(32'hb9e3f216),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d02d6),
	.w1(32'hbca6b566),
	.w2(32'hbd00c67b),
	.w3(32'hbc834b2d),
	.w4(32'hbce33f3f),
	.w5(32'hbd09f92d),
	.w6(32'hbc9e9870),
	.w7(32'hbc6f14aa),
	.w8(32'hb9e064ba),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a921d1a),
	.w1(32'hbac257e3),
	.w2(32'hbbf54e53),
	.w3(32'hbc9187b2),
	.w4(32'hbcc83fcd),
	.w5(32'hbc965401),
	.w6(32'h3ca96ca6),
	.w7(32'h3c033198),
	.w8(32'h3b915d33),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b8c17),
	.w1(32'h3ba6a2fc),
	.w2(32'h3a94b446),
	.w3(32'hbc55cf85),
	.w4(32'hbc5411c3),
	.w5(32'hbc06ae70),
	.w6(32'h3c5acddc),
	.w7(32'h3c41b112),
	.w8(32'h3bd9727e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94540c),
	.w1(32'hbb427fdc),
	.w2(32'hbb990d99),
	.w3(32'hbc37ea5d),
	.w4(32'hbca6fce2),
	.w5(32'hbc2c48a8),
	.w6(32'h3c3dc530),
	.w7(32'h3bb987cc),
	.w8(32'h3d047dc5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc16d8),
	.w1(32'hbbc8b067),
	.w2(32'hbcad23eb),
	.w3(32'hbd0feeaa),
	.w4(32'hbd22382f),
	.w5(32'hbce663b2),
	.w6(32'h3d64abff),
	.w7(32'h3cb71b33),
	.w8(32'h3c19396b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25b7e3),
	.w1(32'hbaf2e89e),
	.w2(32'hbb561b0a),
	.w3(32'hbcaaa7bf),
	.w4(32'hbceef989),
	.w5(32'hbc0ca34c),
	.w6(32'h3d2c1587),
	.w7(32'h3ca678fc),
	.w8(32'h3c8be3ed),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a8798),
	.w1(32'hbbbbd9bd),
	.w2(32'hbab18555),
	.w3(32'hbb49d803),
	.w4(32'hbc1ebeeb),
	.w5(32'h3b1e8df3),
	.w6(32'h3c59c323),
	.w7(32'h3a691ff0),
	.w8(32'h3b9391f1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9e891),
	.w1(32'hbc730f6d),
	.w2(32'hbc9ea3bb),
	.w3(32'hbce1d457),
	.w4(32'hbce792c4),
	.w5(32'hbcded0a2),
	.w6(32'h3bdd2915),
	.w7(32'h3ca31704),
	.w8(32'h3bc5e810),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56a2ae),
	.w1(32'h3a1de49d),
	.w2(32'hbacb5aa5),
	.w3(32'hbc96a79a),
	.w4(32'hbc8cc4ed),
	.w5(32'hbc508a3f),
	.w6(32'h3bbb819c),
	.w7(32'h3c4d915a),
	.w8(32'h3c5aac83),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8428c6),
	.w1(32'hbb8521cf),
	.w2(32'hbc931226),
	.w3(32'hbd3c0e53),
	.w4(32'hbd4f268b),
	.w5(32'hbd2765ab),
	.w6(32'h3bababf0),
	.w7(32'h3b9e497e),
	.w8(32'hbc94698e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd86988a),
	.w1(32'hbc70aab2),
	.w2(32'hbd7a5753),
	.w3(32'hbda26e27),
	.w4(32'hbcb80c99),
	.w5(32'hbd6a6499),
	.w6(32'hbd979eaa),
	.w7(32'hbca886fe),
	.w8(32'hbd35186c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd22229),
	.w1(32'hbb1066b1),
	.w2(32'hbcb2eed4),
	.w3(32'hbd413014),
	.w4(32'hbcc35bca),
	.w5(32'hbd35fb09),
	.w6(32'hbd15f09b),
	.w7(32'hb9ea1c3d),
	.w8(32'hbb3f1a81),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac55f9),
	.w1(32'hbba33d23),
	.w2(32'hbc330e01),
	.w3(32'hbc85fc48),
	.w4(32'hbd0c7338),
	.w5(32'hbccfd25c),
	.w6(32'h3cc29137),
	.w7(32'h3c39292a),
	.w8(32'hbd0805ee),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbede567),
	.w1(32'h3aa4b152),
	.w2(32'hbc041ab9),
	.w3(32'h3cf4ca9b),
	.w4(32'h3d7a67e9),
	.w5(32'h3cd7815a),
	.w6(32'hbd508bed),
	.w7(32'hbcd03332),
	.w8(32'h3c38c0a2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca47e7),
	.w1(32'h3adf7c78),
	.w2(32'h3bd7e292),
	.w3(32'hbc1505e3),
	.w4(32'hbcd5855b),
	.w5(32'hbb6ae96a),
	.w6(32'h3ccd640a),
	.w7(32'h3c1edf6e),
	.w8(32'h3cac5099),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d67fe),
	.w1(32'hba852cc0),
	.w2(32'hbab5b9e7),
	.w3(32'hbc2b9c2e),
	.w4(32'hbc724df6),
	.w5(32'hbc741a6d),
	.w6(32'h3c29d751),
	.w7(32'h3ca0316f),
	.w8(32'hbcdad158),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb32fb2),
	.w1(32'hbaccdc1b),
	.w2(32'hbc1d97e0),
	.w3(32'h3cd15309),
	.w4(32'h3d4f8d85),
	.w5(32'h3c98136d),
	.w6(32'hbd440715),
	.w7(32'hbcef3cdc),
	.w8(32'hbce888dd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc939d49),
	.w1(32'h39abb518),
	.w2(32'hbc6f8c72),
	.w3(32'h3c371f77),
	.w4(32'h3d37ca25),
	.w5(32'h3c3e6217),
	.w6(32'hbd5412df),
	.w7(32'hbccba308),
	.w8(32'h3a5a367b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a868413),
	.w1(32'hb9a46e64),
	.w2(32'hbb7f4c23),
	.w3(32'hbc248747),
	.w4(32'hbbd34642),
	.w5(32'hbc6ee0f6),
	.w6(32'h3b855e1d),
	.w7(32'h3c0ef882),
	.w8(32'h3b858130),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc531fd4),
	.w1(32'h3aff3260),
	.w2(32'h3b0d50f0),
	.w3(32'hbcc390cd),
	.w4(32'hbca970e0),
	.w5(32'hbb82850f),
	.w6(32'h3b83c8c7),
	.w7(32'hbc3409c8),
	.w8(32'hbc36acbc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd8370),
	.w1(32'h3a970f9b),
	.w2(32'hbb3b89c1),
	.w3(32'hbc7c9d31),
	.w4(32'hbc35c3b0),
	.w5(32'hbc30aef0),
	.w6(32'hbadb6c53),
	.w7(32'h3b9333e9),
	.w8(32'hbb85b121),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc353ca),
	.w1(32'h3c9bcabb),
	.w2(32'h3c2c4b9d),
	.w3(32'hbc06dbf6),
	.w4(32'h3a7ceb16),
	.w5(32'hba948bed),
	.w6(32'h3c15fc2e),
	.w7(32'h3b2560d4),
	.w8(32'h3c6d414b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b940f2f),
	.w1(32'h3c8977dd),
	.w2(32'h3c53d254),
	.w3(32'hbcb9edbe),
	.w4(32'hbc37d792),
	.w5(32'hbc85b87b),
	.w6(32'h3b44c77c),
	.w7(32'h3d0358ec),
	.w8(32'hbc015899),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce40d3c),
	.w1(32'hbb687e52),
	.w2(32'hbcedaec6),
	.w3(32'hbcdd0961),
	.w4(32'hbc151527),
	.w5(32'hbc597f68),
	.w6(32'hbc8ca183),
	.w7(32'hbc61b5ff),
	.w8(32'hbcbd3b78),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac12eb9),
	.w1(32'h3bc40197),
	.w2(32'hbaa5bfb5),
	.w3(32'hbc1c7824),
	.w4(32'hbb2da296),
	.w5(32'hbc4fc167),
	.w6(32'h3b1abf3c),
	.w7(32'h3b27efce),
	.w8(32'h3ceb0443),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb5403),
	.w1(32'hbb9ae0cf),
	.w2(32'hbc3ba3cb),
	.w3(32'hbc4a14a3),
	.w4(32'hbcfcb1f5),
	.w5(32'hbc247970),
	.w6(32'h3d9161fa),
	.w7(32'h3cccaccc),
	.w8(32'h3c3b762e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d57f3),
	.w1(32'h3ad3c9ae),
	.w2(32'h3b86ed84),
	.w3(32'hbc089e04),
	.w4(32'hbcd8d706),
	.w5(32'hbbf7859a),
	.w6(32'h3cdd7498),
	.w7(32'h3c51e51c),
	.w8(32'h3ca7d7bd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb808dc5),
	.w1(32'hbc676f65),
	.w2(32'hbc00dbee),
	.w3(32'hbc877dad),
	.w4(32'hbca4bdfe),
	.w5(32'hbcb6dfba),
	.w6(32'h3bdaf115),
	.w7(32'h3caf0591),
	.w8(32'h3c0dbe46),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad76b35),
	.w1(32'hbb5a9c8a),
	.w2(32'hbb233006),
	.w3(32'hbc304f20),
	.w4(32'hbca15b61),
	.w5(32'hbc62f1ba),
	.w6(32'h3c653266),
	.w7(32'h3b60bfc0),
	.w8(32'h3cb2b465),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085ab2),
	.w1(32'h3986fea0),
	.w2(32'hbb8b8ce0),
	.w3(32'hbc91cc25),
	.w4(32'hbd52ac10),
	.w5(32'hbc70dcef),
	.w6(32'h3da15e04),
	.w7(32'h3ce0ff7e),
	.w8(32'h3c5ddf89),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2e240),
	.w1(32'hbab381d6),
	.w2(32'hbc297384),
	.w3(32'hbcfc6a5f),
	.w4(32'hbb8802e8),
	.w5(32'hbc9ee604),
	.w6(32'hbc80ec76),
	.w7(32'h3c33c05b),
	.w8(32'hbc82b79c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc039962),
	.w1(32'h3b93615e),
	.w2(32'hbbadcaf5),
	.w3(32'h3bc300c1),
	.w4(32'h3ce4a2c2),
	.w5(32'h3c04883d),
	.w6(32'hbcdb4a56),
	.w7(32'hbbe0f1f4),
	.w8(32'hbb9fdd92),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc2269),
	.w1(32'hbc0e6ba9),
	.w2(32'h3acb789c),
	.w3(32'hbc936f20),
	.w4(32'hbc36c043),
	.w5(32'hbc0e81b9),
	.w6(32'hbcb93bed),
	.w7(32'hbc426187),
	.w8(32'h3c063419),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc896d3),
	.w1(32'hbd111365),
	.w2(32'h3cb76ab6),
	.w3(32'h3bc31ce4),
	.w4(32'hbd3aea7f),
	.w5(32'h3ba8727c),
	.w6(32'hbc953711),
	.w7(32'h3c4524f9),
	.w8(32'hbb85ba35),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17950a),
	.w1(32'hbbab15eb),
	.w2(32'hba0c090c),
	.w3(32'hbc381910),
	.w4(32'h3c278e3d),
	.w5(32'hbba093ee),
	.w6(32'hbb9492a7),
	.w7(32'h3c0507f4),
	.w8(32'hbb32a0d5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a420e),
	.w1(32'h3a08bacc),
	.w2(32'hbb4309fc),
	.w3(32'h3b6a45e1),
	.w4(32'h3c328728),
	.w5(32'hbb176a0c),
	.w6(32'h39f7026f),
	.w7(32'h3bc0af8f),
	.w8(32'h3bafd8be),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6312e8),
	.w1(32'hbbda3aff),
	.w2(32'h3c3c46d3),
	.w3(32'hbb41b05b),
	.w4(32'hbc17db07),
	.w5(32'hb92e70d4),
	.w6(32'hbb0bf241),
	.w7(32'h3b97d472),
	.w8(32'h3b800559),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4ebfd3),
	.w1(32'hbc06a416),
	.w2(32'h3bae8db6),
	.w3(32'hbd0c1551),
	.w4(32'hbb8d4b9f),
	.w5(32'hbc87d61e),
	.w6(32'hbd340d34),
	.w7(32'h3bfb3849),
	.w8(32'hbbe04fe7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcffd57d),
	.w1(32'hbbd7b812),
	.w2(32'hbb871b4c),
	.w3(32'hbd09af36),
	.w4(32'h3c56a80c),
	.w5(32'h3c4a9772),
	.w6(32'hbceeb64c),
	.w7(32'h3ab46a87),
	.w8(32'hbc8670bc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29d15e),
	.w1(32'h3cbc215d),
	.w2(32'hbbc2fb15),
	.w3(32'hbc1e4ae8),
	.w4(32'h3bd32b58),
	.w5(32'h3b602b64),
	.w6(32'hbc44564b),
	.w7(32'h3ad0ede4),
	.w8(32'h3a93ef98),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5761b2),
	.w1(32'hbc7ef154),
	.w2(32'h3a9d91d6),
	.w3(32'h3b35f603),
	.w4(32'hbb75cf6c),
	.w5(32'h39a4503f),
	.w6(32'h3833abe4),
	.w7(32'h3babef6b),
	.w8(32'hb9cfe202),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3ee74),
	.w1(32'hbc2a050c),
	.w2(32'h3a8df747),
	.w3(32'hbae6b5cb),
	.w4(32'hbbc126d6),
	.w5(32'hbb9d0698),
	.w6(32'hba3f89fc),
	.w7(32'hbaa06b75),
	.w8(32'hbad96b4f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cdb26),
	.w1(32'hbc9e97ba),
	.w2(32'h3a0ffb49),
	.w3(32'hbbeedc3f),
	.w4(32'hbbb0a593),
	.w5(32'hbc1cd7fa),
	.w6(32'h3aa9136f),
	.w7(32'h3b5b1c72),
	.w8(32'h3bcfd67a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc58d41),
	.w1(32'hbd09d89b),
	.w2(32'h3c05ba17),
	.w3(32'h3b6c7273),
	.w4(32'hbcbd1e84),
	.w5(32'hbcb0040d),
	.w6(32'hbcd4596d),
	.w7(32'h3c01c8d7),
	.w8(32'hbba83ff6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7881cd),
	.w1(32'h3c66cf76),
	.w2(32'hba592b89),
	.w3(32'hbca3af23),
	.w4(32'hbbc79559),
	.w5(32'hbc1aecc2),
	.w6(32'hbc4fcfce),
	.w7(32'h3bc41b4b),
	.w8(32'hbcbfb87d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1f8643),
	.w1(32'h3c5622b1),
	.w2(32'h3b1d7a32),
	.w3(32'hbcae184d),
	.w4(32'h3c8b6cf9),
	.w5(32'hbb068426),
	.w6(32'h3ca5bec0),
	.w7(32'hbb9be464),
	.w8(32'hbbe8c969),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb8f89),
	.w1(32'hbb11cbe4),
	.w2(32'hbbf77846),
	.w3(32'h3a0145fe),
	.w4(32'h3b961691),
	.w5(32'h3b69a7eb),
	.w6(32'h3a10d2c8),
	.w7(32'hb926075e),
	.w8(32'hbb59a4b5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ffab2),
	.w1(32'hbbfccfc1),
	.w2(32'hbcee5414),
	.w3(32'hbbd93262),
	.w4(32'hbccf9173),
	.w5(32'hbca87eb7),
	.w6(32'h3bcfb1a6),
	.w7(32'h382afafe),
	.w8(32'h3b641960),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1ceedd),
	.w1(32'hbc8c6dba),
	.w2(32'h3c378843),
	.w3(32'hbc75bade),
	.w4(32'hbd07503d),
	.w5(32'hbc320e74),
	.w6(32'h3b996e5d),
	.w7(32'hbc25476b),
	.w8(32'hbb045383),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af518de),
	.w1(32'hbb5d849d),
	.w2(32'h3a83a265),
	.w3(32'h3a2cc22b),
	.w4(32'h3a0f4e9a),
	.w5(32'hbb7e6227),
	.w6(32'h3b1dfac6),
	.w7(32'h3bb6c93f),
	.w8(32'h3b6d5a87),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04c46c),
	.w1(32'hba16f730),
	.w2(32'hba9fce2e),
	.w3(32'hbc57161f),
	.w4(32'h3aaa2932),
	.w5(32'hbc4a7a3b),
	.w6(32'hbc01efe9),
	.w7(32'hbbba4efe),
	.w8(32'h3c7ddd33),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc105f0b),
	.w1(32'hbc8121c1),
	.w2(32'h3ced77a8),
	.w3(32'hbb903230),
	.w4(32'h38aee3c0),
	.w5(32'h3b9f9788),
	.w6(32'hbc8d1386),
	.w7(32'h3a86e606),
	.w8(32'hbb5fce21),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc3436),
	.w1(32'hbc4f398b),
	.w2(32'h3ca4965a),
	.w3(32'h3b9b7df1),
	.w4(32'hbb78f56c),
	.w5(32'h3c90065d),
	.w6(32'hbbd24b44),
	.w7(32'h3c645a29),
	.w8(32'h3c32184b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23b345),
	.w1(32'hbc7ec706),
	.w2(32'h3bd7cdda),
	.w3(32'hbaf4f2cd),
	.w4(32'hbabea73b),
	.w5(32'h3b28d289),
	.w6(32'hbb403283),
	.w7(32'h3cae4109),
	.w8(32'hbbf60b6a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb090b),
	.w1(32'hbd47e76a),
	.w2(32'h3bf751af),
	.w3(32'h3983d2bf),
	.w4(32'hbc216145),
	.w5(32'hbc994adc),
	.w6(32'h3d06910a),
	.w7(32'h3cacc481),
	.w8(32'h39da87d6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule