module layer_10_featuremap_474(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00b181),
	.w1(32'hbb7d7ef9),
	.w2(32'h3b081a3d),
	.w3(32'hbbbc715f),
	.w4(32'hbaaf114c),
	.w5(32'h3b590f4a),
	.w6(32'h39562c66),
	.w7(32'hbb0ee559),
	.w8(32'hbb84a587),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2bb80),
	.w1(32'h3a665297),
	.w2(32'hbb540edd),
	.w3(32'hbb1fb200),
	.w4(32'hbaa4775b),
	.w5(32'hbb4bb5a4),
	.w6(32'hbbe344f4),
	.w7(32'hbbf16e95),
	.w8(32'hbab9b1e3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc170367),
	.w1(32'h3afb5353),
	.w2(32'h3b2ce926),
	.w3(32'hbb4f0839),
	.w4(32'hbb0c126b),
	.w5(32'h3b4e5ae0),
	.w6(32'h3a0b6c21),
	.w7(32'hbb0f4d3d),
	.w8(32'h3bc11aeb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50d484),
	.w1(32'h3bcc78aa),
	.w2(32'h3b23d7d5),
	.w3(32'h3b8c23d9),
	.w4(32'h39fcaf31),
	.w5(32'h39fc497c),
	.w6(32'h3aa81dbc),
	.w7(32'h3aefa308),
	.w8(32'h3c372804),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff00f0),
	.w1(32'hbba58d9e),
	.w2(32'hbb85a0f3),
	.w3(32'hbb96be12),
	.w4(32'hbbed1ea6),
	.w5(32'hbb9c33bc),
	.w6(32'h3c0255fd),
	.w7(32'hbbb3fa54),
	.w8(32'hbaed5d2d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae6743),
	.w1(32'hbb9ca04f),
	.w2(32'hbbcc54ca),
	.w3(32'hbb866697),
	.w4(32'hbb347e87),
	.w5(32'h3bf67b16),
	.w6(32'hb9e462c0),
	.w7(32'h3bb48fb7),
	.w8(32'hbb501662),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba208f5),
	.w1(32'h3ab22e16),
	.w2(32'h3bcf20ef),
	.w3(32'h3a900d7a),
	.w4(32'hbb65dbec),
	.w5(32'hbbcfc6a6),
	.w6(32'h39606c58),
	.w7(32'hbb0bc542),
	.w8(32'h3aa95766),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e1978),
	.w1(32'hbb978897),
	.w2(32'hbb3b2524),
	.w3(32'hbafe5b50),
	.w4(32'h3bc6700f),
	.w5(32'h3bf99ccf),
	.w6(32'hbb4d89ce),
	.w7(32'h386b7f5e),
	.w8(32'hb71736d1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb235e54),
	.w1(32'h392f066e),
	.w2(32'h3ab6dc66),
	.w3(32'h3c50ada3),
	.w4(32'hb9b3216f),
	.w5(32'hb81063c7),
	.w6(32'hbbebbe97),
	.w7(32'hb42486fa),
	.w8(32'h3b4f9cfe),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad20647),
	.w1(32'hbbbb985f),
	.w2(32'hbc164178),
	.w3(32'hb9dd8dc0),
	.w4(32'hbc3d4fd1),
	.w5(32'h3c063054),
	.w6(32'h3906dc58),
	.w7(32'hbbd694fd),
	.w8(32'h3b1cc020),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0078c1),
	.w1(32'hbb6e29cc),
	.w2(32'hbb8d294c),
	.w3(32'h3aaa1f3d),
	.w4(32'hba18b3cd),
	.w5(32'h3c0c0064),
	.w6(32'hbbb70106),
	.w7(32'h39134d9d),
	.w8(32'hbb8b7885),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90bda8),
	.w1(32'hbb0a23bb),
	.w2(32'hbbd6fd51),
	.w3(32'h3a11ebb9),
	.w4(32'hbb9b7bdc),
	.w5(32'h3a43a0a6),
	.w6(32'h3a7c2824),
	.w7(32'hbb259909),
	.w8(32'hbb138a26),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947d2e),
	.w1(32'hba059788),
	.w2(32'h3a54dadc),
	.w3(32'h3ba2621a),
	.w4(32'hbb86a832),
	.w5(32'h3b3bd820),
	.w6(32'hbbf9be67),
	.w7(32'hb9da6394),
	.w8(32'h3a2f5029),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e41b),
	.w1(32'hbb8a95f7),
	.w2(32'hbad46a75),
	.w3(32'hbb51356e),
	.w4(32'hbb42de6c),
	.w5(32'h3b5317a1),
	.w6(32'h3b09e761),
	.w7(32'h3b244650),
	.w8(32'h3b921bb3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f3246),
	.w1(32'h3b26d476),
	.w2(32'h3bb5a0f7),
	.w3(32'h3b5d8027),
	.w4(32'h3a375298),
	.w5(32'hbb2bd261),
	.w6(32'h3bb02fb3),
	.w7(32'h3adaf446),
	.w8(32'h3b8196b0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d6ce0),
	.w1(32'h39f80a3a),
	.w2(32'h3be806e7),
	.w3(32'h3b8db12d),
	.w4(32'hba1470d1),
	.w5(32'h3b9116cc),
	.w6(32'h3ab5af22),
	.w7(32'h3b46342b),
	.w8(32'hbb89d0b4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17fd50),
	.w1(32'h3b0c8dea),
	.w2(32'h3ba2ef6d),
	.w3(32'h3b0032fc),
	.w4(32'h39e0234e),
	.w5(32'h3a264ddb),
	.w6(32'hb8301a0a),
	.w7(32'hbb842f34),
	.w8(32'h3b0bef2c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e3af),
	.w1(32'hb94246e2),
	.w2(32'h3b227590),
	.w3(32'h39ecba28),
	.w4(32'h39a70ca5),
	.w5(32'h3a203a14),
	.w6(32'h3be730ea),
	.w7(32'hbb291aea),
	.w8(32'hbb709c3a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8328ce),
	.w1(32'h3b40b1e8),
	.w2(32'hb85d6bdb),
	.w3(32'hbb1ac9ba),
	.w4(32'hbac25cd3),
	.w5(32'h3b13b59f),
	.w6(32'hbaf038db),
	.w7(32'h3b5c6f19),
	.w8(32'h3b4aa4c0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66f62c),
	.w1(32'h3c5ba8ed),
	.w2(32'h3c654b44),
	.w3(32'h3c00a280),
	.w4(32'hbb09ab18),
	.w5(32'hbc8ea331),
	.w6(32'hbb8d8274),
	.w7(32'h3ba8381d),
	.w8(32'h3c815ae5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8be646),
	.w1(32'hbbbc6aef),
	.w2(32'hbc3134e1),
	.w3(32'hbbb771d8),
	.w4(32'hbab5a858),
	.w5(32'h3c0cf640),
	.w6(32'hba00e545),
	.w7(32'hb921858d),
	.w8(32'hbb8eb092),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb20e9),
	.w1(32'h3b355e0d),
	.w2(32'hbb1cf1aa),
	.w3(32'h3a1177f5),
	.w4(32'hbbd953d3),
	.w5(32'h3b1a9c1d),
	.w6(32'hbb9b3b00),
	.w7(32'h3c15d2f7),
	.w8(32'h3aa03abd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc36742),
	.w1(32'h3b327225),
	.w2(32'h3bd7211f),
	.w3(32'hbc4d30cd),
	.w4(32'h3b67c72d),
	.w5(32'hbc17633d),
	.w6(32'hbba9f307),
	.w7(32'h3bb79389),
	.w8(32'h3c03f802),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b66b),
	.w1(32'h398fb953),
	.w2(32'h3b5ba867),
	.w3(32'hb9e15af2),
	.w4(32'hbb219245),
	.w5(32'hbbddb5a7),
	.w6(32'h3bb7a4d9),
	.w7(32'hbb9be7d2),
	.w8(32'hbb77dce8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926897),
	.w1(32'h3ac51b2f),
	.w2(32'h3b06b286),
	.w3(32'hbbdf7499),
	.w4(32'h3b95c263),
	.w5(32'h39a3c448),
	.w6(32'hbbae6f25),
	.w7(32'hba9e0336),
	.w8(32'hbbc50443),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21218b),
	.w1(32'hbb9e293e),
	.w2(32'h3a5ca5d1),
	.w3(32'h3bcc4aca),
	.w4(32'h3c0136c0),
	.w5(32'h3be49b85),
	.w6(32'h3b1deb07),
	.w7(32'hbba79a39),
	.w8(32'hbbb50d5f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb740316),
	.w1(32'hbb8d009b),
	.w2(32'hbb6366e4),
	.w3(32'hbb91c8a9),
	.w4(32'hbbc872bb),
	.w5(32'h3c074435),
	.w6(32'hb9ebeadb),
	.w7(32'h3b82966a),
	.w8(32'hba3c823e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e61c9),
	.w1(32'hbb843960),
	.w2(32'hbbc915e2),
	.w3(32'h3a7ca4aa),
	.w4(32'hba819c2e),
	.w5(32'hbbb7acd9),
	.w6(32'hb952c0c2),
	.w7(32'hb9d4f819),
	.w8(32'hbb6696c2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e49b5),
	.w1(32'h3c3b8b2d),
	.w2(32'h3c53f68b),
	.w3(32'h395bb9b4),
	.w4(32'h3bd3b5db),
	.w5(32'hbc23cb6d),
	.w6(32'hbb905d40),
	.w7(32'hba3c4b28),
	.w8(32'hbb4fa77b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c190fd5),
	.w1(32'hbb659697),
	.w2(32'hbb94a740),
	.w3(32'hbb1a58c4),
	.w4(32'hbb33e2a2),
	.w5(32'h3bb270eb),
	.w6(32'h3a6a5b83),
	.w7(32'h3b0f7d09),
	.w8(32'h39f0c6ac),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b503b),
	.w1(32'h3b4a61c0),
	.w2(32'h3c4fcb18),
	.w3(32'h3bd00c30),
	.w4(32'hbbc70266),
	.w5(32'hbc6018ca),
	.w6(32'hbc25cf9e),
	.w7(32'h3a2eec81),
	.w8(32'h3bdcbf65),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57358d),
	.w1(32'h3b6f6cb2),
	.w2(32'hbae70404),
	.w3(32'hbb2defb9),
	.w4(32'h3a7f62c3),
	.w5(32'hba67b778),
	.w6(32'h371d1c6d),
	.w7(32'hbb09eead),
	.w8(32'hba806545),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b809917),
	.w1(32'hbafc84da),
	.w2(32'hbba3cab4),
	.w3(32'h3a64f524),
	.w4(32'hbb557adb),
	.w5(32'hbc0cc744),
	.w6(32'hbb90bacd),
	.w7(32'hbb8075f7),
	.w8(32'hbab72747),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83824f),
	.w1(32'hbb3a23a9),
	.w2(32'hbb169160),
	.w3(32'hbc1a338b),
	.w4(32'h3b8278a8),
	.w5(32'h3a5c94f8),
	.w6(32'hbb521264),
	.w7(32'hb88ddc78),
	.w8(32'hbafd3af1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c92c6),
	.w1(32'h3b6d2440),
	.w2(32'h3c346d3b),
	.w3(32'h3ba807c1),
	.w4(32'h3b4681e8),
	.w5(32'h3b8a7f47),
	.w6(32'hbb3f88cf),
	.w7(32'hba2ebaeb),
	.w8(32'h3a9ba009),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23dfb7),
	.w1(32'h3b95a6f9),
	.w2(32'h3b3e2f7c),
	.w3(32'h3c0797ab),
	.w4(32'h3be6d0ee),
	.w5(32'hbb8f3df7),
	.w6(32'hbbe81a70),
	.w7(32'hbb0decd2),
	.w8(32'h3a3a0652),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9b252),
	.w1(32'hbb31ca4c),
	.w2(32'hbb1984e5),
	.w3(32'hbb22230d),
	.w4(32'h3b8081fd),
	.w5(32'hba15203f),
	.w6(32'h3ba2fc90),
	.w7(32'h3b21919b),
	.w8(32'hbb04a00b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988a074),
	.w1(32'h3a084148),
	.w2(32'hbbdbed8a),
	.w3(32'h3ad6a159),
	.w4(32'hbc0561cd),
	.w5(32'hbc1ed077),
	.w6(32'h3c0b7edd),
	.w7(32'h3ad1e5ba),
	.w8(32'h3be62359),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad051a),
	.w1(32'hbb2a9b50),
	.w2(32'hb99a916e),
	.w3(32'h3a4fecb9),
	.w4(32'hbb8a3441),
	.w5(32'hbb3108ec),
	.w6(32'h3b64aab7),
	.w7(32'hb96f9dee),
	.w8(32'hb99497c7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6756ba),
	.w1(32'hba0f3dbd),
	.w2(32'hbb0c574a),
	.w3(32'h39aae869),
	.w4(32'hbbb9a89a),
	.w5(32'hbb5b7e40),
	.w6(32'h3add124c),
	.w7(32'h39dfa03b),
	.w8(32'hba3edaa5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d2ef2),
	.w1(32'hbab4edbf),
	.w2(32'h3aeecf94),
	.w3(32'hbb6bade9),
	.w4(32'hbc08a774),
	.w5(32'hbc0e2349),
	.w6(32'hbaadc85c),
	.w7(32'h3b5bb1fd),
	.w8(32'h3c5f7527),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1c02f),
	.w1(32'hbb8c11d9),
	.w2(32'hbbbebd3f),
	.w3(32'h3c28c8b5),
	.w4(32'h3a6d77f2),
	.w5(32'h3b07a890),
	.w6(32'h3bd2d537),
	.w7(32'h3b611020),
	.w8(32'h3b2b774c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b406b14),
	.w1(32'hb925483d),
	.w2(32'hbb2a2bf5),
	.w3(32'h3b35049a),
	.w4(32'hba2be5f0),
	.w5(32'hbb7c82ef),
	.w6(32'h3a47d7fd),
	.w7(32'hbb6a69a9),
	.w8(32'h3b3a4625),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e8be0),
	.w1(32'hbb8a4834),
	.w2(32'hbbe7b1ff),
	.w3(32'hbbdc014b),
	.w4(32'hbc12d007),
	.w5(32'h3a3fa99b),
	.w6(32'h3b6976f3),
	.w7(32'hbb0d3549),
	.w8(32'hbb1c485d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a2294),
	.w1(32'hbb3b035a),
	.w2(32'hbbaf8e39),
	.w3(32'hbb56dfbc),
	.w4(32'hbbea9ac3),
	.w5(32'hbba2f8dc),
	.w6(32'hbc09c8b1),
	.w7(32'hba05e531),
	.w8(32'hba9ef9b5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01ac83),
	.w1(32'h3b82972d),
	.w2(32'h3c4d86d5),
	.w3(32'hbaacc5d2),
	.w4(32'h3c0c5ac5),
	.w5(32'h3c66cbf0),
	.w6(32'hbac48cd1),
	.w7(32'h3bc3b468),
	.w8(32'hba605d65),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c0549),
	.w1(32'hbbc93033),
	.w2(32'hbbec5b0f),
	.w3(32'h3ac8884c),
	.w4(32'hbba0b930),
	.w5(32'h3c00b232),
	.w6(32'h3b5b31a9),
	.w7(32'hbc0e7c42),
	.w8(32'hbc053d27),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb466d0b),
	.w1(32'hbb151dde),
	.w2(32'hba5d89f2),
	.w3(32'hbb46bfaa),
	.w4(32'hbb70b294),
	.w5(32'hbb602ad5),
	.w6(32'hba629e85),
	.w7(32'hbb1897fb),
	.w8(32'h394823c1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf768d8),
	.w1(32'h38bc6562),
	.w2(32'hbad78494),
	.w3(32'hbb5a65af),
	.w4(32'h3ac49057),
	.w5(32'hba7ec731),
	.w6(32'h3a7695ba),
	.w7(32'h3b8cafdf),
	.w8(32'h3c0ab162),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb4f03),
	.w1(32'h3c1d3c48),
	.w2(32'hbb5f99bb),
	.w3(32'h3b6a930d),
	.w4(32'h3c17986d),
	.w5(32'hbba0c243),
	.w6(32'h3b18aa54),
	.w7(32'hb9f76f8f),
	.w8(32'hba7e5104),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31a5ce),
	.w1(32'h3be44c07),
	.w2(32'h3a1fc712),
	.w3(32'h392453ca),
	.w4(32'h3bd1bc99),
	.w5(32'hbc0e444c),
	.w6(32'h3b3a2b82),
	.w7(32'h3aaecf14),
	.w8(32'hbc009b91),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2ff32),
	.w1(32'hba0d8ecd),
	.w2(32'hbae4e445),
	.w3(32'hb9b1b10f),
	.w4(32'hbb69d09a),
	.w5(32'hbb2ffc73),
	.w6(32'h3c04e346),
	.w7(32'hbc0d3334),
	.w8(32'hbb209f2d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0165b5),
	.w1(32'h3b385aaf),
	.w2(32'h3b55a208),
	.w3(32'hbbadf751),
	.w4(32'h3a7ed19c),
	.w5(32'hbab23e0e),
	.w6(32'h3b1bb976),
	.w7(32'h3b8944b9),
	.w8(32'hb8a426c9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b172312),
	.w1(32'hbb94cf65),
	.w2(32'hba42cfe0),
	.w3(32'h3bd0941b),
	.w4(32'h3c26ecd8),
	.w5(32'h3bddf47d),
	.w6(32'hbacb683b),
	.w7(32'hbb9b2702),
	.w8(32'hbc111a02),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4cd98),
	.w1(32'h3b5aa4b6),
	.w2(32'h3a8e7064),
	.w3(32'h3bc55f03),
	.w4(32'hbc3a5136),
	.w5(32'hbc1f77e9),
	.w6(32'hbc035aa8),
	.w7(32'hbb422057),
	.w8(32'h38f117f5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e6187),
	.w1(32'hbb3c6cc1),
	.w2(32'h3a12d2cb),
	.w3(32'hbb4ecb57),
	.w4(32'hbbb62cd5),
	.w5(32'hbc0f6b34),
	.w6(32'hbabd06bf),
	.w7(32'hb9ec57b0),
	.w8(32'h3b945bb1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05de2d),
	.w1(32'hbb9ee719),
	.w2(32'hbb2a1a4b),
	.w3(32'hbb60844b),
	.w4(32'h3bbc33f7),
	.w5(32'h3c25c935),
	.w6(32'hba910c0c),
	.w7(32'hbb9298ac),
	.w8(32'hbbe26c85),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dd059),
	.w1(32'hbb27f550),
	.w2(32'hbbef7d2e),
	.w3(32'h3b21c97f),
	.w4(32'hbbac35a5),
	.w5(32'hbc14f962),
	.w6(32'h3b387cd4),
	.w7(32'h3bab2835),
	.w8(32'h3ad59391),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d896da),
	.w1(32'hbbea972f),
	.w2(32'hbb91cc9e),
	.w3(32'hbbe3c6e0),
	.w4(32'hbbf96e73),
	.w5(32'hbb83bd22),
	.w6(32'hbbb41330),
	.w7(32'hbaf7692c),
	.w8(32'h3b57407e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc229a11),
	.w1(32'hbaf6c4d5),
	.w2(32'hbb1ea719),
	.w3(32'hbbaa33e2),
	.w4(32'h3bc8d0b6),
	.w5(32'h3c1c2cbc),
	.w6(32'h3bd684d5),
	.w7(32'hbb30161d),
	.w8(32'hbad2c002),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1e8ec),
	.w1(32'hbc5d786e),
	.w2(32'hbc76830f),
	.w3(32'h3c74c098),
	.w4(32'hbc5f278f),
	.w5(32'h3b542aa7),
	.w6(32'hb9fa950b),
	.w7(32'h3ae78fed),
	.w8(32'h3bce191d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c7e18),
	.w1(32'hbb09c38e),
	.w2(32'h3b3fa086),
	.w3(32'hbc0be75e),
	.w4(32'hbaa87cf7),
	.w5(32'hbc1f6070),
	.w6(32'h3c0904b2),
	.w7(32'h3bcdeab4),
	.w8(32'h3bf1d0f8),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb10c2),
	.w1(32'h3a939b6e),
	.w2(32'h3b690184),
	.w3(32'hba82d9c2),
	.w4(32'hbb1d398f),
	.w5(32'hbc127d24),
	.w6(32'hbb336456),
	.w7(32'hbb62caf7),
	.w8(32'h3a5a99c6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf002),
	.w1(32'h3a837d8c),
	.w2(32'hbb343351),
	.w3(32'h3aa72c03),
	.w4(32'hba9a8e5e),
	.w5(32'hbc27fa13),
	.w6(32'h3c17089e),
	.w7(32'hbbb26394),
	.w8(32'hbb59311b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f16d8),
	.w1(32'h3b3d6dde),
	.w2(32'h3b1c523a),
	.w3(32'hbb49001c),
	.w4(32'h3c075670),
	.w5(32'h3bfd89c6),
	.w6(32'hbbb88664),
	.w7(32'h3b38126a),
	.w8(32'h3b4f729f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf23d50),
	.w1(32'hbbca8860),
	.w2(32'h3b4a4316),
	.w3(32'h3bbfd9c6),
	.w4(32'h3b0fb9e1),
	.w5(32'h3b58be58),
	.w6(32'hba6d29e3),
	.w7(32'h3b4a5071),
	.w8(32'hbb3a7c56),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f6ee9),
	.w1(32'h3b5630b9),
	.w2(32'h388abeb8),
	.w3(32'hbafd6e94),
	.w4(32'h3b50db1d),
	.w5(32'h3bcc1c99),
	.w6(32'h3bafda98),
	.w7(32'hbaa0659c),
	.w8(32'hbb8384f4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4643a),
	.w1(32'hbac46f92),
	.w2(32'h3aeaaed1),
	.w3(32'hba0e95e0),
	.w4(32'h3bff3847),
	.w5(32'hbbb506fe),
	.w6(32'h38b20609),
	.w7(32'h3bd13082),
	.w8(32'h3b36a612),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e3747),
	.w1(32'h3c5651e8),
	.w2(32'h3b06a3c0),
	.w3(32'h3b7c675d),
	.w4(32'hbb7eb9a7),
	.w5(32'hba8ac0b2),
	.w6(32'h3ac20a50),
	.w7(32'hbb643a00),
	.w8(32'hba9ec2fd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb437d29),
	.w1(32'hba9a4273),
	.w2(32'hbc1a27ca),
	.w3(32'h39cc3932),
	.w4(32'hbb8296f3),
	.w5(32'hbc30f5a7),
	.w6(32'h3bd6553c),
	.w7(32'hbb27caf3),
	.w8(32'hbc0ff0cf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad15cb),
	.w1(32'h3ae6a4ad),
	.w2(32'h3baa9e69),
	.w3(32'hbc118268),
	.w4(32'h3b2c36f4),
	.w5(32'h3be2f80b),
	.w6(32'hbbe7eebc),
	.w7(32'h3b53cdfd),
	.w8(32'hbaf23c8f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0d3de),
	.w1(32'h3a6e426d),
	.w2(32'hbbe19c87),
	.w3(32'hba372aba),
	.w4(32'hbbc65879),
	.w5(32'hbad04f2e),
	.w6(32'hbb41f897),
	.w7(32'h3b13d8e2),
	.w8(32'hbb231a58),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b6b39),
	.w1(32'hbb7b16f6),
	.w2(32'hbb9e507f),
	.w3(32'hba12b16d),
	.w4(32'hbbd1b531),
	.w5(32'hbb8e570f),
	.w6(32'hbb2b31fe),
	.w7(32'hbb529420),
	.w8(32'hbb62a79f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba20fe3),
	.w1(32'h3951f173),
	.w2(32'hba844cfb),
	.w3(32'hbba58971),
	.w4(32'h3ba907a4),
	.w5(32'hbc51b03a),
	.w6(32'hbbff80e6),
	.w7(32'h39d1e978),
	.w8(32'h3a0db5b5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905474a),
	.w1(32'hbae9bd0f),
	.w2(32'h3bc64b1a),
	.w3(32'hbb298407),
	.w4(32'hbc12cc4e),
	.w5(32'hbb109f57),
	.w6(32'hbaee7b34),
	.w7(32'h3aac7d21),
	.w8(32'h3bb3d785),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2017c),
	.w1(32'h3b906fd0),
	.w2(32'h3ade88d9),
	.w3(32'h3a9a2a05),
	.w4(32'h3af94aa7),
	.w5(32'hba4a103c),
	.w6(32'h3ba2d9c3),
	.w7(32'hbb28f5ee),
	.w8(32'hb6451959),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ae61b),
	.w1(32'h3993ae47),
	.w2(32'hb922b764),
	.w3(32'hbbb93416),
	.w4(32'hbae9086d),
	.w5(32'h3c0066cf),
	.w6(32'hbb786542),
	.w7(32'hbabddb7a),
	.w8(32'h3b285019),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d70af),
	.w1(32'hbc557215),
	.w2(32'hbc649195),
	.w3(32'h3c495607),
	.w4(32'hb93ee3a8),
	.w5(32'h3b6d48b5),
	.w6(32'h3b9cc5d1),
	.w7(32'hbb972149),
	.w8(32'h39960a7a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc088da4),
	.w1(32'h3bf086cd),
	.w2(32'h3b5f0522),
	.w3(32'hbbc161ca),
	.w4(32'h3c289457),
	.w5(32'h3ccd1208),
	.w6(32'hbc01493c),
	.w7(32'h3a61ae6c),
	.w8(32'h3bb01110),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dec26),
	.w1(32'h3ac947dd),
	.w2(32'hbbb111bd),
	.w3(32'h3bd55f54),
	.w4(32'h3b1b461e),
	.w5(32'h3a68e83c),
	.w6(32'h3b9a124b),
	.w7(32'h3b95ba7a),
	.w8(32'hba908bf5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0db5d1),
	.w1(32'h3b8ac4c0),
	.w2(32'h3baf186d),
	.w3(32'h3bb90c65),
	.w4(32'h3bb241f3),
	.w5(32'h3c361a51),
	.w6(32'h3b1c7296),
	.w7(32'h3ac3e1ce),
	.w8(32'h3c24270c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40dc16),
	.w1(32'hbb88bd4b),
	.w2(32'hbab41e1b),
	.w3(32'h3bb98a48),
	.w4(32'hbb6b90a8),
	.w5(32'hba745645),
	.w6(32'h3bb94203),
	.w7(32'hbb73215c),
	.w8(32'h3a380192),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9a4a0),
	.w1(32'h3bc140d4),
	.w2(32'h3a825981),
	.w3(32'hbb871e76),
	.w4(32'h3c04f575),
	.w5(32'h3bb3c6ee),
	.w6(32'hba94b542),
	.w7(32'h3bfbfd0d),
	.w8(32'hbbe4edae),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10c1ce),
	.w1(32'h3b36bf78),
	.w2(32'hbb11fcd5),
	.w3(32'hbb2ff149),
	.w4(32'hbc1bc434),
	.w5(32'hbb8303fd),
	.w6(32'hbc448dcb),
	.w7(32'hbaf99774),
	.w8(32'h38ca4b70),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f2527),
	.w1(32'h3be8a45f),
	.w2(32'h3b9c254a),
	.w3(32'hbb78c334),
	.w4(32'h3b8e7ae3),
	.w5(32'hba35ab5e),
	.w6(32'h39f1687f),
	.w7(32'h3bc0514d),
	.w8(32'h3c05b9e5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb167e),
	.w1(32'h3ac14a12),
	.w2(32'hbba9158c),
	.w3(32'h3b392eca),
	.w4(32'hbb253b24),
	.w5(32'hbb20e677),
	.w6(32'h3ab012b6),
	.w7(32'h3b3e4d08),
	.w8(32'h3a8ac040),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6553f),
	.w1(32'h399e04ae),
	.w2(32'hbbe181e9),
	.w3(32'h3b3ced9d),
	.w4(32'h3c1a55a3),
	.w5(32'h3a9e6d7c),
	.w6(32'h393810d1),
	.w7(32'h3b9e432f),
	.w8(32'hbb74c419),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a85e6),
	.w1(32'hbb8ed15f),
	.w2(32'hbba50978),
	.w3(32'h3bef6620),
	.w4(32'hbb48c0de),
	.w5(32'hbb8a1b11),
	.w6(32'h3aed5676),
	.w7(32'hbb02a2f8),
	.w8(32'h39f4ca2c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94396c),
	.w1(32'h3ac5046b),
	.w2(32'h3b31a570),
	.w3(32'h3ba8f375),
	.w4(32'hbbb143fc),
	.w5(32'h3b59b14d),
	.w6(32'h3b40b4a2),
	.w7(32'h39a2c2fe),
	.w8(32'h3ad5c750),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a709c),
	.w1(32'hba566518),
	.w2(32'h3b7a2af8),
	.w3(32'h3c12abcf),
	.w4(32'hbb230016),
	.w5(32'h3c1c30c8),
	.w6(32'h3a30aae8),
	.w7(32'hbb9eeb47),
	.w8(32'h3b78ce75),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1c0c3),
	.w1(32'hbb8e45c0),
	.w2(32'h39e24bab),
	.w3(32'h3c014c86),
	.w4(32'hbbf2827e),
	.w5(32'h3aa7b909),
	.w6(32'h3bba45b7),
	.w7(32'hbb3c480c),
	.w8(32'h3b22c871),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7adb79),
	.w1(32'hbb710c6d),
	.w2(32'hbb8582b3),
	.w3(32'hb8dfb259),
	.w4(32'hbab00df5),
	.w5(32'hb9f000e0),
	.w6(32'hbad8127a),
	.w7(32'h3b3d75d3),
	.w8(32'h3a73e140),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9974cfc),
	.w1(32'h396130dd),
	.w2(32'hba4fecea),
	.w3(32'h3a0cdc80),
	.w4(32'h3b1afb25),
	.w5(32'h3b0ce471),
	.w6(32'hb982ae5c),
	.w7(32'h3b1116c5),
	.w8(32'hbaee9815),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfd44a),
	.w1(32'h3bbdb1b0),
	.w2(32'hbae162ba),
	.w3(32'h3c1114a8),
	.w4(32'h3bf38c9e),
	.w5(32'h3b85e09a),
	.w6(32'hbad86102),
	.w7(32'hbafc3cec),
	.w8(32'hba7c5881),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb171319),
	.w1(32'hbad955bc),
	.w2(32'h3a0706bf),
	.w3(32'h3b837b95),
	.w4(32'hbb6eb8db),
	.w5(32'hbb5fad61),
	.w6(32'hba469b31),
	.w7(32'h3bea7a89),
	.w8(32'hba4cd806),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7fdc1),
	.w1(32'hbcd60a26),
	.w2(32'hbc01be7d),
	.w3(32'h399a6af7),
	.w4(32'hbcbe4018),
	.w5(32'hbcadbb62),
	.w6(32'hbbb8b60d),
	.w7(32'hbc8f2a71),
	.w8(32'hbc72100c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb92e88),
	.w1(32'hb82babbf),
	.w2(32'h3b2963b1),
	.w3(32'hbca95df2),
	.w4(32'h3bfcf2fa),
	.w5(32'hbba4db80),
	.w6(32'hbcc7cabd),
	.w7(32'h3b9113da),
	.w8(32'h3bcc81b3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10ffff),
	.w1(32'hbbbbbc02),
	.w2(32'hbb949e91),
	.w3(32'h3b868c0e),
	.w4(32'hbc324eb9),
	.w5(32'hbb3d1e8e),
	.w6(32'hbae0c93b),
	.w7(32'hbb7c6949),
	.w8(32'hbb8ca188),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3846f953),
	.w1(32'hbc25402f),
	.w2(32'hbbc1aab7),
	.w3(32'h3b376166),
	.w4(32'hbc69fae9),
	.w5(32'hbc01a3f7),
	.w6(32'h3b7b3809),
	.w7(32'hbbb8557e),
	.w8(32'h3ab54f03),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb91037),
	.w1(32'h3b992205),
	.w2(32'h3bbde5af),
	.w3(32'hbbff90e5),
	.w4(32'hbbcb18d2),
	.w5(32'hbb8e0bb6),
	.w6(32'hbb8de20b),
	.w7(32'h3b2c5e35),
	.w8(32'h3c2b641d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b5b3c),
	.w1(32'h3b373cfe),
	.w2(32'h3984d648),
	.w3(32'hbb9a7103),
	.w4(32'h3b5323ce),
	.w5(32'h3aa91ca6),
	.w6(32'h3b81e3e7),
	.w7(32'h391d856f),
	.w8(32'h3ad8f928),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002c49),
	.w1(32'hbbbcd82c),
	.w2(32'h398d719c),
	.w3(32'h3b850a9e),
	.w4(32'hbbb8107d),
	.w5(32'hbacbcb7a),
	.w6(32'hbab72e59),
	.w7(32'hbbf89faf),
	.w8(32'hbb71c7ce),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2fa6),
	.w1(32'hbbfdcc03),
	.w2(32'hbbeb9b46),
	.w3(32'h3b6a21ff),
	.w4(32'hbc116549),
	.w5(32'hbc2589be),
	.w6(32'hbbfcf92e),
	.w7(32'hbba08399),
	.w8(32'hbbcc82e0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13fd6a),
	.w1(32'h3b00c7ea),
	.w2(32'h3b592a88),
	.w3(32'hbbbc2380),
	.w4(32'h3a39ef2c),
	.w5(32'h3c931cd2),
	.w6(32'hbb3b9b1a),
	.w7(32'hb9bc2763),
	.w8(32'h3c1b9507),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c0ee1),
	.w1(32'h39811f04),
	.w2(32'h3b2fdee7),
	.w3(32'h3c047c3e),
	.w4(32'hbb3276cb),
	.w5(32'h39b482f5),
	.w6(32'h3b9b4d05),
	.w7(32'hbb92059c),
	.w8(32'hbc2d5b9d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41977c),
	.w1(32'h3949acfb),
	.w2(32'hbb86ce38),
	.w3(32'hbc1092ef),
	.w4(32'hba7e958f),
	.w5(32'h3a7bebb2),
	.w6(32'hbc6e90f7),
	.w7(32'h3b1bb3bd),
	.w8(32'h3b0cc105),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf9ae4),
	.w1(32'h3bfad558),
	.w2(32'hbb0ff546),
	.w3(32'h3b9cd9bd),
	.w4(32'h3c7e7398),
	.w5(32'h3c299f40),
	.w6(32'h3a47d8c2),
	.w7(32'h3b98980b),
	.w8(32'h39883ae0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28d0f8),
	.w1(32'hbae90d9c),
	.w2(32'h3acbf6c0),
	.w3(32'hbc6fd6a6),
	.w4(32'hbb1b2b3f),
	.w5(32'hbc0d54d8),
	.w6(32'hbbf82290),
	.w7(32'h3bbe4c0b),
	.w8(32'hba9fa0f4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbba03c),
	.w1(32'hba37714f),
	.w2(32'hbb038ee2),
	.w3(32'hbc08fc86),
	.w4(32'hbaa226d0),
	.w5(32'hbbcce1f1),
	.w6(32'hbb719e34),
	.w7(32'h3bf581eb),
	.w8(32'hba890e56),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90bffa),
	.w1(32'hbc2979d1),
	.w2(32'hbbade1eb),
	.w3(32'hb9f49829),
	.w4(32'hbc788aca),
	.w5(32'hbbfd5a5f),
	.w6(32'hbc061b31),
	.w7(32'hbc8c2580),
	.w8(32'hbb97f9a7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e8238),
	.w1(32'hbc099c97),
	.w2(32'hbbe2bfb0),
	.w3(32'hbb6a56bd),
	.w4(32'hbbe7b492),
	.w5(32'hbbe09af6),
	.w6(32'hbc1aa9c6),
	.w7(32'hbb94d371),
	.w8(32'h39ec2b73),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38721613),
	.w1(32'hbc224262),
	.w2(32'hbbfeecef),
	.w3(32'hba3fb79c),
	.w4(32'hbc105361),
	.w5(32'hbbc820b5),
	.w6(32'h3b76bbc7),
	.w7(32'hbb9eb91b),
	.w8(32'h38e3f679),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa869de),
	.w1(32'h3730ad15),
	.w2(32'h384e8c7a),
	.w3(32'h3b71150e),
	.w4(32'hbab477d7),
	.w5(32'hbc9e169f),
	.w6(32'h3a30752e),
	.w7(32'hbb7a10b9),
	.w8(32'hb9f4f902),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d3372),
	.w1(32'h39533625),
	.w2(32'hb99d5712),
	.w3(32'h3bbaf6ec),
	.w4(32'h3b572938),
	.w5(32'h3c1acf81),
	.w6(32'h3ae93105),
	.w7(32'h3ba1c2b5),
	.w8(32'h3a90e299),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b402890),
	.w1(32'h3b9b4736),
	.w2(32'hbb0ba076),
	.w3(32'h3b63b9c3),
	.w4(32'h3ba022a3),
	.w5(32'h3c12aa07),
	.w6(32'h39e2964c),
	.w7(32'h3be2fa26),
	.w8(32'h3a768494),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888e0bd),
	.w1(32'h3b2702aa),
	.w2(32'hbb94cda0),
	.w3(32'h3bc374f5),
	.w4(32'hba1a04e1),
	.w5(32'h3a476ab9),
	.w6(32'h3b9c57ed),
	.w7(32'h38a6c3d6),
	.w8(32'hba708a50),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa06b99),
	.w1(32'h3b4d093f),
	.w2(32'h3b387a12),
	.w3(32'h3b52f0ba),
	.w4(32'h3b7b2d3e),
	.w5(32'hbb21787b),
	.w6(32'hbb7e0454),
	.w7(32'hbb00b94c),
	.w8(32'h3b13579a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39a748),
	.w1(32'h3bd04585),
	.w2(32'hbae33ce1),
	.w3(32'hbb9a170e),
	.w4(32'h3bf13c74),
	.w5(32'h3b8e360a),
	.w6(32'hbb95f578),
	.w7(32'h3a59ed71),
	.w8(32'hbb348272),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d7f18),
	.w1(32'hbc1e2f0d),
	.w2(32'h3b0c431c),
	.w3(32'h3b2d50ee),
	.w4(32'h3a8e6708),
	.w5(32'hbbbe8e87),
	.w6(32'hb9f85826),
	.w7(32'h3b8a7d71),
	.w8(32'h3ab91394),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb125a32),
	.w1(32'hbaf2073a),
	.w2(32'hba9aca39),
	.w3(32'hbc182053),
	.w4(32'hbb952dc2),
	.w5(32'hba2cd00a),
	.w6(32'hbbfd6d12),
	.w7(32'hbb62ad08),
	.w8(32'hbac164a7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919d4b),
	.w1(32'h3b5d714c),
	.w2(32'hb8f59b2a),
	.w3(32'hbbcf122c),
	.w4(32'h3b9e5a29),
	.w5(32'h3bf028d3),
	.w6(32'hbb3ce426),
	.w7(32'h39c6000c),
	.w8(32'h3922b766),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831e33),
	.w1(32'h3c0b3d73),
	.w2(32'h3b959fea),
	.w3(32'h3bfbb804),
	.w4(32'hbb07d167),
	.w5(32'hbbc47d42),
	.w6(32'hb9aca5fc),
	.w7(32'hba30dbdb),
	.w8(32'hbaf6260c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57fde6),
	.w1(32'hbb00ad4b),
	.w2(32'hb921fa05),
	.w3(32'h3ad61fc2),
	.w4(32'h36c6b2b4),
	.w5(32'hbb0b2315),
	.w6(32'h3b993ae8),
	.w7(32'h3afc149d),
	.w8(32'h3a68b83d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98d44d),
	.w1(32'hbc090145),
	.w2(32'hbbaab863),
	.w3(32'h3b6ff4ce),
	.w4(32'hbc40ced4),
	.w5(32'hbd0ebcfb),
	.w6(32'hbb4f7bb6),
	.w7(32'hbb87eca3),
	.w8(32'hbc138486),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07b90d),
	.w1(32'h3b992ec2),
	.w2(32'h3a91cc27),
	.w3(32'h3c4545fb),
	.w4(32'hbb6e605d),
	.w5(32'h39f508d2),
	.w6(32'h3bc119c3),
	.w7(32'hbbc4ed03),
	.w8(32'hba7081ab),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e47fe9),
	.w1(32'hbbe15c2d),
	.w2(32'hbc2953d8),
	.w3(32'h3b97e548),
	.w4(32'hbc085ecc),
	.w5(32'h3ad8d4a8),
	.w6(32'h3a64f3a1),
	.w7(32'hbc4a10f0),
	.w8(32'hbc6f6bea),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2da56),
	.w1(32'h3a3661b5),
	.w2(32'h3b8bf384),
	.w3(32'h3a947de0),
	.w4(32'hbb9c659c),
	.w5(32'h3a444e65),
	.w6(32'hbbbf009d),
	.w7(32'hbb3ffcf5),
	.w8(32'h3ad998e2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bc256),
	.w1(32'hbbdac239),
	.w2(32'hbb9215c0),
	.w3(32'hb992bb04),
	.w4(32'hbc13327b),
	.w5(32'hbb838ec0),
	.w6(32'h395a9066),
	.w7(32'h3aa222f7),
	.w8(32'h3b41d3d6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec2815),
	.w1(32'hbc0a5433),
	.w2(32'hbb236fdf),
	.w3(32'hbbc92a5a),
	.w4(32'hbc1d409d),
	.w5(32'hbc1d109a),
	.w6(32'h3b08bf0c),
	.w7(32'hbb3aa25f),
	.w8(32'h3b6abfcc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b525f98),
	.w1(32'hbc43320a),
	.w2(32'hbbdf6507),
	.w3(32'h3aa9404f),
	.w4(32'hbb6687a2),
	.w5(32'h3951cded),
	.w6(32'h3b55fe71),
	.w7(32'hbbfb8e15),
	.w8(32'hbbd8c982),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6082b),
	.w1(32'hbb9d729f),
	.w2(32'hbc1739b9),
	.w3(32'h3c018ef5),
	.w4(32'hbaf42b57),
	.w5(32'hbc139a91),
	.w6(32'h3a84b10a),
	.w7(32'hbbac39d5),
	.w8(32'hbac5ca97),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb775a5),
	.w1(32'h3c30486c),
	.w2(32'h3b96b4bb),
	.w3(32'hbb89e577),
	.w4(32'h3c0e2115),
	.w5(32'h3c3408ca),
	.w6(32'hbbe7614c),
	.w7(32'h3bd8a3ea),
	.w8(32'hbb5fdb5d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c047d63),
	.w1(32'hbb4e72e4),
	.w2(32'h399d7648),
	.w3(32'h3c74a2ff),
	.w4(32'hbb3d0d01),
	.w5(32'hbbddae09),
	.w6(32'h3b8b0a15),
	.w7(32'h3794e5a2),
	.w8(32'hbb3c1ce4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a398d),
	.w1(32'h3bc90830),
	.w2(32'h3b6757ff),
	.w3(32'h3bd19edf),
	.w4(32'h3c45d1d2),
	.w5(32'h3bbda4b9),
	.w6(32'hbaf6e17f),
	.w7(32'h3c27c569),
	.w8(32'h3c131150),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b566d1e),
	.w1(32'hbbd8862e),
	.w2(32'hbad6228f),
	.w3(32'h3bb01e88),
	.w4(32'hbb51de7f),
	.w5(32'hbc0e1f08),
	.w6(32'h3c18880c),
	.w7(32'h3a3fd2f6),
	.w8(32'h3c213b37),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90d2b4),
	.w1(32'hbafb53cc),
	.w2(32'hbbfed92a),
	.w3(32'hbbbe3d94),
	.w4(32'h3b7cf20a),
	.w5(32'hbb265b5b),
	.w6(32'h3a09ba5d),
	.w7(32'hbbe5d08a),
	.w8(32'h3a306166),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc247244),
	.w1(32'h3b67379c),
	.w2(32'hbb816f30),
	.w3(32'hbadcd3b6),
	.w4(32'hb8c16507),
	.w5(32'hbc1baab8),
	.w6(32'hbb9bd719),
	.w7(32'h3a5aa925),
	.w8(32'hbbd7333c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9fd9f),
	.w1(32'h3c1935b3),
	.w2(32'h3bec6506),
	.w3(32'hbc1c87bf),
	.w4(32'h3b73c3c2),
	.w5(32'h3ac8b290),
	.w6(32'hbc056ff6),
	.w7(32'h3b67ffe8),
	.w8(32'hbb967c40),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab08b04),
	.w1(32'h38e5ee48),
	.w2(32'h3b682908),
	.w3(32'hbbee5d8a),
	.w4(32'h39d8dc34),
	.w5(32'hbb92064d),
	.w6(32'hbbd627c6),
	.w7(32'h3b17866a),
	.w8(32'hba9215e1),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97ff1d),
	.w1(32'hbb88ede7),
	.w2(32'h396f71ee),
	.w3(32'hbc1c8ca0),
	.w4(32'hbb810c05),
	.w5(32'h3be4038a),
	.w6(32'hbbd8b7d7),
	.w7(32'hbb9e83af),
	.w8(32'h3b04d810),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8880),
	.w1(32'hbc0562bf),
	.w2(32'hbc45290f),
	.w3(32'h3c122e22),
	.w4(32'hbb146f1b),
	.w5(32'h3cbb3f0c),
	.w6(32'h3bde6039),
	.w7(32'hbc2de4ad),
	.w8(32'hbc4ec17e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085173),
	.w1(32'hbb018e9a),
	.w2(32'hbbbd55b3),
	.w3(32'h3b8e4ff9),
	.w4(32'hbb334ece),
	.w5(32'hbc4e6da6),
	.w6(32'hbc2e429f),
	.w7(32'h3b04a07b),
	.w8(32'hbbe423e0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b450a),
	.w1(32'h3a2a1897),
	.w2(32'h3c228f84),
	.w3(32'hbb2dce97),
	.w4(32'h3bce4d1d),
	.w5(32'hbb174523),
	.w6(32'hbc0b8d14),
	.w7(32'hb9c6cc84),
	.w8(32'h3bb7bf96),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59b905),
	.w1(32'h3b6c26fd),
	.w2(32'h3ad68104),
	.w3(32'hbb9169b6),
	.w4(32'h3bf8a7e0),
	.w5(32'h3b3e38bc),
	.w6(32'hbb92bd7a),
	.w7(32'h3b6ac2e7),
	.w8(32'h3b9dc2ed),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c2aed),
	.w1(32'h39fe813a),
	.w2(32'h3a88e10f),
	.w3(32'hbb8a058b),
	.w4(32'hba94e3b2),
	.w5(32'hbb29c8ed),
	.w6(32'h3832da83),
	.w7(32'hbb25d714),
	.w8(32'hba773077),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff5474),
	.w1(32'hbc195c1c),
	.w2(32'hbb2a9c6a),
	.w3(32'hbbc35cb8),
	.w4(32'hbc3d41c4),
	.w5(32'hbbd56dcc),
	.w6(32'hbb8822f2),
	.w7(32'hbbe66e1a),
	.w8(32'h3a87d6be),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe1fb2),
	.w1(32'h3b75b012),
	.w2(32'hbb9ab959),
	.w3(32'hbb3cd07d),
	.w4(32'h3b941042),
	.w5(32'hbc41ac0b),
	.w6(32'h3a5143d9),
	.w7(32'h3b6e296e),
	.w8(32'hb702e5ac),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06cbf7),
	.w1(32'h3b62576a),
	.w2(32'hba83e635),
	.w3(32'h3b22df50),
	.w4(32'h3a8769d9),
	.w5(32'hbbb2c17c),
	.w6(32'hbb01ad8c),
	.w7(32'h3b1a6274),
	.w8(32'h3bd52926),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9d9cb),
	.w1(32'h3c6335ef),
	.w2(32'h3c000fa1),
	.w3(32'hbb589a7b),
	.w4(32'h3c996512),
	.w5(32'h3c1c8bb4),
	.w6(32'h39ea698c),
	.w7(32'h3c63de4f),
	.w8(32'h3bb27f30),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa569bd),
	.w1(32'hba4b8c20),
	.w2(32'h3b862072),
	.w3(32'hbb12f398),
	.w4(32'h3b05d3f4),
	.w5(32'h3b251bba),
	.w6(32'hba05a2c1),
	.w7(32'hba333a0c),
	.w8(32'h39ab8369),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1def62),
	.w1(32'h3baf9916),
	.w2(32'hbbc82103),
	.w3(32'hb8bad6de),
	.w4(32'hbad22894),
	.w5(32'hbb8b3b44),
	.w6(32'hb913f91e),
	.w7(32'h38b52cbd),
	.w8(32'h3a9318c3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a252e),
	.w1(32'h3b084b79),
	.w2(32'h39fe9c2d),
	.w3(32'h3be05f2a),
	.w4(32'h3c791a64),
	.w5(32'h3b8fbfd2),
	.w6(32'h3b82debe),
	.w7(32'h3b9ec22a),
	.w8(32'h3b6196f4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b663e66),
	.w1(32'h3a9c0a36),
	.w2(32'hbbaef8c3),
	.w3(32'h3c1c6a69),
	.w4(32'h3a896b10),
	.w5(32'hbc246d7d),
	.w6(32'h3b797e0e),
	.w7(32'h3aa66670),
	.w8(32'hbc0333bc),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383a7903),
	.w1(32'h3becd19d),
	.w2(32'h39d54378),
	.w3(32'hbb8873bf),
	.w4(32'h39b46834),
	.w5(32'hbbe2dafc),
	.w6(32'hbbbacf29),
	.w7(32'h3b169bd5),
	.w8(32'hb91cf730),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07eba9),
	.w1(32'hb9fe3833),
	.w2(32'hbaeebe87),
	.w3(32'h3a08f7ce),
	.w4(32'hbb8015e3),
	.w5(32'hba4284c3),
	.w6(32'hbb02425e),
	.w7(32'hb820959d),
	.w8(32'h3a7f6123),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0950c5),
	.w1(32'hbb2381e0),
	.w2(32'hba7a2f62),
	.w3(32'h3a5c0ec0),
	.w4(32'hbbd7b1b4),
	.w5(32'hbb924018),
	.w6(32'h3bd935a8),
	.w7(32'hbb852873),
	.w8(32'h3a81df70),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb384203),
	.w1(32'hbace4976),
	.w2(32'hbba3b8ff),
	.w3(32'hba96c779),
	.w4(32'hbb976fa9),
	.w5(32'hbb8e3aab),
	.w6(32'hbb9b96d3),
	.w7(32'hbb152c08),
	.w8(32'hbb1bf78a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904b8fe),
	.w1(32'hbb12cfd1),
	.w2(32'h3a103fdb),
	.w3(32'h3a1a54d9),
	.w4(32'h3b7f9006),
	.w5(32'h3c695012),
	.w6(32'h3c1658d2),
	.w7(32'h39ef38f2),
	.w8(32'h3b0772cd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3227ca),
	.w1(32'hbac3f716),
	.w2(32'hb97cc796),
	.w3(32'hbafe1445),
	.w4(32'hbb8b60e3),
	.w5(32'h3ab9d47b),
	.w6(32'h3b8c9e49),
	.w7(32'h3ae74c4f),
	.w8(32'h3c3efc52),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5bce7),
	.w1(32'hbbd9ddf0),
	.w2(32'hbb95cf9c),
	.w3(32'h3b7a3839),
	.w4(32'hbaae4884),
	.w5(32'h3c4480ee),
	.w6(32'h3c241f68),
	.w7(32'hbbb9c78c),
	.w8(32'hbb522a4d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38f0b1),
	.w1(32'h3b642b9a),
	.w2(32'h3af05ada),
	.w3(32'hbadb45f4),
	.w4(32'hbab698fc),
	.w5(32'hbb624053),
	.w6(32'hbade8a9e),
	.w7(32'hbb6de68c),
	.w8(32'hbb096e67),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8e0a5),
	.w1(32'hbb9987b0),
	.w2(32'h39d7ed0a),
	.w3(32'hbb7eb93d),
	.w4(32'hbc118d67),
	.w5(32'hbc0aa286),
	.w6(32'hbb7c6925),
	.w7(32'hbb5182b8),
	.w8(32'h3b1223c1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a6486),
	.w1(32'hbb9659d3),
	.w2(32'hbb1873e8),
	.w3(32'h3b76cec6),
	.w4(32'h3a928b39),
	.w5(32'hbaaa7ce1),
	.w6(32'hbac819d0),
	.w7(32'h3ae82ea8),
	.w8(32'hbb8f6dd1),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d82457),
	.w1(32'h3b89a35b),
	.w2(32'h3b9b1197),
	.w3(32'h3c08fdde),
	.w4(32'h3b320c8b),
	.w5(32'h3c82b9c8),
	.w6(32'hbbbc697d),
	.w7(32'h3b1be8b9),
	.w8(32'h3bf2ec92),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3122c),
	.w1(32'hbbc10624),
	.w2(32'hbc039f77),
	.w3(32'h3b83c6ba),
	.w4(32'hbb658f14),
	.w5(32'hbbeeec81),
	.w6(32'h3bd16e10),
	.w7(32'h3b2efe86),
	.w8(32'hbb56bc71),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3957f1),
	.w1(32'hb94f47c9),
	.w2(32'hbc0f265b),
	.w3(32'hbb83c738),
	.w4(32'h3bb41fdc),
	.w5(32'h3cc5e6fc),
	.w6(32'h3b9334ed),
	.w7(32'hbb95f674),
	.w8(32'hba1111ea),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6152c9),
	.w1(32'hbc5e70c9),
	.w2(32'hbbd0dd4d),
	.w3(32'hbc0033b8),
	.w4(32'hbc79c224),
	.w5(32'hbca9a837),
	.w6(32'hbc37e40e),
	.w7(32'hbc19dc40),
	.w8(32'hbbcdee5a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc350f0b),
	.w1(32'h3c49b7bd),
	.w2(32'h3a0dbbc4),
	.w3(32'hbc41c14d),
	.w4(32'h3c8b3ea2),
	.w5(32'h3c231c77),
	.w6(32'hbc2ce5c4),
	.w7(32'h3c48e529),
	.w8(32'h3b6a9142),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923ae6b),
	.w1(32'h3bff384d),
	.w2(32'h3ab1246c),
	.w3(32'h3b255271),
	.w4(32'h3986bd46),
	.w5(32'h3ba34903),
	.w6(32'hbb4f6ffd),
	.w7(32'h3c1bc2e9),
	.w8(32'hbbdf9f12),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59548),
	.w1(32'hbbf7b1c5),
	.w2(32'h3b0a18d4),
	.w3(32'h3b8e4977),
	.w4(32'hbbaa356a),
	.w5(32'h3997473c),
	.w6(32'hbc234088),
	.w7(32'hbba2b52d),
	.w8(32'hbb1471c3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eb7d0),
	.w1(32'hbba6cf38),
	.w2(32'hbb0928c6),
	.w3(32'hbc64cd6a),
	.w4(32'hbaab292e),
	.w5(32'h3c402a9b),
	.w6(32'hbc5677a3),
	.w7(32'hbb62bc19),
	.w8(32'hbc1cb0b2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c07fa),
	.w1(32'hbb816882),
	.w2(32'hbaef917e),
	.w3(32'h3c68c6af),
	.w4(32'hbbbdbb15),
	.w5(32'hbc5e1ae7),
	.w6(32'h3b63caaa),
	.w7(32'hbb50d885),
	.w8(32'hba7ad067),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510fd3),
	.w1(32'h3ba5d658),
	.w2(32'h3b1d0e0c),
	.w3(32'h3aa553e9),
	.w4(32'h3bad1da6),
	.w5(32'hbb1acd64),
	.w6(32'hbb82223f),
	.w7(32'hb9a9b7db),
	.w8(32'h3b88d9b9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac62989),
	.w1(32'h3a6daf46),
	.w2(32'h3bcbde3e),
	.w3(32'h3bbf432e),
	.w4(32'h3a4f7b9d),
	.w5(32'h3bfac68e),
	.w6(32'hbb58dbe6),
	.w7(32'h3afa5b68),
	.w8(32'h3b948b91),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b794c7d),
	.w1(32'h3b7c3a68),
	.w2(32'hba38f897),
	.w3(32'h38e6b298),
	.w4(32'hbb112211),
	.w5(32'hbb58260d),
	.w6(32'h3a9d7ee9),
	.w7(32'hbb24481d),
	.w8(32'hbae27d43),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca739),
	.w1(32'h3b7b3f93),
	.w2(32'h3a8a1f3c),
	.w3(32'hbb739f3b),
	.w4(32'h3a62e114),
	.w5(32'hbb08b8fc),
	.w6(32'hba9590fb),
	.w7(32'h3b47f1b4),
	.w8(32'hb9e20254),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5e2e3),
	.w1(32'h3bf8e02c),
	.w2(32'h3bd43a94),
	.w3(32'hbc304020),
	.w4(32'h3abf6e38),
	.w5(32'hbb9bc0bf),
	.w6(32'hbc1f7c4a),
	.w7(32'h3bc331d3),
	.w8(32'hbabe66cf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053c6c),
	.w1(32'h3b96f714),
	.w2(32'h3c1b0e96),
	.w3(32'h3c35dc46),
	.w4(32'h3b93be0d),
	.w5(32'h3c938a08),
	.w6(32'h3c17a568),
	.w7(32'hb9a221da),
	.w8(32'h3c11e48e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b451c8b),
	.w1(32'h3b7f5de6),
	.w2(32'hbb9b5466),
	.w3(32'h3bda7f4b),
	.w4(32'h3b9cca84),
	.w5(32'hba806600),
	.w6(32'h3be4b0e0),
	.w7(32'h3a31b7e8),
	.w8(32'h3b2fd59c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0861e7),
	.w1(32'hbb50f105),
	.w2(32'hbb193d20),
	.w3(32'h3bbb2f2d),
	.w4(32'hba9a5497),
	.w5(32'hbbed196b),
	.w6(32'hbb15be75),
	.w7(32'h3ad1885b),
	.w8(32'hbb3c0442),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02512a),
	.w1(32'hbbab5d6a),
	.w2(32'hbb407a30),
	.w3(32'hbba3af97),
	.w4(32'hbb1febc9),
	.w5(32'hbba8a12d),
	.w6(32'hbb35260f),
	.w7(32'hbb9fc494),
	.w8(32'h3b0e6365),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb844bde),
	.w1(32'h3bdc69f7),
	.w2(32'hbaa1f554),
	.w3(32'h39dac96a),
	.w4(32'h3be10778),
	.w5(32'h3c3b86c0),
	.w6(32'h3b8c8194),
	.w7(32'h3b6ffc4a),
	.w8(32'h3bcba142),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0c21),
	.w1(32'hbb13726b),
	.w2(32'hbc4051ec),
	.w3(32'h3c65301e),
	.w4(32'h3bc3affb),
	.w5(32'hb8a0aea0),
	.w6(32'h3c5935bd),
	.w7(32'h3bcac9ff),
	.w8(32'hbc103317),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe351a4),
	.w1(32'hbbcaad15),
	.w2(32'hbc7091cb),
	.w3(32'h39c4f163),
	.w4(32'h3adde8af),
	.w5(32'h3ad60df1),
	.w6(32'hbbf242db),
	.w7(32'hbb8bc624),
	.w8(32'hbc81895d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2955f9),
	.w1(32'hbb662908),
	.w2(32'hbb800887),
	.w3(32'hbc0fb0fd),
	.w4(32'hbbc63b70),
	.w5(32'hbb7c1332),
	.w6(32'hbc61c5c1),
	.w7(32'hbbad3f88),
	.w8(32'h3b5146ae),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac32655),
	.w1(32'h3ad7effa),
	.w2(32'h3bd66016),
	.w3(32'hb9b0d1bd),
	.w4(32'h3b8944e2),
	.w5(32'h3b753696),
	.w6(32'h3a1c9fc8),
	.w7(32'h3a56ec15),
	.w8(32'hba4b13d8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d858),
	.w1(32'h39aaf24b),
	.w2(32'hbc27ca42),
	.w3(32'hbb05cd1c),
	.w4(32'h3b050311),
	.w5(32'hbc609816),
	.w6(32'hba9a3fdf),
	.w7(32'h3baa913e),
	.w8(32'hbc2fddc9),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5d1a),
	.w1(32'h3bc0682d),
	.w2(32'hbb8e3a23),
	.w3(32'hbb61a40c),
	.w4(32'h3c1104a9),
	.w5(32'hbb1c533e),
	.w6(32'hbbb2d862),
	.w7(32'h3c6e7118),
	.w8(32'hb9a19e57),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c26a8),
	.w1(32'hbb82fe9b),
	.w2(32'hba9f279d),
	.w3(32'hba704eca),
	.w4(32'hbbda94cb),
	.w5(32'hbb98b857),
	.w6(32'hbb320677),
	.w7(32'hbb662661),
	.w8(32'hba54deb3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843d23),
	.w1(32'hbbb766a1),
	.w2(32'h3b2c577d),
	.w3(32'hbbc746ef),
	.w4(32'hbba5b2cb),
	.w5(32'hbbf681e8),
	.w6(32'hbb1a3816),
	.w7(32'hbbe689c4),
	.w8(32'h3b3de26a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb780193),
	.w1(32'h3b8a6146),
	.w2(32'hbc24767d),
	.w3(32'h39d1977f),
	.w4(32'h3b22deb3),
	.w5(32'hbc90cb48),
	.w6(32'hbb6fa2ad),
	.w7(32'hbb40018f),
	.w8(32'hbc8cd984),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b641baf),
	.w1(32'hba192973),
	.w2(32'hbbc2106c),
	.w3(32'h3c2f2bba),
	.w4(32'hbb16c6e0),
	.w5(32'h3a865d3f),
	.w6(32'h3aff76e3),
	.w7(32'hbb96bd84),
	.w8(32'h3aa93a3b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b220e),
	.w1(32'h3bf87e8d),
	.w2(32'h3b5ba03e),
	.w3(32'h3c4769f3),
	.w4(32'h3c02fd87),
	.w5(32'h3c245423),
	.w6(32'h3923f66b),
	.w7(32'h3b24997a),
	.w8(32'h3ab76ee0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e55f1),
	.w1(32'hbb470dec),
	.w2(32'hbb8abb57),
	.w3(32'hba5e922e),
	.w4(32'hbb06d240),
	.w5(32'hbcbb0e46),
	.w6(32'hbb19c140),
	.w7(32'h3803e43f),
	.w8(32'hbb9fbc2b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc328919),
	.w1(32'h3ad8e87f),
	.w2(32'h3c8636f7),
	.w3(32'hbc48b35d),
	.w4(32'hbbffce64),
	.w5(32'h3c03269f),
	.w6(32'hbba9e4e6),
	.w7(32'hbae6c394),
	.w8(32'h3b6748fa),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c8d6b),
	.w1(32'hbb5279c9),
	.w2(32'h3b97d59f),
	.w3(32'h3b9eb3c2),
	.w4(32'hbc2e0156),
	.w5(32'h3ad87724),
	.w6(32'h3b84c4a6),
	.w7(32'hbb9caa5f),
	.w8(32'hba0b9c59),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24827e),
	.w1(32'hba1832c9),
	.w2(32'hbc137cba),
	.w3(32'h3bc062f5),
	.w4(32'hbbd631f3),
	.w5(32'hbc6e55d4),
	.w6(32'h3b97e410),
	.w7(32'hbbb20b1b),
	.w8(32'hbc50eb7f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e913fc),
	.w1(32'h3a0bacbc),
	.w2(32'h38ae940e),
	.w3(32'hbb2861a0),
	.w4(32'hb9cb2905),
	.w5(32'h3a0e526e),
	.w6(32'hbb3bd02a),
	.w7(32'hb9455494),
	.w8(32'hb913aa2f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a765667),
	.w1(32'hba892cb4),
	.w2(32'hba04d3b2),
	.w3(32'h3aa8f7a7),
	.w4(32'hba8a43b5),
	.w5(32'h38cf6e23),
	.w6(32'h3a8f1433),
	.w7(32'hb9b51ae5),
	.w8(32'h39e5762f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abaaf8),
	.w1(32'hba6cadeb),
	.w2(32'h39a17ea3),
	.w3(32'h398ddc5b),
	.w4(32'hb9f3ec8c),
	.w5(32'hb7c699d6),
	.w6(32'h3a018b91),
	.w7(32'h399ba2a7),
	.w8(32'h3a053c3c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a0a03),
	.w1(32'hba5e3f76),
	.w2(32'h3a232fa4),
	.w3(32'hba055651),
	.w4(32'hba6158bf),
	.w5(32'h3a8c3c7f),
	.w6(32'hba5a1d9e),
	.w7(32'hb815e5db),
	.w8(32'h3a5f21cc),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5a9a8),
	.w1(32'hb9afcbb1),
	.w2(32'hba09117a),
	.w3(32'h3a50fa0f),
	.w4(32'hb8b54dcf),
	.w5(32'hba0cdf4b),
	.w6(32'h3a365503),
	.w7(32'hb92041c0),
	.w8(32'hba7c9d4e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dce958),
	.w1(32'hba2b3be3),
	.w2(32'h3996df2a),
	.w3(32'hba3f9c10),
	.w4(32'hb9d00fd9),
	.w5(32'h39afd0a6),
	.w6(32'hba506b9a),
	.w7(32'hba6d332e),
	.w8(32'h397d6b44),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73dc86),
	.w1(32'hba82573f),
	.w2(32'hbab04abe),
	.w3(32'h3ad93cd3),
	.w4(32'hba0b619e),
	.w5(32'hba157f93),
	.w6(32'h3a41b470),
	.w7(32'hba48f0f5),
	.w8(32'hba12b048),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a2197),
	.w1(32'hba8111b2),
	.w2(32'hbac750d8),
	.w3(32'hba90352f),
	.w4(32'hbac6f8a1),
	.w5(32'hbadf725f),
	.w6(32'hba5537b6),
	.w7(32'hba84d866),
	.w8(32'hbabd230f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0023f0),
	.w1(32'hb9d3e51a),
	.w2(32'hbaf0bda0),
	.w3(32'hbb2f19aa),
	.w4(32'hb91b4e1a),
	.w5(32'hba205fe2),
	.w6(32'hbb1c5061),
	.w7(32'hba9ba8b5),
	.w8(32'hba9847aa),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab289a7),
	.w1(32'hba8d529a),
	.w2(32'hba76c06e),
	.w3(32'hbb0b40ff),
	.w4(32'hba4cc98b),
	.w5(32'hb92b504a),
	.w6(32'hbb3aa18f),
	.w7(32'hbab3d3d6),
	.w8(32'hb9893036),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d2b192),
	.w1(32'hb8c90e34),
	.w2(32'h39003670),
	.w3(32'h3a030190),
	.w4(32'h3892e276),
	.w5(32'h39c06dd5),
	.w6(32'hba15294d),
	.w7(32'hb9187103),
	.w8(32'hba00c22e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba123377),
	.w1(32'h3afd2dfe),
	.w2(32'h3a9766a9),
	.w3(32'hba87a215),
	.w4(32'h3b118392),
	.w5(32'h3a7823c4),
	.w6(32'hba961ae3),
	.w7(32'h3b03dd9b),
	.w8(32'h3a65c9f0),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa083b6),
	.w1(32'h39f3d187),
	.w2(32'h3a005108),
	.w3(32'h3a591209),
	.w4(32'h3a511258),
	.w5(32'h3a85dd19),
	.w6(32'h3a2a282f),
	.w7(32'h3a8dc652),
	.w8(32'h3a4ca692),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19b56f),
	.w1(32'h3a34c72e),
	.w2(32'hb93e9fa1),
	.w3(32'h39805a07),
	.w4(32'h391b3d70),
	.w5(32'hba847e0c),
	.w6(32'h3a154f43),
	.w7(32'hb9154cd9),
	.w8(32'hba5f4872),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d7f78),
	.w1(32'hb930c337),
	.w2(32'hba4c73d8),
	.w3(32'hba9cbc16),
	.w4(32'h3a4e4c75),
	.w5(32'h3a948e8e),
	.w6(32'hbaa7162b),
	.w7(32'h3a2318e6),
	.w8(32'h3ac15a5a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bf80b),
	.w1(32'hb9e624ac),
	.w2(32'h3991b620),
	.w3(32'h39274725),
	.w4(32'h378c1b29),
	.w5(32'h3a2fcb15),
	.w6(32'hba0034e8),
	.w7(32'hb8e4cddc),
	.w8(32'h3a2ff2f9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a508c3f),
	.w1(32'hb7e54169),
	.w2(32'hba5f3906),
	.w3(32'hb8d9f805),
	.w4(32'hbab4a19e),
	.w5(32'h389b0f79),
	.w6(32'h390aa1a9),
	.w7(32'hba9d9171),
	.w8(32'hb9c0be77),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b3729),
	.w1(32'hb9d36e91),
	.w2(32'h36ab8a65),
	.w3(32'hba91800e),
	.w4(32'hba355372),
	.w5(32'hba085ec3),
	.w6(32'hb9273e05),
	.w7(32'hb802581f),
	.w8(32'h389b7119),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933daca),
	.w1(32'h39d4e1f8),
	.w2(32'hb940798a),
	.w3(32'hb951af69),
	.w4(32'hb89fbd5d),
	.w5(32'hba61a9a4),
	.w6(32'hb9e64383),
	.w7(32'h3ae5f2d0),
	.w8(32'h3a352459),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac3a9c),
	.w1(32'h381a85cd),
	.w2(32'hba53c320),
	.w3(32'hb8768504),
	.w4(32'hba44015d),
	.w5(32'hb9815803),
	.w6(32'hba6854be),
	.w7(32'hba6af7dc),
	.w8(32'hb9bb6ada),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f60db6),
	.w1(32'hba94e74f),
	.w2(32'hb99fa5c9),
	.w3(32'h39e6e2b7),
	.w4(32'hba3d1240),
	.w5(32'hba205e79),
	.w6(32'hb91faade),
	.w7(32'hba078fd6),
	.w8(32'hb9c077c1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9181e65),
	.w1(32'h3a477e40),
	.w2(32'h3a2e6cb8),
	.w3(32'hb88f21c2),
	.w4(32'h3a46f151),
	.w5(32'h3a756ad4),
	.w6(32'hb9ebdee5),
	.w7(32'h3a8c5d29),
	.w8(32'h3a31c560),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2bdad),
	.w1(32'hba2388f6),
	.w2(32'hba031240),
	.w3(32'h3a0f388c),
	.w4(32'hbb075847),
	.w5(32'hba6e7a66),
	.w6(32'h3ac62747),
	.w7(32'hbb1cb0dc),
	.w8(32'hbaa15b3f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b00567),
	.w1(32'h3ab41224),
	.w2(32'h3ab5a1f8),
	.w3(32'h3a84866b),
	.w4(32'h3a5cc5e5),
	.w5(32'h3912dbc9),
	.w6(32'hba618ad3),
	.w7(32'h3987d78a),
	.w8(32'h3a005993),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4bf65),
	.w1(32'h3a104047),
	.w2(32'h3a25d643),
	.w3(32'h39603137),
	.w4(32'h3a5c073b),
	.w5(32'h3a98d519),
	.w6(32'h399950bb),
	.w7(32'h3a81f9ee),
	.w8(32'h3a9629fe),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32f3db),
	.w1(32'hb9e729b3),
	.w2(32'hba626694),
	.w3(32'h38781eba),
	.w4(32'hbad1543f),
	.w5(32'h38fe2603),
	.w6(32'hb931a7df),
	.w7(32'hba741628),
	.w8(32'hba080ee6),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabac026),
	.w1(32'hb7a3794e),
	.w2(32'hb9a9efc1),
	.w3(32'hba86dd21),
	.w4(32'hb808a0fe),
	.w5(32'h3a9aea74),
	.w6(32'hba9f9d75),
	.w7(32'hb98721a0),
	.w8(32'h399cbe71),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378d7a2c),
	.w1(32'h3974a086),
	.w2(32'h3a26f04b),
	.w3(32'hb9dbf854),
	.w4(32'h3982632b),
	.w5(32'h3aae449f),
	.w6(32'hb96d2ac4),
	.w7(32'h3a64aca8),
	.w8(32'h39c4dc28),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a814f),
	.w1(32'h3a7e0abe),
	.w2(32'h3aa88633),
	.w3(32'hb9f69c56),
	.w4(32'h3a3fd314),
	.w5(32'h3afcdab0),
	.w6(32'hba25aac3),
	.w7(32'h39e3c697),
	.w8(32'h3aad5591),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba513994),
	.w1(32'hb9f3b896),
	.w2(32'hba4def17),
	.w3(32'hba393b23),
	.w4(32'hba010087),
	.w5(32'hb770f3da),
	.w6(32'hb95a8ea8),
	.w7(32'hba4c01d5),
	.w8(32'hba3a7791),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0e8e3),
	.w1(32'hbb4e7bc2),
	.w2(32'hbb1b4259),
	.w3(32'hb8aa1907),
	.w4(32'hbb300274),
	.w5(32'hbac168c1),
	.w6(32'hb98906bd),
	.w7(32'hbac4697a),
	.w8(32'hba8fde86),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca6ce1),
	.w1(32'hb96d67e1),
	.w2(32'hb996cd25),
	.w3(32'hb9e1b97d),
	.w4(32'hba052628),
	.w5(32'hb9a56e15),
	.w6(32'hbab7d1b7),
	.w7(32'hb90dda0c),
	.w8(32'hba1bb77c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38288a36),
	.w1(32'h3953d47f),
	.w2(32'hb9d15c5f),
	.w3(32'hb76239f2),
	.w4(32'h396d6580),
	.w5(32'h39a4361b),
	.w6(32'hb81f6b2b),
	.w7(32'hb82524cd),
	.w8(32'h3a790d99),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da69ab),
	.w1(32'h39b2f6ec),
	.w2(32'hb8fadfe5),
	.w3(32'hba4a7d54),
	.w4(32'hba0b5dc7),
	.w5(32'h395d9f17),
	.w6(32'h3a1f2ba6),
	.w7(32'hb740b7ca),
	.w8(32'hb9b4c597),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b16e1),
	.w1(32'hba39b8df),
	.w2(32'hb88fc3d1),
	.w3(32'hba167c8d),
	.w4(32'h3939fca8),
	.w5(32'h3a2f17b6),
	.w6(32'hba800601),
	.w7(32'hb864a30f),
	.w8(32'h391aa80b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e2af7),
	.w1(32'h3a0c02c1),
	.w2(32'hba5fcb1f),
	.w3(32'hba1654f5),
	.w4(32'h39c1f1d1),
	.w5(32'hba4e907f),
	.w6(32'hb92ab188),
	.w7(32'hb5cb9b48),
	.w8(32'h390d6006),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a8cd7),
	.w1(32'h3a0a75f1),
	.w2(32'h3a2a27f1),
	.w3(32'hba76c701),
	.w4(32'h3a133500),
	.w5(32'h3a811dee),
	.w6(32'hb91b1da8),
	.w7(32'hb8f9c8ca),
	.w8(32'h3a4a9639),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a89722),
	.w1(32'hba11ede5),
	.w2(32'hba33d8b6),
	.w3(32'h3a2ebc1e),
	.w4(32'h380bd326),
	.w5(32'hba141e25),
	.w6(32'h3a5761a2),
	.w7(32'h391774bb),
	.w8(32'hb75dd53c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e2f2c),
	.w1(32'h39e135cb),
	.w2(32'h39a11741),
	.w3(32'hb98094c7),
	.w4(32'h38c28851),
	.w5(32'h3a6795b3),
	.w6(32'h38bec22c),
	.w7(32'hba079dea),
	.w8(32'hb923d471),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a145b2f),
	.w1(32'h3ac580f8),
	.w2(32'h3a83de17),
	.w3(32'h3a0f0b03),
	.w4(32'h3b07e9d2),
	.w5(32'h3a5e6bd9),
	.w6(32'h3a113f8c),
	.w7(32'h3a479806),
	.w8(32'h3a415281),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16c2ef),
	.w1(32'hba7acfcb),
	.w2(32'hbac8a335),
	.w3(32'h38bc664f),
	.w4(32'hba272f53),
	.w5(32'hba49d604),
	.w6(32'h3aaaf1a6),
	.w7(32'hb990fbeb),
	.w8(32'h39e1788e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19641f),
	.w1(32'hba0a1bb3),
	.w2(32'hb8f324bf),
	.w3(32'hbadff55f),
	.w4(32'hb97f00d8),
	.w5(32'h39b3f740),
	.w6(32'hb8932c1a),
	.w7(32'hba2a0387),
	.w8(32'hba85d3fe),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e908f),
	.w1(32'h3a3e3229),
	.w2(32'h3a4237e8),
	.w3(32'hba82b3df),
	.w4(32'h39d4e876),
	.w5(32'h3a1005e6),
	.w6(32'hbaba796e),
	.w7(32'hb9b3a42d),
	.w8(32'hb9e43d5c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9743376),
	.w1(32'h37dda785),
	.w2(32'h38f1f96d),
	.w3(32'hbaeca811),
	.w4(32'h39faac61),
	.w5(32'h3a478f93),
	.w6(32'hbaea82b4),
	.w7(32'h3a1202c0),
	.w8(32'h394650fd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399552e4),
	.w1(32'hbac98c3d),
	.w2(32'hb9ed92d0),
	.w3(32'hb9cd9192),
	.w4(32'hba1009b1),
	.w5(32'h393ce02e),
	.w6(32'hb8e3adfb),
	.w7(32'hb94f1aa6),
	.w8(32'hba83ca7e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ab08fe),
	.w1(32'hb9df05d4),
	.w2(32'h39fb5c64),
	.w3(32'hba3eb581),
	.w4(32'hb9fbaccf),
	.w5(32'h39aa17a8),
	.w6(32'hb936e98e),
	.w7(32'hba4fb493),
	.w8(32'hb9f16303),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9574fb9),
	.w1(32'h37b9331d),
	.w2(32'hba21e306),
	.w3(32'h39fc9c59),
	.w4(32'hb90e28df),
	.w5(32'h3818b17d),
	.w6(32'h3999cacc),
	.w7(32'hb9fb39f3),
	.w8(32'hb99fa857),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10452f),
	.w1(32'hba06f871),
	.w2(32'hbae030dc),
	.w3(32'hba873967),
	.w4(32'h392973fc),
	.w5(32'hba1ea652),
	.w6(32'hba1e6c6e),
	.w7(32'hb91820cd),
	.w8(32'hb90e5917),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab87219),
	.w1(32'h39fe7bcd),
	.w2(32'h3aa76a4e),
	.w3(32'hbab30c1d),
	.w4(32'h3a647086),
	.w5(32'h39e602ec),
	.w6(32'h390706dc),
	.w7(32'h3a9e98d0),
	.w8(32'h3a792a5e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ef578),
	.w1(32'h39e61e70),
	.w2(32'hb698758e),
	.w3(32'hba73919a),
	.w4(32'h39c0d6da),
	.w5(32'hba2c91e0),
	.w6(32'hb98faf1a),
	.w7(32'h3ac39cec),
	.w8(32'h39f7e238),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884141c),
	.w1(32'h399c3d04),
	.w2(32'hb8c67e5d),
	.w3(32'hba367cfb),
	.w4(32'h39e67c8f),
	.w5(32'h3ada2f73),
	.w6(32'hb9b9c6cb),
	.w7(32'h3a395f0f),
	.w8(32'h3966d1f6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b81ad),
	.w1(32'h3a0a88a5),
	.w2(32'hba29b2bd),
	.w3(32'hba8c1eea),
	.w4(32'hb8a0d368),
	.w5(32'hb9817da6),
	.w6(32'hb93fcc19),
	.w7(32'h3970b074),
	.w8(32'hba1c4781),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e957a),
	.w1(32'hba755662),
	.w2(32'hba5c1c88),
	.w3(32'hba1acb91),
	.w4(32'h39d954c5),
	.w5(32'h39cd538e),
	.w6(32'hb99c04a7),
	.w7(32'hbaa038fb),
	.w8(32'hb9802bd1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9111686),
	.w1(32'h398719a1),
	.w2(32'hb91ad0c4),
	.w3(32'hb966def6),
	.w4(32'hb9dc70d0),
	.w5(32'hb90c2156),
	.w6(32'h39c58fe5),
	.w7(32'h37e7a9f4),
	.w8(32'hba0a4f31),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d2edb),
	.w1(32'hba4dabc4),
	.w2(32'hb984e310),
	.w3(32'hba8fd299),
	.w4(32'hb9d95834),
	.w5(32'h3a70ca2f),
	.w6(32'hbaa8335e),
	.w7(32'hba3e094c),
	.w8(32'hb981a14f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39663b45),
	.w1(32'h3a370b21),
	.w2(32'h3a2a837b),
	.w3(32'h3a759566),
	.w4(32'h39465100),
	.w5(32'hba311d3b),
	.w6(32'hb93a7e40),
	.w7(32'h398a16d3),
	.w8(32'h39c8737d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46ecef),
	.w1(32'hbb1709ec),
	.w2(32'hba05e4df),
	.w3(32'hb984035a),
	.w4(32'hbb10bd6d),
	.w5(32'hb9c57098),
	.w6(32'h3a1aa42b),
	.w7(32'hba80611d),
	.w8(32'hb9d96f08),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01c797),
	.w1(32'hba3f9e53),
	.w2(32'hb9b82e27),
	.w3(32'hba9a94ed),
	.w4(32'hbad22f4b),
	.w5(32'hbb08a543),
	.w6(32'hb9d73270),
	.w7(32'hb9da8fb4),
	.w8(32'hb9ce03dc),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d9104),
	.w1(32'h3a71084b),
	.w2(32'hb93d04f4),
	.w3(32'h3989a3db),
	.w4(32'h39a22489),
	.w5(32'hb93c3756),
	.w6(32'h3a2ddeb1),
	.w7(32'hba515704),
	.w8(32'hb9cb8537),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule