module layer_8_featuremap_229(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24f4d6),
	.w1(32'h3c8c3cf3),
	.w2(32'h3d25c362),
	.w3(32'h3bc4a1ab),
	.w4(32'h3c8b65d1),
	.w5(32'h3c2a28e7),
	.w6(32'h3c5870ec),
	.w7(32'h3c67ea8b),
	.w8(32'h3caff62c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8402fd),
	.w1(32'h3a65052e),
	.w2(32'h3a64b06d),
	.w3(32'hbafe40df),
	.w4(32'hbbb95cfd),
	.w5(32'hbbb3028f),
	.w6(32'h3aca1972),
	.w7(32'hb91900ce),
	.w8(32'hbb35bd6c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadc1bd),
	.w1(32'hbc1dd971),
	.w2(32'hbbb9ebc4),
	.w3(32'hbc11ff35),
	.w4(32'hbbe21373),
	.w5(32'hbc4281c5),
	.w6(32'hbb52d532),
	.w7(32'hbb4b4fb5),
	.w8(32'hbb8b1287),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1e0ba),
	.w1(32'h3bae6f22),
	.w2(32'h3b868ec6),
	.w3(32'hbc6efb09),
	.w4(32'h3a5ad2a7),
	.w5(32'hbbba1ad7),
	.w6(32'h3c390a9c),
	.w7(32'h3bc3de12),
	.w8(32'h3880834c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a0c39),
	.w1(32'h3c1c7931),
	.w2(32'h3ad9199a),
	.w3(32'hbc907222),
	.w4(32'h3bdd9277),
	.w5(32'h3af8ab36),
	.w6(32'h3bb0a378),
	.w7(32'hbbb069a2),
	.w8(32'hbc287298),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01b0a5),
	.w1(32'h3c639e07),
	.w2(32'h3c8fce02),
	.w3(32'hbba5b9b1),
	.w4(32'h3c15a903),
	.w5(32'h3c36c9c5),
	.w6(32'h3c146801),
	.w7(32'h3b5b5476),
	.w8(32'hbabe4544),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c54e4),
	.w1(32'h3a89970d),
	.w2(32'hbbb4e1eb),
	.w3(32'hbb129116),
	.w4(32'h3b457b93),
	.w5(32'hbb446d36),
	.w6(32'h3a181d9e),
	.w7(32'hbb9cf8b1),
	.w8(32'hbbb36015),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe24ca5),
	.w1(32'h3cab0f0a),
	.w2(32'h3c21a05f),
	.w3(32'hbb63ac43),
	.w4(32'h3c51ca10),
	.w5(32'hbbff48b3),
	.w6(32'h3bcee6e2),
	.w7(32'h3b9c1fa6),
	.w8(32'hbb27876a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b1b4c),
	.w1(32'h3c900c42),
	.w2(32'hba86aa7b),
	.w3(32'hbc9fc655),
	.w4(32'h3be07608),
	.w5(32'hbbe3ea2f),
	.w6(32'h3c206cc6),
	.w7(32'hbc0be912),
	.w8(32'hbc4e0892),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e390d),
	.w1(32'h3c9b9978),
	.w2(32'h3cbe1802),
	.w3(32'hbc4ddcd7),
	.w4(32'h3c9d7e55),
	.w5(32'h3c8a712f),
	.w6(32'h3b99e8d4),
	.w7(32'h3ca99c70),
	.w8(32'h39afe676),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c099682),
	.w1(32'hbccf008f),
	.w2(32'hbca54503),
	.w3(32'hb9570d7b),
	.w4(32'hbc9e583f),
	.w5(32'hbcc05fcb),
	.w6(32'hbc1f6a4b),
	.w7(32'hbb73d953),
	.w8(32'h3b84e19b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9e737),
	.w1(32'h3c07a594),
	.w2(32'h3ba96070),
	.w3(32'hbbf5b310),
	.w4(32'h3bebb936),
	.w5(32'hbb04710e),
	.w6(32'h3bb4355a),
	.w7(32'h3b01798c),
	.w8(32'hba244742),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d77af),
	.w1(32'h3bc13581),
	.w2(32'hbac00f7b),
	.w3(32'hbb4f526b),
	.w4(32'hbbc74b4b),
	.w5(32'hbc17deff),
	.w6(32'hbaa77da8),
	.w7(32'hba47053c),
	.w8(32'h3bddc123),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb6071),
	.w1(32'h3beebec1),
	.w2(32'h3c21d8a1),
	.w3(32'hbc0929bf),
	.w4(32'h3c39b19c),
	.w5(32'h3ba1daff),
	.w6(32'h3c7543ca),
	.w7(32'h3b125a76),
	.w8(32'hbb2a049d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2c0ad),
	.w1(32'h3c95f4ba),
	.w2(32'hbb8dfccb),
	.w3(32'h3af85b3a),
	.w4(32'h3c3b92a2),
	.w5(32'hbbc95206),
	.w6(32'h3c4ad31b),
	.w7(32'hbb6cfaf0),
	.w8(32'hbc417f2c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77dc01),
	.w1(32'h3bd9faf9),
	.w2(32'h3bd74ddf),
	.w3(32'hbc7bb7d8),
	.w4(32'h3b6ed477),
	.w5(32'hba8a5f87),
	.w6(32'h3c067efe),
	.w7(32'hbbeb4394),
	.w8(32'h3b3ccf3f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb18468),
	.w1(32'hbbea37d6),
	.w2(32'hbc0c9a88),
	.w3(32'hbb660861),
	.w4(32'hbbc3cdc3),
	.w5(32'hbaf40c99),
	.w6(32'hbc02edd8),
	.w7(32'hbc481629),
	.w8(32'h3bfc00ad),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6031e3),
	.w1(32'hbb4aab6e),
	.w2(32'hb88e2b04),
	.w3(32'h3c1e3d77),
	.w4(32'h3ab6d168),
	.w5(32'hbbef6461),
	.w6(32'hbc12ca76),
	.w7(32'h3a8c8264),
	.w8(32'h3ad32d17),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb829c),
	.w1(32'h3c3ed73e),
	.w2(32'h3c3ed90c),
	.w3(32'hbc0c044b),
	.w4(32'h3c3c4e53),
	.w5(32'h3c4c7826),
	.w6(32'h3c3cda08),
	.w7(32'h3bce41b7),
	.w8(32'h38032ae5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a1483),
	.w1(32'h3a894874),
	.w2(32'hbb89763e),
	.w3(32'h3c31b28d),
	.w4(32'h3b1b6a16),
	.w5(32'hbb6c6e90),
	.w6(32'h3b4531c4),
	.w7(32'h3b2c9cd6),
	.w8(32'h3b2082b4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a577fbb),
	.w1(32'hbd7aae31),
	.w2(32'hbd9f2444),
	.w3(32'hbaa43f95),
	.w4(32'hbd246453),
	.w5(32'hbd6ba9c4),
	.w6(32'hbcdef682),
	.w7(32'hbd0648d6),
	.w8(32'hbc06a0d6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd17a7cd),
	.w1(32'h3c4b6b6a),
	.w2(32'h3c44aaed),
	.w3(32'hbcf56c8b),
	.w4(32'h3c55ee70),
	.w5(32'h3c552f84),
	.w6(32'h3be71b84),
	.w7(32'h3b91b838),
	.w8(32'h3b3cdd44),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65564e),
	.w1(32'hba9e2a3d),
	.w2(32'h3b816c3d),
	.w3(32'h3c1ca1eb),
	.w4(32'hbc08335e),
	.w5(32'h3ae4c863),
	.w6(32'h3b94b40a),
	.w7(32'h3b6a4081),
	.w8(32'hbc0a5132),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4b06),
	.w1(32'h3c5a2855),
	.w2(32'h3c361694),
	.w3(32'h3a1e2642),
	.w4(32'h3b9d2139),
	.w5(32'h3b9e6d57),
	.w6(32'h3a726789),
	.w7(32'h3b0de713),
	.w8(32'h3b29c242),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc01e2a),
	.w1(32'hb9a5f87b),
	.w2(32'hbc62b163),
	.w3(32'h3ba2ec23),
	.w4(32'hbbee501e),
	.w5(32'hbb5c6097),
	.w6(32'h3c828e40),
	.w7(32'h3c3bb448),
	.w8(32'hbb63618c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44bfbc),
	.w1(32'hbcc2f598),
	.w2(32'hbd274348),
	.w3(32'h3b80b6aa),
	.w4(32'hbca24a8c),
	.w5(32'hbcfd251a),
	.w6(32'hbc96d23e),
	.w7(32'hbcd72d40),
	.w8(32'hbbe7d6a1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf5dc6c),
	.w1(32'hbbd05331),
	.w2(32'hbb12136e),
	.w3(32'hbcb985f6),
	.w4(32'h3ba4b59c),
	.w5(32'hbc030aff),
	.w6(32'h395823cd),
	.w7(32'h3b30d0a0),
	.w8(32'h3b376172),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afd051),
	.w1(32'hbcf797c8),
	.w2(32'hbd35487a),
	.w3(32'h3aa090f3),
	.w4(32'hbc9ef491),
	.w5(32'hbcf3240b),
	.w6(32'hbccae7db),
	.w7(32'hbcd8c890),
	.w8(32'hbc927aa7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec4e30),
	.w1(32'h3c8b48fd),
	.w2(32'h3c9af170),
	.w3(32'hbc985868),
	.w4(32'h3c97efd9),
	.w5(32'h3c4218b3),
	.w6(32'h3b4fce96),
	.w7(32'h3c06ee36),
	.w8(32'h3c0ad958),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12e52a),
	.w1(32'h3c493168),
	.w2(32'h3bc54cca),
	.w3(32'hbb88ccfe),
	.w4(32'h3bf48c6b),
	.w5(32'h3b55459b),
	.w6(32'h3ae2ef17),
	.w7(32'h3af69993),
	.w8(32'h3c9242cb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8522a6),
	.w1(32'h3ac5c8df),
	.w2(32'hbb8fe0cd),
	.w3(32'h3c6ed0c8),
	.w4(32'h3c8e9dae),
	.w5(32'h3ba01094),
	.w6(32'hbbe736ee),
	.w7(32'hba8c251c),
	.w8(32'h3bd0aafa),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08885),
	.w1(32'hbcca0f47),
	.w2(32'hbc817b4a),
	.w3(32'hbc11c564),
	.w4(32'hbc614021),
	.w5(32'hbc3d592e),
	.w6(32'hbc5f87de),
	.w7(32'hbc111351),
	.w8(32'hbaf8916e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa74bc),
	.w1(32'h3a51f35b),
	.w2(32'h3c0a6b74),
	.w3(32'hbaab8dce),
	.w4(32'hbb81312e),
	.w5(32'h3b3c4e03),
	.w6(32'h3bab4e4c),
	.w7(32'h3b082e8a),
	.w8(32'hbb979681),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cd9ee),
	.w1(32'h3b75d4dd),
	.w2(32'h3a7aba54),
	.w3(32'hbb7b4249),
	.w4(32'h3abe147c),
	.w5(32'h3bc606d0),
	.w6(32'h3a84ee80),
	.w7(32'h39f4bc4a),
	.w8(32'h3b82414b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd21bb2),
	.w1(32'h3c8ea8ee),
	.w2(32'h3c625841),
	.w3(32'h3ac71fa6),
	.w4(32'hbbe0ca1b),
	.w5(32'h3b89924d),
	.w6(32'h3a336f6e),
	.w7(32'h3bdfe4f1),
	.w8(32'h3bb0b9de),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b745422),
	.w1(32'hbb871cfd),
	.w2(32'hbc12ad4d),
	.w3(32'hbb5866d8),
	.w4(32'hbac95358),
	.w5(32'hbbaec587),
	.w6(32'hb8f9d55c),
	.w7(32'hbbe24ebf),
	.w8(32'hbb85e694),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac87e5c),
	.w1(32'h3a1da033),
	.w2(32'h39843cbc),
	.w3(32'h38e8bd34),
	.w4(32'hbae6c21b),
	.w5(32'hbb0942d1),
	.w6(32'hba8de8ed),
	.w7(32'h3abfeeaa),
	.w8(32'hbad8c71e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e258e),
	.w1(32'h3ccfadc0),
	.w2(32'h3c0dca01),
	.w3(32'h3abb3cc3),
	.w4(32'h3c22dc35),
	.w5(32'h3b6d17a5),
	.w6(32'h3c95d8b0),
	.w7(32'h3b6098b7),
	.w8(32'hbc0c1dfc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7312d),
	.w1(32'h3bd57d6f),
	.w2(32'hbc2e9d89),
	.w3(32'hbbf51b6c),
	.w4(32'h3bb7e9ae),
	.w5(32'hbbf2500c),
	.w6(32'h3b0ec84b),
	.w7(32'hbb881cb4),
	.w8(32'hbbb01952),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cadb2),
	.w1(32'h3b9e9c50),
	.w2(32'h3bf27a29),
	.w3(32'hbbc68062),
	.w4(32'hbb0e9be7),
	.w5(32'h3c5745e2),
	.w6(32'h3b2dd1a3),
	.w7(32'h3aee8ac8),
	.w8(32'h3b92cf22),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3633f1),
	.w1(32'hbbfe29a0),
	.w2(32'hba75de83),
	.w3(32'h3c557a07),
	.w4(32'hbbf4826b),
	.w5(32'hbb23eeb4),
	.w6(32'hbb9a71bc),
	.w7(32'h3ad9a273),
	.w8(32'h3bdd5d5b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc67a93),
	.w1(32'hbcf2062a),
	.w2(32'hbd28c38a),
	.w3(32'h3b7dc232),
	.w4(32'hbc86541c),
	.w5(32'hbcb88aae),
	.w6(32'hbc3f8f1e),
	.w7(32'hbcbd0061),
	.w8(32'hb92cf52c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4527f6),
	.w1(32'h39b56c6f),
	.w2(32'h3c2f0197),
	.w3(32'hbb6872b7),
	.w4(32'hbb9f50a6),
	.w5(32'hba2c631e),
	.w6(32'h3bcda25d),
	.w7(32'h3c8737a8),
	.w8(32'h3b8e9892),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b5a843),
	.w1(32'h3c3c2685),
	.w2(32'h3c8badc6),
	.w3(32'hbb09b335),
	.w4(32'h3c06925e),
	.w5(32'h3c2edaa4),
	.w6(32'h3c70b31f),
	.w7(32'h3c30807b),
	.w8(32'h3c26302a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c5f0d),
	.w1(32'hba124f90),
	.w2(32'h3801016e),
	.w3(32'h3c3c8476),
	.w4(32'hbbe4ad37),
	.w5(32'hbb7f5e64),
	.w6(32'hbab77c5c),
	.w7(32'hbb2d75a1),
	.w8(32'hbb282c3f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b0621),
	.w1(32'h3b372b6e),
	.w2(32'hbbd41848),
	.w3(32'hbc260ce0),
	.w4(32'h3b750ef8),
	.w5(32'hbb9edcd5),
	.w6(32'h3bbb399a),
	.w7(32'h3a27b577),
	.w8(32'h3bb072f9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18ff22),
	.w1(32'h3c285783),
	.w2(32'hbcb23c54),
	.w3(32'hb9a97197),
	.w4(32'h3c5f49f6),
	.w5(32'hbc103b2e),
	.w6(32'h3a4cf2ff),
	.w7(32'hbc9405a2),
	.w8(32'hbcb24055),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01a28e),
	.w1(32'h3bfc371f),
	.w2(32'h3bdf17d7),
	.w3(32'hbcb2f3a2),
	.w4(32'h3b8ab41e),
	.w5(32'h3bc8fda0),
	.w6(32'h3b9d568d),
	.w7(32'h3c202527),
	.w8(32'h3b3982b7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d1c7b0),
	.w1(32'h3c1b0989),
	.w2(32'h3c1f7ab0),
	.w3(32'hbadb8a08),
	.w4(32'h3b97c2ff),
	.w5(32'h3c3c9e20),
	.w6(32'h3baab959),
	.w7(32'h3a436ca2),
	.w8(32'h3c086d3f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f1cf1),
	.w1(32'hbc31b8b3),
	.w2(32'hbcf570a0),
	.w3(32'hb9202493),
	.w4(32'hbb941549),
	.w5(32'hbcc383fb),
	.w6(32'hbc9cffa6),
	.w7(32'hbc974df4),
	.w8(32'hbc4af6ef),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccfddf2),
	.w1(32'hba1b4a61),
	.w2(32'hbbabd430),
	.w3(32'hbca7097e),
	.w4(32'h3b6f73b3),
	.w5(32'hbb3b429f),
	.w6(32'h3b612df7),
	.w7(32'hbb2e8038),
	.w8(32'h3aaf2cd0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2c0ea),
	.w1(32'hbaeec431),
	.w2(32'hbbddd629),
	.w3(32'h3ab5b347),
	.w4(32'h3ab009aa),
	.w5(32'hbb590df1),
	.w6(32'h3b3ea6eb),
	.w7(32'hbac2d001),
	.w8(32'h3bd4f24d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e0eee),
	.w1(32'h3c86f00c),
	.w2(32'h3b9f967d),
	.w3(32'hbaf3837d),
	.w4(32'h3bfa1111),
	.w5(32'h3973e692),
	.w6(32'h3c3f44d5),
	.w7(32'hba9de7b9),
	.w8(32'hbc11327b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28a521),
	.w1(32'hbb48a5ac),
	.w2(32'hbc786c45),
	.w3(32'hbc195931),
	.w4(32'hba9dfe73),
	.w5(32'hbc6732ed),
	.w6(32'hbb63eb9a),
	.w7(32'hbbe8c1df),
	.w8(32'hbb60c93d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02812b),
	.w1(32'h3afe1b06),
	.w2(32'hbc0e2b18),
	.w3(32'hbbcc7afc),
	.w4(32'h3b9ffc22),
	.w5(32'hbbcaaa65),
	.w6(32'hbb485d6d),
	.w7(32'hbc9dd86b),
	.w8(32'hba25cb1e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49c3f6),
	.w1(32'h3bac285a),
	.w2(32'h3c9206c0),
	.w3(32'hbc19baf7),
	.w4(32'h3c6c5f32),
	.w5(32'h3c3b8e07),
	.w6(32'h3c244c04),
	.w7(32'h3b45bf4f),
	.w8(32'h3b7f59fa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd28c05),
	.w1(32'h3d00a2f7),
	.w2(32'h3c80b63b),
	.w3(32'h3c189957),
	.w4(32'h3d1079ed),
	.w5(32'h3bd76e17),
	.w6(32'h3c77fad7),
	.w7(32'h3bb4853d),
	.w8(32'hbc1b9bf9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0fa77),
	.w1(32'hbb8763e4),
	.w2(32'h3c4dce89),
	.w3(32'hbc462587),
	.w4(32'hbbbbc41f),
	.w5(32'h3b8c8c2c),
	.w6(32'hbbdf58bb),
	.w7(32'h3c17a70f),
	.w8(32'h3c21ebdb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26b162),
	.w1(32'h3b557eb9),
	.w2(32'hbbf3e414),
	.w3(32'h3af0e45b),
	.w4(32'h3a5d17f3),
	.w5(32'hbbfe2236),
	.w6(32'hb9d14def),
	.w7(32'hbbc16d18),
	.w8(32'hbbb27e0d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc202538),
	.w1(32'h3c3a5f93),
	.w2(32'h3bd3ff64),
	.w3(32'hbbfeece6),
	.w4(32'h3c11585e),
	.w5(32'h3bc7cc43),
	.w6(32'h3b210dbc),
	.w7(32'h3aaf04cd),
	.w8(32'h38ef6a02),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb5228),
	.w1(32'h3c50656b),
	.w2(32'h3c0cf3ff),
	.w3(32'h3a4f62fd),
	.w4(32'h3b0aab6f),
	.w5(32'hbb0d5644),
	.w6(32'h3cabd04d),
	.w7(32'h3c842dc0),
	.w8(32'h3b9359ce),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c087bbd),
	.w1(32'h3c4edb70),
	.w2(32'h3a41acf8),
	.w3(32'hbb76bcb2),
	.w4(32'hbc0b7dd4),
	.w5(32'hbc5c4254),
	.w6(32'h3c65d442),
	.w7(32'h3bab51db),
	.w8(32'hbb85ca56),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba22fdd),
	.w1(32'hbc0e05a3),
	.w2(32'h3cef54ac),
	.w3(32'h3abfef90),
	.w4(32'hbaa3d96c),
	.w5(32'h3cf4c739),
	.w6(32'hbc0ef287),
	.w7(32'h3c8c4269),
	.w8(32'h3cc534ef),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d41f2ce),
	.w1(32'h3acf1e9f),
	.w2(32'hbbbd7ad1),
	.w3(32'h3d402c8e),
	.w4(32'h3af5d035),
	.w5(32'hbbdb7595),
	.w6(32'h3bbee58c),
	.w7(32'hbaf7d523),
	.w8(32'hbbb55eb4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1262b),
	.w1(32'h3af633bb),
	.w2(32'hbac735b6),
	.w3(32'hbc1b450e),
	.w4(32'h3ae6b813),
	.w5(32'hbb783fec),
	.w6(32'h3ac51146),
	.w7(32'h3a9d7385),
	.w8(32'hbb10d0bd),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac0c7),
	.w1(32'h3b00d96e),
	.w2(32'h3c1a9683),
	.w3(32'hbc11c63c),
	.w4(32'h3b2d1cbb),
	.w5(32'h3c097fb4),
	.w6(32'h3bc54f3a),
	.w7(32'h3beedca7),
	.w8(32'h3b4c916b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00206f),
	.w1(32'h3d02d7c6),
	.w2(32'h3d08479e),
	.w3(32'h3c176a5c),
	.w4(32'h3c92e51b),
	.w5(32'h3c401ee3),
	.w6(32'h3c9ea7a1),
	.w7(32'h3c365d07),
	.w8(32'h3b913c57),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9b463),
	.w1(32'hbd38c622),
	.w2(32'hbd8a76ba),
	.w3(32'h3aa50893),
	.w4(32'hbd03744f),
	.w5(32'hbd411dc1),
	.w6(32'hbd036340),
	.w7(32'hbd2c19bd),
	.w8(32'hbcb14363),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd66d018),
	.w1(32'h3c4504ff),
	.w2(32'h3c21698d),
	.w3(32'hbd2828de),
	.w4(32'h3c9f0b78),
	.w5(32'h3c231067),
	.w6(32'h3b36d3e4),
	.w7(32'h3b1f8cc8),
	.w8(32'hbaff7a6c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d2b89),
	.w1(32'h3a9f31f9),
	.w2(32'hbc132613),
	.w3(32'h3b85f50d),
	.w4(32'hbb67cbb1),
	.w5(32'hbcbfb9c1),
	.w6(32'h3ba2d305),
	.w7(32'hbc01a34f),
	.w8(32'hbc383e9b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8eaebc),
	.w1(32'h3bcafda7),
	.w2(32'hbc9b39b8),
	.w3(32'hbc8a9eb1),
	.w4(32'h3bd54c43),
	.w5(32'hbc222188),
	.w6(32'h3c1ffaf0),
	.w7(32'hbc114486),
	.w8(32'hbbac88e0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc987188),
	.w1(32'h3c8c5185),
	.w2(32'h3c236ec9),
	.w3(32'hbc57d162),
	.w4(32'h3c7e4e61),
	.w5(32'hbb7a4375),
	.w6(32'h3a8093c3),
	.w7(32'h3a8411a4),
	.w8(32'h3a935c99),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacb9fc),
	.w1(32'h3c7148e0),
	.w2(32'h3c45a609),
	.w3(32'hbc261a75),
	.w4(32'h3c51926b),
	.w5(32'h3be45516),
	.w6(32'h3bb5f32c),
	.w7(32'h3c11c1e0),
	.w8(32'h3c3f2463),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac30dcc),
	.w1(32'h3bf3ff10),
	.w2(32'h3b15cf2a),
	.w3(32'h3b5dd301),
	.w4(32'h3ac6b353),
	.w5(32'hbb119b70),
	.w6(32'h3bb83adf),
	.w7(32'hba9e2e0f),
	.w8(32'h3a66393b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2f90a),
	.w1(32'hbba74d7f),
	.w2(32'hbca9a294),
	.w3(32'hbbd37585),
	.w4(32'hbb17aa31),
	.w5(32'hbba9610f),
	.w6(32'h3ac1e980),
	.w7(32'hbb9aa21c),
	.w8(32'h3b80c58f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63a9ea),
	.w1(32'h3c3267fb),
	.w2(32'h3b4b1055),
	.w3(32'h3bef709d),
	.w4(32'h3c190ab6),
	.w5(32'hbc07120c),
	.w6(32'h3bc83377),
	.w7(32'h3999717e),
	.w8(32'hbc0dda97),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5adbaa),
	.w1(32'h3b8acec8),
	.w2(32'h3a7f6955),
	.w3(32'hbc091bb4),
	.w4(32'hbb895600),
	.w5(32'hbb21fbe8),
	.w6(32'h3c0e340e),
	.w7(32'h3bb5cc89),
	.w8(32'hbc225921),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b70b9),
	.w1(32'h3c583398),
	.w2(32'h3b09023f),
	.w3(32'hbc17df09),
	.w4(32'h3bc87291),
	.w5(32'hbac7af3d),
	.w6(32'h3c26f4b3),
	.w7(32'h3c051245),
	.w8(32'hbb8712d7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0804fe),
	.w1(32'h3b5d264d),
	.w2(32'hbc20c83e),
	.w3(32'hbc044e26),
	.w4(32'h3c323221),
	.w5(32'h3bf56ac6),
	.w6(32'h3b815ccb),
	.w7(32'h3bdf0336),
	.w8(32'h3b066d44),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2eaf),
	.w1(32'hbb5aac37),
	.w2(32'h3a9d905e),
	.w3(32'h3acac65b),
	.w4(32'h3a9aea61),
	.w5(32'h3b697bd7),
	.w6(32'h39d7b53a),
	.w7(32'h3b15df15),
	.w8(32'hbb98a971),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5f1dc),
	.w1(32'hbc306711),
	.w2(32'hbc88a148),
	.w3(32'hb9edc604),
	.w4(32'hbc34d57c),
	.w5(32'hbca01026),
	.w6(32'hbbb03c91),
	.w7(32'hbc74ecc5),
	.w8(32'h38153119),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ca949),
	.w1(32'h3bf78bf9),
	.w2(32'h3bd3db86),
	.w3(32'hbc71b1a6),
	.w4(32'h3c837fdb),
	.w5(32'h3c2d8715),
	.w6(32'hba754710),
	.w7(32'h38dcf39d),
	.w8(32'hbb3bd618),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba80f93),
	.w1(32'hbc308df2),
	.w2(32'hbc1eca89),
	.w3(32'h3b5cf40e),
	.w4(32'hbba730d0),
	.w5(32'hbc46ee22),
	.w6(32'hbc0a6a80),
	.w7(32'hbbfd33e5),
	.w8(32'hbbdf14ea),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf97bae),
	.w1(32'h3b4de51b),
	.w2(32'hbd0f5590),
	.w3(32'hbbd88fe8),
	.w4(32'hbc462fc7),
	.w5(32'hbcc3cb88),
	.w6(32'h3bd0e454),
	.w7(32'hbc6d1166),
	.w8(32'hbbdcd72d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc767939),
	.w1(32'hbbe3d95c),
	.w2(32'hbbaa7fb0),
	.w3(32'hbc40a374),
	.w4(32'hbb351eb7),
	.w5(32'hbc090eb1),
	.w6(32'hbc141246),
	.w7(32'hbb946733),
	.w8(32'hbc5e04d1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10d5c0),
	.w1(32'h3c12cbea),
	.w2(32'hba9d205f),
	.w3(32'hbc24654b),
	.w4(32'h3b85bcee),
	.w5(32'hbb6b9fec),
	.w6(32'h393feb4b),
	.w7(32'hbb0e796a),
	.w8(32'hbb7cb24a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac50c87),
	.w1(32'hbc0c10e2),
	.w2(32'hbc4eb2b1),
	.w3(32'hbb0d5da2),
	.w4(32'hbba62a63),
	.w5(32'hbbd2e0ec),
	.w6(32'hbb8b0efe),
	.w7(32'hbb747c47),
	.w8(32'h3aabd6ac),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf7fd7),
	.w1(32'hbc4042f6),
	.w2(32'hbc96a728),
	.w3(32'hbb9f0b85),
	.w4(32'hbc0d1f4a),
	.w5(32'hbc04e517),
	.w6(32'h3c5c13ff),
	.w7(32'h3aa71932),
	.w8(32'hbc3b26f5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03ca0c),
	.w1(32'h3c205115),
	.w2(32'hb885da62),
	.w3(32'h3c49d6e8),
	.w4(32'h3ba4ac5a),
	.w5(32'h3bce2148),
	.w6(32'h3b817ff0),
	.w7(32'h3b03965d),
	.w8(32'h3abb7a15),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8872d5),
	.w1(32'h3c774d9d),
	.w2(32'h3c7479ed),
	.w3(32'hbb415c0f),
	.w4(32'h3c5f9d74),
	.w5(32'h3bbc8d24),
	.w6(32'h3be9a6b2),
	.w7(32'h3c0f425e),
	.w8(32'h3b0c989e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8245b1),
	.w1(32'h3c07c0f8),
	.w2(32'h3b730e15),
	.w3(32'hbbb69c73),
	.w4(32'h3c2b15ed),
	.w5(32'h3b30d3a5),
	.w6(32'h3b0e82a3),
	.w7(32'h3bc2efe9),
	.w8(32'h3bba2fa6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b8f88),
	.w1(32'h3bd418c1),
	.w2(32'h3bd1e809),
	.w3(32'hbb8440a9),
	.w4(32'h3bcf2a76),
	.w5(32'h3bb0d871),
	.w6(32'hbbdcdb47),
	.w7(32'h392fa643),
	.w8(32'h3a9d157c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d2bcd),
	.w1(32'hbc2c1f4d),
	.w2(32'hbbf70b61),
	.w3(32'hbb7feb09),
	.w4(32'hbc1318ac),
	.w5(32'hbbb7cc0d),
	.w6(32'hbbc7daf1),
	.w7(32'hbb1c1ae7),
	.w8(32'h39468d31),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae423c0),
	.w1(32'h3951c174),
	.w2(32'hbafa26a2),
	.w3(32'hba9ba8ff),
	.w4(32'hbaba6076),
	.w5(32'hba892ca4),
	.w6(32'h3ab82365),
	.w7(32'h3a60d846),
	.w8(32'hba0013a0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3350c),
	.w1(32'h3c5c9fab),
	.w2(32'hb9d34c84),
	.w3(32'hbb57c340),
	.w4(32'hb9761bb6),
	.w5(32'hbc87d6d5),
	.w6(32'h3ae9e1fd),
	.w7(32'hbbdc790a),
	.w8(32'h3b09683c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7765a),
	.w1(32'hbb0d51a7),
	.w2(32'hbc20aad1),
	.w3(32'hbc576e2a),
	.w4(32'hbba8dc40),
	.w5(32'hbbf56683),
	.w6(32'h3ab59e67),
	.w7(32'hbbf62906),
	.w8(32'hba126c7e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4b2fe),
	.w1(32'hbc7bffdf),
	.w2(32'hbccf21a3),
	.w3(32'hbc22d189),
	.w4(32'hbbde9374),
	.w5(32'hbcd9bda4),
	.w6(32'hbc0fea58),
	.w7(32'hbc8d9b72),
	.w8(32'hbcce30d2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd46662),
	.w1(32'h3a628be2),
	.w2(32'h3ba4f1d0),
	.w3(32'hbc38b223),
	.w4(32'hba765a2c),
	.w5(32'h3b9a8227),
	.w6(32'h3b8f014f),
	.w7(32'h3bf01083),
	.w8(32'hba9aa8a4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a3e75),
	.w1(32'h3c69a27e),
	.w2(32'h3bc37979),
	.w3(32'hbb76b666),
	.w4(32'h3c2c66b7),
	.w5(32'h3c16ea0d),
	.w6(32'h3bd31d6c),
	.w7(32'h3b9c6521),
	.w8(32'hbb393733),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff06f3),
	.w1(32'h3c4b3c6e),
	.w2(32'h3cafc8a3),
	.w3(32'h3affa640),
	.w4(32'h3be37d71),
	.w5(32'h3ca0bb38),
	.w6(32'h3c2338dd),
	.w7(32'h3bc12d8e),
	.w8(32'h3b3100f6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37baea),
	.w1(32'hbcae55cf),
	.w2(32'hbceb6bfd),
	.w3(32'hba324002),
	.w4(32'h3c08f869),
	.w5(32'hbc6ee7a7),
	.w6(32'hbc00ed24),
	.w7(32'hbc2db87c),
	.w8(32'hbc47e758),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceb9be8),
	.w1(32'h3bda46fb),
	.w2(32'h3c4fa42c),
	.w3(32'hbc825522),
	.w4(32'hbb700678),
	.w5(32'hb90ac153),
	.w6(32'hbb656a62),
	.w7(32'h3c2ecb7d),
	.w8(32'h3c14d80c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c458c0c),
	.w1(32'h3c7fa954),
	.w2(32'h3c442db8),
	.w3(32'h3b1990a9),
	.w4(32'h3c785731),
	.w5(32'h3c4cdfc0),
	.w6(32'h3b1faf94),
	.w7(32'h396f9bd9),
	.w8(32'hb9da3cc9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f654),
	.w1(32'h3ba2f713),
	.w2(32'hb9bfef8a),
	.w3(32'h3b1bd777),
	.w4(32'hbbefaa6e),
	.w5(32'hbc5672f7),
	.w6(32'h3c716e8a),
	.w7(32'h3c14dd5a),
	.w8(32'hbbb0dc11),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25a575),
	.w1(32'hbc943cdf),
	.w2(32'hbc7e273e),
	.w3(32'hbac18bb9),
	.w4(32'hbc8a8517),
	.w5(32'hbc7c55da),
	.w6(32'hbc32e777),
	.w7(32'hbc080d2a),
	.w8(32'hbba6dbec),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0e276),
	.w1(32'h3bac8d38),
	.w2(32'hbc82d9d3),
	.w3(32'h3b762545),
	.w4(32'h3b5a0aad),
	.w5(32'hbc579c9f),
	.w6(32'h3ba72a93),
	.w7(32'hbc19fceb),
	.w8(32'hbbbe7306),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f467d),
	.w1(32'h3c2444d5),
	.w2(32'hbc01a018),
	.w3(32'hbc311b8e),
	.w4(32'h3be7bd97),
	.w5(32'h3bbb251e),
	.w6(32'h3c0975ba),
	.w7(32'h3ac6570e),
	.w8(32'h3ac512f6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba87bf6),
	.w1(32'h3c3f97ff),
	.w2(32'h3a24e512),
	.w3(32'hbbbded55),
	.w4(32'h3950ff08),
	.w5(32'hbb69cf71),
	.w6(32'h3b8a5062),
	.w7(32'h3c231c99),
	.w8(32'h3b428d49),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa00ae2),
	.w1(32'hbbe7f3f7),
	.w2(32'hba8cdd46),
	.w3(32'hbb3999a2),
	.w4(32'hb9b138dd),
	.w5(32'h3c2c2741),
	.w6(32'hbb17355b),
	.w7(32'hb9a767bb),
	.w8(32'h3b969d1d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9766),
	.w1(32'hb9dffe9e),
	.w2(32'h3bae265c),
	.w3(32'h3c02130b),
	.w4(32'h39f04147),
	.w5(32'h3bd2cf8b),
	.w6(32'h3ab164db),
	.w7(32'h3b2098d9),
	.w8(32'h3aafbcb1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6728a),
	.w1(32'h3bfeb69f),
	.w2(32'h3b342c9b),
	.w3(32'h3bbbc0d5),
	.w4(32'h3c3335a3),
	.w5(32'h3ba51814),
	.w6(32'h3b1bb28b),
	.w7(32'h3ad1a1fe),
	.w8(32'h3aea08aa),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a52e4f),
	.w1(32'hbabe4a3e),
	.w2(32'hbbcdffb7),
	.w3(32'hbbe70bab),
	.w4(32'hba2ec04f),
	.w5(32'hbc02d7d0),
	.w6(32'h3b2de5dc),
	.w7(32'h3a9863a4),
	.w8(32'h3b4c7f8d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb890bd2),
	.w1(32'hbae7fef2),
	.w2(32'hbb9baad9),
	.w3(32'hbbe14a51),
	.w4(32'h3b914557),
	.w5(32'hb7ebba7e),
	.w6(32'hbaf2eb63),
	.w7(32'hbb67e5a5),
	.w8(32'h3b5b9f52),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb547653),
	.w1(32'hbb915a1f),
	.w2(32'hbc237c82),
	.w3(32'h3c0397d3),
	.w4(32'h3bd1b6f4),
	.w5(32'h39d52a46),
	.w6(32'h3c7e0589),
	.w7(32'h3afe8834),
	.w8(32'hba66c2d2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f73eb9),
	.w1(32'h39dcdba1),
	.w2(32'hbc66e087),
	.w3(32'hba0d9ca4),
	.w4(32'h3bf9c44f),
	.w5(32'hbae63ca8),
	.w6(32'hbaf3d275),
	.w7(32'hbb8a7725),
	.w8(32'h3c03ba32),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e11814),
	.w1(32'h3b71bb92),
	.w2(32'h3c09ab7d),
	.w3(32'hbb32451b),
	.w4(32'h3b31a328),
	.w5(32'h3bd1c0b6),
	.w6(32'h3b830f5b),
	.w7(32'h3ba86159),
	.w8(32'h3b4d864c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa4835),
	.w1(32'hbbb0df59),
	.w2(32'hbc1d2b40),
	.w3(32'h3b4a2792),
	.w4(32'hbb61c5f0),
	.w5(32'hbbc905fc),
	.w6(32'hba83448e),
	.w7(32'hbb251e6b),
	.w8(32'h3c5aeb9c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c96dc),
	.w1(32'hbb340087),
	.w2(32'h389233d6),
	.w3(32'h3ba9c8a8),
	.w4(32'hba292ab4),
	.w5(32'hbaf1777c),
	.w6(32'h3b3f40c7),
	.w7(32'hbb9aff02),
	.w8(32'h3ab9941d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa1d5f),
	.w1(32'h3c4ed3af),
	.w2(32'h3caeb65c),
	.w3(32'h3b24c20a),
	.w4(32'h3c162e0b),
	.w5(32'h3c30d661),
	.w6(32'h3c56ae66),
	.w7(32'h3ca85fe2),
	.w8(32'h3c265635),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f6f62),
	.w1(32'h3bd59564),
	.w2(32'hbc12c2e4),
	.w3(32'h3ad478a6),
	.w4(32'h3b43f3dd),
	.w5(32'hbacfec88),
	.w6(32'h3bf5b29c),
	.w7(32'hbaa5424c),
	.w8(32'hba77cee0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebce8c),
	.w1(32'h3bf8b3e0),
	.w2(32'h3c565abf),
	.w3(32'hba8070d3),
	.w4(32'h3b47ab55),
	.w5(32'h3bcc2160),
	.w6(32'h3b8ac55d),
	.w7(32'h3c1203d2),
	.w8(32'hb9a1cf8c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3814e2f5),
	.w1(32'h3d07a5e6),
	.w2(32'h3cfc5da7),
	.w3(32'h3c1aa6b4),
	.w4(32'h3cbfc2b0),
	.w5(32'h3c62edcc),
	.w6(32'h3ca1f5eb),
	.w7(32'h3c5d475b),
	.w8(32'h3bbbb983),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abd6f4),
	.w1(32'hbb728402),
	.w2(32'hbbbc44c3),
	.w3(32'hbb96f09d),
	.w4(32'hbbf96957),
	.w5(32'hbbcaba2d),
	.w6(32'hbb4da971),
	.w7(32'h39cc1c29),
	.w8(32'hbaa4964f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac90d8),
	.w1(32'hbb36da72),
	.w2(32'hbb48fcc8),
	.w3(32'hbbfe8b06),
	.w4(32'h3ba3da7e),
	.w5(32'hba72c75c),
	.w6(32'h3b90166a),
	.w7(32'hba23ae92),
	.w8(32'hb9ce558c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5491da),
	.w1(32'h3ca389d1),
	.w2(32'h3bd99e8c),
	.w3(32'h3c349715),
	.w4(32'h3c070bdc),
	.w5(32'hbaf043d1),
	.w6(32'h3c12e4c0),
	.w7(32'h3c1f4435),
	.w8(32'h3b8b540c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39415af0),
	.w1(32'h3c6040be),
	.w2(32'h3bf367b3),
	.w3(32'hbb455b35),
	.w4(32'h3c15c901),
	.w5(32'h3c848c24),
	.w6(32'h3c075fd8),
	.w7(32'h3c0a9488),
	.w8(32'h3bf3e562),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c146b3e),
	.w1(32'h3b28da72),
	.w2(32'hbb1bfa82),
	.w3(32'h3c2669b9),
	.w4(32'hb6f45517),
	.w5(32'hba8ab9ba),
	.w6(32'h3a281f2b),
	.w7(32'hbab9d8a0),
	.w8(32'h3a0e7cf7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6880a5),
	.w1(32'h3cf21894),
	.w2(32'hbcc0b49f),
	.w3(32'h3a455569),
	.w4(32'h3cd20433),
	.w5(32'hbc5f6259),
	.w6(32'h3ca7e256),
	.w7(32'hbca9282d),
	.w8(32'hbbe06bce),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule