module layer_8_featuremap_218(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b956937),
	.w1(32'hbbba4ec3),
	.w2(32'hbba7a0bd),
	.w3(32'hbb95fcc9),
	.w4(32'hbc71f557),
	.w5(32'hbc8a92be),
	.w6(32'hbb6a7050),
	.w7(32'hba8259fc),
	.w8(32'hbaa10ef5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec07d5),
	.w1(32'h3e26a455),
	.w2(32'h3ca01c94),
	.w3(32'hba119711),
	.w4(32'h3dd43fd1),
	.w5(32'h3caa8a72),
	.w6(32'h3d934c70),
	.w7(32'hbc6e35d6),
	.w8(32'hbdb60727),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe108179),
	.w1(32'hba9db6c6),
	.w2(32'h3c011781),
	.w3(32'hbdbd2629),
	.w4(32'h3b0ceee6),
	.w5(32'h3c1081b2),
	.w6(32'h3bbbcf41),
	.w7(32'h3b7b52c2),
	.w8(32'h3ba26139),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d7470),
	.w1(32'hbbe437af),
	.w2(32'hba9722d0),
	.w3(32'hbb8c4843),
	.w4(32'hbbbbb1cf),
	.w5(32'hbc0197aa),
	.w6(32'h39718df2),
	.w7(32'hbb1864b7),
	.w8(32'h3b3c178b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0db4fd),
	.w1(32'h3e09f5ac),
	.w2(32'hbbd8033d),
	.w3(32'h3b81b1fa),
	.w4(32'h3d905d67),
	.w5(32'hbbe26cbf),
	.w6(32'h3d488e54),
	.w7(32'hbcbf5bca),
	.w8(32'hbdbf747b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe11ea33),
	.w1(32'h3c3bc2fe),
	.w2(32'hbbc5e46c),
	.w3(32'hbdb6ed71),
	.w4(32'h3b90b62a),
	.w5(32'hbc820741),
	.w6(32'h3c73da3e),
	.w7(32'hba877c58),
	.w8(32'hbc246790),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ba48d),
	.w1(32'hbdb184ce),
	.w2(32'hbba477ff),
	.w3(32'hbc318562),
	.w4(32'hbd70fc67),
	.w5(32'hbbf786d1),
	.w6(32'hbd22633e),
	.w7(32'h3b20a512),
	.w8(32'h3d2d6d3e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d99ef72),
	.w1(32'h3b60bc0f),
	.w2(32'h3c0ae340),
	.w3(32'h3d3fe595),
	.w4(32'h39996d6d),
	.w5(32'h3b58c257),
	.w6(32'hbbeb9624),
	.w7(32'hbb6ad7f2),
	.w8(32'hbc07a47a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9ee88),
	.w1(32'h3df36328),
	.w2(32'h3c01b618),
	.w3(32'hbb3e7057),
	.w4(32'h3d676a35),
	.w5(32'hb9169815),
	.w6(32'h3d26ee2c),
	.w7(32'hbc72b0f2),
	.w8(32'hbd909648),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbddfbadf),
	.w1(32'hbc4363f8),
	.w2(32'h3c08dddf),
	.w3(32'hbd8548d6),
	.w4(32'hbc4244be),
	.w5(32'h3b5f3d7b),
	.w6(32'h38e340ed),
	.w7(32'hba8cb2ea),
	.w8(32'h3b6b239a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace6a31),
	.w1(32'h3b9c33b7),
	.w2(32'hbbba7bac),
	.w3(32'h3b5d7455),
	.w4(32'hbc486bb0),
	.w5(32'hbaee87e0),
	.w6(32'h3b5ff6a1),
	.w7(32'hbc264c9a),
	.w8(32'hbbe4b2d2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccef10),
	.w1(32'hbb949c5e),
	.w2(32'hbc25c48b),
	.w3(32'hbbfcc8a7),
	.w4(32'hbb5185ad),
	.w5(32'hbc2a6da0),
	.w6(32'h3b417c31),
	.w7(32'hbb2d9aa2),
	.w8(32'hbc0946db),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eaa14),
	.w1(32'hbaf2c8eb),
	.w2(32'hbac82f2d),
	.w3(32'h38c0c146),
	.w4(32'h3b575eab),
	.w5(32'hbb6cebfd),
	.w6(32'hbbdd99eb),
	.w7(32'hbb9c2dfb),
	.w8(32'h3b083458),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae74def),
	.w1(32'hbb668269),
	.w2(32'hbbcc03d3),
	.w3(32'hb9aa7d89),
	.w4(32'hbb3c6011),
	.w5(32'hbc01e0fa),
	.w6(32'h3b4b9856),
	.w7(32'hba85ee35),
	.w8(32'h3ab45cb0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4dfbd),
	.w1(32'hbe0ebdd8),
	.w2(32'hbbc3027f),
	.w3(32'hbbf6730a),
	.w4(32'hbd9c083a),
	.w5(32'hbc163933),
	.w6(32'hbd8e355d),
	.w7(32'h3aa31b59),
	.w8(32'h3d8c71d3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3df71311),
	.w1(32'h3b61426b),
	.w2(32'hbb92f787),
	.w3(32'h3d9c88c0),
	.w4(32'hbb3e73cb),
	.w5(32'h3abb5de3),
	.w6(32'h3c0a2f02),
	.w7(32'h385ce2f5),
	.w8(32'hb951ab2b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee2b4),
	.w1(32'hbaa29a51),
	.w2(32'hbb3b9afa),
	.w3(32'h3bf3a48a),
	.w4(32'h3bddc49d),
	.w5(32'hb8a8a094),
	.w6(32'h3b8f11f3),
	.w7(32'hbc07e7c3),
	.w8(32'hbbd2efb4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc991e6f),
	.w1(32'hbc0fb5c7),
	.w2(32'h3b80cc48),
	.w3(32'hbbc760d6),
	.w4(32'hbb83b542),
	.w5(32'hbc2a3b83),
	.w6(32'hbbbef609),
	.w7(32'h3b485ab5),
	.w8(32'h3be03c86),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be233fb),
	.w1(32'hbc9f897d),
	.w2(32'hbccc412a),
	.w3(32'hbc59bbe8),
	.w4(32'hbd49385d),
	.w5(32'hbd346963),
	.w6(32'hbaffa24f),
	.w7(32'hbc4c028b),
	.w8(32'h3a11097a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eae95),
	.w1(32'hbe39307f),
	.w2(32'hbc9eeb9a),
	.w3(32'h3b228478),
	.w4(32'hbde6f818),
	.w5(32'hbcd451e4),
	.w6(32'hbda04359),
	.w7(32'h3c513962),
	.w8(32'h3db6ed05),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e263799),
	.w1(32'hba4b3249),
	.w2(32'hbbedf6e2),
	.w3(32'h3de16614),
	.w4(32'hbb192002),
	.w5(32'hbc2db5ca),
	.w6(32'h3c0f6a31),
	.w7(32'h3b2b2b6b),
	.w8(32'hbbc5562b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc057bc5),
	.w1(32'hba97c96b),
	.w2(32'h3c218ce1),
	.w3(32'hbada6027),
	.w4(32'h3bbee3ef),
	.w5(32'h3c205659),
	.w6(32'h3b1c6094),
	.w7(32'hb9407c35),
	.w8(32'h3c079b51),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33de40),
	.w1(32'h3ba2cf69),
	.w2(32'h3c9a7a8e),
	.w3(32'hbaabf45c),
	.w4(32'hbcafaa4d),
	.w5(32'hb9becc2b),
	.w6(32'hbbffa151),
	.w7(32'hbc7cb381),
	.w8(32'hbb0a8931),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88a552),
	.w1(32'h3bf664d3),
	.w2(32'h3b3c0ac2),
	.w3(32'h38f77ebe),
	.w4(32'h3c088401),
	.w5(32'hbad1edc5),
	.w6(32'hb7fd928d),
	.w7(32'hbb0dd409),
	.w8(32'hbc3b3f75),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd42998),
	.w1(32'h3ba56a6f),
	.w2(32'h3c12c96a),
	.w3(32'hbba8006f),
	.w4(32'h39bfa09d),
	.w5(32'h3b32b086),
	.w6(32'hbb27a892),
	.w7(32'h3c24d62b),
	.w8(32'h3ba8e891),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ea4cd),
	.w1(32'h3bdc687e),
	.w2(32'h3bc41118),
	.w3(32'hbc4525d3),
	.w4(32'hbc28b9e0),
	.w5(32'hbc59b3ee),
	.w6(32'hbb2e168a),
	.w7(32'hbbb55b4a),
	.w8(32'hbc12f277),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e414f1),
	.w1(32'hbb88219d),
	.w2(32'h3b33be01),
	.w3(32'hba2b87f9),
	.w4(32'hbc0bd1da),
	.w5(32'hbb794afb),
	.w6(32'h3b219a0f),
	.w7(32'h3b7d73bc),
	.w8(32'h3b846190),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e2684),
	.w1(32'hbcd728d5),
	.w2(32'hbbf384fb),
	.w3(32'hbd16c67e),
	.w4(32'hbd5a7397),
	.w5(32'hbdcedfdc),
	.w6(32'hbd2ffc7b),
	.w7(32'hbdc56d2a),
	.w8(32'hbd05d592),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92171f),
	.w1(32'h3b51ace0),
	.w2(32'hbcd64143),
	.w3(32'hbc6d5523),
	.w4(32'hbba93202),
	.w5(32'hbcb54f39),
	.w6(32'h3c1e3477),
	.w7(32'hbc72f275),
	.w8(32'hbc5ebff0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcef6812),
	.w1(32'h3b531164),
	.w2(32'hbb53164d),
	.w3(32'hbc7c844b),
	.w4(32'hbbe8c56a),
	.w5(32'hbc4fa2d0),
	.w6(32'h3b0df29d),
	.w7(32'hbb60f0fa),
	.w8(32'h3c53029c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c312586),
	.w1(32'h3bfd51fe),
	.w2(32'h3bc1d7f2),
	.w3(32'h3beff051),
	.w4(32'hbb88f916),
	.w5(32'hb7a41ac4),
	.w6(32'h3c1a70f8),
	.w7(32'h3c2a5b7b),
	.w8(32'h3b024490),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2217a6),
	.w1(32'h3c5a6816),
	.w2(32'hbbacb9ff),
	.w3(32'hbace1ddd),
	.w4(32'h3c2147d3),
	.w5(32'hba86cb34),
	.w6(32'h3c601403),
	.w7(32'hbbe17cf5),
	.w8(32'hbb90d897),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e87d8),
	.w1(32'h3b87a5d5),
	.w2(32'h3c490134),
	.w3(32'h399b298b),
	.w4(32'hbbcdbb98),
	.w5(32'h3a97a568),
	.w6(32'h3b868148),
	.w7(32'h3b452586),
	.w8(32'h3a87a49d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b13ca),
	.w1(32'h3b797fee),
	.w2(32'hba7e4431),
	.w3(32'h3ba7be5c),
	.w4(32'h3b07c559),
	.w5(32'h3b81d97a),
	.w6(32'h3b989cc0),
	.w7(32'hba59f577),
	.w8(32'hb7a37a38),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b3f27),
	.w1(32'hbb8e5c59),
	.w2(32'hba57376a),
	.w3(32'h3b786fdd),
	.w4(32'h3c6ced77),
	.w5(32'h3c497621),
	.w6(32'h3bc496b7),
	.w7(32'h3c505774),
	.w8(32'h3c9e3cb7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba295f),
	.w1(32'hbbdca537),
	.w2(32'hba0a5318),
	.w3(32'hbbeafaa7),
	.w4(32'hbc860683),
	.w5(32'hbc5af297),
	.w6(32'hbc1c2842),
	.w7(32'hbbca48d2),
	.w8(32'hbb7d986b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfd4bb),
	.w1(32'hbb29768d),
	.w2(32'hbc12105e),
	.w3(32'h3b791e5a),
	.w4(32'hba7bb56d),
	.w5(32'hbc27548f),
	.w6(32'h3a0c40b5),
	.w7(32'hbb0cfa2b),
	.w8(32'h3ba0412d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8caba),
	.w1(32'h3cf58c71),
	.w2(32'h3c0fd1e4),
	.w3(32'hbb58577e),
	.w4(32'h3cda728e),
	.w5(32'h3c0355c5),
	.w6(32'h3c0f688f),
	.w7(32'hbc049261),
	.w8(32'hbcab7db0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd037876),
	.w1(32'hbb5adcc6),
	.w2(32'h3a979c46),
	.w3(32'hbc8ed341),
	.w4(32'hbb19de0d),
	.w5(32'hba974a8d),
	.w6(32'h3882caa5),
	.w7(32'hbabe1579),
	.w8(32'h3ab050aa),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ca711),
	.w1(32'h3b377bcc),
	.w2(32'h3a8af528),
	.w3(32'h3ac0719c),
	.w4(32'h3b04680e),
	.w5(32'h3b6d9297),
	.w6(32'h3badb594),
	.w7(32'hb78e404f),
	.w8(32'h3bb30213),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac853e3),
	.w1(32'hbc0b04f9),
	.w2(32'hbc313760),
	.w3(32'hbca9a3e1),
	.w4(32'hbcb1dfab),
	.w5(32'hbcbbc725),
	.w6(32'hbca0acdc),
	.w7(32'hbc3ea7d2),
	.w8(32'hbc4d4357),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b066a30),
	.w1(32'h3bc060ff),
	.w2(32'hbbde0af2),
	.w3(32'hbab18701),
	.w4(32'h3a484ccd),
	.w5(32'hbb67196d),
	.w6(32'h3c222bed),
	.w7(32'hbb8ed3ea),
	.w8(32'h393398c0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0efd7),
	.w1(32'hbb497961),
	.w2(32'hbc6534df),
	.w3(32'hbb739019),
	.w4(32'hbba9e261),
	.w5(32'hbc5e2d3d),
	.w6(32'h3b077a01),
	.w7(32'hbb456109),
	.w8(32'h3a41851b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab27252),
	.w1(32'hbbbeb8c8),
	.w2(32'hbbed5680),
	.w3(32'hbbf8e4b7),
	.w4(32'hbc9b8c3d),
	.w5(32'hbc641238),
	.w6(32'hbc219972),
	.w7(32'hbc8921ed),
	.w8(32'hbb13f9e2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07a261),
	.w1(32'h3a6ab288),
	.w2(32'hbab078e1),
	.w3(32'h3aa8fb60),
	.w4(32'hbc234718),
	.w5(32'hbbb1e4f8),
	.w6(32'h3bb24b24),
	.w7(32'h3af23916),
	.w8(32'hba0c4229),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2826f5),
	.w1(32'hbde91f2e),
	.w2(32'hbbd7187a),
	.w3(32'h390bd660),
	.w4(32'hbdb4af94),
	.w5(32'hbc8fe7e8),
	.w6(32'hbd6a88d9),
	.w7(32'h3a9f865b),
	.w8(32'h3d78a70c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3de1af87),
	.w1(32'hbb843e22),
	.w2(32'hbb8c87a4),
	.w3(32'h3d86c47d),
	.w4(32'hba2a90d5),
	.w5(32'h3ac5ac2f),
	.w6(32'hbad56c9a),
	.w7(32'hbbaba4cb),
	.w8(32'hbb9127a6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc79194),
	.w1(32'h3b15c256),
	.w2(32'hbc1272fe),
	.w3(32'h3bda933e),
	.w4(32'hbcb22346),
	.w5(32'hbc9fcace),
	.w6(32'h3bf7caff),
	.w7(32'h3a92b945),
	.w8(32'h3b864396),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af95809),
	.w1(32'hbafd1491),
	.w2(32'hba6270ed),
	.w3(32'hbbb2b4b0),
	.w4(32'hbb01af65),
	.w5(32'hbb51eedd),
	.w6(32'h3b4e66f1),
	.w7(32'h3bb36390),
	.w8(32'hbb4bc21c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0952fd),
	.w1(32'hbc18ca07),
	.w2(32'hbc6124d3),
	.w3(32'hbb4f3fbd),
	.w4(32'hbc0c1efe),
	.w5(32'hbc9023eb),
	.w6(32'hbbbad161),
	.w7(32'hbb1ab031),
	.w8(32'hba8fab0a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23f8ee),
	.w1(32'h3c9b8606),
	.w2(32'h3c7455ce),
	.w3(32'h3ac0d71b),
	.w4(32'h3c5d55f9),
	.w5(32'h3c51e2f2),
	.w6(32'h3c384572),
	.w7(32'h3bf54b9d),
	.w8(32'h38fb5a5b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1318c),
	.w1(32'h3cb120dd),
	.w2(32'hb902ca05),
	.w3(32'hbbcc13cb),
	.w4(32'hbc3dcba0),
	.w5(32'hbc038e1b),
	.w6(32'h3ab9019c),
	.w7(32'hbc7a429c),
	.w8(32'hbbf3889f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbea62a),
	.w1(32'h3dd0f416),
	.w2(32'h3bc75448),
	.w3(32'h392ac353),
	.w4(32'h3d5dc0c3),
	.w5(32'hbab5ea74),
	.w6(32'h3d1ccb80),
	.w7(32'hbc52dfa4),
	.w8(32'hbd743b99),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdc3e993),
	.w1(32'hbbda160a),
	.w2(32'hbc5020c6),
	.w3(32'hbd816282),
	.w4(32'hbc27bac0),
	.w5(32'hbb755e3c),
	.w6(32'h3b8254d4),
	.w7(32'h3aea322b),
	.w8(32'h3ba49a4b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b236917),
	.w1(32'h3bfda9ef),
	.w2(32'h3c0143d5),
	.w3(32'h39000074),
	.w4(32'h3b8988df),
	.w5(32'h3c04c2b3),
	.w6(32'h3b9d2f4d),
	.w7(32'h3baaaa06),
	.w8(32'h3acd752d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1e16),
	.w1(32'hbcbef036),
	.w2(32'hbc7442ed),
	.w3(32'hba801fc6),
	.w4(32'hbca58581),
	.w5(32'hbcc01007),
	.w6(32'hbb5e5ae5),
	.w7(32'hbbe0bf1c),
	.w8(32'h3b10844e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a5b6d),
	.w1(32'h3a1adecb),
	.w2(32'hbc2e2194),
	.w3(32'h3b516a5f),
	.w4(32'h3ba66f87),
	.w5(32'h3abd08c3),
	.w6(32'h3c19d154),
	.w7(32'h3b103d9a),
	.w8(32'hba893c8b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e5979),
	.w1(32'hbc106df1),
	.w2(32'hbcba5be3),
	.w3(32'hbc24616c),
	.w4(32'hbc9e62a9),
	.w5(32'hbccfcfed),
	.w6(32'hbc8f41cc),
	.w7(32'hbcdb51e5),
	.w8(32'hbbf179f6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6e402),
	.w1(32'hbb2ea553),
	.w2(32'hbad7e898),
	.w3(32'hbb5d102f),
	.w4(32'hbbed12a3),
	.w5(32'hbbb6e435),
	.w6(32'h3a840081),
	.w7(32'hbc15a2b2),
	.w8(32'hbc77ce2c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28988c),
	.w1(32'hbb02e787),
	.w2(32'h3bc1cbfd),
	.w3(32'h3b95b167),
	.w4(32'hbc0813ba),
	.w5(32'hbb1b511c),
	.w6(32'h3ba2fdde),
	.w7(32'hbb6c37fc),
	.w8(32'hbb0ec980),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b645aa9),
	.w1(32'hb97de081),
	.w2(32'h3ba4d711),
	.w3(32'hbad9d26f),
	.w4(32'hbc29b5bf),
	.w5(32'h3aca647b),
	.w6(32'h3b075227),
	.w7(32'hbac5bbf9),
	.w8(32'hbc05b7cb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2ccda),
	.w1(32'hb9c8050f),
	.w2(32'hbba33b8e),
	.w3(32'h3bb170ed),
	.w4(32'h3bab550a),
	.w5(32'hbc170631),
	.w6(32'h3ab4ceae),
	.w7(32'h3b1ce36e),
	.w8(32'h3b923edd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad263a9),
	.w1(32'hb9a37ee5),
	.w2(32'h38c11587),
	.w3(32'hbcada802),
	.w4(32'hbc807619),
	.w5(32'hbc1e90c4),
	.w6(32'h3bf47da5),
	.w7(32'hbad798b1),
	.w8(32'h3b848cdf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45d547),
	.w1(32'h3b96f73c),
	.w2(32'h3bd12e5f),
	.w3(32'h3c57b1a7),
	.w4(32'h3b8d68e6),
	.w5(32'h3b8bf617),
	.w6(32'h3a886b9f),
	.w7(32'h3a56982f),
	.w8(32'h3abfee15),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1d012),
	.w1(32'hbc8c4674),
	.w2(32'hbc162366),
	.w3(32'h3b8c082e),
	.w4(32'hba843c87),
	.w5(32'hbbf191ad),
	.w6(32'hbbc7f301),
	.w7(32'hbc120dc8),
	.w8(32'hbc380b10),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd48a9c),
	.w1(32'h38e1f20d),
	.w2(32'h3b122db4),
	.w3(32'hbc33348f),
	.w4(32'hbbdb931b),
	.w5(32'hbc0be752),
	.w6(32'hbb62ca1e),
	.w7(32'hbb813bee),
	.w8(32'h3986d500),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b953689),
	.w1(32'h3b7fb25e),
	.w2(32'h3b53195e),
	.w3(32'h3b9d6ca6),
	.w4(32'h3a126b1e),
	.w5(32'h3b112ec2),
	.w6(32'h3b4d88a9),
	.w7(32'h3b3ebd8f),
	.w8(32'hbb14f5a0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53a081),
	.w1(32'hbb5d3804),
	.w2(32'hbbb9f08d),
	.w3(32'h3be3413b),
	.w4(32'hbb1d028e),
	.w5(32'hbb684eb7),
	.w6(32'h3a98c199),
	.w7(32'hbae2360a),
	.w8(32'h3add0433),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baef082),
	.w1(32'h3b84a30e),
	.w2(32'hba7e9a80),
	.w3(32'h3b0367ae),
	.w4(32'hbaca8f91),
	.w5(32'h378e75ab),
	.w6(32'hba65c168),
	.w7(32'h3ae47c12),
	.w8(32'hbaf14e3b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6b0cc),
	.w1(32'h3c18a559),
	.w2(32'hbc32c6c6),
	.w3(32'h3b1e4d83),
	.w4(32'hbcb61b66),
	.w5(32'hbd023ca6),
	.w6(32'hbbf589b9),
	.w7(32'hbcde24c1),
	.w8(32'hbc88d919),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc44e62),
	.w1(32'h3cbeed61),
	.w2(32'h3cd47f99),
	.w3(32'hbb04a4dc),
	.w4(32'h3ca22efd),
	.w5(32'h3cd64e44),
	.w6(32'h3c188dbb),
	.w7(32'h3c334e69),
	.w8(32'h3b86ea38),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda5931),
	.w1(32'h3a23aa03),
	.w2(32'hb98f90c8),
	.w3(32'h3bb942e7),
	.w4(32'hbc000edc),
	.w5(32'hbbb9f178),
	.w6(32'hbb25ad8e),
	.w7(32'hbab65708),
	.w8(32'hbbf37fe1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab8c26),
	.w1(32'hbac547fc),
	.w2(32'hba85e485),
	.w3(32'h3b5c4432),
	.w4(32'hbb4ffb5e),
	.w5(32'hbb95e313),
	.w6(32'h3bbc837c),
	.w7(32'h3b9cb0f4),
	.w8(32'h3b9b9476),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b0811),
	.w1(32'hbc1a17f8),
	.w2(32'hbb9aa3c4),
	.w3(32'hbbb263f2),
	.w4(32'hbbb88cc1),
	.w5(32'hbc023b36),
	.w6(32'hba90274d),
	.w7(32'hbbe18ccb),
	.w8(32'h3b11da24),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b345cce),
	.w1(32'h3be0182e),
	.w2(32'h3b8e1f54),
	.w3(32'h3b0f2f7e),
	.w4(32'h3b9e7950),
	.w5(32'h3b80a55b),
	.w6(32'h3c3c0e3b),
	.w7(32'h3b4013e8),
	.w8(32'h3b5edade),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78d7a8),
	.w1(32'hbc0e2562),
	.w2(32'hbbfbc162),
	.w3(32'h3b71a7cf),
	.w4(32'hbc8414d6),
	.w5(32'hbba924e3),
	.w6(32'hbbbffcf8),
	.w7(32'hbc8e3ab3),
	.w8(32'hbc23809e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f1781),
	.w1(32'hbbb1de0b),
	.w2(32'hbc8462bb),
	.w3(32'hbb6fe132),
	.w4(32'hbc059eba),
	.w5(32'hbb98e9d2),
	.w6(32'h3b484b02),
	.w7(32'hbbce71ab),
	.w8(32'h3c1b2370),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16a7e4),
	.w1(32'hbc488052),
	.w2(32'hbcdaf928),
	.w3(32'hba6e7a72),
	.w4(32'hbcbc68e6),
	.w5(32'hbd157788),
	.w6(32'hbc83005f),
	.w7(32'hbce8f61e),
	.w8(32'h3af0311b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a862),
	.w1(32'hbb2325ac),
	.w2(32'h3b187ffc),
	.w3(32'hbb50159d),
	.w4(32'h391b61c6),
	.w5(32'h3bc7bf04),
	.w6(32'h3a9bba0e),
	.w7(32'hbad407b9),
	.w8(32'h3b8f788f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85edb3),
	.w1(32'h3b1882bb),
	.w2(32'h3b266b09),
	.w3(32'hb9772580),
	.w4(32'h38759277),
	.w5(32'hbaf8f342),
	.w6(32'hbb3aec70),
	.w7(32'hbb577f99),
	.w8(32'h39a785f7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb840fa58),
	.w1(32'h3b598c54),
	.w2(32'hba530b73),
	.w3(32'h3a4dc737),
	.w4(32'h3b1b8f7a),
	.w5(32'h397d79ac),
	.w6(32'h3bf57bd6),
	.w7(32'h3b84d69d),
	.w8(32'h3b253bc7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3b3bd),
	.w1(32'h3b84d36a),
	.w2(32'hbbb82c5a),
	.w3(32'h3a87bb38),
	.w4(32'hbab61b1e),
	.w5(32'hbc20f4e2),
	.w6(32'hbb9953d8),
	.w7(32'hbc2479e0),
	.w8(32'hbbf3fa86),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854751),
	.w1(32'h3bc9e46a),
	.w2(32'h3a31236d),
	.w3(32'hbbbd54f6),
	.w4(32'hbc38941a),
	.w5(32'hbc3b5add),
	.w6(32'hba4cd18d),
	.w7(32'hbbdefb86),
	.w8(32'hbc6a5475),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c3e24),
	.w1(32'hba7e983e),
	.w2(32'hbc3450d1),
	.w3(32'hbd0da311),
	.w4(32'hbc76c763),
	.w5(32'hbc8638e7),
	.w6(32'hbbc8d80d),
	.w7(32'h3bacd083),
	.w8(32'hbb26f82a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d2c3f),
	.w1(32'hbb8e8dde),
	.w2(32'hbbbcf9ce),
	.w3(32'hbcb6ed26),
	.w4(32'hbcff6c71),
	.w5(32'hbccba9ff),
	.w6(32'hbc588e39),
	.w7(32'hbc6d1136),
	.w8(32'hbc24c349),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d958e),
	.w1(32'h3c43dacf),
	.w2(32'hbb352703),
	.w3(32'h3b10be58),
	.w4(32'hbc167861),
	.w5(32'hbc41c58a),
	.w6(32'h3c11cf1c),
	.w7(32'hbc1648c5),
	.w8(32'hbc850829),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46bc59),
	.w1(32'h3c25879b),
	.w2(32'h3bb41a64),
	.w3(32'h3adee9fb),
	.w4(32'h3b5b0b3b),
	.w5(32'hba9dcd23),
	.w6(32'h3b49a965),
	.w7(32'hbb60518f),
	.w8(32'hbbc637fd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95429a),
	.w1(32'h3c92ac6e),
	.w2(32'hba49cae5),
	.w3(32'hba8dbade),
	.w4(32'h3cb717c8),
	.w5(32'h3bc59778),
	.w6(32'h3a6b350a),
	.w7(32'hbb3fcc98),
	.w8(32'h37bd9499),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbee12e),
	.w1(32'hba5dd33e),
	.w2(32'h3ae8f2ac),
	.w3(32'hbba83a92),
	.w4(32'h3b30b477),
	.w5(32'h3b3710d8),
	.w6(32'h3c078374),
	.w7(32'h3ad394f2),
	.w8(32'hbb808864),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9edaa),
	.w1(32'h3b8cda6a),
	.w2(32'h3be52935),
	.w3(32'h3b306cbd),
	.w4(32'h3a5cb3ac),
	.w5(32'h38e0bef4),
	.w6(32'h3b80772e),
	.w7(32'h3baeafdf),
	.w8(32'hbbb3b83c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b290b14),
	.w1(32'hbac48ccd),
	.w2(32'hbb463cda),
	.w3(32'h3baf8893),
	.w4(32'h3a5f2ab4),
	.w5(32'hba85441b),
	.w6(32'h3b30856f),
	.w7(32'h3ab8f766),
	.w8(32'hbb47bc72),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b748c9b),
	.w1(32'h3bbfc952),
	.w2(32'hbb439fd3),
	.w3(32'h3bbd6387),
	.w4(32'h3b7e29e4),
	.w5(32'h3b79764e),
	.w6(32'h3b8925e1),
	.w7(32'hbb18d0b5),
	.w8(32'h36fb1873),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45456b),
	.w1(32'h3d1b9a99),
	.w2(32'h3b9e045a),
	.w3(32'h3b866297),
	.w4(32'h3cc7b491),
	.w5(32'h3bd83d68),
	.w6(32'h3c881f48),
	.w7(32'hba049e14),
	.w8(32'hbc8b5e92),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc900839),
	.w1(32'h3d97dd0d),
	.w2(32'h3ba007dc),
	.w3(32'hbc70d3a0),
	.w4(32'h3d274496),
	.w5(32'h3b901d79),
	.w6(32'h3d0f6007),
	.w7(32'hbb79cb0c),
	.w8(32'hbd147512),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd717a1c),
	.w1(32'hbb9c4a80),
	.w2(32'hbc9e410d),
	.w3(32'hbd0abbf9),
	.w4(32'h3ac5fd3e),
	.w5(32'hbbadbab6),
	.w6(32'h3c0f6da9),
	.w7(32'h3b811a19),
	.w8(32'hb9881d54),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1e000),
	.w1(32'hbaee3dd6),
	.w2(32'hbc77b8ff),
	.w3(32'hbb057b1f),
	.w4(32'hbc4a70dc),
	.w5(32'hbc8c13ff),
	.w6(32'h3b878c27),
	.w7(32'hbc143b88),
	.w8(32'hbb9a5b89),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983db5),
	.w1(32'h3b05dcc0),
	.w2(32'h3b769857),
	.w3(32'hbbd73e43),
	.w4(32'hbc38a8e2),
	.w5(32'hbc49ef4e),
	.w6(32'h3bbcb560),
	.w7(32'hbb3d5f47),
	.w8(32'hbb926acc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4075),
	.w1(32'hbb0557fd),
	.w2(32'h3908065b),
	.w3(32'hbbc7eab9),
	.w4(32'hba5146ae),
	.w5(32'hbb2a739f),
	.w6(32'hba34f9a8),
	.w7(32'hbbc7ada7),
	.w8(32'h3b41e592),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad88b19),
	.w1(32'hbc033a9a),
	.w2(32'hbb0cf6fa),
	.w3(32'hbb0750c8),
	.w4(32'hbbf5922e),
	.w5(32'hbc454d09),
	.w6(32'hbb6fe441),
	.w7(32'hbb1b1aeb),
	.w8(32'h3bac75d9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b825ce7),
	.w1(32'hbb1aea37),
	.w2(32'h3a7ad87f),
	.w3(32'hbbd70cb5),
	.w4(32'hbbf00b4e),
	.w5(32'h3b05c79c),
	.w6(32'hbab3663d),
	.w7(32'h3b8a8a13),
	.w8(32'hb9b6d396),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a2899),
	.w1(32'h3b8c2bc7),
	.w2(32'h3ba0658e),
	.w3(32'h3b3088d5),
	.w4(32'h3b8389e3),
	.w5(32'hbae24e2b),
	.w6(32'h3a0a714d),
	.w7(32'h3b4fd0ea),
	.w8(32'hbb301980),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8f648),
	.w1(32'h3aba969d),
	.w2(32'h3a948b36),
	.w3(32'hbb8eb407),
	.w4(32'hbb8a01bb),
	.w5(32'h3af07669),
	.w6(32'h3b466a81),
	.w7(32'hbba95f3d),
	.w8(32'hbb9bcdb2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb943a12),
	.w1(32'hb9eb08f2),
	.w2(32'hbbc105a9),
	.w3(32'hbad03f47),
	.w4(32'hbb87d4e5),
	.w5(32'hbbc563b3),
	.w6(32'h3a326959),
	.w7(32'h3adc01ad),
	.w8(32'hbb524ae8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc280fb5),
	.w1(32'hba38386b),
	.w2(32'hbc1881fd),
	.w3(32'h3a409e9d),
	.w4(32'hbbe48379),
	.w5(32'h3ac90f5c),
	.w6(32'h3b44159b),
	.w7(32'hba916d17),
	.w8(32'hbbb11447),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf809f),
	.w1(32'hbac041a0),
	.w2(32'hb8d650da),
	.w3(32'h39bc1a8b),
	.w4(32'hbb22d943),
	.w5(32'h3ab2060a),
	.w6(32'hbac9e811),
	.w7(32'hba954aa2),
	.w8(32'hbbbc2932),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95be885),
	.w1(32'hbdb37337),
	.w2(32'hbb1f16fa),
	.w3(32'hbb0f46b0),
	.w4(32'hbd6d7630),
	.w5(32'hbcd188b6),
	.w6(32'hbd46d3e5),
	.w7(32'hbc2d8fa9),
	.w8(32'h3cf507f1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dafefcf),
	.w1(32'hbb24a2a1),
	.w2(32'hbb94678e),
	.w3(32'h3d357aaa),
	.w4(32'hbc0588bf),
	.w5(32'hbb8ae602),
	.w6(32'hbbbf56ef),
	.w7(32'hbc4a1566),
	.w8(32'hbc65cf11),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c2fab),
	.w1(32'hbbb770e0),
	.w2(32'hbc11b15e),
	.w3(32'h3bf795e1),
	.w4(32'h3bcd8b83),
	.w5(32'hbba3eb05),
	.w6(32'hbb85dabc),
	.w7(32'hbabcd18a),
	.w8(32'h3afb50f3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1feb7),
	.w1(32'h3bea8bbc),
	.w2(32'h3b033587),
	.w3(32'h3bb5bff0),
	.w4(32'h3c592fea),
	.w5(32'h3ae1009a),
	.w6(32'h3b5fb73c),
	.w7(32'hbb627dc7),
	.w8(32'hbabe4be8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70ec24),
	.w1(32'h3dd9b9c5),
	.w2(32'h3c73c569),
	.w3(32'hbc2d2c60),
	.w4(32'h3d833797),
	.w5(32'h3c72851f),
	.w6(32'h3d515805),
	.w7(32'hbc493712),
	.w8(32'hbd804bae),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdba3dfc),
	.w1(32'h39594c7f),
	.w2(32'hb922bfa5),
	.w3(32'hbd753995),
	.w4(32'hbb84e29e),
	.w5(32'hbc058cef),
	.w6(32'h3be5a37a),
	.w7(32'h3ba09588),
	.w8(32'hbaf5c4eb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba380531),
	.w1(32'hbd171f41),
	.w2(32'hbc30c5a0),
	.w3(32'hbae4025f),
	.w4(32'hbcc8eda7),
	.w5(32'hbc4d4280),
	.w6(32'hbc9c120f),
	.w7(32'hb8450855),
	.w8(32'h3ca31ebd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf50175),
	.w1(32'h3b2c0744),
	.w2(32'hbb4f3f5d),
	.w3(32'h3c9afab7),
	.w4(32'h3be51b7d),
	.w5(32'hbb44b496),
	.w6(32'hba040c0e),
	.w7(32'h3b8edf7a),
	.w8(32'h3b383f93),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33b5aa),
	.w1(32'hbad4f306),
	.w2(32'h3b7624c1),
	.w3(32'hbc2aa7b9),
	.w4(32'hbabd9331),
	.w5(32'hbb48c5a3),
	.w6(32'hbac1753f),
	.w7(32'h39d99b77),
	.w8(32'h3b6a7ef9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392990),
	.w1(32'h3bd3890e),
	.w2(32'h3c496476),
	.w3(32'hbb24b3ce),
	.w4(32'h3c14e3bb),
	.w5(32'h3c158d42),
	.w6(32'h3ba941b5),
	.w7(32'h3ba2b4a2),
	.w8(32'hb98147f1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c149190),
	.w1(32'h3d922c59),
	.w2(32'h3bf55f72),
	.w3(32'h3c4256fd),
	.w4(32'h3d517a77),
	.w5(32'h3c19d768),
	.w6(32'h3d10b63f),
	.w7(32'hbbd5579b),
	.w8(32'hbd309e0b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8219aa),
	.w1(32'h3b64060c),
	.w2(32'hbb202a0e),
	.w3(32'hbd1ed2fa),
	.w4(32'hbb8f4321),
	.w5(32'hbc158520),
	.w6(32'h3c04a80a),
	.w7(32'hbad6b501),
	.w8(32'h3bb3b51b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c046887),
	.w1(32'hb9ec8482),
	.w2(32'hbc1d77e2),
	.w3(32'hbacf3c2c),
	.w4(32'hbc558038),
	.w5(32'hbc8a76b9),
	.w6(32'hbba9c300),
	.w7(32'hbb95e7eb),
	.w8(32'hbc347a17),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc297c15),
	.w1(32'hbb2af7b3),
	.w2(32'hbbb3d795),
	.w3(32'hbc16b8ba),
	.w4(32'hbbba9c7d),
	.w5(32'hbb88ee6c),
	.w6(32'hbaea0d75),
	.w7(32'h3afc52a3),
	.w8(32'h3a81c1ee),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1887d2),
	.w1(32'h3b4fa1c1),
	.w2(32'h3b2aec61),
	.w3(32'hbc094b8d),
	.w4(32'hb994e2f6),
	.w5(32'h3b682417),
	.w6(32'h3c0157a6),
	.w7(32'h3b0a4d5a),
	.w8(32'h39132355),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d79ad),
	.w1(32'hbb1abb4a),
	.w2(32'hbb53fde5),
	.w3(32'h3bb69dac),
	.w4(32'h3acfa625),
	.w5(32'h3c10db71),
	.w6(32'h3ba1bf6b),
	.w7(32'hbbc8eaeb),
	.w8(32'hbb48a6be),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91cd3ab),
	.w1(32'hbb6b2470),
	.w2(32'hbb17dc7c),
	.w3(32'hbb90e04d),
	.w4(32'hbba7749c),
	.w5(32'h3b1a3d45),
	.w6(32'h3b3aaae0),
	.w7(32'h3bd922c0),
	.w8(32'h3bb1b942),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c93cc),
	.w1(32'h3dad236b),
	.w2(32'h3bb1d817),
	.w3(32'h3b80c936),
	.w4(32'h3d356115),
	.w5(32'h3b9fdcf4),
	.w6(32'h3d037952),
	.w7(32'hbbe9aeb7),
	.w8(32'hbd2647fa),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd91e252),
	.w1(32'h3bfcc51f),
	.w2(32'hbbade03c),
	.w3(32'hbd2c8549),
	.w4(32'h3a7a89c6),
	.w5(32'hbba283f3),
	.w6(32'h3b83ad9c),
	.w7(32'hbb107eb1),
	.w8(32'hb9e13233),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71128),
	.w1(32'h3b143f62),
	.w2(32'h3c138c7f),
	.w3(32'h3a008ef8),
	.w4(32'h3a2cb4e9),
	.w5(32'hb9bc8653),
	.w6(32'h3c0f068f),
	.w7(32'h3a6aaa30),
	.w8(32'h3c063c5b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd774a7),
	.w1(32'h3b1360d3),
	.w2(32'hbac6ada1),
	.w3(32'h3babac2d),
	.w4(32'hbc051472),
	.w5(32'hbb8da093),
	.w6(32'h3b08a804),
	.w7(32'hbbac7536),
	.w8(32'h3b8c7046),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae837d4),
	.w1(32'hb9d06032),
	.w2(32'h3a93f298),
	.w3(32'hbb3eec9a),
	.w4(32'h39ba9d2d),
	.w5(32'h3b754f45),
	.w6(32'h3a862399),
	.w7(32'h3b663672),
	.w8(32'h3ab210f6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f719a),
	.w1(32'h3c6beb85),
	.w2(32'h3b588689),
	.w3(32'h3b2aac24),
	.w4(32'hbc0f694a),
	.w5(32'hbcc889b5),
	.w6(32'h3c4aca75),
	.w7(32'h3cd3b2b9),
	.w8(32'h3caa19f7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule