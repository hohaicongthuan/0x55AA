module layer_10_featuremap_467(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea3617),
	.w1(32'h3b2589d8),
	.w2(32'h3b28ef94),
	.w3(32'hbadc938d),
	.w4(32'h3b2ea1f2),
	.w5(32'h3b5431ef),
	.w6(32'hba816d74),
	.w7(32'h3b0e3f72),
	.w8(32'h3b0a1105),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a58f9),
	.w1(32'hbb6d1f2f),
	.w2(32'hbb8232be),
	.w3(32'h3b1ec9f0),
	.w4(32'hbbcf770f),
	.w5(32'hbbe405b9),
	.w6(32'h3b11f79c),
	.w7(32'hbb8e6cc3),
	.w8(32'hbbe1a56d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbe611),
	.w1(32'hbadf9385),
	.w2(32'hbb45826e),
	.w3(32'h3a83d088),
	.w4(32'h39f4c1b8),
	.w5(32'hba8a58eb),
	.w6(32'hb9ce7f29),
	.w7(32'hba889074),
	.w8(32'hbadaae16),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1db1),
	.w1(32'h3a9305d5),
	.w2(32'h3add3d10),
	.w3(32'hbab9e61c),
	.w4(32'hb9df04f2),
	.w5(32'hbaacfd2a),
	.w6(32'hbaeb3d6d),
	.w7(32'hb950e1bf),
	.w8(32'hbb1f3eac),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28840e),
	.w1(32'h38d050d0),
	.w2(32'h3a2957a8),
	.w3(32'hbac9847b),
	.w4(32'h39589519),
	.w5(32'h3a9cf5a8),
	.w6(32'hbb2d32b0),
	.w7(32'h38db3e57),
	.w8(32'h3a33cffe),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09a2db),
	.w1(32'hb961b5b1),
	.w2(32'hba935312),
	.w3(32'hb9c8a003),
	.w4(32'h37bdf779),
	.w5(32'hbad32e49),
	.w6(32'h390a933b),
	.w7(32'hb9a456be),
	.w8(32'hb95985d9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba94f03),
	.w1(32'h3c9cc84a),
	.w2(32'h3b69d071),
	.w3(32'hbaf0af13),
	.w4(32'h3c9323b8),
	.w5(32'h3b228d6a),
	.w6(32'h3c22c65e),
	.w7(32'h3c22918b),
	.w8(32'hba92be6b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a6272),
	.w1(32'h3c116f35),
	.w2(32'hbc99ce68),
	.w3(32'h3b8a5c26),
	.w4(32'h3b42796d),
	.w5(32'hba7a086f),
	.w6(32'hbc7b9477),
	.w7(32'h3aabae67),
	.w8(32'hbc9135e1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae260be),
	.w1(32'hba5cceb7),
	.w2(32'hbaa4ee17),
	.w3(32'h3abb9169),
	.w4(32'hba22a295),
	.w5(32'hb99bb6ec),
	.w6(32'h38d56e24),
	.w7(32'hb9d8b919),
	.w8(32'hba4a7e4c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bd43c),
	.w1(32'h3680aa22),
	.w2(32'hbc877537),
	.w3(32'hbbe42aaf),
	.w4(32'h3c0a088c),
	.w5(32'hbc21883c),
	.w6(32'h3aab8e8a),
	.w7(32'h3c0d4547),
	.w8(32'hbb937b89),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dc678),
	.w1(32'hbb26a5c6),
	.w2(32'hba761ca5),
	.w3(32'hb9d87a6f),
	.w4(32'hbaec73d1),
	.w5(32'h37e7b012),
	.w6(32'hba3de9d5),
	.w7(32'hbb481d37),
	.w8(32'hbb3a3234),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c6fbd),
	.w1(32'h3c828acd),
	.w2(32'h3c229a38),
	.w3(32'hbc4670a4),
	.w4(32'h3cbcc84c),
	.w5(32'h3bb828d3),
	.w6(32'hbb820050),
	.w7(32'h3ca7c035),
	.w8(32'hbbb20c6b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd01179),
	.w1(32'h3b9c0668),
	.w2(32'hbc6c1b82),
	.w3(32'hbb0d51c7),
	.w4(32'h3bea5fba),
	.w5(32'hbc36b33e),
	.w6(32'hbafa6b22),
	.w7(32'h3b51a883),
	.w8(32'hbc03f483),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68b9ae),
	.w1(32'hbb1cfcbe),
	.w2(32'hbc21df41),
	.w3(32'h3c2dc394),
	.w4(32'hbb77f85c),
	.w5(32'hbb9aed87),
	.w6(32'h3b7b1e46),
	.w7(32'hbbb1a0c4),
	.w8(32'hbbffc1de),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf786f5),
	.w1(32'hbb66e3b3),
	.w2(32'hbba15733),
	.w3(32'hbbc08898),
	.w4(32'hbbc78f5c),
	.w5(32'hbbb1f0d8),
	.w6(32'hbaa765c6),
	.w7(32'hbb048724),
	.w8(32'hbbbf90c0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ef2a4),
	.w1(32'hbc1bcc8e),
	.w2(32'hbcc98274),
	.w3(32'h3bf3c025),
	.w4(32'hbb012cf5),
	.w5(32'hbcdaa2f8),
	.w6(32'h3a27e5f0),
	.w7(32'hbc09f098),
	.w8(32'hbc653596),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d051c),
	.w1(32'h3a573225),
	.w2(32'h3a920a24),
	.w3(32'hbb23c579),
	.w4(32'h39f95995),
	.w5(32'h3aef6668),
	.w6(32'hba371ea2),
	.w7(32'h3b20dda9),
	.w8(32'h3b28bf2c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da2c1),
	.w1(32'h3c463ab3),
	.w2(32'hbcd6702b),
	.w3(32'h3c5c71e0),
	.w4(32'h3c900934),
	.w5(32'hbc32b02a),
	.w6(32'h3a8e82ec),
	.w7(32'h3bd39366),
	.w8(32'hbc3bd89a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb57b6),
	.w1(32'h3b8e3118),
	.w2(32'hbc6f1677),
	.w3(32'h3bc41653),
	.w4(32'h3bc7dd91),
	.w5(32'hbc0c910c),
	.w6(32'h3afa3b11),
	.w7(32'h3aae76bf),
	.w8(32'hbc033fdd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372f926e),
	.w1(32'hbab10c27),
	.w2(32'hb9b9292a),
	.w3(32'hba81cf5b),
	.w4(32'hbb0743f6),
	.w5(32'hba084840),
	.w6(32'h38fa966d),
	.w7(32'hbb046e16),
	.w8(32'hbb72cd91),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd6682),
	.w1(32'h3aef7076),
	.w2(32'h3a19f68b),
	.w3(32'hba2bfcbb),
	.w4(32'h3992d159),
	.w5(32'hbaa09624),
	.w6(32'hba5560d8),
	.w7(32'hb8b161f1),
	.w8(32'hbaa243b3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e386f),
	.w1(32'h3a4711a6),
	.w2(32'h3a3186b1),
	.w3(32'hbb97a8fd),
	.w4(32'hbad0e88d),
	.w5(32'hbb118fc6),
	.w6(32'hbb2140be),
	.w7(32'hba1214f4),
	.w8(32'hbb60a4f2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c4ff6),
	.w1(32'h3c2a75a9),
	.w2(32'hbc0da1e0),
	.w3(32'h39b8a4af),
	.w4(32'h3cc64566),
	.w5(32'hbc5d0fac),
	.w6(32'h3c0d9d8e),
	.w7(32'h3ca22a04),
	.w8(32'hb8cfd117),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e0968),
	.w1(32'hbb2e2ffb),
	.w2(32'hbc23fc68),
	.w3(32'hbba04870),
	.w4(32'hb9852a4d),
	.w5(32'hbc10c43c),
	.w6(32'hbb4feac7),
	.w7(32'h3b74fed5),
	.w8(32'hbb868cd0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b5201),
	.w1(32'hbb8a5c33),
	.w2(32'hba8f64f5),
	.w3(32'hbc8ea140),
	.w4(32'hbc3c0faf),
	.w5(32'hbc3dc63b),
	.w6(32'hbc2b06ef),
	.w7(32'hbb8c5c71),
	.w8(32'hbc522452),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace7ecf),
	.w1(32'h3adb2797),
	.w2(32'h3a987862),
	.w3(32'h3934603a),
	.w4(32'h3aa9f497),
	.w5(32'hb6b7eb24),
	.w6(32'hba999ad5),
	.w7(32'h3aec12f8),
	.w8(32'h3a42bc63),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56e3fd),
	.w1(32'h3a9b1c8c),
	.w2(32'h3b0d2416),
	.w3(32'hb9dae7c4),
	.w4(32'hb8bba278),
	.w5(32'h3a090858),
	.w6(32'hb9e9c49e),
	.w7(32'hb9f9ef4d),
	.w8(32'h3a89742b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4bf20),
	.w1(32'h3c02f8b3),
	.w2(32'hbb8e29c8),
	.w3(32'hbc4454bd),
	.w4(32'h3bacb613),
	.w5(32'hbc193a5b),
	.w6(32'h39c739d6),
	.w7(32'h3c986c1d),
	.w8(32'hbbf85a87),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5338e),
	.w1(32'h39ef56a9),
	.w2(32'h3ac22fc4),
	.w3(32'hbba6a949),
	.w4(32'hb8ab640d),
	.w5(32'h3b53e228),
	.w6(32'hbba63ebd),
	.w7(32'h3a766408),
	.w8(32'h3b56373d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebd69e),
	.w1(32'h3bee8a96),
	.w2(32'hbba6d645),
	.w3(32'hbc0bc996),
	.w4(32'h3b333c2a),
	.w5(32'hbc2b2013),
	.w6(32'hb8be0100),
	.w7(32'h3c65eb65),
	.w8(32'hbc2cb527),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a119a67),
	.w1(32'hb86577bb),
	.w2(32'hba12aead),
	.w3(32'h3a230d6a),
	.w4(32'hbaf948b8),
	.w5(32'hbb0340e0),
	.w6(32'h3a0dce90),
	.w7(32'hbae583ad),
	.w8(32'hbb21fa22),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8e76f),
	.w1(32'hbb02366b),
	.w2(32'hbb05d776),
	.w3(32'hba967538),
	.w4(32'hbaad57c8),
	.w5(32'hbadadaf6),
	.w6(32'hbae6371f),
	.w7(32'hba8cde8f),
	.w8(32'hba5b23be),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bcdd6),
	.w1(32'h3986966d),
	.w2(32'hbbf1b166),
	.w3(32'hba90abb1),
	.w4(32'h3b5e046a),
	.w5(32'hbb57c5e6),
	.w6(32'hba9e4c0e),
	.w7(32'h3b47eb1f),
	.w8(32'hbb28b9c0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2857e2),
	.w1(32'h39fb3ad7),
	.w2(32'h3aeaf838),
	.w3(32'hbba6475a),
	.w4(32'hbb69dae3),
	.w5(32'hbb0f4325),
	.w6(32'hbb0952a5),
	.w7(32'hba2e364e),
	.w8(32'hbae06291),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d4790),
	.w1(32'hb8c8516a),
	.w2(32'hba827b58),
	.w3(32'hbab8206f),
	.w4(32'h3acac214),
	.w5(32'hbb0e1848),
	.w6(32'h3b4b2141),
	.w7(32'h3990dd92),
	.w8(32'hbb70ab85),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fbccf),
	.w1(32'h3c07bd29),
	.w2(32'h3bc9efc4),
	.w3(32'hbb8c16b5),
	.w4(32'h3c0b14a1),
	.w5(32'h3b358db4),
	.w6(32'hbb868dde),
	.w7(32'h3b505f91),
	.w8(32'hbb63a3f8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ebae2),
	.w1(32'h3ca04439),
	.w2(32'h3d2efd3a),
	.w3(32'hbd25fcfc),
	.w4(32'h3cfe88b5),
	.w5(32'h3d39e6ed),
	.w6(32'h3953639e),
	.w7(32'h3d3304bf),
	.w8(32'h3c135781),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc997ce0),
	.w1(32'h3c129e82),
	.w2(32'h3bb8e60b),
	.w3(32'hbc9ae632),
	.w4(32'hbb223454),
	.w5(32'hbb81b8f5),
	.w6(32'hbb4427ec),
	.w7(32'h3c4dafc0),
	.w8(32'hbc472f1d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ff34e),
	.w1(32'h3c4150eb),
	.w2(32'h3b62321d),
	.w3(32'hbc8d3d6e),
	.w4(32'h3bb47f19),
	.w5(32'hbbb27238),
	.w6(32'hbbeb0fea),
	.w7(32'h3cbc1729),
	.w8(32'hbb51eda8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5ac3c),
	.w1(32'h3b10cd77),
	.w2(32'h3887a03c),
	.w3(32'hbb2742dc),
	.w4(32'h37c5f0d1),
	.w5(32'hba486ccb),
	.w6(32'hba5f9cc0),
	.w7(32'h399ad42a),
	.w8(32'hbb97f6a6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9580e77),
	.w1(32'hba33072a),
	.w2(32'h37293c2f),
	.w3(32'hb9cea94b),
	.w4(32'hb7dba6c0),
	.w5(32'hba6f382d),
	.w6(32'hba7c7f46),
	.w7(32'hba6ae12b),
	.w8(32'h3a036904),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d76ff),
	.w1(32'hba723281),
	.w2(32'hb94ada84),
	.w3(32'hba39328e),
	.w4(32'hbafabbd7),
	.w5(32'hbab81c42),
	.w6(32'h39bdb947),
	.w7(32'hbafcbdd2),
	.w8(32'hbab2b35c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb512c),
	.w1(32'hb9e3076e),
	.w2(32'hb9cedf63),
	.w3(32'hbae81ceb),
	.w4(32'hba6dd978),
	.w5(32'hbb0413ab),
	.w6(32'hba52cb56),
	.w7(32'hb99e71b6),
	.w8(32'hba87bc55),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc684f4d),
	.w1(32'h3b3efc0f),
	.w2(32'hbcb4edc0),
	.w3(32'hbbabbcbe),
	.w4(32'h3be02580),
	.w5(32'hbc6c909b),
	.w6(32'hbc2e5bf0),
	.w7(32'hba16b8a6),
	.w8(32'hbbd66991),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22dd89),
	.w1(32'hbb57ce7c),
	.w2(32'hbb247c7d),
	.w3(32'hbc1a6ef7),
	.w4(32'hbb8edf6e),
	.w5(32'hbb38f34f),
	.w6(32'hbb0fa222),
	.w7(32'h3b9e022b),
	.w8(32'h3b08ec21),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75e03d),
	.w1(32'hbabddc1a),
	.w2(32'hbc218821),
	.w3(32'hbc69cbcb),
	.w4(32'hbbf21578),
	.w5(32'hbc1c3686),
	.w6(32'hbc31970a),
	.w7(32'hbb3e4bec),
	.w8(32'hbc313c50),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b1395),
	.w1(32'hbbcd382e),
	.w2(32'hbbfa90a6),
	.w3(32'hbc340d59),
	.w4(32'hbb2cba50),
	.w5(32'hbbaa21f9),
	.w6(32'hbb795744),
	.w7(32'h3a9f13a9),
	.w8(32'hbab25646),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9109e0),
	.w1(32'h3c4f4d75),
	.w2(32'hbc6f36e8),
	.w3(32'h3b849f08),
	.w4(32'h3cafaefb),
	.w5(32'hbbe6cd83),
	.w6(32'h3b8f240f),
	.w7(32'h3c8dd4a2),
	.w8(32'hbc3faf72),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f42ef),
	.w1(32'h3889cd98),
	.w2(32'h3a308280),
	.w3(32'hb9fd9ddf),
	.w4(32'h39dc11f2),
	.w5(32'h3a2defbc),
	.w6(32'hb7bc088c),
	.w7(32'hba0d8f6e),
	.w8(32'h3a64fa94),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aa210),
	.w1(32'h3b1329b6),
	.w2(32'h39cc14fa),
	.w3(32'hbadca9ef),
	.w4(32'h3b4e973b),
	.w5(32'hbab4d4b2),
	.w6(32'hba717690),
	.w7(32'h3b0a0111),
	.w8(32'hb9a78182),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30d189),
	.w1(32'h3a0eb798),
	.w2(32'h38fcb0f8),
	.w3(32'hba62e6c4),
	.w4(32'h3a68bfe3),
	.w5(32'h399b50d1),
	.w6(32'hbad86fe7),
	.w7(32'h3a6af319),
	.w8(32'h3a5f8903),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52ed4),
	.w1(32'hbb581171),
	.w2(32'hbb8cf490),
	.w3(32'hbb0413dc),
	.w4(32'hbb1261af),
	.w5(32'hbbf7c6e6),
	.w6(32'hbab05b94),
	.w7(32'hbb1d9b3f),
	.w8(32'hba913a45),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39540802),
	.w1(32'h3b3fc0af),
	.w2(32'h3a50763c),
	.w3(32'h39aa9350),
	.w4(32'h3b14f5a3),
	.w5(32'hb9b60097),
	.w6(32'hbb4c0b29),
	.w7(32'h3a527998),
	.w8(32'hb7cadc23),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf630da),
	.w1(32'h3c61eb13),
	.w2(32'hbc9e02f7),
	.w3(32'h3b3449f5),
	.w4(32'h3ca643eb),
	.w5(32'hbbb365c1),
	.w6(32'h3c29afad),
	.w7(32'h3c746e94),
	.w8(32'hbbd82747),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac76c25),
	.w1(32'h3ba9d543),
	.w2(32'hb985b2d4),
	.w3(32'hbb0ed376),
	.w4(32'h38a12875),
	.w5(32'h37fbd1e9),
	.w6(32'hbbbbf9b0),
	.w7(32'hb9fcdad0),
	.w8(32'hba3c8056),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeeec80),
	.w1(32'h3aa92572),
	.w2(32'h3a428718),
	.w3(32'hb9afa83b),
	.w4(32'hba678a63),
	.w5(32'h398827b2),
	.w6(32'hb9b98ece),
	.w7(32'h3a3a0f8f),
	.w8(32'hb90832a6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb0d2f),
	.w1(32'h3a967560),
	.w2(32'h3b00a699),
	.w3(32'h39b1bc81),
	.w4(32'h399d139c),
	.w5(32'h3a45d26d),
	.w6(32'h39a14a51),
	.w7(32'h399c8a9f),
	.w8(32'h3a9306e7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11c1af),
	.w1(32'hbb27e3ec),
	.w2(32'hbb44c84c),
	.w3(32'h3af70dcb),
	.w4(32'hbac4a368),
	.w5(32'hbad65e8c),
	.w6(32'h3b397b18),
	.w7(32'h3a07da0f),
	.w8(32'hbafd4ea9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4007e6),
	.w1(32'h3b575e20),
	.w2(32'h3b2a7586),
	.w3(32'hbb8220b4),
	.w4(32'h3b497047),
	.w5(32'h3b133c42),
	.w6(32'hbb27f5e4),
	.w7(32'h3ade0065),
	.w8(32'h39b90496),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a8c27),
	.w1(32'h3aba53c4),
	.w2(32'hba778b79),
	.w3(32'h3b0ebcac),
	.w4(32'h3ab4d4d2),
	.w5(32'hbad99e69),
	.w6(32'h3b875473),
	.w7(32'h3a71715f),
	.w8(32'hbac9445e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06bd16),
	.w1(32'h3ba035cc),
	.w2(32'hbbb22f12),
	.w3(32'hbafe4b61),
	.w4(32'h3b5b70f2),
	.w5(32'hbbe1cab0),
	.w6(32'hbb86b062),
	.w7(32'h3abd5e43),
	.w8(32'hbb164e20),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadf7e3),
	.w1(32'hbb591093),
	.w2(32'hbc19cc8b),
	.w3(32'hba3cefb1),
	.w4(32'hbb99e87d),
	.w5(32'hbc1695a7),
	.w6(32'hbbe19200),
	.w7(32'hbc019fd7),
	.w8(32'hbb98d4be),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98418b9),
	.w1(32'h39b2f6f8),
	.w2(32'hbab985ac),
	.w3(32'hba75024c),
	.w4(32'h3a9f5349),
	.w5(32'hbad9845c),
	.w6(32'hba6f35e0),
	.w7(32'h3a98c0a8),
	.w8(32'hbb3274ce),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad22bb7),
	.w1(32'h39c5b429),
	.w2(32'h3a437947),
	.w3(32'hbab9c73a),
	.w4(32'h3a5afc1e),
	.w5(32'hb9004354),
	.w6(32'hbb13c005),
	.w7(32'h3a52529b),
	.w8(32'h3ab1ec9a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7c878),
	.w1(32'h3b403c4b),
	.w2(32'h3b3e6cd1),
	.w3(32'h3ae85bda),
	.w4(32'h3af20221),
	.w5(32'h3ad087ca),
	.w6(32'h3b66dd0a),
	.w7(32'h3b249876),
	.w8(32'h3afff714),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b6222),
	.w1(32'hba89388c),
	.w2(32'hb96f2fda),
	.w3(32'h3abea3f1),
	.w4(32'hba2de306),
	.w5(32'hba00ab7a),
	.w6(32'h3a99da3f),
	.w7(32'hbaa1efd6),
	.w8(32'hba3c49e5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6842e3),
	.w1(32'hbc37be8e),
	.w2(32'hbd22cf38),
	.w3(32'h3c19542e),
	.w4(32'h3c963a53),
	.w5(32'hbc922432),
	.w6(32'h3cab324e),
	.w7(32'h3c479322),
	.w8(32'hbc3fb0ab),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5134c),
	.w1(32'h3c881c3f),
	.w2(32'h3afb72cc),
	.w3(32'hbbd79155),
	.w4(32'h3ad41929),
	.w5(32'hbc2ec262),
	.w6(32'hbcfefd74),
	.w7(32'hbc88a494),
	.w8(32'hbcac28ce),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b720b),
	.w1(32'h3bb9c49f),
	.w2(32'hbbe61d31),
	.w3(32'hbb6297bc),
	.w4(32'h3bafa12b),
	.w5(32'hbc0fafc4),
	.w6(32'hbc5b1124),
	.w7(32'hbb17f034),
	.w8(32'hbb260d1f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93ee52),
	.w1(32'h3b62a296),
	.w2(32'h3af7b499),
	.w3(32'hbcb67cbd),
	.w4(32'hbc0cfe07),
	.w5(32'hbbff5d84),
	.w6(32'hbc122668),
	.w7(32'h3bddca10),
	.w8(32'hbc11c1e2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e0af3),
	.w1(32'hbac0b0ef),
	.w2(32'hba795449),
	.w3(32'hbb3090df),
	.w4(32'hbb012a1e),
	.w5(32'h3a912131),
	.w6(32'hbab0295e),
	.w7(32'h3959c6f3),
	.w8(32'h3a99c6b8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a439057),
	.w1(32'hbaf422f0),
	.w2(32'h3a166c68),
	.w3(32'h3ab52196),
	.w4(32'hba8427f7),
	.w5(32'h3b42375f),
	.w6(32'h399265db),
	.w7(32'hb9ca17bb),
	.w8(32'h39f3ca2a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87a666),
	.w1(32'hba916be1),
	.w2(32'h3b358600),
	.w3(32'hb96690e2),
	.w4(32'hbb01199a),
	.w5(32'h3b83b436),
	.w6(32'h3b073370),
	.w7(32'hbb23ab03),
	.w8(32'h3b382faa),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3729f9de),
	.w1(32'h3afcf164),
	.w2(32'hbbb47d12),
	.w3(32'h3abab110),
	.w4(32'h3ae9febe),
	.w5(32'hbb2d1d08),
	.w6(32'hbb486fb7),
	.w7(32'hbad46f8a),
	.w8(32'hbbaaa8dd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a756a),
	.w1(32'h3982cbe7),
	.w2(32'h3a45f15a),
	.w3(32'hbafbb09f),
	.w4(32'h3af2cc36),
	.w5(32'h3b0d5fe5),
	.w6(32'hba5422fd),
	.w7(32'h3ae42d95),
	.w8(32'h3b2ff609),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb18619),
	.w1(32'h3b21a288),
	.w2(32'hbb9432cc),
	.w3(32'hbb2affce),
	.w4(32'h3c3db715),
	.w5(32'h3b4cd35a),
	.w6(32'h3c1600f8),
	.w7(32'h3c471125),
	.w8(32'h3b145e9c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb628ecd),
	.w1(32'h3b949c0b),
	.w2(32'hbb0c7594),
	.w3(32'hbb3ecdfc),
	.w4(32'h3c005cdd),
	.w5(32'hbb4db80a),
	.w6(32'hbc066b9a),
	.w7(32'h3bd97003),
	.w8(32'hbc4cacbc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc210adf),
	.w1(32'hbc139343),
	.w2(32'hbc1bdd13),
	.w3(32'hbc5380ee),
	.w4(32'hbc3adeed),
	.w5(32'hbc33c8ae),
	.w6(32'hbbc22a2c),
	.w7(32'hbb6776ec),
	.w8(32'hbc220976),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb218561),
	.w1(32'h39e04b7a),
	.w2(32'hbc0cfd7d),
	.w3(32'h3a305e79),
	.w4(32'h3b8c39dc),
	.w5(32'hbb8f53d6),
	.w6(32'hbaccf17a),
	.w7(32'h3af0c024),
	.w8(32'hbb223c19),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be08d),
	.w1(32'h3a1613e3),
	.w2(32'hbc19e6aa),
	.w3(32'h38fa0cfb),
	.w4(32'h3c19659c),
	.w5(32'hbb940f75),
	.w6(32'h3c4a53e2),
	.w7(32'h3c28b8be),
	.w8(32'hbb7ec0a1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3f81e),
	.w1(32'hba236a7d),
	.w2(32'h3b2e0338),
	.w3(32'hbbcf3cf9),
	.w4(32'h3ad7111b),
	.w5(32'hbaa6683d),
	.w6(32'hbb8ff0e9),
	.w7(32'h3bd01351),
	.w8(32'h3bec34ff),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac293c0),
	.w1(32'h3bccd859),
	.w2(32'hbb1548bd),
	.w3(32'h3ba53ce3),
	.w4(32'h3c0d906d),
	.w5(32'hba54e5d3),
	.w6(32'h3bdd86eb),
	.w7(32'h3bf195ec),
	.w8(32'hba9a3058),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaad0c),
	.w1(32'hb730dc17),
	.w2(32'hb738e6cb),
	.w3(32'h3ab964aa),
	.w4(32'hb98c9fd9),
	.w5(32'hba646cf7),
	.w6(32'h3a311702),
	.w7(32'hba88336d),
	.w8(32'hb9d97cdf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af03095),
	.w1(32'h38d52d1d),
	.w2(32'h39c10e6c),
	.w3(32'h3b592fb8),
	.w4(32'h3a914cab),
	.w5(32'h3b18847a),
	.w6(32'h3b4084a3),
	.w7(32'h3aa9e9f2),
	.w8(32'h3a617631),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba996717),
	.w1(32'hb9c9a881),
	.w2(32'h3a134cc9),
	.w3(32'hbac411f9),
	.w4(32'hbace5cf7),
	.w5(32'h3ad1ad0b),
	.w6(32'h3a05dd27),
	.w7(32'hbb168b21),
	.w8(32'hb9bc069d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ce82f),
	.w1(32'hb9fbf285),
	.w2(32'hbb1aef2d),
	.w3(32'h3aa8ef9c),
	.w4(32'h3a9a54d4),
	.w5(32'h3a4afb84),
	.w6(32'h3a564325),
	.w7(32'h393845c4),
	.w8(32'hbaa4b2d0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3a5b),
	.w1(32'hbba4317e),
	.w2(32'h3b791d09),
	.w3(32'hbc716060),
	.w4(32'hbbf2de09),
	.w5(32'h3b0bcf21),
	.w6(32'hbbbaf689),
	.w7(32'h3b48deb8),
	.w8(32'h3b6c60cc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff1348),
	.w1(32'hbb586c06),
	.w2(32'hbac118a5),
	.w3(32'hbb855b49),
	.w4(32'hbb40cf1a),
	.w5(32'hbb4ac040),
	.w6(32'hbb47e43f),
	.w7(32'hbb6a1a7f),
	.w8(32'hbaa01635),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a995),
	.w1(32'hbb05dd1c),
	.w2(32'h39c81a35),
	.w3(32'hbc2b5641),
	.w4(32'hbb337cdb),
	.w5(32'hbb6864b8),
	.w6(32'hbb973553),
	.w7(32'hbb394e72),
	.w8(32'hbb20d08a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d7fe2),
	.w1(32'h3b9a4a3b),
	.w2(32'hbc5b9287),
	.w3(32'hbb028108),
	.w4(32'h3c12ded7),
	.w5(32'hbbc70d16),
	.w6(32'hbaf8ba05),
	.w7(32'h3b9bc180),
	.w8(32'hbc1510ab),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a483a),
	.w1(32'h3bb77560),
	.w2(32'hb8300651),
	.w3(32'hbc230541),
	.w4(32'h3b6f6f1e),
	.w5(32'h3b658505),
	.w6(32'hbb2bd82f),
	.w7(32'h3c292b89),
	.w8(32'h3b805d0b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dab69),
	.w1(32'h3c1d829e),
	.w2(32'hbbf11cea),
	.w3(32'hbb8c83ce),
	.w4(32'h3cd691b9),
	.w5(32'hbbdcd20d),
	.w6(32'h3c6d04c0),
	.w7(32'h3cdc8a9f),
	.w8(32'hb9e96d82),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd8f10),
	.w1(32'h3b99e764),
	.w2(32'h3a305bc2),
	.w3(32'hbb65bb9d),
	.w4(32'h3b5c7aeb),
	.w5(32'hba99b656),
	.w6(32'h3b20d717),
	.w7(32'h3c04e8ce),
	.w8(32'h3bb4dc28),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948303),
	.w1(32'h3ae12edc),
	.w2(32'hbccacef7),
	.w3(32'h3c5fd8c1),
	.w4(32'h3b486b0f),
	.w5(32'hbcab1869),
	.w6(32'h3bdaf9ec),
	.w7(32'h3ab66a35),
	.w8(32'hbc6bc322),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66f7ab),
	.w1(32'h3b2e962c),
	.w2(32'hbb496cb2),
	.w3(32'h3af902d1),
	.w4(32'h3b4e71b9),
	.w5(32'hbb6b173f),
	.w6(32'h3c3869a9),
	.w7(32'h3c15a3ec),
	.w8(32'h3b6869bb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0d90f),
	.w1(32'hbb8f8d1f),
	.w2(32'hbc141cba),
	.w3(32'hba7d5e67),
	.w4(32'hbbae8a36),
	.w5(32'hbc328ede),
	.w6(32'hbb95c6b6),
	.w7(32'hba84749e),
	.w8(32'hbc2a469f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0e08a),
	.w1(32'hba86b321),
	.w2(32'hbb01d33b),
	.w3(32'hbbad23f8),
	.w4(32'hbb6e8942),
	.w5(32'h398ab28e),
	.w6(32'hbb1a2c11),
	.w7(32'hbb32b3ad),
	.w8(32'h3a762bc4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba6b65),
	.w1(32'h3bf7d935),
	.w2(32'hbc7cccb3),
	.w3(32'h3a5ce2cd),
	.w4(32'h3c3be647),
	.w5(32'hbbba8c66),
	.w6(32'hba4b6642),
	.w7(32'h3bdb5fe4),
	.w8(32'hbbf0542e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce14c64),
	.w1(32'h3bb8e2f0),
	.w2(32'hbb1c74a9),
	.w3(32'hbc5889be),
	.w4(32'h3c8ff950),
	.w5(32'h3bc8dd07),
	.w6(32'h3c404e7e),
	.w7(32'h3cdf1248),
	.w8(32'h3c85128e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98ca27),
	.w1(32'h3c89719b),
	.w2(32'h3d090206),
	.w3(32'hbcbada2c),
	.w4(32'h3c9c032b),
	.w5(32'h3c57f07a),
	.w6(32'hbc90233b),
	.w7(32'h3b9403e3),
	.w8(32'hbbacfd48),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07499d),
	.w1(32'h3c7519cf),
	.w2(32'h3c6a25c7),
	.w3(32'hbc3a016d),
	.w4(32'h3c14b2f4),
	.w5(32'h3c308373),
	.w6(32'h37e657a8),
	.w7(32'h3c0601c7),
	.w8(32'hbbcb1f3c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc008f2e),
	.w1(32'hbaaa7193),
	.w2(32'hbbb3c8e9),
	.w3(32'hbc141322),
	.w4(32'hbbe29cd8),
	.w5(32'hbbbd69db),
	.w6(32'hbb708906),
	.w7(32'hb96ded56),
	.w8(32'hbbaa57d8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca57605),
	.w1(32'h3c2e65a4),
	.w2(32'h3bd25b02),
	.w3(32'hbc2a2908),
	.w4(32'h3cdc56fc),
	.w5(32'h3c54a5a2),
	.w6(32'h3b4e63bb),
	.w7(32'h3ccc5e54),
	.w8(32'h3be112ac),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab56347),
	.w1(32'hbacb3ee8),
	.w2(32'h39c4fb0b),
	.w3(32'h3b517daf),
	.w4(32'hbb3378a5),
	.w5(32'h3ac859c0),
	.w6(32'h3a1c0834),
	.w7(32'hbaca8186),
	.w8(32'hba15ee25),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc465a66),
	.w1(32'h3adbddbf),
	.w2(32'h3c42f155),
	.w3(32'hbc4be705),
	.w4(32'h3c933558),
	.w5(32'h3c8d108f),
	.w6(32'hbc81d190),
	.w7(32'h3c61bc4c),
	.w8(32'hbba62134),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35c979),
	.w1(32'h3aedc47e),
	.w2(32'h3c84741c),
	.w3(32'hbbedf498),
	.w4(32'h3bdff53a),
	.w5(32'h3c5b3d61),
	.w6(32'hbbf78d32),
	.w7(32'h3c3d10fc),
	.w8(32'h3c4212ae),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2b314),
	.w1(32'h39ba3ce0),
	.w2(32'hb97c26ab),
	.w3(32'h38f0f4df),
	.w4(32'h3a31f725),
	.w5(32'hbac13484),
	.w6(32'h3987d64a),
	.w7(32'h3a46b462),
	.w8(32'hbad4c335),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f8cea),
	.w1(32'hbb2e3567),
	.w2(32'hbb8c1b6e),
	.w3(32'h3b628906),
	.w4(32'hba70e172),
	.w5(32'hbbffd783),
	.w6(32'h3bbc81e2),
	.w7(32'h3aa33f64),
	.w8(32'hbb89960d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb495382),
	.w1(32'h3abf2ff4),
	.w2(32'hbc4cf431),
	.w3(32'hba5c92c3),
	.w4(32'h3bc61659),
	.w5(32'hbc1d3042),
	.w6(32'hbb090eed),
	.w7(32'h3af218f8),
	.w8(32'hbc18ec05),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9c29),
	.w1(32'h3af2ce66),
	.w2(32'h38be36a5),
	.w3(32'hbb794ec3),
	.w4(32'hbaa44d87),
	.w5(32'hbb767554),
	.w6(32'h3a546360),
	.w7(32'h3b26ba0f),
	.w8(32'hbb157265),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb992d3b),
	.w1(32'h39c179ab),
	.w2(32'hbc14186b),
	.w3(32'hba11d243),
	.w4(32'h3b90872b),
	.w5(32'hbbb17aa0),
	.w6(32'h3ba90216),
	.w7(32'h3c25031a),
	.w8(32'hbbaad7f0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc85c7),
	.w1(32'hbb0a9149),
	.w2(32'hbb1b8a55),
	.w3(32'hbc15c668),
	.w4(32'hbbbc810c),
	.w5(32'hbb49bab4),
	.w6(32'hbb450e61),
	.w7(32'hba602a3d),
	.w8(32'hbb78a788),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc208d5d),
	.w1(32'h3c027bd9),
	.w2(32'h3c1a15de),
	.w3(32'hbc60eadc),
	.w4(32'h3b8e58e9),
	.w5(32'hbb692ede),
	.w6(32'hbc9783d0),
	.w7(32'hbbb90f1a),
	.w8(32'hbc3bd894),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d4509),
	.w1(32'hbaea9963),
	.w2(32'hbca75042),
	.w3(32'h3c38d5cc),
	.w4(32'h3b8502d7),
	.w5(32'hbcaadce1),
	.w6(32'h3b31eda8),
	.w7(32'h3b09e261),
	.w8(32'hbc1720d3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8dc61),
	.w1(32'hb9c4b16b),
	.w2(32'hbaaaa67b),
	.w3(32'hbb200781),
	.w4(32'hba953576),
	.w5(32'hbb2551b5),
	.w6(32'hb9f89db8),
	.w7(32'h3b429681),
	.w8(32'hbae99025),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b033621),
	.w1(32'hb9a4daf9),
	.w2(32'h38245d24),
	.w3(32'h3a37cb9f),
	.w4(32'hba943ab1),
	.w5(32'h399168e9),
	.w6(32'h3aa06347),
	.w7(32'hb9e32880),
	.w8(32'h38181846),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35fa6c),
	.w1(32'h396fd4a5),
	.w2(32'hbaca39ea),
	.w3(32'h3adec3a5),
	.w4(32'h3b0e128e),
	.w5(32'h3a6bcf4d),
	.w6(32'hba81a781),
	.w7(32'h3a447492),
	.w8(32'h3a08884c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c16fa),
	.w1(32'h3aa03be8),
	.w2(32'h39e322ac),
	.w3(32'h3ae6476f),
	.w4(32'h38d09ba1),
	.w5(32'hbac02327),
	.w6(32'h3aa79ace),
	.w7(32'h3aaf873e),
	.w8(32'hbacebd30),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a275b9),
	.w1(32'hbb3b4d37),
	.w2(32'hba48a8ae),
	.w3(32'hba7a26a7),
	.w4(32'hbac3d842),
	.w5(32'h3a7ff271),
	.w6(32'h3a576cfd),
	.w7(32'hbab66d26),
	.w8(32'hb88f7c6f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cbd2e),
	.w1(32'hbb1825d6),
	.w2(32'hb9d21722),
	.w3(32'hbc090a4c),
	.w4(32'hbba1438e),
	.w5(32'h3a3e94f6),
	.w6(32'hbba3803d),
	.w7(32'hba797c27),
	.w8(32'h3b0199ca),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b219286),
	.w1(32'hba97165f),
	.w2(32'hba1d5976),
	.w3(32'h3b1227b0),
	.w4(32'hba28e9c0),
	.w5(32'hba7a0eb9),
	.w6(32'h3a8ec998),
	.w7(32'hba24670a),
	.w8(32'h396f061f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac78118),
	.w1(32'h3bb94672),
	.w2(32'hbb8786df),
	.w3(32'h3a69b40c),
	.w4(32'h3bc978af),
	.w5(32'hbb09b78b),
	.w6(32'h3b9fe90f),
	.w7(32'h3bc3718a),
	.w8(32'hbb03c2bf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc17e4f),
	.w1(32'hbae42e73),
	.w2(32'hbbc8abcd),
	.w3(32'hbbaa6bea),
	.w4(32'hbc2a35fb),
	.w5(32'hbc3d7c76),
	.w6(32'hbb5f8b2a),
	.w7(32'hbb956479),
	.w8(32'hbc476807),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cfb66),
	.w1(32'h3b18e149),
	.w2(32'h3a88754b),
	.w3(32'h3b0e308e),
	.w4(32'h3aa8286c),
	.w5(32'h3afecbcc),
	.w6(32'h3b1e9223),
	.w7(32'h3a01b97d),
	.w8(32'h3b2d76f4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ef95a),
	.w1(32'hbab67d4c),
	.w2(32'h3b02a6b1),
	.w3(32'h3af4207d),
	.w4(32'hba935850),
	.w5(32'h39f24b18),
	.w6(32'h3a7609c8),
	.w7(32'hba06ff53),
	.w8(32'h3992a808),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf7bf7),
	.w1(32'h3a0e899b),
	.w2(32'hb8c3f2bf),
	.w3(32'hba4dd576),
	.w4(32'h3aa800db),
	.w5(32'hba204c35),
	.w6(32'hb9b0b255),
	.w7(32'hb81950e9),
	.w8(32'hbafeb84f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aced682),
	.w1(32'h3b2e8fe0),
	.w2(32'hba99b9aa),
	.w3(32'h38718f6a),
	.w4(32'h397a6b02),
	.w5(32'hbb15607e),
	.w6(32'h3a9c6b1e),
	.w7(32'h3b01a9d2),
	.w8(32'hbb65c117),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc313a78),
	.w1(32'h3c96211d),
	.w2(32'h3ba6d3c2),
	.w3(32'hbb6ef7c1),
	.w4(32'h3c5ba363),
	.w5(32'hbc458480),
	.w6(32'hbca85da5),
	.w7(32'hbc0a08b6),
	.w8(32'hbc9d6b5e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc025c61),
	.w1(32'h3b6abd4a),
	.w2(32'hbc9eb4e4),
	.w3(32'h3b243893),
	.w4(32'h3c422115),
	.w5(32'hbc380ab5),
	.w6(32'h3b897dde),
	.w7(32'h3bc42593),
	.w8(32'hbc02d6ef),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d9bf3),
	.w1(32'hbad4e691),
	.w2(32'hbb974a03),
	.w3(32'hbb040d2e),
	.w4(32'h3a017ba0),
	.w5(32'hbb24b35c),
	.w6(32'h3a09b299),
	.w7(32'h3aafb42e),
	.w8(32'hbb91a24c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb069e9b),
	.w1(32'h3b8266f3),
	.w2(32'hba5e51f6),
	.w3(32'hbb863274),
	.w4(32'h3b58035e),
	.w5(32'hba826ffa),
	.w6(32'hbbea7a41),
	.w7(32'hbb08f5c4),
	.w8(32'hbb2a04e4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef86d7),
	.w1(32'hbaa2a7a4),
	.w2(32'hbb50b56a),
	.w3(32'hbb7184ee),
	.w4(32'hbac97b63),
	.w5(32'hba1200df),
	.w6(32'hba5517b6),
	.w7(32'h3a7eb218),
	.w8(32'h38080d1a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad27b44),
	.w1(32'h3a8e425d),
	.w2(32'hbc0dee39),
	.w3(32'h3a6f30c4),
	.w4(32'hb9095406),
	.w5(32'hbb89fe15),
	.w6(32'hbacdbbfd),
	.w7(32'hbb488223),
	.w8(32'hbb600c53),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8928f6),
	.w1(32'h3a3a19ac),
	.w2(32'hbb900281),
	.w3(32'h3b19302d),
	.w4(32'h3ae6cff5),
	.w5(32'hbc0a6a9e),
	.w6(32'h3baabebb),
	.w7(32'h3b96d9c0),
	.w8(32'h393672fa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb3a46),
	.w1(32'h3bdd7ed2),
	.w2(32'hbc999c24),
	.w3(32'h3c12e8e1),
	.w4(32'h3ca003c1),
	.w5(32'hbbf62f2a),
	.w6(32'h3bf865cf),
	.w7(32'h3c52335a),
	.w8(32'hbbaa24be),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78c61d),
	.w1(32'hbb040269),
	.w2(32'hba3313aa),
	.w3(32'hbba099fd),
	.w4(32'hbbcfba88),
	.w5(32'hbb662faa),
	.w6(32'hbac338c8),
	.w7(32'hbad46065),
	.w8(32'hbbd37d31),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29f807),
	.w1(32'hbaadf019),
	.w2(32'hbc04505e),
	.w3(32'h3b8208a6),
	.w4(32'h3bf2109d),
	.w5(32'hbb98730c),
	.w6(32'h3bad3379),
	.w7(32'h3bf4a95f),
	.w8(32'hbb895bd8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b9de),
	.w1(32'h3c2dffda),
	.w2(32'hbbb7a2f3),
	.w3(32'hb825fa0f),
	.w4(32'h3c872624),
	.w5(32'hbb108cf7),
	.w6(32'h3bce9b6b),
	.w7(32'h3c2f4452),
	.w8(32'hbb7b0399),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc137aa),
	.w1(32'hb9211474),
	.w2(32'h3b823e9e),
	.w3(32'hbbd16514),
	.w4(32'hbb1b1c0e),
	.w5(32'hb83dfcf9),
	.w6(32'hbbcc29f6),
	.w7(32'hbb6872c6),
	.w8(32'hbb88cd46),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d8c70),
	.w1(32'h3904c0cf),
	.w2(32'hbc051f4f),
	.w3(32'h3b215cc3),
	.w4(32'h3c0eb310),
	.w5(32'hbb800843),
	.w6(32'h3bf0fc5e),
	.w7(32'h3be64ad8),
	.w8(32'hbb038541),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb140e08),
	.w1(32'hba03aa68),
	.w2(32'hbb8714bd),
	.w3(32'hba6835bd),
	.w4(32'hbb16ebfd),
	.w5(32'hbb86fb78),
	.w6(32'hba7bfd09),
	.w7(32'hbab229f1),
	.w8(32'hbb9423c6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99aee1),
	.w1(32'h3c84f06b),
	.w2(32'hbb981f0d),
	.w3(32'hba2273ac),
	.w4(32'h3c08fad6),
	.w5(32'hbc1dc394),
	.w6(32'hb903a89c),
	.w7(32'h3c035a68),
	.w8(32'hbc923197),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1778c2),
	.w1(32'h3b15377f),
	.w2(32'h3b1862c9),
	.w3(32'h39e699d8),
	.w4(32'h3a88de49),
	.w5(32'h3b8898a7),
	.w6(32'h3a5c886d),
	.w7(32'h3b0c33c1),
	.w8(32'h3b018d3f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c412),
	.w1(32'hbace3129),
	.w2(32'h3a137fb0),
	.w3(32'h3b5fe44f),
	.w4(32'hbafa6135),
	.w5(32'h3adc9970),
	.w6(32'h3a84e35b),
	.w7(32'hbab3bb25),
	.w8(32'h3a454d1b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81a35e),
	.w1(32'hb9977927),
	.w2(32'h3aaa1fa3),
	.w3(32'h3b09100c),
	.w4(32'h3a8c4f97),
	.w5(32'h3aae6272),
	.w6(32'h3ac4d473),
	.w7(32'hb9bce1d2),
	.w8(32'hbac9c4a6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fb0d9),
	.w1(32'hbace1293),
	.w2(32'h3b0309ad),
	.w3(32'hb95f5dee),
	.w4(32'h39efe6a2),
	.w5(32'h3b03f238),
	.w6(32'hbab3701d),
	.w7(32'h3b159360),
	.w8(32'hb9cc898f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc153d79),
	.w1(32'h3aba745c),
	.w2(32'h3afa49c0),
	.w3(32'hbc13f720),
	.w4(32'hbb12bc54),
	.w5(32'h3ace9809),
	.w6(32'hb8991cca),
	.w7(32'h3bb4f49a),
	.w8(32'h3a3778b9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01af10),
	.w1(32'hba8fd32d),
	.w2(32'hbc0886be),
	.w3(32'hbc01ae59),
	.w4(32'hb9c0d67d),
	.w5(32'hbbb5d78e),
	.w6(32'hbc1c708e),
	.w7(32'hbb53732f),
	.w8(32'hbc193e83),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc49d6),
	.w1(32'h3a14cfe4),
	.w2(32'h38fc8a77),
	.w3(32'hbb36632e),
	.w4(32'h38e196bc),
	.w5(32'hbabedad2),
	.w6(32'hbb49b5e4),
	.w7(32'hbacb365e),
	.w8(32'hba889780),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea32d8),
	.w1(32'h3a327239),
	.w2(32'hbc42640f),
	.w3(32'hbb1b15d2),
	.w4(32'h3bb120fa),
	.w5(32'hbb6b25b4),
	.w6(32'h3a19f49b),
	.w7(32'h3bf58a2b),
	.w8(32'hbb597b38),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b6351),
	.w1(32'h382828e6),
	.w2(32'hbba3d4e8),
	.w3(32'hbb0e7aff),
	.w4(32'hba851729),
	.w5(32'hbb7085de),
	.w6(32'hbb5de7fd),
	.w7(32'h39376907),
	.w8(32'hbb8c3bfe),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb191d1),
	.w1(32'h3b7643d1),
	.w2(32'hbc6e44a4),
	.w3(32'h3b63451f),
	.w4(32'h3c639abd),
	.w5(32'hbc12eb6d),
	.w6(32'h3c46240b),
	.w7(32'h3c706101),
	.w8(32'hbbbab7ba),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f4dec),
	.w1(32'hbb1c35db),
	.w2(32'hbc02e571),
	.w3(32'hbc90e1c5),
	.w4(32'hbc24feb8),
	.w5(32'hbbf7a6d6),
	.w6(32'hbab786b5),
	.w7(32'h3c99c31b),
	.w8(32'hbb2791c0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e0a0a),
	.w1(32'h3b8fbbaf),
	.w2(32'h3b8ee618),
	.w3(32'h3b0ca66d),
	.w4(32'hba656eac),
	.w5(32'hbbca1891),
	.w6(32'h3a34e528),
	.w7(32'hbb1faa21),
	.w8(32'hbbbb8202),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81e622),
	.w1(32'h38d005f8),
	.w2(32'h3983c043),
	.w3(32'hba666ef9),
	.w4(32'h3a023fd0),
	.w5(32'h3a332938),
	.w6(32'h374910aa),
	.w7(32'hbaafa510),
	.w8(32'hbb0217c3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aefc1),
	.w1(32'h3a72288c),
	.w2(32'h3a21471f),
	.w3(32'hbc4f16f5),
	.w4(32'hbb6814cf),
	.w5(32'h3a932b51),
	.w6(32'hbc0ef871),
	.w7(32'h3aa21d33),
	.w8(32'h3b5d694a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb790449),
	.w1(32'h3b8a93f3),
	.w2(32'h3bcc7050),
	.w3(32'hbbc072ac),
	.w4(32'h3b4cfa1e),
	.w5(32'h3ba83c82),
	.w6(32'hb9488e81),
	.w7(32'h3bd55c57),
	.w8(32'hba14d221),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ccce8),
	.w1(32'h3a7f2f9d),
	.w2(32'h3b94a5c7),
	.w3(32'hbc279ae7),
	.w4(32'hbb10c4fe),
	.w5(32'hbaa96b26),
	.w6(32'hbbf24c1f),
	.w7(32'hba342ce4),
	.w8(32'hbb7ebfcd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf473f1),
	.w1(32'h3b630ed2),
	.w2(32'h3b4885ce),
	.w3(32'h3a48d1d0),
	.w4(32'h3bd1b1b4),
	.w5(32'h3b62d51c),
	.w6(32'h3b68f203),
	.w7(32'h3b96195e),
	.w8(32'hbaa10568),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b315b8a),
	.w1(32'hba7e8952),
	.w2(32'hb9310c17),
	.w3(32'h39f48261),
	.w4(32'hbb2e93d9),
	.w5(32'hba88c132),
	.w6(32'h3a97dbc8),
	.w7(32'hbb33d220),
	.w8(32'hba1f487f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefe7aa),
	.w1(32'hba88a90c),
	.w2(32'hbc230ade),
	.w3(32'h3a65c4bc),
	.w4(32'h3c018aca),
	.w5(32'hbbc31085),
	.w6(32'h3a95ad35),
	.w7(32'hbab185bf),
	.w8(32'hbc180880),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2711c2),
	.w1(32'h3b092da6),
	.w2(32'hba981c32),
	.w3(32'hbb7e7eaa),
	.w4(32'h3b2c2e6b),
	.w5(32'h39fb8f37),
	.w6(32'h3a61f5b6),
	.w7(32'h3b001f89),
	.w8(32'hb8ccacb4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4d3f),
	.w1(32'h3a6b6f70),
	.w2(32'h3b1cff28),
	.w3(32'hbb99be53),
	.w4(32'hbb806d6c),
	.w5(32'hbb2f746b),
	.w6(32'hbb1041e5),
	.w7(32'hba79e74e),
	.w8(32'h3a294f41),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01991a),
	.w1(32'h3aa46a32),
	.w2(32'h3ace7e49),
	.w3(32'h3a929202),
	.w4(32'h3aefc265),
	.w5(32'h3aba2b92),
	.w6(32'h3b7040b7),
	.w7(32'h3b680572),
	.w8(32'h3ab6a2c0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25baf6),
	.w1(32'h3a4e729d),
	.w2(32'hbb653f51),
	.w3(32'hbc1595c2),
	.w4(32'hba80bcd5),
	.w5(32'hbbf09ce7),
	.w6(32'hbc40cfa3),
	.w7(32'hbba4e36c),
	.w8(32'hbc339803),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8ce2a),
	.w1(32'h38651f82),
	.w2(32'hbb2b4956),
	.w3(32'hba0b41de),
	.w4(32'h3a7406ef),
	.w5(32'hba6e8213),
	.w6(32'hbac46332),
	.w7(32'h3a272c56),
	.w8(32'hbb086918),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a888591),
	.w1(32'h389a119c),
	.w2(32'hbabf95a5),
	.w3(32'h3a1c6d78),
	.w4(32'hbad31b85),
	.w5(32'hb8bd0c11),
	.w6(32'hb94380a4),
	.w7(32'h3a261f53),
	.w8(32'h3adfd3ac),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae63425),
	.w1(32'hbae6fbd0),
	.w2(32'hbb8685f8),
	.w3(32'hbb10be11),
	.w4(32'hbaab047a),
	.w5(32'hbb44e477),
	.w6(32'h39e555a9),
	.w7(32'h3a417324),
	.w8(32'hbb570450),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b37c1),
	.w1(32'h3bfed436),
	.w2(32'h3b9fecbc),
	.w3(32'hbbbe817e),
	.w4(32'h3c5262a8),
	.w5(32'hba011c1a),
	.w6(32'hbc38a927),
	.w7(32'h3c0a2621),
	.w8(32'hbc1a47aa),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb723c22),
	.w1(32'h3a3d0054),
	.w2(32'h39a967b2),
	.w3(32'hbae27aef),
	.w4(32'hb9061152),
	.w5(32'h3b05b1f8),
	.w6(32'hbbadb158),
	.w7(32'hbab7bcad),
	.w8(32'h3a9b2e75),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e9288),
	.w1(32'hb8832f5a),
	.w2(32'hbb921169),
	.w3(32'hba8fcbb7),
	.w4(32'hbb40fd92),
	.w5(32'hbba32fc2),
	.w6(32'hbb07837b),
	.w7(32'hb9b5b717),
	.w8(32'hbbceae4e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45f942),
	.w1(32'hbb2175db),
	.w2(32'hbb681a84),
	.w3(32'hbb130917),
	.w4(32'hbb0585ea),
	.w5(32'hbace383b),
	.w6(32'hba974b6b),
	.w7(32'h3afbc458),
	.w8(32'h39976f1e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8859d8),
	.w1(32'hbb076b77),
	.w2(32'hbc8b8cad),
	.w3(32'hbb194642),
	.w4(32'h3b1fb8a2),
	.w5(32'hbc47d029),
	.w6(32'hbbce4b16),
	.w7(32'h3b5e0507),
	.w8(32'hbaeaef9b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b916a),
	.w1(32'hbad11a4c),
	.w2(32'hbbbca0af),
	.w3(32'h3aabb641),
	.w4(32'h39222f94),
	.w5(32'hb9ca9d36),
	.w6(32'hbac5c370),
	.w7(32'h3b35df68),
	.w8(32'hbb026725),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb96b4),
	.w1(32'h3bf8251d),
	.w2(32'hbc4c9d96),
	.w3(32'h3b5c5b19),
	.w4(32'h3c354e78),
	.w5(32'hbc24a7cc),
	.w6(32'h3b90e60b),
	.w7(32'h3bbc0a6e),
	.w8(32'hbbc7b894),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d6002),
	.w1(32'hbb086b87),
	.w2(32'h39b34fb9),
	.w3(32'hba10b9ab),
	.w4(32'hbb03b72f),
	.w5(32'h3b5acb52),
	.w6(32'h3984ea25),
	.w7(32'hba488436),
	.w8(32'h3b134f97),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a485c73),
	.w1(32'hb90b5033),
	.w2(32'hbbf5e9f0),
	.w3(32'h3ada0625),
	.w4(32'h3ad5574d),
	.w5(32'hbc10fa2e),
	.w6(32'h3b516eaa),
	.w7(32'h3b4983ef),
	.w8(32'hbb4482c4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39317f70),
	.w1(32'hba87ad6f),
	.w2(32'h3ab21509),
	.w3(32'hbab91137),
	.w4(32'h390a964c),
	.w5(32'h3ac3918a),
	.w6(32'hb9a214e3),
	.w7(32'hbad60850),
	.w8(32'h3b71a954),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b7c47),
	.w1(32'h3a954282),
	.w2(32'hba819e67),
	.w3(32'h3b538e6c),
	.w4(32'h3add6382),
	.w5(32'h3a6028ff),
	.w6(32'h3b57b2f3),
	.w7(32'h3b706e4e),
	.w8(32'h3a5e4f8d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4244b),
	.w1(32'hbaf30e52),
	.w2(32'hba877f93),
	.w3(32'h3a2de497),
	.w4(32'hbb2dc13f),
	.w5(32'hbab679ef),
	.w6(32'h3a646776),
	.w7(32'hbb027be0),
	.w8(32'hbb33d10f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb153c8),
	.w1(32'hbafa62b2),
	.w2(32'hbc56fe1f),
	.w3(32'h39bdf789),
	.w4(32'h384eba78),
	.w5(32'hbc326334),
	.w6(32'hbb2d68ba),
	.w7(32'h39a48ece),
	.w8(32'hbbdd479e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af14e20),
	.w1(32'h3a17a67f),
	.w2(32'h3af64e7e),
	.w3(32'h3a727afe),
	.w4(32'h3a43ffbd),
	.w5(32'h3a9c5de9),
	.w6(32'h3a524ad1),
	.w7(32'h3ad87b27),
	.w8(32'h3aae6f1b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f4ce4),
	.w1(32'hb9a3147c),
	.w2(32'hbaa2e5fe),
	.w3(32'h39374402),
	.w4(32'hba1011e3),
	.w5(32'h39d437ea),
	.w6(32'h3abfec1f),
	.w7(32'hbb104345),
	.w8(32'hbb17dad9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1df3b1),
	.w1(32'hbac486d8),
	.w2(32'hbb1323c0),
	.w3(32'hbb9073af),
	.w4(32'hbb5d9257),
	.w5(32'hbb193592),
	.w6(32'hbbcd614e),
	.w7(32'hbb02ea8d),
	.w8(32'hbbccf98c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d101e),
	.w1(32'hb62688a5),
	.w2(32'hbb20d9e3),
	.w3(32'hbbe319c9),
	.w4(32'h3c4bc9d2),
	.w5(32'hba125a5d),
	.w6(32'hba6ea733),
	.w7(32'h3c6d93a1),
	.w8(32'h3bf5084a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22dbda),
	.w1(32'h3ba3b5cd),
	.w2(32'h3c910dc4),
	.w3(32'hbc1e498c),
	.w4(32'h3c2b24f6),
	.w5(32'h3cb839ea),
	.w6(32'hbb888c47),
	.w7(32'h3c50e2bf),
	.w8(32'h3b08f7fa),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba936a4f),
	.w1(32'hb9bb6f70),
	.w2(32'hbb6e64b7),
	.w3(32'hbb1d6266),
	.w4(32'hba354b5d),
	.w5(32'hbb3432f1),
	.w6(32'hbb9d4d89),
	.w7(32'hbab27cca),
	.w8(32'hbb644008),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e0f9b),
	.w1(32'h3a2a4e26),
	.w2(32'hbceaf18d),
	.w3(32'hba126018),
	.w4(32'h3b0d0dab),
	.w5(32'hbcfae098),
	.w6(32'hbc2eb968),
	.w7(32'hbb9d4e55),
	.w8(32'hbcb6f58d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73248f),
	.w1(32'hbc28108f),
	.w2(32'hbab419d4),
	.w3(32'hbbe3af31),
	.w4(32'h3b2cc7da),
	.w5(32'hbb952505),
	.w6(32'h3c13c053),
	.w7(32'h3c8589be),
	.w8(32'h3b99ebe6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b979),
	.w1(32'h3b1debed),
	.w2(32'h3ad4aa1e),
	.w3(32'hbbb2eef7),
	.w4(32'h3b8c8081),
	.w5(32'h3b644745),
	.w6(32'h3a80f481),
	.w7(32'h3be122f3),
	.w8(32'h3b3e578e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdb4de),
	.w1(32'hbaf7d2cb),
	.w2(32'hbaf8bb66),
	.w3(32'h39e81eed),
	.w4(32'hbb8550b1),
	.w5(32'h3a7e1601),
	.w6(32'hb9a4d240),
	.w7(32'hbb5ba0e4),
	.w8(32'hb9fff3ca),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3c4e8),
	.w1(32'h3b1d6286),
	.w2(32'h3ac4d6ac),
	.w3(32'hbaaf2d5c),
	.w4(32'h3b02fecf),
	.w5(32'h399b6f51),
	.w6(32'hba9a29bd),
	.w7(32'h3af3552b),
	.w8(32'h3aea8500),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3f10e),
	.w1(32'h3acebb1d),
	.w2(32'h3b0de253),
	.w3(32'h3ab01634),
	.w4(32'h3af26808),
	.w5(32'hb9803811),
	.w6(32'h39f152db),
	.w7(32'h3b1a83f2),
	.w8(32'h3aff0be3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9050ac),
	.w1(32'h3bd85b30),
	.w2(32'h3bb06198),
	.w3(32'h3b58619e),
	.w4(32'h3c554d4f),
	.w5(32'h3ba35028),
	.w6(32'h3be5c892),
	.w7(32'h3c2d79f5),
	.w8(32'hba0cd9c8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f965f),
	.w1(32'h3bc3d628),
	.w2(32'h3b05865c),
	.w3(32'h39af7462),
	.w4(32'h3bf1cec1),
	.w5(32'h3a900780),
	.w6(32'hbacad783),
	.w7(32'h3b7a37d8),
	.w8(32'hbb308833),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc289de8),
	.w1(32'hbbe1c817),
	.w2(32'hbbcbdee5),
	.w3(32'hbc3c3ce2),
	.w4(32'hbc3f8b87),
	.w5(32'hbbd2af96),
	.w6(32'hbc1b9125),
	.w7(32'hbbafdd2f),
	.w8(32'hbbc0b918),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbada3de),
	.w1(32'hbb323d22),
	.w2(32'hbb0a2e3e),
	.w3(32'hbbf33ed0),
	.w4(32'hbba23b94),
	.w5(32'hb94d9bc2),
	.w6(32'hbb85520e),
	.w7(32'hbb6dbca9),
	.w8(32'hbb69716a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20fcc4),
	.w1(32'h3a8226bd),
	.w2(32'hbc4acf68),
	.w3(32'hbb86bad6),
	.w4(32'h3c210f01),
	.w5(32'hbc15e293),
	.w6(32'hbb386f05),
	.w7(32'h3bb31074),
	.w8(32'hbba0ab65),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8caf00),
	.w1(32'hbab85fb1),
	.w2(32'h3bc9d535),
	.w3(32'hbc017fb6),
	.w4(32'hbb6cb243),
	.w5(32'h3bda2188),
	.w6(32'hbba2a6ac),
	.w7(32'hba8d5951),
	.w8(32'h3b0db9e8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75c54d),
	.w1(32'hba68a748),
	.w2(32'hbabdb1c7),
	.w3(32'hbadd5dd1),
	.w4(32'hb9af0615),
	.w5(32'hb9a5583a),
	.w6(32'hbafae9f8),
	.w7(32'h3a29f744),
	.w8(32'hb9cbe43a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcc7b6),
	.w1(32'hb98f8747),
	.w2(32'hbb467a8e),
	.w3(32'h3bc16ee5),
	.w4(32'h3b4213d5),
	.w5(32'hbb866b03),
	.w6(32'hbacd44f8),
	.w7(32'h3ad21259),
	.w8(32'hbb507937),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a1f1d),
	.w1(32'hb982daea),
	.w2(32'hba7d585f),
	.w3(32'h3a67dbb8),
	.w4(32'hbae042f8),
	.w5(32'hbb17d70b),
	.w6(32'h3a36a8e5),
	.w7(32'hbb25d03e),
	.w8(32'hbb1c512d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17068d),
	.w1(32'h3b56ed9f),
	.w2(32'hb9c536ea),
	.w3(32'hbba2f98b),
	.w4(32'h3ba1b8c2),
	.w5(32'hba359a84),
	.w6(32'hbbb5acfe),
	.w7(32'h3b3bb9a0),
	.w8(32'h3a2d8aaa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaccede),
	.w1(32'hbacc11b5),
	.w2(32'h3b99c53d),
	.w3(32'hbbd0a2bc),
	.w4(32'hbb9041ca),
	.w5(32'hb97c45b1),
	.w6(32'h3adfcc5d),
	.w7(32'h3b634e50),
	.w8(32'h3a778c4d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eca58),
	.w1(32'hbaf6486b),
	.w2(32'hbb3a5cda),
	.w3(32'hbbb3ff1b),
	.w4(32'hbaa125b5),
	.w5(32'hbb343fc7),
	.w6(32'hbb181ae5),
	.w7(32'h3b0376c4),
	.w8(32'h3a2312e4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188132),
	.w1(32'h389dc4a5),
	.w2(32'h3a09693b),
	.w3(32'hbb0015c3),
	.w4(32'hba8f2987),
	.w5(32'hbad1591b),
	.w6(32'hba4a708f),
	.w7(32'hbaba13ac),
	.w8(32'hba789d26),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934b35),
	.w1(32'hbb8047bb),
	.w2(32'hbba76fd5),
	.w3(32'hbbe7b71d),
	.w4(32'hbbc809ed),
	.w5(32'hbba79c91),
	.w6(32'hbbc0ef7d),
	.w7(32'hba5412ed),
	.w8(32'hb963bf82),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8077ad),
	.w1(32'hbac0e1b9),
	.w2(32'hbc023714),
	.w3(32'hba1f05f8),
	.w4(32'h3b943e8b),
	.w5(32'hbbcd34ee),
	.w6(32'hba9505b1),
	.w7(32'h3b57c7c2),
	.w8(32'hbb5cc10c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc664ef4),
	.w1(32'h3bb761b9),
	.w2(32'hbb8b6d67),
	.w3(32'hbc4539b2),
	.w4(32'h3b54748d),
	.w5(32'hbb658cc4),
	.w6(32'hbc4a3247),
	.w7(32'h3b06cff4),
	.w8(32'hbb93fd2d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73f797),
	.w1(32'hba1d07b5),
	.w2(32'hba35bada),
	.w3(32'h3b5f0bc8),
	.w4(32'hba1384a1),
	.w5(32'hba01c1c3),
	.w6(32'h3b7dabe4),
	.w7(32'hb92a80ca),
	.w8(32'hb94cbb39),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a7f02),
	.w1(32'h3a8f3843),
	.w2(32'hba401433),
	.w3(32'hbaa535bc),
	.w4(32'hba07e9ca),
	.w5(32'hba86df31),
	.w6(32'h3863fb6b),
	.w7(32'hb983315a),
	.w8(32'hba9af4c9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dc64c),
	.w1(32'h3be5253b),
	.w2(32'h3bb77930),
	.w3(32'hbc84e248),
	.w4(32'h3b01df4f),
	.w5(32'h3b576489),
	.w6(32'hbc7c368d),
	.w7(32'hbbf88a9a),
	.w8(32'hbc859c45),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b9bb),
	.w1(32'h3bc587d2),
	.w2(32'hbb409cba),
	.w3(32'h3b1d4207),
	.w4(32'h3bd754a8),
	.w5(32'hbbf29e99),
	.w6(32'hbbfc6355),
	.w7(32'hbaa4afbc),
	.w8(32'hbc0163f5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09c215),
	.w1(32'hbb6174be),
	.w2(32'hbbf3772a),
	.w3(32'hbc297161),
	.w4(32'hbbd5a4a2),
	.w5(32'hbb944ebc),
	.w6(32'hbbddfddf),
	.w7(32'h3afecaf0),
	.w8(32'hbb35dcee),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc988541),
	.w1(32'h3c1f14a5),
	.w2(32'hbc025f74),
	.w3(32'hba3d0328),
	.w4(32'h3cb8dd2f),
	.w5(32'hbb8ecb0c),
	.w6(32'h3ca97fce),
	.w7(32'h3cc53740),
	.w8(32'hbb482ef4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac99210),
	.w1(32'h3a5701dd),
	.w2(32'hbb4456bd),
	.w3(32'h3b8a0a6a),
	.w4(32'h3a94993d),
	.w5(32'hbb7bca34),
	.w6(32'h3b03c7ec),
	.w7(32'hbb5520e4),
	.w8(32'hbb7984c5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba38c78),
	.w1(32'h3b9a3210),
	.w2(32'hba83d411),
	.w3(32'h3b6b07fe),
	.w4(32'h3a95ca27),
	.w5(32'hbb0c13b9),
	.w6(32'hbab80c7e),
	.w7(32'hbacb3666),
	.w8(32'hbb37d808),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc965931),
	.w1(32'h3cbea9b6),
	.w2(32'h3d0fdfc8),
	.w3(32'hbcb5fdf4),
	.w4(32'h3cd7eb35),
	.w5(32'h3c8e7de2),
	.w6(32'hbc6f6788),
	.w7(32'h3cae7304),
	.w8(32'hbc5707fe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ac7ba),
	.w1(32'h3bb8cc95),
	.w2(32'hbc9b3553),
	.w3(32'hbad9f38a),
	.w4(32'h3bef12ea),
	.w5(32'hbc884fb6),
	.w6(32'hbc1c4d9e),
	.w7(32'hbae6e499),
	.w8(32'hbc562f45),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8afc06),
	.w1(32'h3b62360e),
	.w2(32'h3b21f98d),
	.w3(32'hbb00fa68),
	.w4(32'h3c673323),
	.w5(32'h3b85a104),
	.w6(32'h3baf9496),
	.w7(32'h3c6cf2a4),
	.w8(32'h38ae74a4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f3f82),
	.w1(32'h3c00485a),
	.w2(32'h3b9de760),
	.w3(32'hbbd1df93),
	.w4(32'h3a178dff),
	.w5(32'h39cae1d6),
	.w6(32'h3a95edc1),
	.w7(32'h3bd817f8),
	.w8(32'hbb39265a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08a02b),
	.w1(32'hbb6e53c9),
	.w2(32'hbb936520),
	.w3(32'hbc04366f),
	.w4(32'hbbc1901a),
	.w5(32'hbc02cc13),
	.w6(32'hbb07b29b),
	.w7(32'h3b31e5f6),
	.w8(32'hbba88b17),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a283e10),
	.w1(32'h39801796),
	.w2(32'h3a68b697),
	.w3(32'h3a3bc3e5),
	.w4(32'h39946b8d),
	.w5(32'h3a805251),
	.w6(32'h3a1e7464),
	.w7(32'h3af75d52),
	.w8(32'h3b0ea6b7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9fa00),
	.w1(32'hbad6e7e5),
	.w2(32'h3a235244),
	.w3(32'h3b675435),
	.w4(32'hbae9c257),
	.w5(32'hbb1ba59d),
	.w6(32'h3b60bb7e),
	.w7(32'hbb167493),
	.w8(32'hbacf597b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb838b69),
	.w1(32'hba9fe055),
	.w2(32'hbb8e9fc6),
	.w3(32'hbb23ca47),
	.w4(32'h3a49c78e),
	.w5(32'hbbba708d),
	.w6(32'hbb21f5d7),
	.w7(32'hbbe62c31),
	.w8(32'hbbf01875),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac190bc),
	.w1(32'h3a8114d8),
	.w2(32'h3afde10a),
	.w3(32'hbb0fa6f9),
	.w4(32'h3ae094b4),
	.w5(32'h3a8ad288),
	.w6(32'hbb0a1509),
	.w7(32'h3afdada0),
	.w8(32'h3a8399bb),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a28c),
	.w1(32'h3b688ca6),
	.w2(32'h39bae2ef),
	.w3(32'h3a9a1ea3),
	.w4(32'h3b994342),
	.w5(32'h3a9a9897),
	.w6(32'hbb550d4c),
	.w7(32'h3b44f7ee),
	.w8(32'hbb3845fc),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f920d),
	.w1(32'h3c6747f4),
	.w2(32'h3a85e77b),
	.w3(32'h3b4e84ec),
	.w4(32'h3c2a8ff8),
	.w5(32'hbc33d53a),
	.w6(32'hbbe13779),
	.w7(32'hbb2d1f14),
	.w8(32'hbc1555b9),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab363bb),
	.w1(32'hbaace45b),
	.w2(32'hbb8f50f2),
	.w3(32'hbb15a623),
	.w4(32'hbaee1841),
	.w5(32'hbb8e8d7c),
	.w6(32'hbaa05117),
	.w7(32'h398987e8),
	.w8(32'hbb1f9b07),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f1a45),
	.w1(32'hbae1a5bd),
	.w2(32'hbaed2647),
	.w3(32'hba5303f4),
	.w4(32'hbac5f708),
	.w5(32'hbb3b6161),
	.w6(32'hba831083),
	.w7(32'hba3886d2),
	.w8(32'hbb06e319),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc366490),
	.w1(32'h3c1a71bd),
	.w2(32'h3be8241a),
	.w3(32'hbc331fbe),
	.w4(32'h3c9de081),
	.w5(32'h3b9695fa),
	.w6(32'hb9b0c3fd),
	.w7(32'h3c9023ce),
	.w8(32'hbbee2bce),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4942f7),
	.w1(32'h3b502935),
	.w2(32'hbba19f4e),
	.w3(32'h3b5037ed),
	.w4(32'h3baffbeb),
	.w5(32'hbb75e474),
	.w6(32'h3ab95732),
	.w7(32'h3b4eef66),
	.w8(32'hbb9edf2e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad96156),
	.w1(32'hba2c9c35),
	.w2(32'hbad468ba),
	.w3(32'hb895e52e),
	.w4(32'hbabf00da),
	.w5(32'hba3c4398),
	.w6(32'h3960760e),
	.w7(32'hbacd9fbd),
	.w8(32'hbb08637c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7888d1),
	.w1(32'h3bb4d3e9),
	.w2(32'hbb7dee77),
	.w3(32'h3a3d1aa4),
	.w4(32'h3c0da992),
	.w5(32'hba24eaec),
	.w6(32'hba193052),
	.w7(32'h3bbc150f),
	.w8(32'hbb8a47ad),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5baf5),
	.w1(32'h380881e2),
	.w2(32'hb863546d),
	.w3(32'hb9e3914c),
	.w4(32'hba6a0111),
	.w5(32'hba1af657),
	.w6(32'hb9cb9e72),
	.w7(32'hba4b5ec5),
	.w8(32'hba4ecf1f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91a415),
	.w1(32'hb98cc381),
	.w2(32'hbb0f1d45),
	.w3(32'hbacbacd9),
	.w4(32'h38b72e0c),
	.w5(32'hbb0a124c),
	.w6(32'hbaebf574),
	.w7(32'hb9d88c2c),
	.w8(32'hbb4eb389),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de2397),
	.w1(32'h39b178d0),
	.w2(32'h3a5fb83a),
	.w3(32'hba967c80),
	.w4(32'h3a5e1a48),
	.w5(32'h3ab3cceb),
	.w6(32'hbb00a8c7),
	.w7(32'h3a9e52f6),
	.w8(32'h3a8e409d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d33059),
	.w1(32'hba995d5e),
	.w2(32'hbaa4c7c7),
	.w3(32'h3abbe4e1),
	.w4(32'hbb1b9176),
	.w5(32'hbb78c21e),
	.w6(32'h3a61ce11),
	.w7(32'hba6cec64),
	.w8(32'hbb87cd0a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dcb7c),
	.w1(32'h3a89ce9a),
	.w2(32'h3b3c6b6e),
	.w3(32'hbba509d0),
	.w4(32'hbab53410),
	.w5(32'h3af42aa1),
	.w6(32'hbbaac148),
	.w7(32'hba0aef72),
	.w8(32'h39d91cb4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53a5fb),
	.w1(32'hbb3453ce),
	.w2(32'hbcc8d524),
	.w3(32'h3b721409),
	.w4(32'h3c327ddb),
	.w5(32'hbc50c4f0),
	.w6(32'h3c723f59),
	.w7(32'h3c78ce73),
	.w8(32'hba279b10),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8208b6),
	.w1(32'h3b95b2c4),
	.w2(32'hbc2dcfa3),
	.w3(32'h3a280c3e),
	.w4(32'h3bf781f2),
	.w5(32'hbb9a340d),
	.w6(32'h3a8ba8c8),
	.w7(32'h3b5059ac),
	.w8(32'hbba4f922),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc566626),
	.w1(32'hb9997623),
	.w2(32'hbc9c6327),
	.w3(32'h399a8dac),
	.w4(32'h3bc5237f),
	.w5(32'hbc7db7d7),
	.w6(32'h3b9d699d),
	.w7(32'h3b3b0cc4),
	.w8(32'hbc059a27),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44e79c),
	.w1(32'h3b097a82),
	.w2(32'h3ae7bd4d),
	.w3(32'hba955ecd),
	.w4(32'h3a16fb42),
	.w5(32'h3aa52db6),
	.w6(32'hba8a9c2c),
	.w7(32'h3a0390a7),
	.w8(32'h39430b38),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaffe0),
	.w1(32'hba995293),
	.w2(32'hbb2bb118),
	.w3(32'h3aac67b4),
	.w4(32'h39ed59e2),
	.w5(32'hba76c669),
	.w6(32'hbabee055),
	.w7(32'hba2682fe),
	.w8(32'hbade1ac6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb115254),
	.w1(32'h3a1066ef),
	.w2(32'h3af6fd18),
	.w3(32'hbab78a10),
	.w4(32'h3a22cb79),
	.w5(32'hb9c1157f),
	.w6(32'hba67bf84),
	.w7(32'hb9a93e91),
	.w8(32'hb917c01f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11c167),
	.w1(32'h3a22eae0),
	.w2(32'hba7412e6),
	.w3(32'h3a2a7629),
	.w4(32'h3a17bc97),
	.w5(32'h381a75fd),
	.w6(32'h39dd00f5),
	.w7(32'h3a3026d3),
	.w8(32'hba33378b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8a03a),
	.w1(32'hbab3865e),
	.w2(32'hbc93c482),
	.w3(32'h3bc1362b),
	.w4(32'hbb42ed7d),
	.w5(32'hbc5eeb14),
	.w6(32'h3ac177ff),
	.w7(32'hbc098dc3),
	.w8(32'hbc129ab6),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2a4fd),
	.w1(32'h383ac00f),
	.w2(32'h36886b68),
	.w3(32'hbaee1323),
	.w4(32'h3a18b6d4),
	.w5(32'h3a08647d),
	.w6(32'hbb283b19),
	.w7(32'h3a303dcf),
	.w8(32'h3a2bb76b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa860c),
	.w1(32'h3b30a565),
	.w2(32'h3b3e6876),
	.w3(32'hbb0db362),
	.w4(32'h3a231de1),
	.w5(32'h3aeaea35),
	.w6(32'hbb5b4072),
	.w7(32'h3a29f0f1),
	.w8(32'h3b1ebb80),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fcae0),
	.w1(32'h3abb2727),
	.w2(32'h3b834b1e),
	.w3(32'h3a678533),
	.w4(32'h3ab1a48b),
	.w5(32'h3ae83450),
	.w6(32'hbaf1d6d2),
	.w7(32'h388de64c),
	.w8(32'h3adf06ed),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c7005),
	.w1(32'hb9ee5ab4),
	.w2(32'hbaa49479),
	.w3(32'h3a377999),
	.w4(32'hb9a07a18),
	.w5(32'hb92e3742),
	.w6(32'h3af7ecf9),
	.w7(32'hba3273a9),
	.w8(32'hba3a16e4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae08877),
	.w1(32'h3b16d2d5),
	.w2(32'hbb0377dc),
	.w3(32'hba1d1738),
	.w4(32'h3b3e15fc),
	.w5(32'hbac5261d),
	.w6(32'hba4667af),
	.w7(32'h3b1f1205),
	.w8(32'hba281511),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c251a),
	.w1(32'hba985fe8),
	.w2(32'hbb0b303b),
	.w3(32'h3af224ee),
	.w4(32'h3a7a841a),
	.w5(32'hba19679b),
	.w6(32'h3b51a71b),
	.w7(32'h3a979a66),
	.w8(32'hb906d380),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc290c86),
	.w1(32'hbc14fc8f),
	.w2(32'hbd0d6b52),
	.w3(32'h3c30e257),
	.w4(32'h3b9de5eb),
	.w5(32'hbcf07e52),
	.w6(32'h3ba0c44d),
	.w7(32'hbb79931a),
	.w8(32'hbc36a61d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba893c19),
	.w1(32'hb9c003be),
	.w2(32'hba8e4f80),
	.w3(32'hba983c59),
	.w4(32'hba957064),
	.w5(32'hbabc14a6),
	.w6(32'hbb058e8d),
	.w7(32'hbacdff06),
	.w8(32'hba10a89d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030b15),
	.w1(32'h3c209d43),
	.w2(32'h3c1d9ba7),
	.w3(32'hbc53b85c),
	.w4(32'h3b4b5291),
	.w5(32'h3beb8184),
	.w6(32'hbbf0711b),
	.w7(32'hbaf80435),
	.w8(32'hbb633f98),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule