module layer_8_featuremap_33(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b746d6a),
	.w1(32'h3ba06205),
	.w2(32'h3b8db27f),
	.w3(32'h3b714f28),
	.w4(32'h3ba1145f),
	.w5(32'h3b87efdb),
	.w6(32'h3ae2bd06),
	.w7(32'h3a9cb247),
	.w8(32'h3b0453f6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f859c),
	.w1(32'hbb0e1b32),
	.w2(32'hbb2289a1),
	.w3(32'hbb34d6dc),
	.w4(32'hbb3fe3c0),
	.w5(32'hbb4e7da2),
	.w6(32'hbb63dac6),
	.w7(32'hbb6911f2),
	.w8(32'hbb4a50aa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b66de),
	.w1(32'hbb061e2e),
	.w2(32'hbae5fb18),
	.w3(32'hbb2daf45),
	.w4(32'hbb41d89a),
	.w5(32'hbb1c3168),
	.w6(32'hbb55c7b0),
	.w7(32'hbb54f3dc),
	.w8(32'hbb11ef7d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a7a63),
	.w1(32'h3b451a90),
	.w2(32'h3b38f1ce),
	.w3(32'h3adc823f),
	.w4(32'h3b19e177),
	.w5(32'h3b266c3c),
	.w6(32'h3b2e4375),
	.w7(32'h3b4c0a52),
	.w8(32'h3b3b9531),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad70f81),
	.w1(32'hbad14978),
	.w2(32'hb9c3e732),
	.w3(32'hbaee019e),
	.w4(32'hbadfbfef),
	.w5(32'hba1f47f2),
	.w6(32'hbb647f77),
	.w7(32'hbb2c4b68),
	.w8(32'hbaf5d81a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb829aaa),
	.w1(32'hbb8b1d56),
	.w2(32'hbb5e66c6),
	.w3(32'hbb61c208),
	.w4(32'hbb0e5555),
	.w5(32'hba813228),
	.w6(32'hbaffe7a1),
	.w7(32'hb9210e60),
	.w8(32'hbb0e8e6d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914c802),
	.w1(32'h3900129d),
	.w2(32'h380f0ea8),
	.w3(32'hb2ae0afa),
	.w4(32'h38d0aa52),
	.w5(32'hb66e1707),
	.w6(32'h382d1c35),
	.w7(32'h37c368af),
	.w8(32'h35261a4b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0927d5),
	.w1(32'hbb222307),
	.w2(32'hbabdaabe),
	.w3(32'hbaf582e7),
	.w4(32'hbb181af1),
	.w5(32'hbaf55baa),
	.w6(32'hbba4ff74),
	.w7(32'hbb88e4ff),
	.w8(32'hbb62614b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba982f72),
	.w1(32'hbaeb4bae),
	.w2(32'hba9e0db1),
	.w3(32'hbb3594a9),
	.w4(32'hbb370146),
	.w5(32'hba94da77),
	.w6(32'hbb745a17),
	.w7(32'hbb1e3287),
	.w8(32'hba733393),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49048c),
	.w1(32'h3a269e57),
	.w2(32'hba52fef0),
	.w3(32'hbac67575),
	.w4(32'hba50f443),
	.w5(32'hba772967),
	.w6(32'hbb87345a),
	.w7(32'hbb794155),
	.w8(32'hbb4f6bc3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7840ce),
	.w1(32'h3ba3e221),
	.w2(32'h3b772f37),
	.w3(32'h3b2deecc),
	.w4(32'h3b84b5e2),
	.w5(32'h3b0c7fce),
	.w6(32'h3a55117a),
	.w7(32'h3aba0e15),
	.w8(32'hb634b4e0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eda35),
	.w1(32'hbaa59897),
	.w2(32'hba9f7c9c),
	.w3(32'hb9052b20),
	.w4(32'h3aa79562),
	.w5(32'h3a02b12c),
	.w6(32'hbb1785a9),
	.w7(32'hbaa702dc),
	.w8(32'hba28861d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb578a35),
	.w1(32'hbb4da5de),
	.w2(32'hbb810941),
	.w3(32'hbb6f3f86),
	.w4(32'hbb2e3b10),
	.w5(32'hbb381ef3),
	.w6(32'hbb9bfa8d),
	.w7(32'hbb848a8c),
	.w8(32'hbb7e1b65),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ff69af),
	.w1(32'hb8051123),
	.w2(32'hb8f7d023),
	.w3(32'hb9d326dd),
	.w4(32'hb96a81e6),
	.w5(32'hb8a41251),
	.w6(32'hb95a3199),
	.w7(32'hb9fa2eff),
	.w8(32'hb8a61202),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a8c4de),
	.w1(32'hb78712e1),
	.w2(32'hb80f39c5),
	.w3(32'hb83db229),
	.w4(32'hb7f798fa),
	.w5(32'hb8282944),
	.w6(32'hb8039bf6),
	.w7(32'hb85ae5e4),
	.w8(32'hb7fe1aab),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e15ec1),
	.w1(32'hb553e119),
	.w2(32'h39795dfb),
	.w3(32'hb8882968),
	.w4(32'hb934119c),
	.w5(32'h38eea0ac),
	.w6(32'hb93e7b9c),
	.w7(32'hb8358190),
	.w8(32'h393e17a4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39113d51),
	.w1(32'h3a644689),
	.w2(32'h3a0f9f04),
	.w3(32'h3a864616),
	.w4(32'h3ac02149),
	.w5(32'h3a580111),
	.w6(32'h3a5fc16d),
	.w7(32'h3ab4752c),
	.w8(32'h3a328496),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb802638b),
	.w1(32'hb9bd4ed4),
	.w2(32'hba9a60c9),
	.w3(32'hba2a0f68),
	.w4(32'hba50960c),
	.w5(32'hbacb3aab),
	.w6(32'hbb264ce0),
	.w7(32'hbb44868a),
	.w8(32'hbb0eb773),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb858c1),
	.w1(32'h3c140aa2),
	.w2(32'h3bfd3c16),
	.w3(32'h3c1280bf),
	.w4(32'h3c35b53a),
	.w5(32'h3be59382),
	.w6(32'hb94b40a8),
	.w7(32'hbb58cebc),
	.w8(32'hbb9934e7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e06d4),
	.w1(32'h3b8c20db),
	.w2(32'h3b78b193),
	.w3(32'h3a89095a),
	.w4(32'h39f093ce),
	.w5(32'hb982c968),
	.w6(32'hbb00dd81),
	.w7(32'hbb0da163),
	.w8(32'hbad3a7b2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cc70e),
	.w1(32'hb9a67a7e),
	.w2(32'hbace3308),
	.w3(32'hbac01b03),
	.w4(32'h3b4c7513),
	.w5(32'h380bb326),
	.w6(32'h39364b62),
	.w7(32'h3b015552),
	.w8(32'hbabfa502),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941354),
	.w1(32'hbb8a0e38),
	.w2(32'hbbc006f9),
	.w3(32'hbbe0fec9),
	.w4(32'hbbff8daa),
	.w5(32'hbc0cb639),
	.w6(32'hbbb4fecd),
	.w7(32'hbbff0a60),
	.w8(32'hbc12a8a3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b22b7),
	.w1(32'h3c17e60e),
	.w2(32'h3bf343f5),
	.w3(32'h3b8b3fa4),
	.w4(32'h3bfe8ec3),
	.w5(32'h3c024629),
	.w6(32'h39eb245b),
	.w7(32'h3b7c3ab5),
	.w8(32'h3b93ccb3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca1173),
	.w1(32'h3a191388),
	.w2(32'h3a2737ee),
	.w3(32'hba9ebcf2),
	.w4(32'hbadad23b),
	.w5(32'hbb039bc1),
	.w6(32'hba6498d9),
	.w7(32'hba92c0e2),
	.w8(32'hb8d8ac14),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc2e8),
	.w1(32'hb9d08788),
	.w2(32'h39a2f507),
	.w3(32'h397e0b68),
	.w4(32'hb9edc17d),
	.w5(32'hb9862670),
	.w6(32'hb91e0d77),
	.w7(32'hb9263a2c),
	.w8(32'h3a880839),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ea3b1),
	.w1(32'h3a8872b8),
	.w2(32'h39d6f3e5),
	.w3(32'h39aa7f4e),
	.w4(32'h3b14d38e),
	.w5(32'h3b2e97c7),
	.w6(32'hba1a7b6e),
	.w7(32'h39269866),
	.w8(32'h3a1672a7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f7248),
	.w1(32'h38185c6f),
	.w2(32'h3836f066),
	.w3(32'h3982596c),
	.w4(32'h399275b9),
	.w5(32'h39389f42),
	.w6(32'h3959f8b2),
	.w7(32'h39521337),
	.w8(32'h3922e79f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5393d),
	.w1(32'h3c6bea9c),
	.w2(32'h3c5393e9),
	.w3(32'h3a66f027),
	.w4(32'h3c1455e2),
	.w5(32'h3c9216ef),
	.w6(32'hbbc78d59),
	.w7(32'h3bb612af),
	.w8(32'hbbf312f6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e1c3c),
	.w1(32'h3a9072bc),
	.w2(32'h39e96e90),
	.w3(32'h3861af42),
	.w4(32'h3af86440),
	.w5(32'h3a7fe41e),
	.w6(32'hba2e6309),
	.w7(32'h3a291769),
	.w8(32'h3a45296f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba616483),
	.w1(32'hba3b80fa),
	.w2(32'hba3a59e0),
	.w3(32'hba7ddcdd),
	.w4(32'hba61d47c),
	.w5(32'hba78508a),
	.w6(32'hba849fcc),
	.w7(32'hba512358),
	.w8(32'hba9f8883),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a65c56),
	.w1(32'h3a1121bb),
	.w2(32'hba762600),
	.w3(32'h3aadd775),
	.w4(32'h3aaf279f),
	.w5(32'hb8dbf6ab),
	.w6(32'h3a0d3507),
	.w7(32'h3888f7dc),
	.w8(32'hba052fd6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d3e53),
	.w1(32'hbb2b0d5d),
	.w2(32'hbb06ae53),
	.w3(32'hbb419c46),
	.w4(32'hbb2b3776),
	.w5(32'hbabcb9db),
	.w6(32'hbb41f6c3),
	.w7(32'hbb1b50c3),
	.w8(32'hbb2a3e81),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901d74a),
	.w1(32'h38de0c12),
	.w2(32'h38c5e613),
	.w3(32'h3817328d),
	.w4(32'h3717f1bd),
	.w5(32'h379d3870),
	.w6(32'h384e1b4a),
	.w7(32'h3815f69f),
	.w8(32'h38531dc2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea8c44),
	.w1(32'h37aa6bf6),
	.w2(32'h37c835b8),
	.w3(32'hb7297ef9),
	.w4(32'hb805b9c6),
	.w5(32'hb7f5b49f),
	.w6(32'h381add7e),
	.w7(32'h373180f7),
	.w8(32'h37866a9c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b44a),
	.w1(32'hbb4f07bf),
	.w2(32'hbb3a0c78),
	.w3(32'hbb15fb53),
	.w4(32'hbb6404c0),
	.w5(32'hbb613f5c),
	.w6(32'hbb37d61c),
	.w7(32'hbb78e8de),
	.w8(32'hbb87646b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0256cb),
	.w1(32'h3b10ab36),
	.w2(32'h39472178),
	.w3(32'h3b63f0d0),
	.w4(32'h3b52eae0),
	.w5(32'h39d3ccb6),
	.w6(32'h3a13bb5f),
	.w7(32'hb9804a9f),
	.w8(32'hbb042037),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e9a5ce),
	.w1(32'hb976f4e7),
	.w2(32'h390ee915),
	.w3(32'hb76ca7e6),
	.w4(32'hb9565502),
	.w5(32'h3955635f),
	.w6(32'hb64e3fd5),
	.w7(32'hb8bfcb3f),
	.w8(32'h397b5aa4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1e5a4),
	.w1(32'hbad0b6b3),
	.w2(32'hba894a8c),
	.w3(32'hbb161350),
	.w4(32'hbb07cc48),
	.w5(32'hbad03cd3),
	.w6(32'hbb245d71),
	.w7(32'hbb008147),
	.w8(32'hbab9965b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a06b46),
	.w1(32'h3902a73e),
	.w2(32'h38ec8ba3),
	.w3(32'h383ac88b),
	.w4(32'hb9186b1c),
	.w5(32'hb95d820f),
	.w6(32'hb930f8b0),
	.w7(32'hb90e9970),
	.w8(32'hb9a26ca0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb808bf6c),
	.w1(32'h37f382e5),
	.w2(32'hb8c21d3f),
	.w3(32'hb921d370),
	.w4(32'hb9438c3a),
	.w5(32'hb9c1049a),
	.w6(32'h39452190),
	.w7(32'h382fd4dd),
	.w8(32'hb935d87c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca22a0),
	.w1(32'hbb9c82dd),
	.w2(32'hbb599f44),
	.w3(32'hbaa80266),
	.w4(32'h39e6829d),
	.w5(32'h3b3460d4),
	.w6(32'hba8bf285),
	.w7(32'h379582c4),
	.w8(32'h3b8fa14b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd12e9),
	.w1(32'hb78f353f),
	.w2(32'h3b005b44),
	.w3(32'h3958f987),
	.w4(32'h39367649),
	.w5(32'hbacff7ac),
	.w6(32'hba909693),
	.w7(32'hba76102b),
	.w8(32'hbb8586f3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97ac46),
	.w1(32'hbb2a7920),
	.w2(32'h3b19e51a),
	.w3(32'h3a207562),
	.w4(32'hbab394c6),
	.w5(32'h3b5e5747),
	.w6(32'hbabfc757),
	.w7(32'hbb6b20f6),
	.w8(32'hba2a68ea),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0496c7),
	.w1(32'h3acbdc8a),
	.w2(32'h3b01ebcb),
	.w3(32'h3aa4074b),
	.w4(32'h3b334914),
	.w5(32'h39955f55),
	.w6(32'h3ac0aa5a),
	.w7(32'h3af710c8),
	.w8(32'h3a75cdd6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948ba59),
	.w1(32'h3b7df041),
	.w2(32'h3b7d88de),
	.w3(32'h3b2e60d3),
	.w4(32'h3b973c41),
	.w5(32'h3ad4324a),
	.w6(32'hbb00e495),
	.w7(32'hba931cde),
	.w8(32'hbb902f80),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa110ac),
	.w1(32'h3b02d609),
	.w2(32'hba19e945),
	.w3(32'h3b038ec1),
	.w4(32'h3ad76c73),
	.w5(32'h3818aa69),
	.w6(32'hba8db395),
	.w7(32'hba7affaf),
	.w8(32'hbc708eb9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c669d),
	.w1(32'h3b75c186),
	.w2(32'hbb65a4f4),
	.w3(32'h3ac11f6a),
	.w4(32'hbaffe383),
	.w5(32'h3a337004),
	.w6(32'hbbe64e2b),
	.w7(32'hbb20d595),
	.w8(32'hba24d027),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb572e51),
	.w1(32'hbadc89c2),
	.w2(32'h3ba5e0b7),
	.w3(32'hba901c80),
	.w4(32'h3aebd4ba),
	.w5(32'h3b47ea2b),
	.w6(32'hbb8ee2f7),
	.w7(32'hbb482e4c),
	.w8(32'hbb3e231b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa599b4),
	.w1(32'hb8e2b606),
	.w2(32'hb9a894f8),
	.w3(32'h3ad05b68),
	.w4(32'h3af4670b),
	.w5(32'h3ba579af),
	.w6(32'h3a50754c),
	.w7(32'h3ac6a59c),
	.w8(32'hb9caee2c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bc865),
	.w1(32'h3a99ead6),
	.w2(32'h3ae61808),
	.w3(32'hba22e3b9),
	.w4(32'h3ad6c2c6),
	.w5(32'h3b08c78d),
	.w6(32'h3919c79f),
	.w7(32'h3b275546),
	.w8(32'h3a18ec1f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3823b2),
	.w1(32'hbc52e549),
	.w2(32'hbc35e3b1),
	.w3(32'hbc34f392),
	.w4(32'hbc391411),
	.w5(32'hbc2174f4),
	.w6(32'hbc340c26),
	.w7(32'hbc1941dc),
	.w8(32'hbbeb7e14),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be9b7),
	.w1(32'hb846aaef),
	.w2(32'h3b8d36d7),
	.w3(32'h3b4652eb),
	.w4(32'h3b99b9eb),
	.w5(32'h3b4c1fdf),
	.w6(32'hbb05e407),
	.w7(32'hba7ae480),
	.w8(32'hba9230a0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc87703),
	.w1(32'h3a9219b0),
	.w2(32'h397a6c48),
	.w3(32'h3a62fbbe),
	.w4(32'hbb037cf0),
	.w5(32'h3a9ffb97),
	.w6(32'hbafe9ff6),
	.w7(32'hb8bd322e),
	.w8(32'h3a833464),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c76eaa),
	.w1(32'h3b01df56),
	.w2(32'h395e32ba),
	.w3(32'hb9cfdb37),
	.w4(32'h398cce44),
	.w5(32'h3a6b0996),
	.w6(32'hbab545d1),
	.w7(32'hbb27ab7f),
	.w8(32'hbc109bbb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bee67),
	.w1(32'h3890124c),
	.w2(32'hbb321312),
	.w3(32'hbb55efec),
	.w4(32'h3b3245e8),
	.w5(32'h3b69f36a),
	.w6(32'h3b16ea2e),
	.w7(32'hbbc15a80),
	.w8(32'h378393ff),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1819e),
	.w1(32'h3a4bee28),
	.w2(32'hbb91142a),
	.w3(32'h3abb08f4),
	.w4(32'h3b16b624),
	.w5(32'hba7433c7),
	.w6(32'hbbc94af2),
	.w7(32'hbbbc8cf0),
	.w8(32'hbb0bc7da),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33c2ea),
	.w1(32'h3bc769cc),
	.w2(32'hbb401540),
	.w3(32'h3abeba53),
	.w4(32'hb9d7e37a),
	.w5(32'hbb4033ee),
	.w6(32'h3b1fcd5a),
	.w7(32'h3aeeecfa),
	.w8(32'hbaa71355),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd13a21),
	.w1(32'hbb0ecd9b),
	.w2(32'h3af5875f),
	.w3(32'h3b0d1c91),
	.w4(32'h3b8bc681),
	.w5(32'h3b693adb),
	.w6(32'hbb9a6ee0),
	.w7(32'hbbf30e13),
	.w8(32'h3a2bf631),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b505201),
	.w1(32'h3b1fedc0),
	.w2(32'h3b79d8a8),
	.w3(32'h3b6bda8d),
	.w4(32'h3b9baa50),
	.w5(32'h3b3d0ee3),
	.w6(32'h3b4612b0),
	.w7(32'h3b90311a),
	.w8(32'hbac7a84f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84810c),
	.w1(32'h3af28d19),
	.w2(32'hbb039355),
	.w3(32'hbb7bbf4a),
	.w4(32'hbab672ba),
	.w5(32'hb9e4ed08),
	.w6(32'hbaaa2cf7),
	.w7(32'hbb0bcd67),
	.w8(32'h3af994da),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d3c1b),
	.w1(32'h3b6e89a0),
	.w2(32'h3ba1af03),
	.w3(32'h3b3e387b),
	.w4(32'h3bab9eb0),
	.w5(32'hba64505c),
	.w6(32'hbc2f6690),
	.w7(32'h3a824ecd),
	.w8(32'hbb0efbfa),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b39df),
	.w1(32'hbb39a260),
	.w2(32'hba90558c),
	.w3(32'hbae00bba),
	.w4(32'hba753ecf),
	.w5(32'h39f41323),
	.w6(32'hbaf47a64),
	.w7(32'hba92d76f),
	.w8(32'h3b1eee53),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb6a4),
	.w1(32'hbb8618df),
	.w2(32'hbb4d1425),
	.w3(32'h3b63d230),
	.w4(32'h3b018b33),
	.w5(32'hba2aa827),
	.w6(32'hbb10526b),
	.w7(32'h39614213),
	.w8(32'hb9e2fbae),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb815d0),
	.w1(32'h3a2f37d2),
	.w2(32'h3ae245cf),
	.w3(32'hbbb74cf5),
	.w4(32'hbbaa3507),
	.w5(32'hbb18adcf),
	.w6(32'h3b923031),
	.w7(32'hbba4c48a),
	.w8(32'h39e22297),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a071454),
	.w1(32'h3a9627dd),
	.w2(32'h3a9fb095),
	.w3(32'h3ae7c182),
	.w4(32'h3b1c287e),
	.w5(32'h37ecc86e),
	.w6(32'h3ab9e14e),
	.w7(32'h3b1aaccd),
	.w8(32'h3a825c8e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01ad4a),
	.w1(32'hb87591ac),
	.w2(32'hba449f38),
	.w3(32'h39c9fcf1),
	.w4(32'h39b47abb),
	.w5(32'hba98df2e),
	.w6(32'hbb1be178),
	.w7(32'hbadf4312),
	.w8(32'hbade935e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad78f4),
	.w1(32'hbba812aa),
	.w2(32'hbb756f5d),
	.w3(32'hbb764dc5),
	.w4(32'hbb7eb294),
	.w5(32'hbb791250),
	.w6(32'hbb918315),
	.w7(32'hbb5c5797),
	.w8(32'hbb41b85d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc04a28),
	.w1(32'hbbc780c6),
	.w2(32'hbb7e2824),
	.w3(32'hbbe59401),
	.w4(32'hbb72a4e2),
	.w5(32'hba0aaa71),
	.w6(32'hbbc5b13c),
	.w7(32'hbc1ba773),
	.w8(32'hbad73aab),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f463ea),
	.w1(32'hb9b1e71a),
	.w2(32'h3a813e4b),
	.w3(32'hb8dc763f),
	.w4(32'h3a280019),
	.w5(32'h3a4f40f5),
	.w6(32'hba419d8a),
	.w7(32'h3a5a58c4),
	.w8(32'h3bbc71dc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6af0b),
	.w1(32'h3c184b95),
	.w2(32'h3c407862),
	.w3(32'h3c0e542d),
	.w4(32'h3c5001d5),
	.w5(32'h3b963d43),
	.w6(32'h3bf47065),
	.w7(32'h3c0a8504),
	.w8(32'h3ac21302),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7a7bf),
	.w1(32'h38ec5778),
	.w2(32'h3a97f3f0),
	.w3(32'h3a58670f),
	.w4(32'h3aa7048c),
	.w5(32'hb9f7ed63),
	.w6(32'h38e6deed),
	.w7(32'h3ac1eb62),
	.w8(32'h39a913e1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ca12e),
	.w1(32'hbb04a3bb),
	.w2(32'h393b41bb),
	.w3(32'hbb586a28),
	.w4(32'hbab2221c),
	.w5(32'hb9de9c05),
	.w6(32'hbb9c4b75),
	.w7(32'hbb1f70d0),
	.w8(32'hbac755e3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3380c),
	.w1(32'h38feaa81),
	.w2(32'h3a46eece),
	.w3(32'h3ae8f477),
	.w4(32'h3a979fd6),
	.w5(32'hba641a3f),
	.w6(32'hb9e14fe7),
	.w7(32'h3a93d0ad),
	.w8(32'hbaf8cde2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd40853),
	.w1(32'hbb229ef5),
	.w2(32'hbb0a6c2c),
	.w3(32'hbc4c8850),
	.w4(32'hbb79b23a),
	.w5(32'h3b1bd42f),
	.w6(32'hbb2f8c88),
	.w7(32'hbc0780e2),
	.w8(32'hbb4dd4c1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74d87f),
	.w1(32'hb9ef81b9),
	.w2(32'hb86b8906),
	.w3(32'hba8d5071),
	.w4(32'h39856391),
	.w5(32'hbb06f5ad),
	.w6(32'hba696fb7),
	.w7(32'hbad27237),
	.w8(32'h3953ef80),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26dbf9),
	.w1(32'hbad40073),
	.w2(32'hb929bd3f),
	.w3(32'hbae7b877),
	.w4(32'h39903ed4),
	.w5(32'hba811945),
	.w6(32'hbb39f9e2),
	.w7(32'h37d125db),
	.w8(32'hb9a4cccc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c1b65f),
	.w1(32'hb9a6215b),
	.w2(32'h39a34e06),
	.w3(32'h321bf215),
	.w4(32'h3a2afd96),
	.w5(32'hba4aad25),
	.w6(32'hba0aef1f),
	.w7(32'h38b71d3d),
	.w8(32'h3bcbbeab),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8a4d1),
	.w1(32'h3ac1222f),
	.w2(32'h3b1bef9b),
	.w3(32'h3ba106c1),
	.w4(32'h3b9fc388),
	.w5(32'hbabc32ac),
	.w6(32'h3b0513c2),
	.w7(32'h3b7732ba),
	.w8(32'h3b86d167),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e9b55),
	.w1(32'h395ceb8f),
	.w2(32'h3a9fb11f),
	.w3(32'h3b3ebf7e),
	.w4(32'h3b0d80c2),
	.w5(32'hbacda1d8),
	.w6(32'hbaa19d39),
	.w7(32'hb97d2401),
	.w8(32'hbada029c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6426f),
	.w1(32'h397ce241),
	.w2(32'h398a3fbe),
	.w3(32'hbac0af27),
	.w4(32'h38fd2245),
	.w5(32'hba1b0675),
	.w6(32'hba795c12),
	.w7(32'hbad5f9ce),
	.w8(32'hb9d64792),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd4cb5),
	.w1(32'hbc0b5363),
	.w2(32'hbc3a7599),
	.w3(32'hbb6bf9a6),
	.w4(32'h3948991f),
	.w5(32'h3a3506b7),
	.w6(32'hbb425db8),
	.w7(32'hbb97a28d),
	.w8(32'hba598c8b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b5047),
	.w1(32'h3ab60183),
	.w2(32'h3af1e0a2),
	.w3(32'hb9bded65),
	.w4(32'h3b113713),
	.w5(32'h3a8505a7),
	.w6(32'h39a5bd7c),
	.w7(32'h3ae76929),
	.w8(32'hba56a401),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb449bfb),
	.w1(32'h3a4ed77c),
	.w2(32'hba5e5e93),
	.w3(32'hb9eac25b),
	.w4(32'h3b0d4acc),
	.w5(32'hba43b869),
	.w6(32'hbb28a79a),
	.w7(32'hbb01e18f),
	.w8(32'h3bab9a15),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c5a76),
	.w1(32'hbc8023be),
	.w2(32'hbca5f533),
	.w3(32'hbc074dcf),
	.w4(32'hbbf0d789),
	.w5(32'hbb7f3850),
	.w6(32'hb9375599),
	.w7(32'hbbce7cd1),
	.w8(32'hba916f23),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa1f11),
	.w1(32'h3bd3e023),
	.w2(32'h3bb53153),
	.w3(32'h3b66b594),
	.w4(32'h3bce17fe),
	.w5(32'h3bd00c17),
	.w6(32'h3a84ef83),
	.w7(32'h3b8604ff),
	.w8(32'h3a933894),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbd483),
	.w1(32'h3bc1f055),
	.w2(32'h3bac3c69),
	.w3(32'h3b1a2c5f),
	.w4(32'h3bb60ba9),
	.w5(32'h3bc861bb),
	.w6(32'h3b73c9ff),
	.w7(32'h3bc5a0c3),
	.w8(32'h3bdc0bc5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06b174),
	.w1(32'hba18e407),
	.w2(32'h3a214035),
	.w3(32'h3af7a4d8),
	.w4(32'h3a8e4a0a),
	.w5(32'h3bcfa4c5),
	.w6(32'h3b10647e),
	.w7(32'h3b0d1bed),
	.w8(32'h3b152054),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b9b4e),
	.w1(32'hba5fbc51),
	.w2(32'h38b59494),
	.w3(32'hba13b2d3),
	.w4(32'h3b02da7f),
	.w5(32'hb91f6ff1),
	.w6(32'h3960a188),
	.w7(32'h39bb6aa7),
	.w8(32'hbb9d27b0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc8764),
	.w1(32'h3a60f99b),
	.w2(32'hba6acfec),
	.w3(32'hbb7e4d11),
	.w4(32'hb9fb4c20),
	.w5(32'h3a9b5a43),
	.w6(32'hbaadca2c),
	.w7(32'hbb927ed0),
	.w8(32'h3a448b2d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef9001),
	.w1(32'hba4f3fc7),
	.w2(32'hb9460e70),
	.w3(32'h3b26ccb5),
	.w4(32'h3ad06668),
	.w5(32'h3bbb4985),
	.w6(32'h3b13b43c),
	.w7(32'h3b0d6a7d),
	.w8(32'h3a378b6a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b660c),
	.w1(32'hba6fe984),
	.w2(32'hb9f897fc),
	.w3(32'h3a6faa96),
	.w4(32'h3afd1ae9),
	.w5(32'h3bb71bb0),
	.w6(32'h3a88a8ec),
	.w7(32'h3b2054fa),
	.w8(32'hbb310328),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84b63a),
	.w1(32'hb94b7095),
	.w2(32'hb90c3b24),
	.w3(32'hba95a1cd),
	.w4(32'hbaba8f82),
	.w5(32'h39b80b4c),
	.w6(32'hb9f7b0d5),
	.w7(32'h3a7ce335),
	.w8(32'h3c0050da),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994c8d),
	.w1(32'hbb86cd74),
	.w2(32'hbaae00d3),
	.w3(32'hbba54cec),
	.w4(32'hbb4792c7),
	.w5(32'hbb1bdb35),
	.w6(32'h3b8d4d2e),
	.w7(32'hba1554a2),
	.w8(32'hbb0634ac),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b8cf1),
	.w1(32'hba16c908),
	.w2(32'hb9a3ad35),
	.w3(32'hba55f033),
	.w4(32'hba907cb3),
	.w5(32'hbaf569f9),
	.w6(32'hbb066516),
	.w7(32'hbb0299cd),
	.w8(32'h3b5a2f35),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b5fcb),
	.w1(32'hbb995821),
	.w2(32'hbbfef8c6),
	.w3(32'hbbc28f41),
	.w4(32'hbc232b4c),
	.w5(32'hbbe1d6db),
	.w6(32'hbb6e313d),
	.w7(32'hbc206a37),
	.w8(32'hbbcb5e20),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9b5e4),
	.w1(32'h3b72da95),
	.w2(32'hb9b8261b),
	.w3(32'h3acc6243),
	.w4(32'h3aa887f4),
	.w5(32'h3ac38a4a),
	.w6(32'h3b77fbf4),
	.w7(32'h3a830d45),
	.w8(32'h3b842b15),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa203f0),
	.w1(32'hba8d82e8),
	.w2(32'h3b360efc),
	.w3(32'hbb70003b),
	.w4(32'hba7a39f6),
	.w5(32'hb8e9b17c),
	.w6(32'hb9896328),
	.w7(32'hbabc2016),
	.w8(32'h3bc9b312),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8588b7),
	.w1(32'hbb799187),
	.w2(32'hbb9ba133),
	.w3(32'hbb4e27e0),
	.w4(32'hbb8d32f4),
	.w5(32'hbb22b332),
	.w6(32'h3be00355),
	.w7(32'hbab62c99),
	.w8(32'h3bb1d748),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6587b5),
	.w1(32'hb9a4cdf0),
	.w2(32'h3a984d68),
	.w3(32'h3b08f1f9),
	.w4(32'h3afce7d6),
	.w5(32'hbb5ad591),
	.w6(32'h3ac7124b),
	.w7(32'h3b067167),
	.w8(32'h3a22a42a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848f66b),
	.w1(32'h39e52d74),
	.w2(32'hb6c0a6ee),
	.w3(32'h38d4b654),
	.w4(32'h3acc01cd),
	.w5(32'hba0da964),
	.w6(32'hb9d120d5),
	.w7(32'h39a51aa6),
	.w8(32'hb98f9908),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15c7f5),
	.w1(32'h3b0c0a14),
	.w2(32'hbab3759c),
	.w3(32'hbb07ea1a),
	.w4(32'h399d549b),
	.w5(32'hba914390),
	.w6(32'hba92b8c7),
	.w7(32'hbb073fa7),
	.w8(32'hb9245a5d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7127),
	.w1(32'hbb354c62),
	.w2(32'hba92774b),
	.w3(32'hbb661837),
	.w4(32'hbb5994e9),
	.w5(32'hbb587888),
	.w6(32'hbb87651a),
	.w7(32'hbb2edf53),
	.w8(32'h3b8fa3bc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b415e0d),
	.w1(32'h37fb795e),
	.w2(32'h3b866760),
	.w3(32'h3b56a587),
	.w4(32'h3b423442),
	.w5(32'h39248f00),
	.w6(32'h3ab17933),
	.w7(32'h3b915a9f),
	.w8(32'hbad0565c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aa7cb),
	.w1(32'h39b172bb),
	.w2(32'h3a85f3e1),
	.w3(32'hbbaffcab),
	.w4(32'hbb6cd807),
	.w5(32'hbab3848f),
	.w6(32'hbb699636),
	.w7(32'hbb2c98cf),
	.w8(32'hbb499b67),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812383a),
	.w1(32'hba689049),
	.w2(32'hba607d0d),
	.w3(32'h39aa378f),
	.w4(32'hb8d5cb98),
	.w5(32'h3ae798e9),
	.w6(32'h39bc3623),
	.w7(32'h39bec753),
	.w8(32'hba4d43aa),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66b9f3),
	.w1(32'h3bbf7143),
	.w2(32'h3c0c2cff),
	.w3(32'h3b76293d),
	.w4(32'h3bc7002a),
	.w5(32'h3be20a10),
	.w6(32'h3afaf799),
	.w7(32'h3b88a1e3),
	.w8(32'h3b3fd9b8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b004147),
	.w1(32'h3abe7c31),
	.w2(32'h3b1b922f),
	.w3(32'h397ccf2e),
	.w4(32'hb9dd94df),
	.w5(32'h3a421dbc),
	.w6(32'h3a9015fb),
	.w7(32'h3a10f833),
	.w8(32'h3a6196c0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98de89),
	.w1(32'hbab8c153),
	.w2(32'hbaa338eb),
	.w3(32'hbac26ba7),
	.w4(32'hbae97bbb),
	.w5(32'hbaf1c980),
	.w6(32'hbaa07005),
	.w7(32'hbab67d01),
	.w8(32'hbae2c9da),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b4be8),
	.w1(32'hba34d92b),
	.w2(32'hbae34f3a),
	.w3(32'hb93ea7ec),
	.w4(32'hb9602600),
	.w5(32'hbaaa7ac0),
	.w6(32'hba3b0d19),
	.w7(32'hba604f67),
	.w8(32'hbab7a768),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacafcda),
	.w1(32'hbac9c155),
	.w2(32'hbab957f2),
	.w3(32'hbb4cf7f6),
	.w4(32'hbb41ce13),
	.w5(32'hbad5e53e),
	.w6(32'hbb09b6d0),
	.w7(32'hbae4138e),
	.w8(32'hba1b07be),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45487d),
	.w1(32'hbb712b2d),
	.w2(32'hbb8d4d4e),
	.w3(32'hbabd1606),
	.w4(32'hbacdb9e3),
	.w5(32'hbb256557),
	.w6(32'hbb85858b),
	.w7(32'hbb8d0a78),
	.w8(32'hbba3dee3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56e9b6),
	.w1(32'hbb03f7ba),
	.w2(32'hbb15c5a9),
	.w3(32'hbb21bb7d),
	.w4(32'hba6d1179),
	.w5(32'hba317d4c),
	.w6(32'hbb5df367),
	.w7(32'hbb109c8f),
	.w8(32'hbb3ff617),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39017c66),
	.w1(32'hba20466b),
	.w2(32'hba183993),
	.w3(32'h3a7eca47),
	.w4(32'h37d3d828),
	.w5(32'hb9e2bccc),
	.w6(32'h39cbccde),
	.w7(32'hb548f2ec),
	.w8(32'hba33a1c6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3833773e),
	.w1(32'h38ca38e8),
	.w2(32'h397a4de0),
	.w3(32'h369ff24d),
	.w4(32'h380407f1),
	.w5(32'h3936a759),
	.w6(32'h3922e1e7),
	.w7(32'h38da39e3),
	.w8(32'h39ad1bdb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5d0c6),
	.w1(32'h39bbdff4),
	.w2(32'h3a4ae6a8),
	.w3(32'hb97e3330),
	.w4(32'h392f4690),
	.w5(32'h3a0f02a9),
	.w6(32'h3a4d2775),
	.w7(32'h397f8508),
	.w8(32'h3a45f585),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3957634f),
	.w1(32'h39b82e70),
	.w2(32'h38862619),
	.w3(32'h3984904e),
	.w4(32'h3a2d10e2),
	.w5(32'h3a788b7d),
	.w6(32'hb9109c3f),
	.w7(32'h39ff99a5),
	.w8(32'h39995b0d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaf952),
	.w1(32'hba2b402e),
	.w2(32'hbae36a57),
	.w3(32'hba74db67),
	.w4(32'h398c8fdf),
	.w5(32'hba025587),
	.w6(32'hbabf5089),
	.w7(32'hb96c0e5e),
	.w8(32'hbaac9a81),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba838206),
	.w1(32'h39434cc1),
	.w2(32'hb9412de0),
	.w3(32'h3a253883),
	.w4(32'h3b2eb7a1),
	.w5(32'h3b046f31),
	.w6(32'hb8859fa2),
	.w7(32'h3aa21996),
	.w8(32'h3a12253a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a6ef4c),
	.w1(32'h37400ab7),
	.w2(32'h37be852b),
	.w3(32'h372093a4),
	.w4(32'hb69d97c9),
	.w5(32'h36eb9f6e),
	.w6(32'h3798ddc4),
	.w7(32'h36f5c5f7),
	.w8(32'h378bd06a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c00d6),
	.w1(32'hb7e63683),
	.w2(32'hb6f11002),
	.w3(32'h38c77343),
	.w4(32'h37909dc4),
	.w5(32'hb93986b8),
	.w6(32'hb987b7ab),
	.w7(32'hb9e4cda0),
	.w8(32'hb9c898e5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0b599),
	.w1(32'hba809037),
	.w2(32'hbb0cc9c3),
	.w3(32'hbad827d6),
	.w4(32'hb9da7a7d),
	.w5(32'hbac5b778),
	.w6(32'hbad5ad31),
	.w7(32'hb9e8a5da),
	.w8(32'hb831f70f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39284eea),
	.w1(32'h3a9f7aec),
	.w2(32'h3ad275f6),
	.w3(32'hb8968fdd),
	.w4(32'h3a0d4f98),
	.w5(32'h3a8db4c5),
	.w6(32'h394a614e),
	.w7(32'h3a6ef918),
	.w8(32'h3aaf142f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfd960),
	.w1(32'hba4c95e0),
	.w2(32'hb9d14d2c),
	.w3(32'hba25a82e),
	.w4(32'hb9f5cfb0),
	.w5(32'hb971d02d),
	.w6(32'hba2e7558),
	.w7(32'hba1e6b02),
	.w8(32'hba0f7ff3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9603f),
	.w1(32'hb9485154),
	.w2(32'hb95cbc3a),
	.w3(32'h3972c0b6),
	.w4(32'h3a3c9a0c),
	.w5(32'h3a04ed42),
	.w6(32'hb87818f0),
	.w7(32'h384f5b6e),
	.w8(32'hb99c105e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d640e),
	.w1(32'hbab50f26),
	.w2(32'hba30fc5c),
	.w3(32'hbadb98ea),
	.w4(32'hbada7335),
	.w5(32'hba9b33e5),
	.w6(32'hba98cd70),
	.w7(32'hbaa615f7),
	.w8(32'hba6fa6eb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11f413),
	.w1(32'hbabb51e8),
	.w2(32'hba93c703),
	.w3(32'hbadcaf62),
	.w4(32'hbac64b4f),
	.w5(32'hbaa26964),
	.w6(32'hbae796a2),
	.w7(32'hbb08d5b9),
	.w8(32'hbb30d382),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a479fd),
	.w1(32'hba9a498a),
	.w2(32'hba8158e7),
	.w3(32'hba1b2e4c),
	.w4(32'hbac2ae06),
	.w5(32'hba374ae6),
	.w6(32'hbaf1b232),
	.w7(32'hbb209e41),
	.w8(32'hbac09c4d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6e66d),
	.w1(32'h3a90b84d),
	.w2(32'h38c73be1),
	.w3(32'h3a995662),
	.w4(32'h3a8698c4),
	.w5(32'hb9b885f1),
	.w6(32'h3ab64e11),
	.w7(32'h3a07e88e),
	.w8(32'hba91fd7a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule