module layer_10_featuremap_432(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18b3cf),
	.w1(32'h398f5f42),
	.w2(32'hbb222627),
	.w3(32'hbbd93bb7),
	.w4(32'hbb1b5bba),
	.w5(32'h3a426533),
	.w6(32'hbbe614b1),
	.w7(32'hbaa15388),
	.w8(32'hba9343db),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb98ba),
	.w1(32'h3bd7a790),
	.w2(32'hba2f51e9),
	.w3(32'hbb5fdaba),
	.w4(32'h3ae2ef37),
	.w5(32'h3ba00d3e),
	.w6(32'hba75b7da),
	.w7(32'hbb6f17f1),
	.w8(32'h3bed98b1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe4fca),
	.w1(32'h3b73e50d),
	.w2(32'hbb556d9d),
	.w3(32'hbaad3a30),
	.w4(32'h3c003007),
	.w5(32'hbc01693c),
	.w6(32'hba08d1dd),
	.w7(32'h3bba14c7),
	.w8(32'h3b0a9d09),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0302ad),
	.w1(32'hbbc23086),
	.w2(32'hbb57d729),
	.w3(32'hbb97f4d8),
	.w4(32'hbba0efe8),
	.w5(32'hbb4baa73),
	.w6(32'h3aa1760c),
	.w7(32'h391f0c82),
	.w8(32'h39b4829b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a125284),
	.w1(32'hbb27e49e),
	.w2(32'h3b12ca7a),
	.w3(32'h3b12d2df),
	.w4(32'hbb3c02ab),
	.w5(32'h3b24c86d),
	.w6(32'h3b0e56ca),
	.w7(32'h3a2ef53e),
	.w8(32'hba8df045),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dd02c),
	.w1(32'hbb117d3b),
	.w2(32'hb732b68e),
	.w3(32'h3ae9031e),
	.w4(32'h39122035),
	.w5(32'h39a6830c),
	.w6(32'h3b407687),
	.w7(32'hbadc990a),
	.w8(32'hbbea29b5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd98cf),
	.w1(32'h3b8c0148),
	.w2(32'hbb39bf9a),
	.w3(32'h3b67368d),
	.w4(32'h3beddb50),
	.w5(32'hbbfce2b1),
	.w6(32'h3b9e1bd1),
	.w7(32'h38970861),
	.w8(32'hbb9904f5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc21b1),
	.w1(32'h3b1fa37e),
	.w2(32'hbba17729),
	.w3(32'hbbeab2dc),
	.w4(32'h3a5909b7),
	.w5(32'h39894cf7),
	.w6(32'hbc186b59),
	.w7(32'hbbbb9844),
	.w8(32'hbb87d8ad),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaf4a7),
	.w1(32'hbb07ecd9),
	.w2(32'h3af0a30a),
	.w3(32'hbc04b1b2),
	.w4(32'h3aa685e7),
	.w5(32'hbbd6e11b),
	.w6(32'hbc343d64),
	.w7(32'h39618878),
	.w8(32'hbbe39bac),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07314f),
	.w1(32'hbbc7c6bf),
	.w2(32'hbba028aa),
	.w3(32'h3c2c7442),
	.w4(32'hbb97183a),
	.w5(32'hbc28d907),
	.w6(32'h3af1e699),
	.w7(32'h3baf3743),
	.w8(32'hbb028393),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94503d),
	.w1(32'hbb7b5edd),
	.w2(32'hbb3d2bdb),
	.w3(32'hbab7fa8d),
	.w4(32'hbb5ccac4),
	.w5(32'hbb3a872e),
	.w6(32'hba91ce5f),
	.w7(32'hbb2f61f6),
	.w8(32'hbbb4ec4b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ccf50),
	.w1(32'h3ad226c3),
	.w2(32'h3899ca8a),
	.w3(32'h3bd9cdf8),
	.w4(32'h3b2b1e33),
	.w5(32'h3b260e53),
	.w6(32'h3badec17),
	.w7(32'h3af1a22e),
	.w8(32'h3a10ac04),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a7de5),
	.w1(32'hbaa73000),
	.w2(32'hbb0ea5f8),
	.w3(32'hba889957),
	.w4(32'h3b31a557),
	.w5(32'hba834769),
	.w6(32'h3b810c5e),
	.w7(32'h3bbc7555),
	.w8(32'h3c2f1b66),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb213e58),
	.w1(32'hba19a64a),
	.w2(32'h3bbe04d2),
	.w3(32'hbb58991d),
	.w4(32'hba9ed335),
	.w5(32'h3ad8e1c6),
	.w6(32'h3a062377),
	.w7(32'h3b8413a8),
	.w8(32'h38b082e2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3931e842),
	.w1(32'hbb047785),
	.w2(32'h3b04b4d7),
	.w3(32'h3c1405f1),
	.w4(32'h3b8d4673),
	.w5(32'h3b982c07),
	.w6(32'h3c448b66),
	.w7(32'h3b5630cb),
	.w8(32'hbad4a278),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4c2ad),
	.w1(32'h3b437ace),
	.w2(32'hbb6166ea),
	.w3(32'hbb6ce3a4),
	.w4(32'h3c23fdfd),
	.w5(32'hbb0b82c9),
	.w6(32'hba06477a),
	.w7(32'h3b97e745),
	.w8(32'hbaa8e04b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb508937),
	.w1(32'h3b08865e),
	.w2(32'h3b36c42f),
	.w3(32'hbaa87ff5),
	.w4(32'hbadf931e),
	.w5(32'hbb5a45a6),
	.w6(32'hbba164c8),
	.w7(32'hb9c81d93),
	.w8(32'hbb816b20),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27d2b7),
	.w1(32'hbc20df60),
	.w2(32'hbc30af6f),
	.w3(32'hbc34fed0),
	.w4(32'hbbaf4044),
	.w5(32'hbbacb3b6),
	.w6(32'hbb99660a),
	.w7(32'hbba09461),
	.w8(32'hbbe2be0e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe288cd),
	.w1(32'hbc0b93bf),
	.w2(32'hba9edcfb),
	.w3(32'hbc0dcc24),
	.w4(32'hbb7c4871),
	.w5(32'hbba0d7a0),
	.w6(32'hbb5d4277),
	.w7(32'hbb01594f),
	.w8(32'hbbc3cd5b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8f963),
	.w1(32'hbb5f2fdd),
	.w2(32'h3b158a50),
	.w3(32'h3ace41e8),
	.w4(32'hbaaa0f58),
	.w5(32'hba22ba93),
	.w6(32'h3a591f20),
	.w7(32'hba8052c1),
	.w8(32'hbb1b54f0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6d04a),
	.w1(32'hb99dd862),
	.w2(32'h3a1cb12a),
	.w3(32'h39b07b81),
	.w4(32'h3a32f617),
	.w5(32'h3928984e),
	.w6(32'h3bb97c80),
	.w7(32'hb89eccfe),
	.w8(32'hbb498b18),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8f07c),
	.w1(32'hbb4b1d47),
	.w2(32'h39d5435b),
	.w3(32'h3c039dc2),
	.w4(32'hbb49cd3b),
	.w5(32'h38c69c20),
	.w6(32'h3b5a9b48),
	.w7(32'hba4104a9),
	.w8(32'hba5b87e7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40b84f),
	.w1(32'hbc4c0e18),
	.w2(32'hbc122972),
	.w3(32'hbc209ddc),
	.w4(32'hbb21c4e4),
	.w5(32'hbc29cb3b),
	.w6(32'hbc368bb8),
	.w7(32'hba9b0e7c),
	.w8(32'hbc021567),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3862cf),
	.w1(32'hbb56655a),
	.w2(32'hbaf750cd),
	.w3(32'h3b4c99ca),
	.w4(32'h3b075bd1),
	.w5(32'hbb175c58),
	.w6(32'hbab55ed9),
	.w7(32'hb9f8d753),
	.w8(32'hbb55ceec),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d8985),
	.w1(32'h3bcf64e8),
	.w2(32'hbc0be596),
	.w3(32'h3b937cac),
	.w4(32'h3befa9ff),
	.w5(32'hbbbe3b23),
	.w6(32'hbb0b3785),
	.w7(32'h3b797f36),
	.w8(32'hb9e9b106),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d9c95),
	.w1(32'hbaabf8f3),
	.w2(32'hba8ffad8),
	.w3(32'h3aa55e26),
	.w4(32'hba6cbe52),
	.w5(32'h3b35e8bc),
	.w6(32'hbada7918),
	.w7(32'h39f98ea5),
	.w8(32'hbb1a752d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f7815),
	.w1(32'hbbbadd16),
	.w2(32'hbb4b494a),
	.w3(32'h3ad8df6f),
	.w4(32'hbaf41f0b),
	.w5(32'hbc08bf79),
	.w6(32'h3aa352a0),
	.w7(32'h3ad1f32c),
	.w8(32'hbc0037d4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88cea4),
	.w1(32'h3bc13f1d),
	.w2(32'h3c00b218),
	.w3(32'hbb3666d8),
	.w4(32'h3b7e5fb5),
	.w5(32'h3b049cb5),
	.w6(32'hbc130c2d),
	.w7(32'hbb075e77),
	.w8(32'hbb949aef),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8b7be),
	.w1(32'hbb2eee85),
	.w2(32'hbbc7654b),
	.w3(32'h3b8560e4),
	.w4(32'hbbc09984),
	.w5(32'hbc01d753),
	.w6(32'h3b70f290),
	.w7(32'hba3f2ce3),
	.w8(32'hbba46100),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc1c4e),
	.w1(32'h3b3ba86f),
	.w2(32'h3a7dd27a),
	.w3(32'hbab46418),
	.w4(32'h3b9dd0bf),
	.w5(32'h3b0b99a9),
	.w6(32'hbb2672e3),
	.w7(32'h3a8d6cfe),
	.w8(32'hbb9a52c1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39c00e),
	.w1(32'h3ab5ef1b),
	.w2(32'hbad36b38),
	.w3(32'hbb6e5364),
	.w4(32'h3bbc7b50),
	.w5(32'h3b3b5326),
	.w6(32'hbb7d7553),
	.w7(32'h3b012df7),
	.w8(32'hbaab372e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ba989),
	.w1(32'h3c0446bb),
	.w2(32'hbb09c7dd),
	.w3(32'hbb10d46d),
	.w4(32'h3c3b1be5),
	.w5(32'h3a8e58f0),
	.w6(32'h3acc61e2),
	.w7(32'h3bc3879c),
	.w8(32'h3b859580),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08fc77),
	.w1(32'h3ba50c9c),
	.w2(32'hba1d7c83),
	.w3(32'hbb8c26bf),
	.w4(32'h3b7c5756),
	.w5(32'hbbce4610),
	.w6(32'hbb911f39),
	.w7(32'h3b8dc9c0),
	.w8(32'h3ba9b348),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f63c8),
	.w1(32'h3b84d58f),
	.w2(32'h3aebcded),
	.w3(32'h3ad01f9e),
	.w4(32'h3b7ce314),
	.w5(32'hbc123e9f),
	.w6(32'hbb8575e7),
	.w7(32'h38ae5788),
	.w8(32'hbb9fc179),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ced678),
	.w1(32'hbb3f40df),
	.w2(32'hbb329286),
	.w3(32'h3b7d229b),
	.w4(32'hbb07e373),
	.w5(32'hbab91cab),
	.w6(32'hbb1c2209),
	.w7(32'h3ae6132d),
	.w8(32'hba2c1783),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab037cb),
	.w1(32'hbb74cf57),
	.w2(32'hbbee395d),
	.w3(32'h38f8a3c9),
	.w4(32'h3ac49fee),
	.w5(32'hba196473),
	.w6(32'h3b916513),
	.w7(32'h3a7b0a3d),
	.w8(32'h3acfdcf1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73a8c),
	.w1(32'hbbb7fd53),
	.w2(32'h3b054789),
	.w3(32'h3b927e47),
	.w4(32'hbb4aff1d),
	.w5(32'h3b0c7050),
	.w6(32'h3b2a9dcf),
	.w7(32'h3ba70599),
	.w8(32'h3b0bedbb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc19061),
	.w1(32'h3c716797),
	.w2(32'hbb08fc52),
	.w3(32'h3c5a9e78),
	.w4(32'h3ca585af),
	.w5(32'h3c3a74f7),
	.w6(32'h3c23e8d6),
	.w7(32'h3a6f1734),
	.w8(32'h3c3f18f7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb263dd),
	.w1(32'h3c396453),
	.w2(32'h3c3a1443),
	.w3(32'h3b92f3ee),
	.w4(32'h3bf27699),
	.w5(32'h3bfe1c4b),
	.w6(32'h3bd0a0cf),
	.w7(32'h3b2fa666),
	.w8(32'hbab81f9b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b984ced),
	.w1(32'hbad0aa30),
	.w2(32'hbb117d40),
	.w3(32'h3bbd61e0),
	.w4(32'h3adb0a53),
	.w5(32'h3a833bbb),
	.w6(32'h3bc1f37c),
	.w7(32'hbb351bd5),
	.w8(32'h390da9d3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9671cd),
	.w1(32'hba90333f),
	.w2(32'h3c40f9e2),
	.w3(32'hbb876488),
	.w4(32'hbbd5ef6e),
	.w5(32'h3c8d94c3),
	.w6(32'hbb5eb6a8),
	.w7(32'hbbb171e6),
	.w8(32'h3c49445d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba98f46),
	.w1(32'hbb06afaf),
	.w2(32'h3ba13834),
	.w3(32'hbb48049f),
	.w4(32'hbb006512),
	.w5(32'h3a40b644),
	.w6(32'h3b388721),
	.w7(32'hbadd46aa),
	.w8(32'hbb132a4f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b099fdb),
	.w1(32'h3ab9488f),
	.w2(32'hbbb2809d),
	.w3(32'h3b4b98fe),
	.w4(32'h3be015db),
	.w5(32'h3af472e3),
	.w6(32'h3b28955f),
	.w7(32'h3bb86c5d),
	.w8(32'h3bf853f6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba32629),
	.w1(32'h3b2e83dc),
	.w2(32'h3b821176),
	.w3(32'hbc222e41),
	.w4(32'hbacc723f),
	.w5(32'h3c16708f),
	.w6(32'hbb6e0f57),
	.w7(32'hbab2e5e3),
	.w8(32'hba327af1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45ecd7),
	.w1(32'h3a8ab0b1),
	.w2(32'hb8a45cc6),
	.w3(32'h3b045ea7),
	.w4(32'hbac2011e),
	.w5(32'hbbafc70b),
	.w6(32'hb9d62040),
	.w7(32'h3b786003),
	.w8(32'h3a18937f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ac3aa),
	.w1(32'hbaffc69e),
	.w2(32'hbb93addb),
	.w3(32'h3b8a2f79),
	.w4(32'h3c0d5e7c),
	.w5(32'hbb50a66f),
	.w6(32'h3b6b349e),
	.w7(32'h3bb17c83),
	.w8(32'hba467549),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb432bad),
	.w1(32'hbba1b8e7),
	.w2(32'hbaeb9c66),
	.w3(32'hbad4cdc7),
	.w4(32'hbb487799),
	.w5(32'hbb6509df),
	.w6(32'hbc35b0f3),
	.w7(32'h3a1fae44),
	.w8(32'hbaadbeb0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac21c95),
	.w1(32'hbc1862ea),
	.w2(32'hbbc96f78),
	.w3(32'h39e38d01),
	.w4(32'hbbb2558f),
	.w5(32'hbbb6a2ff),
	.w6(32'h3b98aa4f),
	.w7(32'hbb6ebb89),
	.w8(32'hbbfeed72),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfb5a0),
	.w1(32'hbbc8fa94),
	.w2(32'h3b9a4abf),
	.w3(32'h3b045cb6),
	.w4(32'hbb696fa6),
	.w5(32'h3a50390e),
	.w6(32'h39861e8a),
	.w7(32'hbbb5bee1),
	.w8(32'hbbbd91b2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba243b8),
	.w1(32'h3b4d4c6a),
	.w2(32'h39851d70),
	.w3(32'h3bc7ec90),
	.w4(32'h3ba2d050),
	.w5(32'h3bcd12cd),
	.w6(32'h3a83000e),
	.w7(32'h39d89781),
	.w8(32'h3bc5c773),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e8b28),
	.w1(32'h3a290c5d),
	.w2(32'hbb182a4f),
	.w3(32'hbae487e0),
	.w4(32'hba2850f8),
	.w5(32'hb9e8fa44),
	.w6(32'hbbaf6612),
	.w7(32'hbb597451),
	.w8(32'h3b2cb63f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacd2c8),
	.w1(32'h3a9409d5),
	.w2(32'hbb15f31f),
	.w3(32'h3a3647d9),
	.w4(32'h3ba1657b),
	.w5(32'hbaba367c),
	.w6(32'hba90acfb),
	.w7(32'h3a8efee0),
	.w8(32'hbad99d55),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e3557),
	.w1(32'h3b06b40e),
	.w2(32'h3a98e00d),
	.w3(32'h3a0e0129),
	.w4(32'h3b81b6af),
	.w5(32'hba7ec5ad),
	.w6(32'hba4efb29),
	.w7(32'hbb566c64),
	.w8(32'hbbfa65c5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f1573),
	.w1(32'hbb36d80b),
	.w2(32'hbc026d51),
	.w3(32'hbc2dba53),
	.w4(32'h3a4c2f6a),
	.w5(32'hbbce3fcf),
	.w6(32'hbbf91ed5),
	.w7(32'hbb88965d),
	.w8(32'hbb92f3b2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88199b),
	.w1(32'h399fa5b3),
	.w2(32'hbb5c3a06),
	.w3(32'hbab319c6),
	.w4(32'h3b539c04),
	.w5(32'hba3eea92),
	.w6(32'hbbd5a827),
	.w7(32'hbb20f893),
	.w8(32'h3adc0c7c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddde2a),
	.w1(32'h3aa6dde2),
	.w2(32'hbb03cbb5),
	.w3(32'hbad57f26),
	.w4(32'h3c0532e5),
	.w5(32'hbad28660),
	.w6(32'hbb27e1a6),
	.w7(32'h39ce06fb),
	.w8(32'h3b927d85),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05d08c),
	.w1(32'h3a7c8dd3),
	.w2(32'h396f73b3),
	.w3(32'hbb633586),
	.w4(32'h3a2edd25),
	.w5(32'h3916e60b),
	.w6(32'hbb022e81),
	.w7(32'h3abb7c20),
	.w8(32'h3adf2b54),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9750b),
	.w1(32'hbaed2c6b),
	.w2(32'h3b440c68),
	.w3(32'hbad3b077),
	.w4(32'hbbb2eaa0),
	.w5(32'h3af44266),
	.w6(32'h3a8fa66e),
	.w7(32'hbb2f21e5),
	.w8(32'hbb292f2b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf955fd),
	.w1(32'h3a5184f1),
	.w2(32'h3b09f671),
	.w3(32'h3aebed0c),
	.w4(32'hbba46a91),
	.w5(32'h3b70ae83),
	.w6(32'hbad5b08a),
	.w7(32'hbbd3c633),
	.w8(32'h3a452ba6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ae44),
	.w1(32'hb9a74b39),
	.w2(32'hbb5a32f0),
	.w3(32'hb922f125),
	.w4(32'hb9197071),
	.w5(32'h3a2e8fac),
	.w6(32'h3b31b150),
	.w7(32'hbb1166f6),
	.w8(32'hbac0124c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88846c),
	.w1(32'hbbe72e0b),
	.w2(32'hbb9afead),
	.w3(32'hbb9f2fe9),
	.w4(32'hbbd66396),
	.w5(32'hbbbe82fb),
	.w6(32'hbb73c00c),
	.w7(32'hba32bebe),
	.w8(32'hbc321e9c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf883df),
	.w1(32'hbaa2c6f8),
	.w2(32'h3bc53ba9),
	.w3(32'hbc0fd6e2),
	.w4(32'hbb51182e),
	.w5(32'h3b073c2a),
	.w6(32'hbbe61345),
	.w7(32'hbb383c0f),
	.w8(32'hbaaf8550),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3d1f3),
	.w1(32'h3a463688),
	.w2(32'hbb7560f5),
	.w3(32'h3b9ae73d),
	.w4(32'h3a902671),
	.w5(32'hba9a2a2d),
	.w6(32'h3b80f2a4),
	.w7(32'h3a6f0930),
	.w8(32'h3beada02),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83c75d),
	.w1(32'h3a9b6205),
	.w2(32'hba0b90a9),
	.w3(32'hbba42e53),
	.w4(32'hb9e823f6),
	.w5(32'hbb20ca8e),
	.w6(32'hbb9095d9),
	.w7(32'hb909e00c),
	.w8(32'hb9a9dbba),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a6419),
	.w1(32'h3b895cd8),
	.w2(32'h3ae4c83b),
	.w3(32'hbb51589b),
	.w4(32'h3b7c43ba),
	.w5(32'h3b07eabc),
	.w6(32'hb933a4bb),
	.w7(32'h3adbe089),
	.w8(32'h3b34469c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5c28d),
	.w1(32'hb8b1c54c),
	.w2(32'h3bb977e2),
	.w3(32'hbac1d562),
	.w4(32'hba438aac),
	.w5(32'h3b4f2416),
	.w6(32'hba753224),
	.w7(32'hba82e32b),
	.w8(32'hbaac0989),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c6eeed),
	.w1(32'hbb74c964),
	.w2(32'hb9c851e5),
	.w3(32'h3a3f51a9),
	.w4(32'hbbc73bc1),
	.w5(32'hba9d6ea4),
	.w6(32'h3b1f8dc7),
	.w7(32'hbbbe0f4b),
	.w8(32'hbbfb700e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb930d81),
	.w1(32'hbb55d12d),
	.w2(32'hbb474f1f),
	.w3(32'h3b71e6fd),
	.w4(32'h3a936908),
	.w5(32'hba8115bc),
	.w6(32'hbb7e02d9),
	.w7(32'h39d5679f),
	.w8(32'hbacc6c20),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6053cd),
	.w1(32'hbc35b25e),
	.w2(32'hbbba34b4),
	.w3(32'hba47ea4d),
	.w4(32'hbbd541aa),
	.w5(32'hbadff0e7),
	.w6(32'hbbee88ea),
	.w7(32'hbc1e83a4),
	.w8(32'hbbb1a05c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c42e5),
	.w1(32'h3af7a6c6),
	.w2(32'h38af931b),
	.w3(32'h3bc9b1c8),
	.w4(32'h3bf39fc1),
	.w5(32'h39cc86f0),
	.w6(32'hbb603cfc),
	.w7(32'h3a06deac),
	.w8(32'hb9f1b1f0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a9b388),
	.w1(32'hb790d80d),
	.w2(32'h382a0390),
	.w3(32'h369316cd),
	.w4(32'hb6d922f7),
	.w5(32'h381bf9f1),
	.w6(32'hb79d67ff),
	.w7(32'h3798c2b4),
	.w8(32'h385aee36),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c5411c),
	.w1(32'h3732020c),
	.w2(32'h3886917a),
	.w3(32'hb769d1dc),
	.w4(32'hb82d2bee),
	.w5(32'h37c3c6c4),
	.w6(32'h37b92a28),
	.w7(32'h382382d7),
	.w8(32'h38e62854),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb791e881),
	.w1(32'hb872c7fb),
	.w2(32'h37a1184c),
	.w3(32'hb836432b),
	.w4(32'hb814b1c0),
	.w5(32'hb6dc12b7),
	.w6(32'h384185b2),
	.w7(32'hb8443294),
	.w8(32'hb7ab734d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5523e0),
	.w1(32'hbaae1c2d),
	.w2(32'hba7b93ef),
	.w3(32'hba0ac6f6),
	.w4(32'hba8b0042),
	.w5(32'hb9befacf),
	.w6(32'h38e948fa),
	.w7(32'hba83da64),
	.w8(32'hbaa36599),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370f951e),
	.w1(32'h36bcc2dd),
	.w2(32'h3860aa0d),
	.w3(32'hb5e5c868),
	.w4(32'hb7e34586),
	.w5(32'h3831024a),
	.w6(32'h38272b80),
	.w7(32'hb71db5e1),
	.w8(32'h380c4ee9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee4c3),
	.w1(32'hbbce029f),
	.w2(32'hbb2e6615),
	.w3(32'hbb61edd6),
	.w4(32'hbb442fa5),
	.w5(32'h39fde432),
	.w6(32'hba8f8ce9),
	.w7(32'hbac4d115),
	.w8(32'hbadfe2a2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad34cb6),
	.w1(32'hbc160001),
	.w2(32'hbbad89f5),
	.w3(32'hbb7e83cc),
	.w4(32'hbbd0e3a5),
	.w5(32'hbb2a543a),
	.w6(32'hbb44fba9),
	.w7(32'hbbc273d7),
	.w8(32'hbb9f2f2f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a404781),
	.w1(32'h3aefca5a),
	.w2(32'hba36b653),
	.w3(32'h3b199fa0),
	.w4(32'h3b33b3ae),
	.w5(32'hbaaa3982),
	.w6(32'h3b341c16),
	.w7(32'h3af85f17),
	.w8(32'hba3d4a7e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb116c80),
	.w1(32'hbada03d3),
	.w2(32'hba8d4d5b),
	.w3(32'hbab26d77),
	.w4(32'hba9cdc0c),
	.w5(32'hb99c04eb),
	.w6(32'hba560665),
	.w7(32'hba86829b),
	.w8(32'hbaf34170),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803b78),
	.w1(32'hbb7bee81),
	.w2(32'h38b2ef76),
	.w3(32'hbaa92bc5),
	.w4(32'hba8afbcb),
	.w5(32'h3a9f3bac),
	.w6(32'hb9efdfea),
	.w7(32'hba8f28f8),
	.w8(32'hbac3d71c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2540f3),
	.w1(32'h3a79bbee),
	.w2(32'hb9f6bbb4),
	.w3(32'hb7fb7283),
	.w4(32'h3a8d8951),
	.w5(32'hb9ceb18c),
	.w6(32'hb90b61e3),
	.w7(32'h39b3d0a9),
	.w8(32'hba75111c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb009f7f),
	.w1(32'hbb22442f),
	.w2(32'hbac0e50f),
	.w3(32'hbab64adc),
	.w4(32'hbacf052e),
	.w5(32'hba087f25),
	.w6(32'hba6825ff),
	.w7(32'hba4e9805),
	.w8(32'hbacd974e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a3f63),
	.w1(32'hb7f503fe),
	.w2(32'h3732d871),
	.w3(32'hb8444837),
	.w4(32'hb7e11720),
	.w5(32'h379949d5),
	.w6(32'hb7e0804f),
	.w7(32'h370d84be),
	.w8(32'h388cf930),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385ac9e7),
	.w1(32'hb742dc66),
	.w2(32'h3683e1ba),
	.w3(32'h38284e55),
	.w4(32'hb82032fa),
	.w5(32'hb7d4309b),
	.w6(32'h3792fc98),
	.w7(32'hb74a7373),
	.w8(32'hb6b3e733),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b961ce),
	.w1(32'h38c1c3d2),
	.w2(32'h39370b91),
	.w3(32'h3914a287),
	.w4(32'h38c7fef8),
	.w5(32'h3907a510),
	.w6(32'h39aa61e0),
	.w7(32'h390c86b3),
	.w8(32'h393f5d03),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a046aa3),
	.w1(32'h39d735a6),
	.w2(32'h39be2f22),
	.w3(32'h39e7e1a1),
	.w4(32'h39bb5797),
	.w5(32'h399d71cd),
	.w6(32'h39a9b65a),
	.w7(32'h38baf5c0),
	.w8(32'h385a1da0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a823e),
	.w1(32'h3a04f601),
	.w2(32'hb8f4f742),
	.w3(32'h3ad401f9),
	.w4(32'h3ad7761c),
	.w5(32'h3ad435b5),
	.w6(32'hba09f83a),
	.w7(32'hba9fab2c),
	.w8(32'h39513e86),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999db16),
	.w1(32'h397ac8fe),
	.w2(32'h39dc1092),
	.w3(32'h38b06e0d),
	.w4(32'h38d01bd7),
	.w5(32'h39f7e82a),
	.w6(32'hb5daefb6),
	.w7(32'hb86ea2bd),
	.w8(32'h39025a18),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ed2f),
	.w1(32'hbb4141c2),
	.w2(32'hba884a89),
	.w3(32'hb87a110f),
	.w4(32'h3a2e1e1d),
	.w5(32'hb95571b7),
	.w6(32'hb9bce931),
	.w7(32'h3acfa496),
	.w8(32'h3a66e047),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd8324),
	.w1(32'hbbe73333),
	.w2(32'hba7f4d5b),
	.w3(32'hbc05a3d6),
	.w4(32'hbb905f21),
	.w5(32'h3a94fbd7),
	.w6(32'hbbc8e29e),
	.w7(32'hbbcfd3be),
	.w8(32'hbb0ce993),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00315c),
	.w1(32'h3b786bd8),
	.w2(32'h3b2456af),
	.w3(32'h3ad9d58c),
	.w4(32'h3b4eff71),
	.w5(32'h3b2a09c1),
	.w6(32'h3a47f565),
	.w7(32'h3a1d3d0f),
	.w8(32'h39703005),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb056c6),
	.w1(32'hbb9bfa80),
	.w2(32'hbb2be0b8),
	.w3(32'hbb940ed8),
	.w4(32'hba0250d1),
	.w5(32'h3a893f0a),
	.w6(32'hb9d0dd2b),
	.w7(32'h3b88456d),
	.w8(32'h3ac52e3d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8071c),
	.w1(32'h3b184ee7),
	.w2(32'h3b0aa480),
	.w3(32'h3b5f7468),
	.w4(32'h3b6e3693),
	.w5(32'h3ac61ac1),
	.w6(32'h3ad3adc6),
	.w7(32'h3aaf447d),
	.w8(32'h3a485d88),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc99350),
	.w1(32'hbbb1384b),
	.w2(32'hbb80902d),
	.w3(32'hbb97fef4),
	.w4(32'hbb7dea4c),
	.w5(32'hba960076),
	.w6(32'hbabd6c78),
	.w7(32'hba462364),
	.w8(32'hbb0cd053),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9af7a),
	.w1(32'h3a13a270),
	.w2(32'h3ad96038),
	.w3(32'hb9427800),
	.w4(32'h3b051346),
	.w5(32'h3b227ef9),
	.w6(32'h3ac16878),
	.w7(32'h3a8613ee),
	.w8(32'h3a4f0d08),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a289a71),
	.w1(32'h3b1fb172),
	.w2(32'hbaa09b74),
	.w3(32'h3ada61f1),
	.w4(32'h3b4f6924),
	.w5(32'h3abd4189),
	.w6(32'hb73abe3a),
	.w7(32'h386799cf),
	.w8(32'h3a2f999a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a092789),
	.w1(32'h39c9a719),
	.w2(32'h393e39c6),
	.w3(32'h3a46eb92),
	.w4(32'h35f1571a),
	.w5(32'hb92ba18a),
	.w6(32'h39f46617),
	.w7(32'h38aa2385),
	.w8(32'hb90bd6cf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb271),
	.w1(32'hbb732d14),
	.w2(32'hbb3769f7),
	.w3(32'hbb2d129c),
	.w4(32'hba7bdd3d),
	.w5(32'hba6999c2),
	.w6(32'hb9d962e6),
	.w7(32'h3a08b710),
	.w8(32'hba9634e6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba74d4),
	.w1(32'hbb5ad800),
	.w2(32'h3b07bff5),
	.w3(32'hbb9524be),
	.w4(32'hb8bc3120),
	.w5(32'h3b4456e8),
	.w6(32'hbab3e223),
	.w7(32'h3a529fed),
	.w8(32'h3b061399),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a326670),
	.w1(32'hbc0f7d13),
	.w2(32'hbc0058dd),
	.w3(32'hba672faf),
	.w4(32'hbb0a1c98),
	.w5(32'hbb239684),
	.w6(32'hbbad1e56),
	.w7(32'hba492f74),
	.w8(32'hbb1dbb37),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02f667),
	.w1(32'h3b30561a),
	.w2(32'hba76da94),
	.w3(32'h3b14c6e6),
	.w4(32'h3b839767),
	.w5(32'h3a9c2e46),
	.w6(32'h39577aaf),
	.w7(32'h3b294d92),
	.w8(32'h3b0e7e91),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992332d),
	.w1(32'h3a88099f),
	.w2(32'h3affd474),
	.w3(32'h3b4b705a),
	.w4(32'h3b986a27),
	.w5(32'h3a06dda3),
	.w6(32'h3b03e019),
	.w7(32'h3b403a48),
	.w8(32'h3ab6c34b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed31af),
	.w1(32'hbb730a1d),
	.w2(32'hba9a3c1c),
	.w3(32'hbae54093),
	.w4(32'h3ad7bc75),
	.w5(32'h38d54e2a),
	.w6(32'hb91cbe6e),
	.w7(32'h3b869e00),
	.w8(32'hb8d24346),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a4c5c),
	.w1(32'h39c89677),
	.w2(32'h3a64ae54),
	.w3(32'hba619f8a),
	.w4(32'h397c8d5d),
	.w5(32'h3a7e3635),
	.w6(32'hba1a19b4),
	.w7(32'h3a130628),
	.w8(32'h3a81299a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc044ce),
	.w1(32'hbc72ddb1),
	.w2(32'hbc61f931),
	.w3(32'hbba30159),
	.w4(32'hbbb66e82),
	.w5(32'hbb79a004),
	.w6(32'hbb423129),
	.w7(32'hbb7eb8fd),
	.w8(32'hbba316e0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89384a),
	.w1(32'hb9a0a32a),
	.w2(32'h3761e5e7),
	.w3(32'h3b013227),
	.w4(32'h3a7a7dcf),
	.w5(32'hbabbbef3),
	.w6(32'h3b0e116a),
	.w7(32'h3b3409d1),
	.w8(32'h38e78dbd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddfa28),
	.w1(32'h398ca352),
	.w2(32'h38ddda6b),
	.w3(32'h39d7f0bf),
	.w4(32'h39598b16),
	.w5(32'h381530f6),
	.w6(32'h39f5d9c8),
	.w7(32'h391215d0),
	.w8(32'h39017d1e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba611e12),
	.w1(32'h38c887cb),
	.w2(32'hba643328),
	.w3(32'hb9e660f9),
	.w4(32'h3a3c4caf),
	.w5(32'hb8a90acb),
	.w6(32'hbaa40f5d),
	.w7(32'hba7b083d),
	.w8(32'hba23f292),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b0377),
	.w1(32'hb9089f13),
	.w2(32'h3a4e415f),
	.w3(32'h39fface4),
	.w4(32'h39536178),
	.w5(32'hba87e2ea),
	.w6(32'h3b0f444b),
	.w7(32'h3b0bf83d),
	.w8(32'h39650b51),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13907c),
	.w1(32'h3b029a99),
	.w2(32'h3a514c91),
	.w3(32'h3b26834b),
	.w4(32'h3b597335),
	.w5(32'h3a1dd731),
	.w6(32'h3b0f8e53),
	.w7(32'h3b58fbb0),
	.w8(32'h3ab275f3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394eaf89),
	.w1(32'h3b358de2),
	.w2(32'hb9ca54d3),
	.w3(32'h39dce2e8),
	.w4(32'h3a918fbb),
	.w5(32'hb7b10c2f),
	.w6(32'h3ac494e0),
	.w7(32'hb9b15e2f),
	.w8(32'hba8289bf),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac564b6),
	.w1(32'h38bbf33c),
	.w2(32'hba18ca50),
	.w3(32'hb7630606),
	.w4(32'h3a50eaf4),
	.w5(32'hba028a01),
	.w6(32'hb9f7afc9),
	.w7(32'h38c839cc),
	.w8(32'hbaa9f064),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb800b3e),
	.w1(32'hbad1ec0f),
	.w2(32'h3b260a99),
	.w3(32'hba6c6920),
	.w4(32'h3b3c5dd1),
	.w5(32'h3b89a686),
	.w6(32'hbad443d8),
	.w7(32'h3b834d61),
	.w8(32'h3b9fdb36),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcbf44),
	.w1(32'hba8ce5d7),
	.w2(32'hba37d22c),
	.w3(32'hbb3f880a),
	.w4(32'hb9a7d4f0),
	.w5(32'hba6ca6f1),
	.w6(32'hba986406),
	.w7(32'hba8a1ca7),
	.w8(32'hbb0869cc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3830e563),
	.w1(32'h388b97f0),
	.w2(32'h3a473cd7),
	.w3(32'h3a802a04),
	.w4(32'h3aaa1672),
	.w5(32'h377a1935),
	.w6(32'h3afd00cc),
	.w7(32'h3ad171d4),
	.w8(32'h3a168457),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916b447),
	.w1(32'hb8ff3f81),
	.w2(32'hb8a34c7d),
	.w3(32'hb9841ba4),
	.w4(32'hb94308b2),
	.w5(32'hb941cc7a),
	.w6(32'hb980d69a),
	.w7(32'hb948ca6e),
	.w8(32'hb916b933),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866019d),
	.w1(32'hb7b36dc0),
	.w2(32'hb90c872c),
	.w3(32'h390b2553),
	.w4(32'hb8e709fc),
	.w5(32'h372f8577),
	.w6(32'h378b9a48),
	.w7(32'h38d7bffe),
	.w8(32'hb9a91ca0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b8712),
	.w1(32'h37bc200e),
	.w2(32'h3698d29f),
	.w3(32'h37194148),
	.w4(32'h376f6c16),
	.w5(32'h366a0743),
	.w6(32'h36392f54),
	.w7(32'h37ad57d5),
	.w8(32'h37eb64f3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd940a),
	.w1(32'h39d7f1a6),
	.w2(32'h3a0f7b75),
	.w3(32'h3a3273e0),
	.w4(32'h3a1b9415),
	.w5(32'h3a0d2bc7),
	.w6(32'h3a305709),
	.w7(32'h3988e461),
	.w8(32'hb98c4f51),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961b4b0),
	.w1(32'h3a9cc531),
	.w2(32'h3a31e3f1),
	.w3(32'h3aae1105),
	.w4(32'h3b19a181),
	.w5(32'h39191dcc),
	.w6(32'h3ae832c8),
	.w7(32'h3b1c99f0),
	.w8(32'h3a7c234e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39583378),
	.w1(32'h38072b55),
	.w2(32'hba0e39a0),
	.w3(32'hb5fc7596),
	.w4(32'h3996da91),
	.w5(32'hb989d525),
	.w6(32'h3a0f43f9),
	.w7(32'h39fb2cf1),
	.w8(32'hb955dd5a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04cc49),
	.w1(32'hbb2edee4),
	.w2(32'hba02c87d),
	.w3(32'hbaf28956),
	.w4(32'hba74564d),
	.w5(32'h38244c12),
	.w6(32'hbabe9ab9),
	.w7(32'h39dac220),
	.w8(32'hb93f1ce7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f48abf),
	.w1(32'h3b4ee684),
	.w2(32'h3a12aaae),
	.w3(32'h3b797080),
	.w4(32'h3b863f1d),
	.w5(32'h39fdfb97),
	.w6(32'h3b74b78b),
	.w7(32'h3a546737),
	.w8(32'hba595ffa),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391df6b4),
	.w1(32'h39474e11),
	.w2(32'h37f0c6d7),
	.w3(32'h39096a67),
	.w4(32'h38638ba8),
	.w5(32'hb7eec961),
	.w6(32'h38adfa28),
	.w7(32'hb808f0ce),
	.w8(32'h38283e42),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d028f),
	.w1(32'h39715dd2),
	.w2(32'h3937f4f5),
	.w3(32'h39822219),
	.w4(32'h38f85d24),
	.w5(32'hb7c598f6),
	.w6(32'h3940a2a8),
	.w7(32'h38fcde21),
	.w8(32'h381e105d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dca04d),
	.w1(32'h36d4ae8c),
	.w2(32'h37ba0050),
	.w3(32'h377cc47c),
	.w4(32'h3790d4bc),
	.w5(32'h37b5bfa3),
	.w6(32'h3816c9a9),
	.w7(32'h38301a6b),
	.w8(32'h38123d9d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dda5f3),
	.w1(32'h3993eea6),
	.w2(32'h38d72837),
	.w3(32'h3a800639),
	.w4(32'h3a445b3c),
	.w5(32'h393c6c1c),
	.w6(32'h3a800de1),
	.w7(32'h3a50a795),
	.w8(32'h3a197969),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba650c7a),
	.w1(32'hbb8005f9),
	.w2(32'hbaaeeb4a),
	.w3(32'h3b17d285),
	.w4(32'hbae104a2),
	.w5(32'hbafede42),
	.w6(32'hb9b92eef),
	.w7(32'h3a4f2efa),
	.w8(32'h393548f7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c986d),
	.w1(32'hbb3a3cc5),
	.w2(32'hba98879d),
	.w3(32'hbb4d0652),
	.w4(32'hbb3962a3),
	.w5(32'hba8f7e0f),
	.w6(32'hb99c4e2a),
	.w7(32'hba416560),
	.w8(32'hbab1c75d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1a21b),
	.w1(32'hba859927),
	.w2(32'hba53c86d),
	.w3(32'hb9f985f0),
	.w4(32'hb9e9cd82),
	.w5(32'hb9bea56e),
	.w6(32'hb98163fd),
	.w7(32'hb9a84e33),
	.w8(32'hba18d468),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2146e0),
	.w1(32'hbb1668cb),
	.w2(32'hb9f2ca81),
	.w3(32'hba3d1f3f),
	.w4(32'hba5010b2),
	.w5(32'h38f8c505),
	.w6(32'hbab0eb4f),
	.w7(32'hba845f7e),
	.w8(32'hba5b156f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0242ad),
	.w1(32'h3a1e9877),
	.w2(32'h395f40ad),
	.w3(32'h3a817e2c),
	.w4(32'h3a5e3a17),
	.w5(32'h3a168d38),
	.w6(32'h3a6f9f9e),
	.w7(32'h3a03471f),
	.w8(32'h39b34863),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae67089),
	.w1(32'hba37f2da),
	.w2(32'h3951e6ba),
	.w3(32'hbaaa5f48),
	.w4(32'hba6fb92a),
	.w5(32'h39f3096b),
	.w6(32'hb8f7ca27),
	.w7(32'hb8f51517),
	.w8(32'h398a9ac6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b5c23),
	.w1(32'h3a2660a2),
	.w2(32'h3b281f6c),
	.w3(32'hba883a81),
	.w4(32'h3adb120c),
	.w5(32'h3b463627),
	.w6(32'h3a2fdd72),
	.w7(32'h3a8e8541),
	.w8(32'h3adf3312),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe72e4a),
	.w1(32'hbbed86e8),
	.w2(32'hbb8c054f),
	.w3(32'hbbb287fe),
	.w4(32'hbb637f07),
	.w5(32'hba5d6fdd),
	.w6(32'hbb7df2f3),
	.w7(32'hbb4c9e39),
	.w8(32'hbb833593),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b836e),
	.w1(32'h3a972f45),
	.w2(32'hba919746),
	.w3(32'h3b158332),
	.w4(32'h3ab672e3),
	.w5(32'hba76d1f6),
	.w6(32'h3ab9ef82),
	.w7(32'h3a08d5be),
	.w8(32'hba4f5849),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d033c),
	.w1(32'hbb1c3c42),
	.w2(32'hbad1b411),
	.w3(32'hbb128ae5),
	.w4(32'hb9cc4914),
	.w5(32'hb92118fb),
	.w6(32'hba9ffafb),
	.w7(32'h3a582ce6),
	.w8(32'h3a140359),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0aaa6),
	.w1(32'hbb9ff4ad),
	.w2(32'hba93d1f1),
	.w3(32'hbb87a27f),
	.w4(32'hba20116f),
	.w5(32'h3aba4924),
	.w6(32'hba1cc272),
	.w7(32'h39af5823),
	.w8(32'h39285d00),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdf646),
	.w1(32'hba5924ac),
	.w2(32'h37e0bc7f),
	.w3(32'h3a7cee30),
	.w4(32'h3af153a9),
	.w5(32'h39955641),
	.w6(32'hba5622cb),
	.w7(32'h3a2fb5c5),
	.w8(32'h3aa17f66),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac05e6d),
	.w1(32'hbb0bc6ac),
	.w2(32'hba94fd87),
	.w3(32'hbabd82d2),
	.w4(32'hba9db5e6),
	.w5(32'hba96c02b),
	.w6(32'hb8e4a891),
	.w7(32'h3a1c3846),
	.w8(32'hbacb0fdb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913a198),
	.w1(32'h3781798a),
	.w2(32'hb9492a17),
	.w3(32'h37720e21),
	.w4(32'h39486d3b),
	.w5(32'hb98ff905),
	.w6(32'h392e134d),
	.w7(32'h3a074a9d),
	.w8(32'hb927cf50),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b49c8),
	.w1(32'h3a09428c),
	.w2(32'hb9e9d3db),
	.w3(32'h3b9de745),
	.w4(32'h3b8b4ef2),
	.w5(32'h399ff585),
	.w6(32'h3b409978),
	.w7(32'h3b013266),
	.w8(32'hbaa66d80),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafafa22),
	.w1(32'hba96b8d8),
	.w2(32'hba1bf5dc),
	.w3(32'hbb0213a0),
	.w4(32'hb9f6c397),
	.w5(32'h3a15f3a3),
	.w6(32'hbb311c06),
	.w7(32'hb8dd3902),
	.w8(32'h37abb5ba),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb852cbc6),
	.w1(32'hb88f6efe),
	.w2(32'h388c738d),
	.w3(32'hb846187b),
	.w4(32'hb798f233),
	.w5(32'h3833bf36),
	.w6(32'hb8215b2a),
	.w7(32'h382b7a59),
	.w8(32'h38e679c9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8351a30),
	.w1(32'hb864e005),
	.w2(32'h363aa403),
	.w3(32'h36f74cdc),
	.w4(32'h351a5bb0),
	.w5(32'h36e57727),
	.w6(32'h37220298),
	.w7(32'hb84d80f8),
	.w8(32'hb50e6597),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97bafd),
	.w1(32'hbab31d47),
	.w2(32'hba15d1ad),
	.w3(32'hba327417),
	.w4(32'hba7b83f2),
	.w5(32'hba9c8fcb),
	.w6(32'h39106aae),
	.w7(32'h38b0e1ab),
	.w8(32'hb96c3016),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf8df7),
	.w1(32'hba885013),
	.w2(32'hbb6ccdaf),
	.w3(32'hb99eb377),
	.w4(32'hb9cb73e6),
	.w5(32'hbb08d9c3),
	.w6(32'hbaeb3034),
	.w7(32'hbb14d7dc),
	.w8(32'hba9b4669),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845f25),
	.w1(32'hba4863f2),
	.w2(32'h394d7f82),
	.w3(32'h3a0af840),
	.w4(32'hb9f9ceb5),
	.w5(32'hbaa65447),
	.w6(32'h3b333ccb),
	.w7(32'h3a34f5a2),
	.w8(32'hba15bd69),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86dc625),
	.w1(32'hb846bd59),
	.w2(32'hb65ff00e),
	.w3(32'hb8002dc7),
	.w4(32'hb7cc5338),
	.w5(32'h3637ae47),
	.w6(32'h36502ffc),
	.w7(32'hb7cedc27),
	.w8(32'hb7cd5833),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd66d7),
	.w1(32'hbb098e03),
	.w2(32'hba533458),
	.w3(32'hbac72d71),
	.w4(32'hbb0d3c5c),
	.w5(32'hbad668cd),
	.w6(32'h3a2c6225),
	.w7(32'h3a160cf3),
	.w8(32'hbaf393c4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e00f1c),
	.w1(32'hba2cd869),
	.w2(32'h382aefb3),
	.w3(32'h3a525b65),
	.w4(32'hb9181265),
	.w5(32'hbadbe543),
	.w6(32'h3a95c319),
	.w7(32'h3aa4d5e2),
	.w8(32'hba648b4d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb630d0c),
	.w1(32'hbb7ba58b),
	.w2(32'hbb335ffc),
	.w3(32'hbab93358),
	.w4(32'hba3e60a8),
	.w5(32'hbad1d4a5),
	.w6(32'hb96b369a),
	.w7(32'h3a3fe16c),
	.w8(32'hba2323c2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68fffa),
	.w1(32'h3b188883),
	.w2(32'h3aa03d86),
	.w3(32'hba664339),
	.w4(32'h3b0c2bb5),
	.w5(32'h3a9fd423),
	.w6(32'h3a92b9b7),
	.w7(32'hb91e5285),
	.w8(32'hb9c5d0c1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948ca7e),
	.w1(32'h3a202cd7),
	.w2(32'hb8f98a2f),
	.w3(32'h38d5ca33),
	.w4(32'h3a56b1cc),
	.w5(32'h3a450dbb),
	.w6(32'h3993dcf4),
	.w7(32'hb94206d6),
	.w8(32'h38fe71ac),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba0152),
	.w1(32'h3a051162),
	.w2(32'h3a3d3d15),
	.w3(32'h39d5c450),
	.w4(32'h3a364b3a),
	.w5(32'h3a51c78f),
	.w6(32'h39f0336d),
	.w7(32'h3a1c9713),
	.w8(32'h3a46dbd7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2a51c),
	.w1(32'hb7d50292),
	.w2(32'hb952145e),
	.w3(32'h3a7e5945),
	.w4(32'h3af34465),
	.w5(32'hb94d15ab),
	.w6(32'h38592338),
	.w7(32'h3b07c54d),
	.w8(32'h3a59f3a9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3609ac),
	.w1(32'hb979f7fb),
	.w2(32'h38fa50fd),
	.w3(32'hba91b17b),
	.w4(32'h3916d496),
	.w5(32'h3a1d53cf),
	.w6(32'h38ed98f4),
	.w7(32'hba5ec7a8),
	.w8(32'hb952ea57),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b102fc0),
	.w1(32'h3b1d90f7),
	.w2(32'h3a9dbe23),
	.w3(32'h3b2b0155),
	.w4(32'h3b183637),
	.w5(32'h3acc6fe1),
	.w6(32'h3ae82aab),
	.w7(32'h3a52df14),
	.w8(32'h3989095f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb7e13),
	.w1(32'hbad95353),
	.w2(32'hba28e13a),
	.w3(32'hbad1ac32),
	.w4(32'hba822060),
	.w5(32'h38e118e3),
	.w6(32'hba803204),
	.w7(32'hb9d00833),
	.w8(32'h38887781),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933c7d0),
	.w1(32'h393c5014),
	.w2(32'hb6f47bdd),
	.w3(32'h39f76269),
	.w4(32'h3a0e20e1),
	.w5(32'h398c862b),
	.w6(32'h39d24030),
	.w7(32'h39dcb07a),
	.w8(32'h38a5db01),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45b045),
	.w1(32'hbba03a8e),
	.w2(32'hbafa3b58),
	.w3(32'hbb370071),
	.w4(32'hbb162d7b),
	.w5(32'h398a7df1),
	.w6(32'hbaaef92c),
	.w7(32'h39d723ea),
	.w8(32'h3a34efdf),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394054f5),
	.w1(32'hb8899bbb),
	.w2(32'hb913597b),
	.w3(32'h380d2511),
	.w4(32'h38ed6d21),
	.w5(32'hb982144f),
	.w6(32'h393d3af4),
	.w7(32'h3a01fef0),
	.w8(32'h398f12ae),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d0cf),
	.w1(32'hba82db9e),
	.w2(32'hba035de0),
	.w3(32'hba31b053),
	.w4(32'h3aa7d568),
	.w5(32'h3963f8b9),
	.w6(32'hba637c29),
	.w7(32'h3aee5c7b),
	.w8(32'h3a303c78),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39975993),
	.w1(32'h39aefad5),
	.w2(32'h393d8655),
	.w3(32'h3963157c),
	.w4(32'h38c3ee94),
	.w5(32'h39013132),
	.w6(32'h393cdf9b),
	.w7(32'h391b4462),
	.w8(32'h39213a90),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ce1f2),
	.w1(32'h39e46b8e),
	.w2(32'h3a912dfa),
	.w3(32'h3b96dbfe),
	.w4(32'h3aaf24c5),
	.w5(32'h3a5d1fb5),
	.w6(32'h3b5f56c6),
	.w7(32'hb9b110e8),
	.w8(32'hba882ce4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895a8e5),
	.w1(32'hb857ac4e),
	.w2(32'hb92397b5),
	.w3(32'hb8c3b02c),
	.w4(32'hb8ed9fa5),
	.w5(32'hb9603607),
	.w6(32'hb840d4b4),
	.w7(32'h3839f150),
	.w8(32'hb8c02b80),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39450425),
	.w1(32'hb98417bc),
	.w2(32'hba286169),
	.w3(32'h380b239f),
	.w4(32'hb9b2059b),
	.w5(32'hba49075b),
	.w6(32'h391befd5),
	.w7(32'hb9d53064),
	.w8(32'hba73f178),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1947e3),
	.w1(32'h3a541e27),
	.w2(32'hbabba68b),
	.w3(32'h3a4a6be8),
	.w4(32'h3a9cfa60),
	.w5(32'hba79e9cc),
	.w6(32'hb8f07b75),
	.w7(32'h3a27008b),
	.w8(32'h39854638),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc0eb),
	.w1(32'hbb07f9d2),
	.w2(32'hba669953),
	.w3(32'hba8afad7),
	.w4(32'hba835321),
	.w5(32'hba42d150),
	.w6(32'hbb93d693),
	.w7(32'hba983972),
	.w8(32'hbb15a70d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa06eb),
	.w1(32'h3aa7c052),
	.w2(32'h3aa9d0cb),
	.w3(32'h3aad9139),
	.w4(32'h3a8316a0),
	.w5(32'h3a965dfe),
	.w6(32'h3a5e1014),
	.w7(32'h3a03711c),
	.w8(32'h39d0e2f3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97223da),
	.w1(32'h3ad587aa),
	.w2(32'hba3dbde4),
	.w3(32'h3acc8f59),
	.w4(32'h3b1bef67),
	.w5(32'hbadc1c23),
	.w6(32'h3b33c826),
	.w7(32'h3b27561b),
	.w8(32'hba0093ce),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f31e25),
	.w1(32'h3abb3f8b),
	.w2(32'h3a382af8),
	.w3(32'hb8c4b0ed),
	.w4(32'hb88c79ba),
	.w5(32'h39b1c905),
	.w6(32'hb917d328),
	.w7(32'hba5b0824),
	.w8(32'hba3583fc),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc985ce),
	.w1(32'h3907cf3c),
	.w2(32'h399d8507),
	.w3(32'hbb106b10),
	.w4(32'h3a9bf340),
	.w5(32'hba040750),
	.w6(32'h39b050f5),
	.w7(32'hba0f1521),
	.w8(32'hbb3bc1b8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5dd7e),
	.w1(32'hbb10a131),
	.w2(32'hbab8a212),
	.w3(32'hba887887),
	.w4(32'hbaae11b9),
	.w5(32'hb9b09bff),
	.w6(32'hb8d19721),
	.w7(32'h392b6237),
	.w8(32'hb9443121),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd17f3),
	.w1(32'hbb5f404e),
	.w2(32'hbaf7deaa),
	.w3(32'hbb91a871),
	.w4(32'hbb02044d),
	.w5(32'hbac39eb7),
	.w6(32'hbae9f1f3),
	.w7(32'h3a017ac9),
	.w8(32'hbaf09e3b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e7227),
	.w1(32'h391071e6),
	.w2(32'hb80115aa),
	.w3(32'hb7b1527d),
	.w4(32'h38c43c48),
	.w5(32'h39a99f05),
	.w6(32'hba1390ff),
	.w7(32'hb8d47a98),
	.w8(32'h39d69b4b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c041),
	.w1(32'hba98d7a7),
	.w2(32'hba7e32be),
	.w3(32'hbb36b2e8),
	.w4(32'hb9b9b5e4),
	.w5(32'hba4871c2),
	.w6(32'hba9bd68f),
	.w7(32'h388dfa09),
	.w8(32'hbad08983),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3725d1c5),
	.w1(32'hb6ec353e),
	.w2(32'h38ac05ec),
	.w3(32'h37b4f1f8),
	.w4(32'h36832e8d),
	.w5(32'h3886c019),
	.w6(32'h38187f36),
	.w7(32'h37836272),
	.w8(32'h38927078),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c9d3b),
	.w1(32'hb88e0406),
	.w2(32'h3a0a7c8e),
	.w3(32'hba290d44),
	.w4(32'h367c550b),
	.w5(32'h39f77f78),
	.w6(32'hb9a7a079),
	.w7(32'hb7e397cf),
	.w8(32'h396bb933),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba348d8e),
	.w1(32'hb9b7cc6b),
	.w2(32'hb9c939e8),
	.w3(32'h393fb781),
	.w4(32'h38e8d50c),
	.w5(32'hb99a70c1),
	.w6(32'h36ca5c6a),
	.w7(32'hb9882ed3),
	.w8(32'hba032885),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c9d43),
	.w1(32'hba927234),
	.w2(32'hba9f9137),
	.w3(32'hbb13b0c9),
	.w4(32'hba85b25d),
	.w5(32'hbaa0d1fd),
	.w6(32'hb981b7df),
	.w7(32'hbae77ae7),
	.w8(32'hbb144141),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8007c23),
	.w1(32'hb74ad80b),
	.w2(32'hb73d288a),
	.w3(32'hb74d2705),
	.w4(32'h369cf8f0),
	.w5(32'h3777370a),
	.w6(32'h36a63380),
	.w7(32'hb782a997),
	.w8(32'h35f29f2a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ef9de),
	.w1(32'hb9872495),
	.w2(32'hb99c1533),
	.w3(32'hb9897b7d),
	.w4(32'hb8ba9528),
	.w5(32'hb89071d9),
	.w6(32'hb95db1bd),
	.w7(32'h3713b3bc),
	.w8(32'h3637b98d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d5e91),
	.w1(32'h384f1541),
	.w2(32'h3a11b50a),
	.w3(32'h3a45f9c6),
	.w4(32'h3abe16ec),
	.w5(32'h3a240080),
	.w6(32'hb9f52bfc),
	.w7(32'h399aa2d7),
	.w8(32'hb9a473ca),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1321b),
	.w1(32'hbb2b3109),
	.w2(32'hbb0041b1),
	.w3(32'h3b41a47c),
	.w4(32'h3a74bb9e),
	.w5(32'h39d7f867),
	.w6(32'h3a305327),
	.w7(32'hbae563bf),
	.w8(32'hbb447df4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cddf2),
	.w1(32'hb926f554),
	.w2(32'h383c963c),
	.w3(32'hbaad8d56),
	.w4(32'h39cb65a3),
	.w5(32'h38789ab5),
	.w6(32'hb8889255),
	.w7(32'h3ac5cd0a),
	.w8(32'hb9421eb5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce7d3b),
	.w1(32'hba683925),
	.w2(32'hba030a49),
	.w3(32'hb9ec8749),
	.w4(32'hb95f2252),
	.w5(32'hb9d110df),
	.w6(32'hba77977a),
	.w7(32'hba1c3d55),
	.w8(32'hba70828a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc313112),
	.w1(32'hbc2a0c8f),
	.w2(32'hbbc51d5e),
	.w3(32'hbb506021),
	.w4(32'hbb5ef7b0),
	.w5(32'hbbccdfea),
	.w6(32'h38f024b0),
	.w7(32'hb8927be6),
	.w8(32'hbbde2b78),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57d267),
	.w1(32'h3b4efed9),
	.w2(32'h3b2354fa),
	.w3(32'hbae877ab),
	.w4(32'h3b7b0f1e),
	.w5(32'h3b4273f4),
	.w6(32'h3a9d0583),
	.w7(32'h3b2e8ecb),
	.w8(32'h38f9c602),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ac698),
	.w1(32'hb8ec2f58),
	.w2(32'h3a1c09b8),
	.w3(32'h39b93066),
	.w4(32'hb912699b),
	.w5(32'hb50f9902),
	.w6(32'h3a875bee),
	.w7(32'h3a15b683),
	.w8(32'hb9a89b15),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810e366),
	.w1(32'hb7adb5fa),
	.w2(32'hb706a1a3),
	.w3(32'hb8710afb),
	.w4(32'hb7f90bef),
	.w5(32'hb823cfb2),
	.w6(32'hb807a182),
	.w7(32'hb7afbb9b),
	.w8(32'hb8889638),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96751aa),
	.w1(32'hb881c656),
	.w2(32'hb8f9fb85),
	.w3(32'hb995af46),
	.w4(32'h378f31e7),
	.w5(32'hb890d83f),
	.w6(32'hb98b449e),
	.w7(32'h382d084f),
	.w8(32'h383367de),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c571cd),
	.w1(32'h371a262f),
	.w2(32'h372f44e6),
	.w3(32'h375f9cea),
	.w4(32'h370ff256),
	.w5(32'hb6a40ecc),
	.w6(32'h37ab3956),
	.w7(32'h377fbae8),
	.w8(32'h36d57441),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b0f91),
	.w1(32'h3a3ce89a),
	.w2(32'h3a76c6e3),
	.w3(32'h3ac1c01e),
	.w4(32'h3aab61b0),
	.w5(32'h39f8e347),
	.w6(32'h3a6a3c8e),
	.w7(32'h3af92a2f),
	.w8(32'hb808a588),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6b1a7),
	.w1(32'hba5b2e32),
	.w2(32'hba5272da),
	.w3(32'hb97c0a1c),
	.w4(32'hb99c72a5),
	.w5(32'h3a702b4f),
	.w6(32'hba92e361),
	.w7(32'hbac5c8bf),
	.w8(32'hba5413ab),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad53d75),
	.w1(32'h3abb455e),
	.w2(32'hb9913e03),
	.w3(32'h3b347047),
	.w4(32'h3b0650d4),
	.w5(32'hba1fa4f8),
	.w6(32'h3b0ef594),
	.w7(32'h3a8addea),
	.w8(32'hb92a70a3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931cad2),
	.w1(32'hba012d2a),
	.w2(32'h37da9b3d),
	.w3(32'h39ab53a8),
	.w4(32'h399f3b35),
	.w5(32'h39830334),
	.w6(32'hba0b7898),
	.w7(32'hb90f0aa3),
	.w8(32'hb8a47a8d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2f98a),
	.w1(32'hbc031375),
	.w2(32'hbc11aa91),
	.w3(32'h3909ec59),
	.w4(32'hb98ab30c),
	.w5(32'hbc4c94d5),
	.w6(32'h3b1393fb),
	.w7(32'h3aab4ba5),
	.w8(32'hbc3a9ef8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95ced9),
	.w1(32'h3a1cbbd1),
	.w2(32'h3915c2d4),
	.w3(32'hbbabbd56),
	.w4(32'hb97aab1d),
	.w5(32'hbbf7a137),
	.w6(32'hbbc024b4),
	.w7(32'hbabc5048),
	.w8(32'hbb15e74a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab656c4),
	.w1(32'hbbc63daf),
	.w2(32'hbb0342cf),
	.w3(32'h3b286b28),
	.w4(32'hba12b7bc),
	.w5(32'hbb980be8),
	.w6(32'h3bdb268e),
	.w7(32'hbbc665b6),
	.w8(32'hbba969e8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1cd5f),
	.w1(32'hbb269adf),
	.w2(32'hbb01df38),
	.w3(32'hbaa30daa),
	.w4(32'hbbea8681),
	.w5(32'h39b9e237),
	.w6(32'hbba61f1e),
	.w7(32'hbb89e6f8),
	.w8(32'hbba5c80e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf563fa),
	.w1(32'hbbdc07cb),
	.w2(32'hba72bc18),
	.w3(32'hbb75105c),
	.w4(32'hba3a6bcc),
	.w5(32'h3b2ba057),
	.w6(32'hbb6b65de),
	.w7(32'hbacb069e),
	.w8(32'h3b11840a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b09af),
	.w1(32'h3a8095a8),
	.w2(32'hbbb5ee63),
	.w3(32'h3b86edd5),
	.w4(32'h3a9394e7),
	.w5(32'hbb6933e0),
	.w6(32'hbac2b528),
	.w7(32'hbbbfc818),
	.w8(32'hbc28eb9d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef0634),
	.w1(32'hbad85a5e),
	.w2(32'h3a518f7c),
	.w3(32'h3b3ebf65),
	.w4(32'h3b137501),
	.w5(32'hb88942ce),
	.w6(32'hbae2f839),
	.w7(32'hbb1deb3c),
	.w8(32'hbbbb47b6),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b5d15),
	.w1(32'hbb3c5fe9),
	.w2(32'hbaabef51),
	.w3(32'h3b9d3820),
	.w4(32'hbb9e3cab),
	.w5(32'hba9365f2),
	.w6(32'h3b14f090),
	.w7(32'hbba417a5),
	.w8(32'hbb94dc42),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98bf51),
	.w1(32'h3b100c5b),
	.w2(32'hbbc8cafb),
	.w3(32'hbb0ebfbd),
	.w4(32'hbb1af28c),
	.w5(32'hbbd57860),
	.w6(32'hbaeb65ba),
	.w7(32'h3aa46fb7),
	.w8(32'hbc143cfd),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c99fa),
	.w1(32'h3b71fff9),
	.w2(32'h3b19efef),
	.w3(32'h3aab646a),
	.w4(32'h3b8ef60f),
	.w5(32'h3b8903af),
	.w6(32'hbb127ec3),
	.w7(32'h3b930d97),
	.w8(32'h3ba48948),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b1684),
	.w1(32'hbb8721ac),
	.w2(32'h3aa75805),
	.w3(32'hbc3575db),
	.w4(32'hbb7c9059),
	.w5(32'hbbf2626e),
	.w6(32'hbbecab8d),
	.w7(32'hba855910),
	.w8(32'hbb8cd776),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19c5bd),
	.w1(32'hbb765259),
	.w2(32'h3b5c4fb8),
	.w3(32'hba3062d2),
	.w4(32'h3b6d29f1),
	.w5(32'h3c6d3834),
	.w6(32'h3b453541),
	.w7(32'h3880dae4),
	.w8(32'h3b24f59e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bac57),
	.w1(32'hbad53bc0),
	.w2(32'hba59925d),
	.w3(32'hbaa796c1),
	.w4(32'hbb285cec),
	.w5(32'hbb507a0e),
	.w6(32'hbb1d3364),
	.w7(32'hbaa5432d),
	.w8(32'hbbb226f5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf2ed5),
	.w1(32'h3a62c90e),
	.w2(32'hbb419c3e),
	.w3(32'h3afcee09),
	.w4(32'h3b103686),
	.w5(32'h3aec2e8b),
	.w6(32'h3b1409ab),
	.w7(32'hbb036d19),
	.w8(32'hbb23b95d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb913fba),
	.w1(32'hbba7c533),
	.w2(32'hb9be277a),
	.w3(32'h3b99f5e2),
	.w4(32'h3baa07f9),
	.w5(32'hbb9c50bc),
	.w6(32'hba38fe48),
	.w7(32'hbb2ae5e3),
	.w8(32'hbac144db),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f420a),
	.w1(32'hbbae591f),
	.w2(32'hbbd04059),
	.w3(32'hbc0cbd89),
	.w4(32'hbaea427c),
	.w5(32'h3aaf60eb),
	.w6(32'hbc5ddece),
	.w7(32'h39099f5f),
	.w8(32'hbbc078d5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9331972),
	.w1(32'hbbb0bcf6),
	.w2(32'hbc0ece3d),
	.w3(32'h3b0704b5),
	.w4(32'hbbda876f),
	.w5(32'hbb930974),
	.w6(32'h3aa46912),
	.w7(32'hbac7ab86),
	.w8(32'h3a6c1085),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aa118),
	.w1(32'hbb0fce40),
	.w2(32'hb9b76f99),
	.w3(32'h3b6207f8),
	.w4(32'h3be8f069),
	.w5(32'h3c4b13ab),
	.w6(32'h3b6de564),
	.w7(32'hbb94ce3f),
	.w8(32'hba687cd1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72218c),
	.w1(32'hb986bff5),
	.w2(32'hbbab3f4b),
	.w3(32'hbb961aca),
	.w4(32'h3bdbd4c5),
	.w5(32'h3abcdab0),
	.w6(32'h3a262591),
	.w7(32'hb94f2d70),
	.w8(32'h3a0667f5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5300ea),
	.w1(32'hbb12486b),
	.w2(32'hb9aeedde),
	.w3(32'h3b916bd4),
	.w4(32'h398b58f8),
	.w5(32'hbbfa9354),
	.w6(32'h3b9aa96f),
	.w7(32'hbbdc5127),
	.w8(32'hbb946ccd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf4e38),
	.w1(32'h3be3f506),
	.w2(32'h3b8928f1),
	.w3(32'h3a28fa4c),
	.w4(32'h3aff305a),
	.w5(32'hbb4f8799),
	.w6(32'h3b4fa203),
	.w7(32'h3bf2f4f4),
	.w8(32'h3b141f49),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe36ef6),
	.w1(32'hbbd30ac8),
	.w2(32'hbba86e57),
	.w3(32'hbbc05692),
	.w4(32'h3b33089f),
	.w5(32'hbad11158),
	.w6(32'h3b27154a),
	.w7(32'hbaba1d15),
	.w8(32'hbb121e9f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f49d6b),
	.w1(32'hbb82763f),
	.w2(32'hba49c001),
	.w3(32'h39ae8d80),
	.w4(32'hbb61ae83),
	.w5(32'hbba1eedc),
	.w6(32'h3b6cabe6),
	.w7(32'h3a5dd8a7),
	.w8(32'hba4eba52),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf375d),
	.w1(32'h3a7caf93),
	.w2(32'hbac144ca),
	.w3(32'hbab5cbac),
	.w4(32'h3bd3386f),
	.w5(32'h3c0fc033),
	.w6(32'hbb829911),
	.w7(32'hbbc98ae8),
	.w8(32'hbb1a27c5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0252f),
	.w1(32'hbb258e07),
	.w2(32'hbb8bb8c4),
	.w3(32'h3bb08622),
	.w4(32'h3b202d63),
	.w5(32'h3b4c377f),
	.w6(32'hbb7c0694),
	.w7(32'hb9ec58d6),
	.w8(32'hbb6239b2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc65a0),
	.w1(32'h3be828f8),
	.w2(32'h3af11fe9),
	.w3(32'h3b001e5c),
	.w4(32'h3b021bb5),
	.w5(32'hbbb9a8bd),
	.w6(32'hba0fd3d4),
	.w7(32'hbb551239),
	.w8(32'hbbe018a6),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe00df0),
	.w1(32'hbb703a5c),
	.w2(32'hba9523b7),
	.w3(32'h3b3d0070),
	.w4(32'hbba7623c),
	.w5(32'h3b653572),
	.w6(32'hbbc4e6cf),
	.w7(32'hbbcda11f),
	.w8(32'h3bcd93f9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96166f),
	.w1(32'hbb6db76f),
	.w2(32'hb9db9f5c),
	.w3(32'h3b89b8c0),
	.w4(32'hba999ff6),
	.w5(32'hbbb73234),
	.w6(32'hb93ee33e),
	.w7(32'hbb88d03b),
	.w8(32'hbb0dcdff),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7faf2e),
	.w1(32'h3be7ec5c),
	.w2(32'h3b8ce5d3),
	.w3(32'h3b409665),
	.w4(32'h3be4fbdd),
	.w5(32'h3b5bb32f),
	.w6(32'hbac48126),
	.w7(32'h3b6578fb),
	.w8(32'h3c00b1d0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd1f60),
	.w1(32'hba0a039c),
	.w2(32'h3afcb210),
	.w3(32'hbc3bab0e),
	.w4(32'hbac9615f),
	.w5(32'hbc0e3b63),
	.w6(32'hb99356fe),
	.w7(32'h3ba0c9db),
	.w8(32'h3bd398d2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ec7b3),
	.w1(32'hbb884d31),
	.w2(32'hbb0d58ed),
	.w3(32'h38e4e2ef),
	.w4(32'hba26515f),
	.w5(32'hbc482e22),
	.w6(32'h3b8fda42),
	.w7(32'h3bedf453),
	.w8(32'h3b042d94),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998d5a5),
	.w1(32'hbb289cec),
	.w2(32'hbaaa997f),
	.w3(32'hbb4c79a0),
	.w4(32'h3b69b4f3),
	.w5(32'hbb56fc28),
	.w6(32'h3a78076c),
	.w7(32'hba958a1a),
	.w8(32'hbb59b5e9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1c23),
	.w1(32'hbb81467f),
	.w2(32'h3b606bfe),
	.w3(32'h3b81c418),
	.w4(32'hbb350e58),
	.w5(32'h3bbf2a51),
	.w6(32'hbb6c15d7),
	.w7(32'hbb75ee47),
	.w8(32'h3b699e96),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95f279),
	.w1(32'hbc1a0381),
	.w2(32'hbb7efa4b),
	.w3(32'h3b8864bf),
	.w4(32'hbb8308cd),
	.w5(32'hbb9db9dc),
	.w6(32'h3ab40541),
	.w7(32'hbad07893),
	.w8(32'hbc0bb55d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffd429),
	.w1(32'h399ec717),
	.w2(32'h3b17d7f8),
	.w3(32'hbae1cced),
	.w4(32'hbb1ed1b7),
	.w5(32'h3b970cb1),
	.w6(32'hbb71dbd9),
	.w7(32'hbb8d64a3),
	.w8(32'h3bdd257b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba54119),
	.w1(32'h3b497f08),
	.w2(32'h3b785159),
	.w3(32'hbb645641),
	.w4(32'h3b401f10),
	.w5(32'hba649cdc),
	.w6(32'hbb136bf4),
	.w7(32'hbb6b1f96),
	.w8(32'hbb2ecadf),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ddf19),
	.w1(32'hbbd13917),
	.w2(32'hbb260871),
	.w3(32'hbb54f0d5),
	.w4(32'hba0f3e4f),
	.w5(32'hba92aa9e),
	.w6(32'hbb2cf8c2),
	.w7(32'hba0f9bef),
	.w8(32'hba19b31f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e71c2),
	.w1(32'h3aaac103),
	.w2(32'hbb539cfd),
	.w3(32'hbab0b472),
	.w4(32'hbb373df6),
	.w5(32'hba842a9f),
	.w6(32'hba3c34df),
	.w7(32'hb9892556),
	.w8(32'hbb9f46d2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba006c5),
	.w1(32'hbaae049e),
	.w2(32'hbb44fb25),
	.w3(32'h3b9f7eac),
	.w4(32'h3b4c7102),
	.w5(32'hbb813ed5),
	.w6(32'h3be95f2d),
	.w7(32'hbadcda1e),
	.w8(32'hbae45f4f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38081bb2),
	.w1(32'hbb218b9b),
	.w2(32'hbac0259c),
	.w3(32'h3a91e9f5),
	.w4(32'h3ae14927),
	.w5(32'h3c26b195),
	.w6(32'hba413188),
	.w7(32'hbb643a96),
	.w8(32'hba89bc95),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ea41),
	.w1(32'hbab1f15c),
	.w2(32'hbaedb176),
	.w3(32'h39cf4cba),
	.w4(32'hbb309ebe),
	.w5(32'h3b959e43),
	.w6(32'hbb39cb97),
	.w7(32'hbbbace21),
	.w8(32'hba8a5778),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807616),
	.w1(32'hba056dba),
	.w2(32'hba3ec016),
	.w3(32'h3b22aa8e),
	.w4(32'hbb7a3af0),
	.w5(32'hba9dea41),
	.w6(32'hbb870dc8),
	.w7(32'hbad21d45),
	.w8(32'h3b585e08),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb2f8),
	.w1(32'hbb97fa1b),
	.w2(32'h39890054),
	.w3(32'hbbde11e7),
	.w4(32'hbba8b9b3),
	.w5(32'hbbcd27cb),
	.w6(32'hbb0e0a6c),
	.w7(32'hba98564b),
	.w8(32'hba3ba923),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943452f),
	.w1(32'hbbed9a5f),
	.w2(32'hbaebefd0),
	.w3(32'h3b5e66e5),
	.w4(32'hba905766),
	.w5(32'hb96cd960),
	.w6(32'h3bce5536),
	.w7(32'h3b33c795),
	.w8(32'h3b7b1cc7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4062f9),
	.w1(32'hbc28a636),
	.w2(32'hbbc9c708),
	.w3(32'h3ad8de27),
	.w4(32'hbc2ec3c8),
	.w5(32'hbb309c2c),
	.w6(32'hbb204526),
	.w7(32'hbbee4f07),
	.w8(32'hbbc2de0a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba428f9),
	.w1(32'hbaffde52),
	.w2(32'hbb3489df),
	.w3(32'hb9823bc4),
	.w4(32'h3aab1715),
	.w5(32'h3aa956c3),
	.w6(32'hbc120f36),
	.w7(32'hba5b4ef0),
	.w8(32'h3b88ce7a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe87a7e),
	.w1(32'hbb41234e),
	.w2(32'hbaa1ab15),
	.w3(32'hbc102ce2),
	.w4(32'hbad6f702),
	.w5(32'hbba24ba9),
	.w6(32'hbc25b3ca),
	.w7(32'hba9c8102),
	.w8(32'hbbd9c9c6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ce115),
	.w1(32'hbb32a796),
	.w2(32'hbb45c172),
	.w3(32'hbbbbbc21),
	.w4(32'hbb1a6a6c),
	.w5(32'h3b8793e1),
	.w6(32'hbbff8572),
	.w7(32'hbb8ff5c2),
	.w8(32'hbae670af),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba949227),
	.w1(32'hbb9e9741),
	.w2(32'hbb8541f0),
	.w3(32'hbac50ae6),
	.w4(32'h3ae22fc7),
	.w5(32'h3b954298),
	.w6(32'hbb8ca6b6),
	.w7(32'h3a38fc18),
	.w8(32'hbaa5c6c9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c7f1a),
	.w1(32'hbba9d8ea),
	.w2(32'hbba0906d),
	.w3(32'h3a9bcab6),
	.w4(32'hbb3fd74e),
	.w5(32'hbb5fe93d),
	.w6(32'h39975ec2),
	.w7(32'hbb06ca1c),
	.w8(32'hbb9006c8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e1638),
	.w1(32'hbb478180),
	.w2(32'h39c69ab9),
	.w3(32'h3ae73041),
	.w4(32'h3a725fef),
	.w5(32'hb8e69e19),
	.w6(32'hbbc899d1),
	.w7(32'h3b00d1e1),
	.w8(32'h3b2f64a7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39802565),
	.w1(32'h3a3adf11),
	.w2(32'h3b1d15b1),
	.w3(32'h3a58d940),
	.w4(32'h3a83dcf7),
	.w5(32'h3b10f5f8),
	.w6(32'hbb03a97f),
	.w7(32'hbb08b728),
	.w8(32'hba911da0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b067886),
	.w1(32'hbaa5819a),
	.w2(32'hbb3d754e),
	.w3(32'hbb302f56),
	.w4(32'hbadcffc4),
	.w5(32'hbba300bc),
	.w6(32'hbb028141),
	.w7(32'h3b2696a9),
	.w8(32'hbbb58fc6),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4aa6f),
	.w1(32'hbb320c04),
	.w2(32'hbb26a136),
	.w3(32'hbb93d2ad),
	.w4(32'h3a565e4f),
	.w5(32'hbb2d1445),
	.w6(32'hbbb0540b),
	.w7(32'h3a616bb5),
	.w8(32'h3a9055b3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d22d),
	.w1(32'hbb998eea),
	.w2(32'h3bb4f435),
	.w3(32'h3c33e6dc),
	.w4(32'hbb86b046),
	.w5(32'h3b186d93),
	.w6(32'h3bc362b6),
	.w7(32'h398a4d0a),
	.w8(32'h3b7751a3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be976ad),
	.w1(32'hbbb5567f),
	.w2(32'hba1bf29f),
	.w3(32'h3bec1b0d),
	.w4(32'h3bb35b7c),
	.w5(32'h3b548cfe),
	.w6(32'h3b35fcc1),
	.w7(32'hbb674d7f),
	.w8(32'hbc027dd4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcbe62),
	.w1(32'hbb9942f3),
	.w2(32'hbb3f6336),
	.w3(32'h3b94bfa3),
	.w4(32'hbbb018e4),
	.w5(32'hbb937a35),
	.w6(32'hbb368017),
	.w7(32'hbb8500b6),
	.w8(32'hbb0a018e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb55635),
	.w1(32'hb9821ec0),
	.w2(32'hbb3e7bab),
	.w3(32'hbae52b11),
	.w4(32'hbbc47269),
	.w5(32'hbc6c355d),
	.w6(32'hbbf6deb9),
	.w7(32'h39ea0d7d),
	.w8(32'hbbc2cefb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5deb1),
	.w1(32'hbb42e02b),
	.w2(32'h397f68c4),
	.w3(32'hbb9e60d6),
	.w4(32'hbafe9a85),
	.w5(32'hbb29a0f2),
	.w6(32'hbba57e32),
	.w7(32'hbb4d8a8d),
	.w8(32'hbb7484d8),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule