module layer_10_featuremap_132(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d42b8),
	.w1(32'h3bbd10f7),
	.w2(32'h3af6e86d),
	.w3(32'hbadeebfc),
	.w4(32'h3c174b8b),
	.w5(32'h3c420f8a),
	.w6(32'h3b232c6c),
	.w7(32'h39a15ca8),
	.w8(32'hbb2d445f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc22bdd),
	.w1(32'h3c16b7e9),
	.w2(32'h3c961e3e),
	.w3(32'h3b9ec2e5),
	.w4(32'h3b253faa),
	.w5(32'h3c1ca098),
	.w6(32'h3899fb66),
	.w7(32'h3bd3bb0c),
	.w8(32'h3a8da4b1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2be0ec),
	.w1(32'h3a7ec686),
	.w2(32'h3c1feb21),
	.w3(32'h3b17075b),
	.w4(32'hbb98e0bd),
	.w5(32'h3aaf3716),
	.w6(32'hbb9fc869),
	.w7(32'h3aabdf40),
	.w8(32'hbb088316),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71f2d5),
	.w1(32'hbbb23a03),
	.w2(32'hbb8d091d),
	.w3(32'hbb527ad6),
	.w4(32'hbc07b1ee),
	.w5(32'hbc151012),
	.w6(32'h39be43c5),
	.w7(32'h3b2fd9a4),
	.w8(32'h3b12e1ec),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4d2c),
	.w1(32'hbb87ca56),
	.w2(32'hbafe816c),
	.w3(32'hbbc66843),
	.w4(32'hbb0ae95c),
	.w5(32'hbb358fc1),
	.w6(32'hbb0c68ae),
	.w7(32'hb9b15632),
	.w8(32'h3bdba8dc),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f43e3),
	.w1(32'hbc146aab),
	.w2(32'hbbff6fce),
	.w3(32'h3b89aa10),
	.w4(32'hbc04db6e),
	.w5(32'hbbe3c394),
	.w6(32'hbbd7ab7c),
	.w7(32'hbbdc3e88),
	.w8(32'hbb80ae4c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e42d),
	.w1(32'h3babc22c),
	.w2(32'h3c6dceae),
	.w3(32'hbb26d5a5),
	.w4(32'hbad1ae19),
	.w5(32'h3b97098b),
	.w6(32'hbb5095b1),
	.w7(32'h3b5f9125),
	.w8(32'hbacfff39),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20d224),
	.w1(32'hbc02575f),
	.w2(32'hbc13cd3b),
	.w3(32'hba243839),
	.w4(32'hbba509c2),
	.w5(32'hbbe4fd1c),
	.w6(32'hbba8fe57),
	.w7(32'hbbda0e30),
	.w8(32'hbb8406d4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce3200),
	.w1(32'h3a4f5343),
	.w2(32'h3ae44cb9),
	.w3(32'hbb4aa7e0),
	.w4(32'h3a792da7),
	.w5(32'h3b06370f),
	.w6(32'h3a66c12d),
	.w7(32'h3a88a706),
	.w8(32'h3aaf38f9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea437a),
	.w1(32'h3baea666),
	.w2(32'h3c686db9),
	.w3(32'h3b29e04e),
	.w4(32'h391b568a),
	.w5(32'h3be5872f),
	.w6(32'hbacec27d),
	.w7(32'h3b7aeb85),
	.w8(32'h39da526a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b6bd7),
	.w1(32'hbb4788d2),
	.w2(32'hbb355626),
	.w3(32'h3ad75943),
	.w4(32'hbb647eff),
	.w5(32'hbb779132),
	.w6(32'hbb2f2d8f),
	.w7(32'hbb09431d),
	.w8(32'hbaf4c81f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95ff3a),
	.w1(32'hbaea8e5a),
	.w2(32'hbb245e8d),
	.w3(32'hba0fe00d),
	.w4(32'hbadaab9f),
	.w5(32'hbb5392c0),
	.w6(32'hba29a6d8),
	.w7(32'h39090793),
	.w8(32'h39e87cf8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a7948),
	.w1(32'h390fd047),
	.w2(32'hb927352c),
	.w3(32'hbab7f46c),
	.w4(32'h3a9047a8),
	.w5(32'h3ab7169d),
	.w6(32'h3a6cc828),
	.w7(32'h3a7f8fe2),
	.w8(32'h3a79333c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac59bf4),
	.w1(32'hbcb4f129),
	.w2(32'hbcf38837),
	.w3(32'h3b28adf8),
	.w4(32'hbc81e182),
	.w5(32'hbcab7956),
	.w6(32'hbc75fdc4),
	.w7(32'hbca33ddd),
	.w8(32'hbc86f50a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb9bb4),
	.w1(32'h3a2f0f6e),
	.w2(32'h3b3258f7),
	.w3(32'hbc821540),
	.w4(32'hbad067cf),
	.w5(32'hbb98ed02),
	.w6(32'h3b128ef4),
	.w7(32'h3bb747ca),
	.w8(32'h3b9db042),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a3f8c),
	.w1(32'h3a2a0d33),
	.w2(32'h3b96119b),
	.w3(32'hbb5b022b),
	.w4(32'hb7e9ee8e),
	.w5(32'h3b67cb2b),
	.w6(32'h39d319c4),
	.w7(32'h3b13de24),
	.w8(32'h3b117788),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fa9ad),
	.w1(32'hbba45419),
	.w2(32'hbbcd0c57),
	.w3(32'h3b82fd7a),
	.w4(32'hbb85452b),
	.w5(32'hbb6ec7af),
	.w6(32'hbb874b49),
	.w7(32'hbba745c1),
	.w8(32'hbb033815),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3edf92),
	.w1(32'h3c492cda),
	.w2(32'h3cd1a98e),
	.w3(32'hbaecf1f6),
	.w4(32'h3b7084e9),
	.w5(32'h3c5938cb),
	.w6(32'h3b2a7af4),
	.w7(32'h3c2f2754),
	.w8(32'h3b8df96f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c2840),
	.w1(32'hb8885ed3),
	.w2(32'h3bf490a4),
	.w3(32'h3bc164b3),
	.w4(32'hbb426582),
	.w5(32'h3b5d9377),
	.w6(32'hbb7cc99a),
	.w7(32'hb88ec80a),
	.w8(32'hbb98df6d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11d88d),
	.w1(32'h3a8a6f5b),
	.w2(32'h3a91f3dc),
	.w3(32'hbad9b095),
	.w4(32'h3aa4c661),
	.w5(32'h3ac9b05c),
	.w6(32'h3a1a12e9),
	.w7(32'h3a05403d),
	.w8(32'h39e7a424),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5da09c),
	.w1(32'hba843a09),
	.w2(32'hbb211609),
	.w3(32'h3ac031ec),
	.w4(32'h3847ba4b),
	.w5(32'hba8c2a26),
	.w6(32'h3905e0e7),
	.w7(32'hba52e818),
	.w8(32'h390e3e8e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4009d),
	.w1(32'h3b039baf),
	.w2(32'h3b9e92bb),
	.w3(32'h392fd4de),
	.w4(32'h3bbf2a53),
	.w5(32'h3c263999),
	.w6(32'hbab7a4f0),
	.w7(32'h3b230e8c),
	.w8(32'h3b26fb80),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c2620),
	.w1(32'h398835af),
	.w2(32'h396057e4),
	.w3(32'h3bfca6e0),
	.w4(32'h3a46d8a5),
	.w5(32'h3b226593),
	.w6(32'hb9347a2f),
	.w7(32'hb9e1acf4),
	.w8(32'hbb01a888),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e079cc),
	.w1(32'hbbc971d8),
	.w2(32'hbbee00f5),
	.w3(32'h3a6eabe8),
	.w4(32'hbb8cde7f),
	.w5(32'hbbafc3b8),
	.w6(32'hbb896023),
	.w7(32'hbbac50a8),
	.w8(32'hbb8b9952),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4d43c),
	.w1(32'hbabc9574),
	.w2(32'h3b156929),
	.w3(32'hbb6c4085),
	.w4(32'hbb89d08d),
	.w5(32'hbb4a0ef9),
	.w6(32'hbb870312),
	.w7(32'hbac5a053),
	.w8(32'hbb84e3fc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80176e),
	.w1(32'h3ad7693c),
	.w2(32'h3ace6219),
	.w3(32'hbbd91c61),
	.w4(32'h3b1d3d52),
	.w5(32'h3b5b9496),
	.w6(32'h3ac13bf6),
	.w7(32'hbab1f434),
	.w8(32'h39cc8945),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b1543),
	.w1(32'h38f9326b),
	.w2(32'h36ffafbd),
	.w3(32'h3b344b5a),
	.w4(32'h39988178),
	.w5(32'h39b282a1),
	.w6(32'hb832b537),
	.w7(32'h37da0bb8),
	.w8(32'h38d3d6e7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efe33f),
	.w1(32'hbb8f0027),
	.w2(32'h3b11cdb0),
	.w3(32'h3a06dd31),
	.w4(32'hbba9cb6a),
	.w5(32'hbb142ce3),
	.w6(32'hbbf8f3d0),
	.w7(32'hbb91c869),
	.w8(32'hbbbb6b83),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833ae3),
	.w1(32'hbbbb323a),
	.w2(32'hbb8df8ad),
	.w3(32'hbbbff9ba),
	.w4(32'hbb858be9),
	.w5(32'hbb3111d5),
	.w6(32'hbbe4f3e0),
	.w7(32'hbbe03dd9),
	.w8(32'hbb752451),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29a41),
	.w1(32'hbb4831d4),
	.w2(32'hbb5509fa),
	.w3(32'h3a6158c5),
	.w4(32'hbb3baef0),
	.w5(32'hbb643da3),
	.w6(32'hbb0fdbcd),
	.w7(32'hbb108b09),
	.w8(32'hbb179608),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eaa51),
	.w1(32'hba8c1466),
	.w2(32'hbae779fc),
	.w3(32'hbb7b6c90),
	.w4(32'hb975c78e),
	.w5(32'hba501cea),
	.w6(32'hb9cd4b71),
	.w7(32'hba7b66ea),
	.w8(32'hb9d67061),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba719d4d),
	.w1(32'h3a12786f),
	.w2(32'h3a09bdf8),
	.w3(32'hb899e227),
	.w4(32'h3ab9a977),
	.w5(32'h3ae2a928),
	.w6(32'h3a23a54f),
	.w7(32'h3a797668),
	.w8(32'h3aa119c2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf7bca),
	.w1(32'hbb26288a),
	.w2(32'hba6e2488),
	.w3(32'h3b1ffd79),
	.w4(32'hba24281d),
	.w5(32'h3890e58e),
	.w6(32'hbb8837fe),
	.w7(32'hbb6ff41a),
	.w8(32'h3b823e4b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf5bce),
	.w1(32'h3b176d6b),
	.w2(32'hbb16917a),
	.w3(32'h3bab2966),
	.w4(32'h3af48ac5),
	.w5(32'h3ab98830),
	.w6(32'h3b2d7da7),
	.w7(32'hbb0e5171),
	.w8(32'hbbb3f9c6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6bb15),
	.w1(32'h3c12a94a),
	.w2(32'h3c99b106),
	.w3(32'h398046bb),
	.w4(32'h3b02735f),
	.w5(32'h3c1cf90b),
	.w6(32'hb998facf),
	.w7(32'h3ba432d2),
	.w8(32'hba7b662b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20e6ab),
	.w1(32'hba52cf9a),
	.w2(32'hba7a593f),
	.w3(32'h3b2186ec),
	.w4(32'h386de98a),
	.w5(32'hb91b9691),
	.w6(32'hba51a2f2),
	.w7(32'hb97b2e4e),
	.w8(32'hb9984330),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27651f),
	.w1(32'h3c11ae5d),
	.w2(32'h3c885b92),
	.w3(32'h3a6d1654),
	.w4(32'h3b0ca6a4),
	.w5(32'h3be3c39f),
	.w6(32'h3a48da10),
	.w7(32'h3b87aeba),
	.w8(32'hb9f88aa9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38fe31),
	.w1(32'h3c07cb91),
	.w2(32'h3c8277b1),
	.w3(32'h3b1b713e),
	.w4(32'h3b118f37),
	.w5(32'h3c04a814),
	.w6(32'h3a8497fd),
	.w7(32'h3bd00edd),
	.w8(32'h3aa085d5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17369c),
	.w1(32'hbb75328d),
	.w2(32'hbb5569f4),
	.w3(32'h3b37f730),
	.w4(32'hbaef4ee6),
	.w5(32'hbae8b8d2),
	.w6(32'hbaea8c3c),
	.w7(32'hbaef9d44),
	.w8(32'hbab37e47),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dec2b),
	.w1(32'h3a86e1c8),
	.w2(32'h3bf58894),
	.w3(32'hba8474b8),
	.w4(32'hbae962e1),
	.w5(32'h3b2c4258),
	.w6(32'hbba4451a),
	.w7(32'hba1fc382),
	.w8(32'hbb977b2e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cbca3),
	.w1(32'hba2447b6),
	.w2(32'hb9d27175),
	.w3(32'hbb10dba8),
	.w4(32'hb9a705f4),
	.w5(32'hb9d72040),
	.w6(32'hba764b89),
	.w7(32'hba268e22),
	.w8(32'hbb0b5833),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51c7d6),
	.w1(32'h3abf53c8),
	.w2(32'h3c295e74),
	.w3(32'hbb190df6),
	.w4(32'hbb8f5fbb),
	.w5(32'h3ac60858),
	.w6(32'hbb8cee69),
	.w7(32'h3aa4ee6f),
	.w8(32'hbb48b47c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8e33b),
	.w1(32'h3a85a330),
	.w2(32'h3a6efe3d),
	.w3(32'hba2a8d17),
	.w4(32'h3aeca101),
	.w5(32'h3b16774b),
	.w6(32'h3ab5f84f),
	.w7(32'h3ac11709),
	.w8(32'h3b00b90e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec1824),
	.w1(32'h3bf21a0c),
	.w2(32'h3c7ea3ad),
	.w3(32'h3b37d433),
	.w4(32'h3b0ecf9a),
	.w5(32'h3c0877c7),
	.w6(32'h3b058b2e),
	.w7(32'h3bbc4ac7),
	.w8(32'h3b53583a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3571a5),
	.w1(32'hbab11d47),
	.w2(32'h3afe57ec),
	.w3(32'h3b795e3a),
	.w4(32'hbb823bd9),
	.w5(32'hba5b7334),
	.w6(32'hbaec8eee),
	.w7(32'h3b0a31c5),
	.w8(32'h3a6ae5ec),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72be90),
	.w1(32'hbb691177),
	.w2(32'h39e35b33),
	.w3(32'hbb0b616e),
	.w4(32'hbb89d870),
	.w5(32'hbaa3d4a7),
	.w6(32'hbbfb0db8),
	.w7(32'hbb8d9ec8),
	.w8(32'hbbe0dcce),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fefb4),
	.w1(32'hb8a6f113),
	.w2(32'h3ba1c595),
	.w3(32'hbbada37f),
	.w4(32'hbb06b175),
	.w5(32'hb8b54fbc),
	.w6(32'h3b73aee2),
	.w7(32'h3c2b973c),
	.w8(32'h3c28a55b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc734f9),
	.w1(32'hbb0c9e3d),
	.w2(32'hbb3ee854),
	.w3(32'h3ac1ae3e),
	.w4(32'hba4b46ee),
	.w5(32'hba486f38),
	.w6(32'hbab185a1),
	.w7(32'hbb64cac4),
	.w8(32'hbb472fbd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe111c),
	.w1(32'h3949c0c4),
	.w2(32'h3946c4a8),
	.w3(32'h3a79b69d),
	.w4(32'h3a99acd5),
	.w5(32'h3ad2be22),
	.w6(32'h3931cffb),
	.w7(32'h3a279d6f),
	.w8(32'h39f11685),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987152a),
	.w1(32'hbbaba6a0),
	.w2(32'hbbecd6a1),
	.w3(32'h3aa01a48),
	.w4(32'hbb1c0051),
	.w5(32'hbb7cf2d4),
	.w6(32'hbb31020a),
	.w7(32'hbb73901b),
	.w8(32'hbb15f900),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4e6c8),
	.w1(32'hbb701bc5),
	.w2(32'hb96fcd7b),
	.w3(32'hbb1991d5),
	.w4(32'hbbde1e01),
	.w5(32'hbb5cddbd),
	.w6(32'hbc05ef82),
	.w7(32'hbbbb3999),
	.w8(32'hbc1ca13b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f9dba),
	.w1(32'h3bf8a905),
	.w2(32'h3bc55b62),
	.w3(32'hbbfc9944),
	.w4(32'h3a587b80),
	.w5(32'hbb48cf63),
	.w6(32'h394e080d),
	.w7(32'h3b03f5b7),
	.w8(32'hbb13abed),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1c875),
	.w1(32'hb9d533b3),
	.w2(32'h3b602bbc),
	.w3(32'hbb9bcf81),
	.w4(32'hbaf8ea59),
	.w5(32'h3a9b7100),
	.w6(32'hba125211),
	.w7(32'h3a95e8b9),
	.w8(32'h3aa183de),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7377ac),
	.w1(32'hbc175296),
	.w2(32'hbbc9de0e),
	.w3(32'h3afabd53),
	.w4(32'hbc18147b),
	.w5(32'hbc018f5f),
	.w6(32'hbbd8a4cd),
	.w7(32'hbbace3d0),
	.w8(32'hbb27097a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d9cac),
	.w1(32'hbb7ac021),
	.w2(32'hbb0c4c9d),
	.w3(32'hbbaa2954),
	.w4(32'hbba98e9f),
	.w5(32'hbb29e34c),
	.w6(32'hbbabf639),
	.w7(32'hbb892136),
	.w8(32'hbb58b74a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee3d9c),
	.w1(32'h3a6b55bc),
	.w2(32'h3b1f9d0b),
	.w3(32'hbb1f5d41),
	.w4(32'h3ace5836),
	.w5(32'h3ac53b6b),
	.w6(32'hb9c9887b),
	.w7(32'h3a669899),
	.w8(32'hb99b177f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2ae18),
	.w1(32'hbbd96142),
	.w2(32'hbb571118),
	.w3(32'h3a041a1c),
	.w4(32'hbc2e418f),
	.w5(32'hbbcf4314),
	.w6(32'hbc291ee2),
	.w7(32'hbc016bf5),
	.w8(32'hbc4967bd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc011b2a),
	.w1(32'h3a8545cd),
	.w2(32'hbae4591e),
	.w3(32'hbc1888ef),
	.w4(32'h3b7e151e),
	.w5(32'h3aa78500),
	.w6(32'hba78787f),
	.w7(32'hbac74a8f),
	.w8(32'h39888d89),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a771c),
	.w1(32'h3b0c02b9),
	.w2(32'h3c1c9866),
	.w3(32'h3a8df50c),
	.w4(32'hbbe149c4),
	.w5(32'hba861b66),
	.w6(32'hbbcbcf0c),
	.w7(32'hbaf94ce6),
	.w8(32'hbc0d4fd3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23b1c2),
	.w1(32'hbb997eca),
	.w2(32'hbba012a9),
	.w3(32'hbc0ca6e5),
	.w4(32'hbb48847c),
	.w5(32'hbb5e15c1),
	.w6(32'hbb59711e),
	.w7(32'hbb76f755),
	.w8(32'hbb5b0e34),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c34f),
	.w1(32'hbb1281ae),
	.w2(32'h3c400aae),
	.w3(32'hbb24e29a),
	.w4(32'hbbcf4b5b),
	.w5(32'h3b52458c),
	.w6(32'hbc146afd),
	.w7(32'h3a8887e1),
	.w8(32'hbb67895a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba03e99),
	.w1(32'hbb9b747e),
	.w2(32'hbbc6e8ee),
	.w3(32'hbb28f21c),
	.w4(32'hbb1da1c2),
	.w5(32'hbb339967),
	.w6(32'hbb5c2034),
	.w7(32'hbb9b5017),
	.w8(32'hbb666ab2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922e2f),
	.w1(32'hbb17d84b),
	.w2(32'hba68b840),
	.w3(32'hbacee7d6),
	.w4(32'hbae1084a),
	.w5(32'hba3edfcd),
	.w6(32'hbb642b6a),
	.w7(32'h3941e4b7),
	.w8(32'h3bcba76b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5035c),
	.w1(32'h3bc9e987),
	.w2(32'h3c410a50),
	.w3(32'h3baa6a4a),
	.w4(32'h3af4484d),
	.w5(32'h3bc0ee79),
	.w6(32'h3a94ecc5),
	.w7(32'h3b9cbf9e),
	.w8(32'h3b1829c6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf84fd5),
	.w1(32'hbb55cc56),
	.w2(32'h3ba121d7),
	.w3(32'h3ae43596),
	.w4(32'hbbcb6ba2),
	.w5(32'hb98943b7),
	.w6(32'hbbb88fc9),
	.w7(32'h3a98fc35),
	.w8(32'h3a0b9d24),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99db9e),
	.w1(32'h3bb6b5f7),
	.w2(32'h3a1e55ed),
	.w3(32'hbad9dd51),
	.w4(32'h3c00aa8b),
	.w5(32'h3ba5c7a7),
	.w6(32'h3ba657fc),
	.w7(32'h3ab31b53),
	.w8(32'h3b5d9415),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5332bd),
	.w1(32'h385ab5e0),
	.w2(32'h3aa98ab3),
	.w3(32'h3b9fac56),
	.w4(32'hba0e9ea5),
	.w5(32'h39df897b),
	.w6(32'h3b14ffa1),
	.w7(32'h3aadf14b),
	.w8(32'hb91dcbe2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c6858),
	.w1(32'hba556047),
	.w2(32'hb89331d1),
	.w3(32'h39a49024),
	.w4(32'hbaa7fda3),
	.w5(32'hb9737a28),
	.w6(32'hba4c9dde),
	.w7(32'hba70a658),
	.w8(32'hba43b6f9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4197a),
	.w1(32'hb8264e3a),
	.w2(32'h3b2cb2c2),
	.w3(32'h389ce1e3),
	.w4(32'hb9c04cc5),
	.w5(32'h3adf924b),
	.w6(32'hb98c9c0d),
	.w7(32'h3a8617a0),
	.w8(32'h3acc94de),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b557c15),
	.w1(32'hbbda4218),
	.w2(32'hbbf28011),
	.w3(32'h3b506697),
	.w4(32'hbb7585ac),
	.w5(32'hbbb8084e),
	.w6(32'hbbfb766a),
	.w7(32'hbbef78d5),
	.w8(32'hbc126909),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc149ab1),
	.w1(32'h3c26c55a),
	.w2(32'h3c99d935),
	.w3(32'hbc2377eb),
	.w4(32'h3b1ce2e8),
	.w5(32'h3c0366e9),
	.w6(32'h3b2978ae),
	.w7(32'h3bffea36),
	.w8(32'h3aa3daf2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1197a5),
	.w1(32'hbb4173c1),
	.w2(32'hbb5d5d76),
	.w3(32'h3a6e2f22),
	.w4(32'hbae358ef),
	.w5(32'hbb26ffe5),
	.w6(32'hbb191acc),
	.w7(32'hbb23a427),
	.w8(32'hbac94cfd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040899),
	.w1(32'hbb55ad9f),
	.w2(32'hbb38f28d),
	.w3(32'hba88abf1),
	.w4(32'hbb0b3de9),
	.w5(32'hbb0aff6e),
	.w6(32'hbb1190ef),
	.w7(32'hbb13820c),
	.w8(32'hbaee4436),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300572),
	.w1(32'hb92a53f2),
	.w2(32'h3912817d),
	.w3(32'hbaaabe50),
	.w4(32'h3a8ad2ae),
	.w5(32'h3abdd1ac),
	.w6(32'h39909140),
	.w7(32'h3a63bafa),
	.w8(32'h3a851b6a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bbd25),
	.w1(32'h3a538d6e),
	.w2(32'h3c22e1e1),
	.w3(32'h3aedc3ec),
	.w4(32'hbbdb396e),
	.w5(32'h390e041e),
	.w6(32'hbbce4ced),
	.w7(32'h3a8be73b),
	.w8(32'hbb3fd816),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82db7b),
	.w1(32'h3b89ecf5),
	.w2(32'h3c0b6d75),
	.w3(32'hbb939917),
	.w4(32'h3b84260e),
	.w5(32'h3c1a5cb6),
	.w6(32'h3a4023de),
	.w7(32'h3b036963),
	.w8(32'h3b29a530),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dd0c0),
	.w1(32'hbc17966b),
	.w2(32'hbc79b93c),
	.w3(32'h3c42e003),
	.w4(32'hbb3c4d78),
	.w5(32'hbbe7998e),
	.w6(32'hbb195bf9),
	.w7(32'hbbee0f42),
	.w8(32'hbb2290d2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07140f),
	.w1(32'hbb50d446),
	.w2(32'h3beaebfb),
	.w3(32'hba68423d),
	.w4(32'hbc129c90),
	.w5(32'h39437710),
	.w6(32'hbc053a07),
	.w7(32'hbac21fbb),
	.w8(32'hbbc4a5ce),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f46df),
	.w1(32'hbad4d74d),
	.w2(32'hba1945fc),
	.w3(32'hbb6bd6f1),
	.w4(32'h388ed438),
	.w5(32'h3b4e4028),
	.w6(32'hba723f2b),
	.w7(32'hbaa334d6),
	.w8(32'h3b85d43a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b860b1c),
	.w1(32'hbab1db39),
	.w2(32'hbb35fa64),
	.w3(32'h3b91dcfe),
	.w4(32'hba0fe078),
	.w5(32'hbab56843),
	.w6(32'h38a8c46c),
	.w7(32'hbab15ad1),
	.w8(32'hb9e1b3d3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8433b6),
	.w1(32'h3a532889),
	.w2(32'h3b145cc4),
	.w3(32'h38d64064),
	.w4(32'h390c8b62),
	.w5(32'h3af5a718),
	.w6(32'h3a012520),
	.w7(32'h3ad76f30),
	.w8(32'h394a8b91),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61fecd),
	.w1(32'hbb05150f),
	.w2(32'h3bc9890b),
	.w3(32'h3acbd89d),
	.w4(32'hbc146a96),
	.w5(32'hbada1b2c),
	.w6(32'hbc06448c),
	.w7(32'hbb5a6395),
	.w8(32'hbc17f36e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06a762),
	.w1(32'h3b393442),
	.w2(32'h3b8db281),
	.w3(32'hbbe01101),
	.w4(32'h3a2efaa9),
	.w5(32'h3a465379),
	.w6(32'h3ae540c3),
	.w7(32'h3b12cf93),
	.w8(32'hba67ea08),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71602d),
	.w1(32'hba715754),
	.w2(32'h3bb3927b),
	.w3(32'hbb0fe12c),
	.w4(32'hbbcf76c3),
	.w5(32'hb95c08b2),
	.w6(32'hbbf2e550),
	.w7(32'hbb1d7b63),
	.w8(32'hbbd97952),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b82f3b),
	.w1(32'hb946ef83),
	.w2(32'hbb23c9ea),
	.w3(32'hbbab387d),
	.w4(32'hba563e27),
	.w5(32'hbabc9756),
	.w6(32'h3b7e1652),
	.w7(32'h3add400d),
	.w8(32'h3af46140),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba641f77),
	.w1(32'hbb1a148f),
	.w2(32'h37e74fa8),
	.w3(32'h3a5ff744),
	.w4(32'hbbaa5241),
	.w5(32'hbb3824a0),
	.w6(32'hbb7945a5),
	.w7(32'hbb3e9b0b),
	.w8(32'hbbc4ab5b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500402),
	.w1(32'hbb254ce0),
	.w2(32'hbb36fb44),
	.w3(32'hbbb24fe0),
	.w4(32'hbb326954),
	.w5(32'hbaa99c42),
	.w6(32'hbbc6ded8),
	.w7(32'hbc010064),
	.w8(32'hbc4dab4b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c92cb),
	.w1(32'hba1443e1),
	.w2(32'hbaabb5ce),
	.w3(32'hbb9cb5f3),
	.w4(32'h38eff3ec),
	.w5(32'hb9f56d7c),
	.w6(32'h38e643d8),
	.w7(32'hb9deb908),
	.w8(32'h37ee27ac),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3da630),
	.w1(32'hbb9affd2),
	.w2(32'hbb705f4e),
	.w3(32'h391ae5e0),
	.w4(32'hbbe295d1),
	.w5(32'hbbba9abc),
	.w6(32'hbbd565eb),
	.w7(32'hbbd7d012),
	.w8(32'hbbe7a6b9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cd696),
	.w1(32'hb88fd4a9),
	.w2(32'hba6aa1c6),
	.w3(32'hbbd38a4b),
	.w4(32'h3a740fe4),
	.w5(32'h398d49f9),
	.w6(32'h3a87251f),
	.w7(32'h388692d2),
	.w8(32'h3a3fda49),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15b8e7),
	.w1(32'hb9dd568f),
	.w2(32'hba81a0b4),
	.w3(32'h3afd9946),
	.w4(32'h3a66ffea),
	.w5(32'h39b7f01a),
	.w6(32'hb94fe46d),
	.w7(32'hb9445dc6),
	.w8(32'hb99515b0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d891e6),
	.w1(32'h3bcc14a6),
	.w2(32'h3c45e8df),
	.w3(32'h3a5f5603),
	.w4(32'hb9ed9d8a),
	.w5(32'h3bc429ca),
	.w6(32'h3b15072d),
	.w7(32'h3bdd36be),
	.w8(32'h3b6d3269),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c343891),
	.w1(32'h3b639c13),
	.w2(32'h3bf64355),
	.w3(32'h3b704abd),
	.w4(32'h37f4b912),
	.w5(32'h3b8f6842),
	.w6(32'h39d3d489),
	.w7(32'h3b6173b3),
	.w8(32'h3b1263a6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5e95d),
	.w1(32'hba34b329),
	.w2(32'h3a9fb8b7),
	.w3(32'h3b503eef),
	.w4(32'hba0ca33d),
	.w5(32'h3ac88d74),
	.w6(32'hbaf62131),
	.w7(32'hb9bfbaaf),
	.w8(32'hba084a5c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec5c28),
	.w1(32'h3b783006),
	.w2(32'h3c30e090),
	.w3(32'h3a8f4d45),
	.w4(32'hb98063d5),
	.w5(32'h3ba0a00b),
	.w6(32'hbb4e1eb3),
	.w7(32'h3a91bf38),
	.w8(32'hbb24f127),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b744),
	.w1(32'hbbb28576),
	.w2(32'hbb65c127),
	.w3(32'h3a96c80e),
	.w4(32'h3a22e057),
	.w5(32'h3ba8469e),
	.w6(32'hbbbbd109),
	.w7(32'hbbc3923a),
	.w8(32'hbb684649),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e4558),
	.w1(32'h3b44827d),
	.w2(32'h3bda5623),
	.w3(32'h3bbcb886),
	.w4(32'h3b13f441),
	.w5(32'h3bbf839f),
	.w6(32'h3a447235),
	.w7(32'h3b4b27d1),
	.w8(32'h3aee2cfb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ea757),
	.w1(32'h3a8ef53b),
	.w2(32'hbb5609de),
	.w3(32'h3b856f72),
	.w4(32'h3a890b0b),
	.w5(32'hbb5205ae),
	.w6(32'h3b030376),
	.w7(32'hbad63600),
	.w8(32'hbbbb89a1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1269ee),
	.w1(32'h3a8af554),
	.w2(32'h3c5d6ef8),
	.w3(32'hbbebda36),
	.w4(32'hbc0200a4),
	.w5(32'h3b6a68bb),
	.w6(32'hbbb1941f),
	.w7(32'h3b687749),
	.w8(32'hbb708316),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2d150),
	.w1(32'h3a6d3575),
	.w2(32'h3b1c8cde),
	.w3(32'hbaff8926),
	.w4(32'hbb0aa54f),
	.w5(32'hbac6d80c),
	.w6(32'hb909120d),
	.w7(32'hbad9147d),
	.w8(32'hbb5169b4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4812bf),
	.w1(32'h3c063698),
	.w2(32'h3c4a9aa1),
	.w3(32'hbaef3e56),
	.w4(32'h3c135de2),
	.w5(32'h3c490158),
	.w6(32'h3b1fef0a),
	.w7(32'h3c0d4089),
	.w8(32'h3bdbcd61),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6803eb),
	.w1(32'hbbbd17be),
	.w2(32'hbbcbca2b),
	.w3(32'h3c1fa0eb),
	.w4(32'h3b0e8b90),
	.w5(32'h3b712329),
	.w6(32'hbadc1337),
	.w7(32'hbb0d9261),
	.w8(32'h3ba7b01b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8b3e7),
	.w1(32'hbc59fbfe),
	.w2(32'hbcbcebe2),
	.w3(32'h3c188c3b),
	.w4(32'hbb744c64),
	.w5(32'hbc2b7705),
	.w6(32'hbb559bfc),
	.w7(32'hbc31156c),
	.w8(32'hbb780cf2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d2f58),
	.w1(32'hbab1c93f),
	.w2(32'hbaf0e195),
	.w3(32'hbadf6da9),
	.w4(32'hba114c8d),
	.w5(32'hbaba0645),
	.w6(32'hba993e31),
	.w7(32'hbacd5d89),
	.w8(32'hb9ac5d61),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89508d1),
	.w1(32'hbbd3e9f7),
	.w2(32'hbc3688e2),
	.w3(32'hba0bef85),
	.w4(32'hbad95fca),
	.w5(32'hbbaf771c),
	.w6(32'hba8baa55),
	.w7(32'hbb9b9328),
	.w8(32'hbb139c5f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb94e7d),
	.w1(32'h3a5680c2),
	.w2(32'hb948a000),
	.w3(32'hb968b872),
	.w4(32'h3aae25bf),
	.w5(32'h398726bd),
	.w6(32'h3a210927),
	.w7(32'hb8d802ab),
	.w8(32'hb8fff7df),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e4555),
	.w1(32'h3a8de605),
	.w2(32'h3c16d71d),
	.w3(32'h3a47efae),
	.w4(32'hbbd1ec30),
	.w5(32'hb9899826),
	.w6(32'hbb8c3061),
	.w7(32'h3b2c168c),
	.w8(32'hba6f1e69),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2b87f),
	.w1(32'hbabf2ab6),
	.w2(32'hbb2699fa),
	.w3(32'hbb17ab7c),
	.w4(32'hb994ef3c),
	.w5(32'hba93d5fb),
	.w6(32'hba1231af),
	.w7(32'hbaadb5e3),
	.w8(32'hba7e6e9c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1397c6),
	.w1(32'hbc077661),
	.w2(32'hbc518ca5),
	.w3(32'hba233945),
	.w4(32'hbb46929f),
	.w5(32'hbbc0427c),
	.w6(32'hbb36012b),
	.w7(32'hbbd4d8f0),
	.w8(32'hbb195062),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56052),
	.w1(32'hbbd37c18),
	.w2(32'h39b2af80),
	.w3(32'hbabce93c),
	.w4(32'hbc31d8f4),
	.w5(32'hbba643a0),
	.w6(32'hbc32698d),
	.w7(32'hbbb8984b),
	.w8(32'hbbf11757),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac61f05),
	.w1(32'h3abf6bc0),
	.w2(32'h3b747f12),
	.w3(32'hbc05a3ed),
	.w4(32'h3aa15d13),
	.w5(32'h3b273b79),
	.w6(32'h3a3a542d),
	.w7(32'h3b4d5e25),
	.w8(32'h3b45fe3a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40dc33),
	.w1(32'h3923bb7d),
	.w2(32'hbae322fa),
	.w3(32'h3b662c3e),
	.w4(32'hb8b6ab1d),
	.w5(32'hbb00d9fe),
	.w6(32'h3a87893f),
	.w7(32'h3a06b634),
	.w8(32'h3b0de4f4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93f1e4),
	.w1(32'hbab72018),
	.w2(32'h3b0a07a8),
	.w3(32'h3ae5f03a),
	.w4(32'hbb0c6b04),
	.w5(32'hba4af2f8),
	.w6(32'hbafdd838),
	.w7(32'h39cfda32),
	.w8(32'h3a3cf67e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea9f64),
	.w1(32'h3b24a0ae),
	.w2(32'h3c0622ae),
	.w3(32'h38fc87cc),
	.w4(32'hbbcd3317),
	.w5(32'hbb523538),
	.w6(32'hbb7ea974),
	.w7(32'hb9aac8ef),
	.w8(32'hbc025a2a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3114),
	.w1(32'hbb453693),
	.w2(32'hbb79811b),
	.w3(32'hbc1bfc5b),
	.w4(32'hbb00f518),
	.w5(32'hbade1dea),
	.w6(32'hbaf7a150),
	.w7(32'hbb31bbd9),
	.w8(32'hbadff9c7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa6b7c),
	.w1(32'hbc25d7ac),
	.w2(32'hbc896f56),
	.w3(32'hb9887315),
	.w4(32'hbb3b04f9),
	.w5(32'hbbf4dac6),
	.w6(32'hbb379ba7),
	.w7(32'hbbffffca),
	.w8(32'hbb0e7799),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1445c9),
	.w1(32'hbbaebe94),
	.w2(32'hbbcba2d5),
	.w3(32'hba5c5f56),
	.w4(32'hbb713f01),
	.w5(32'hbb9b0dae),
	.w6(32'hbb27b651),
	.w7(32'hbb644268),
	.w8(32'hbad0f320),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e46e3),
	.w1(32'hbbdaaf30),
	.w2(32'hbbee8971),
	.w3(32'hbad972a9),
	.w4(32'hbb832221),
	.w5(32'hbb9a8a60),
	.w6(32'hbb5dd952),
	.w7(32'hbb82a237),
	.w8(32'hba54f6f1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407c8a),
	.w1(32'hbb53f529),
	.w2(32'hbb570cd1),
	.w3(32'hba047fa0),
	.w4(32'h3a2b3e6a),
	.w5(32'h3a2444cb),
	.w6(32'hbae84d41),
	.w7(32'hb96f0850),
	.w8(32'h3ac615ec),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee95b4),
	.w1(32'h3be87c8b),
	.w2(32'h3c41676e),
	.w3(32'h3b095b0e),
	.w4(32'h3b88b959),
	.w5(32'h3be8492b),
	.w6(32'h3adf5d46),
	.w7(32'h3b98183a),
	.w8(32'hbb121979),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5335d3),
	.w1(32'hb958b104),
	.w2(32'h3afd757f),
	.w3(32'hbaf6d44e),
	.w4(32'hba133cff),
	.w5(32'h3a02e5e9),
	.w6(32'hb9db0d45),
	.w7(32'h3b06a717),
	.w8(32'h3b157f58),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95619f),
	.w1(32'h398be877),
	.w2(32'h3b3dad2f),
	.w3(32'h3b076c74),
	.w4(32'hba0f4725),
	.w5(32'h3b1dd885),
	.w6(32'hba9c88f0),
	.w7(32'h3a41a023),
	.w8(32'hba97e1c1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23c1f5),
	.w1(32'hbbb9108e),
	.w2(32'hbbd496d6),
	.w3(32'h3ac46c99),
	.w4(32'hbb752bcf),
	.w5(32'hbb946b20),
	.w6(32'hbb8013ec),
	.w7(32'hbb971192),
	.w8(32'hbb776272),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd9c3f),
	.w1(32'hba9292b6),
	.w2(32'hbaf0338e),
	.w3(32'hbb5b036e),
	.w4(32'h3bc5a0e0),
	.w5(32'h3bff8612),
	.w6(32'h3b086fdc),
	.w7(32'h3a7e06c5),
	.w8(32'h3b80b6ec),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953808f),
	.w1(32'hbb80c2d8),
	.w2(32'hba44040e),
	.w3(32'h3bd900e1),
	.w4(32'hbb932b6c),
	.w5(32'hba6a57a4),
	.w6(32'hbb312623),
	.w7(32'hbad749fe),
	.w8(32'hba6421ba),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d1f9e),
	.w1(32'hba92124d),
	.w2(32'hbaf21e8f),
	.w3(32'h3ae0e0fd),
	.w4(32'h37f0756c),
	.w5(32'hba32fc24),
	.w6(32'hba10be83),
	.w7(32'hba82f97d),
	.w8(32'hba2d8405),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5c78c),
	.w1(32'hb80874bc),
	.w2(32'hb8115873),
	.w3(32'hb8ccacf3),
	.w4(32'hb8032106),
	.w5(32'hb7051980),
	.w6(32'hb8798c74),
	.w7(32'hb843edf2),
	.w8(32'hb73d6329),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82daff7),
	.w1(32'hb91cc42a),
	.w2(32'hb98537b9),
	.w3(32'h39812a11),
	.w4(32'h38949570),
	.w5(32'h384722ee),
	.w6(32'h3891b650),
	.w7(32'hba357c6b),
	.w8(32'hba12b8d9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bfebf),
	.w1(32'hba14e942),
	.w2(32'hb9f5efcd),
	.w3(32'hb8fdf948),
	.w4(32'hb9f0a57b),
	.w5(32'hb993d7e9),
	.w6(32'hb879cb51),
	.w7(32'hba0edb58),
	.w8(32'hb9e7b32b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367cdc38),
	.w1(32'hb7e1f505),
	.w2(32'hb894d9bf),
	.w3(32'hb72006c0),
	.w4(32'hb8801c2d),
	.w5(32'hb85946a5),
	.w6(32'h37ab59f2),
	.w7(32'hb81226dd),
	.w8(32'hb8eb0aff),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b656ba),
	.w1(32'hb91b992b),
	.w2(32'hb763010c),
	.w3(32'h37c558fa),
	.w4(32'hb6bad8ed),
	.w5(32'hb8d17c38),
	.w6(32'hb92bd323),
	.w7(32'hb9297682),
	.w8(32'hb81a42b1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c5a175),
	.w1(32'h3825ce9e),
	.w2(32'h385ed629),
	.w3(32'h36e9e5ed),
	.w4(32'h3794bd42),
	.w5(32'h37acb7d1),
	.w6(32'h36873b3c),
	.w7(32'h37dc07bd),
	.w8(32'hb7c784ce),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb713e46e),
	.w1(32'hb8a26991),
	.w2(32'h389b419c),
	.w3(32'hb8852338),
	.w4(32'hb8b73ee9),
	.w5(32'hb6fd757e),
	.w6(32'hb95ba4e7),
	.w7(32'hb90d5fb4),
	.w8(32'hb86408fe),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828c6d7),
	.w1(32'hb8e6aa63),
	.w2(32'h38f4c6f8),
	.w3(32'hb830a521),
	.w4(32'hb98a0412),
	.w5(32'hb72fca93),
	.w6(32'hb97beebe),
	.w7(32'hb9922aa6),
	.w8(32'hb991f81c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8196f20),
	.w1(32'hba084d18),
	.w2(32'hba44ba0b),
	.w3(32'hb8e60d9c),
	.w4(32'hba22b87a),
	.w5(32'hba080615),
	.w6(32'h383f73bf),
	.w7(32'hba389bcd),
	.w8(32'hba3f5c3a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f81fc8),
	.w1(32'h39396464),
	.w2(32'h39160612),
	.w3(32'h38a44a29),
	.w4(32'h392e3787),
	.w5(32'h3894b689),
	.w6(32'h38ee8eab),
	.w7(32'h3942930f),
	.w8(32'h3895fb9e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3896396d),
	.w1(32'hb867c3d9),
	.w2(32'hb8e1d860),
	.w3(32'hb8a9f429),
	.w4(32'hb8fb101d),
	.w5(32'h3682ccaa),
	.w6(32'hb7a1be47),
	.w7(32'hb8da17dc),
	.w8(32'hb96cb2b4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985e1c5),
	.w1(32'hb98977f7),
	.w2(32'hb9e6a48f),
	.w3(32'h3761b906),
	.w4(32'hb98213f7),
	.w5(32'hb9a1bc9e),
	.w6(32'h3848665f),
	.w7(32'hb9a12f88),
	.w8(32'hba084f44),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0bdab),
	.w1(32'h38e3db3b),
	.w2(32'h392b6817),
	.w3(32'h38c8d741),
	.w4(32'h39580674),
	.w5(32'h39287494),
	.w6(32'h39235ab6),
	.w7(32'h38dc37b8),
	.w8(32'h3909ca04),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942237b),
	.w1(32'h376fb51e),
	.w2(32'hb8b39eb6),
	.w3(32'h37ca8468),
	.w4(32'hb9079f3c),
	.w5(32'hb91e9155),
	.w6(32'h397db1db),
	.w7(32'hb8de1781),
	.w8(32'hb97bf36c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f34c08),
	.w1(32'hb8388dd4),
	.w2(32'hb8048553),
	.w3(32'h383d7bf6),
	.w4(32'hb7272f38),
	.w5(32'h34880e2a),
	.w6(32'h3799dd60),
	.w7(32'h371001f8),
	.w8(32'h375c0836),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399283b5),
	.w1(32'h3a03bb9f),
	.w2(32'h39989b99),
	.w3(32'h3a044870),
	.w4(32'h39ed9fdd),
	.w5(32'h3993c383),
	.w6(32'h3a05a65a),
	.w7(32'h39cfea79),
	.w8(32'h3961b37b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38495218),
	.w1(32'hb7f27886),
	.w2(32'h385d08eb),
	.w3(32'h382efd38),
	.w4(32'h3763bf35),
	.w5(32'hb850d60c),
	.w6(32'hb8902e32),
	.w7(32'h361f72a2),
	.w8(32'hb870064c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360f54da),
	.w1(32'hb7f866af),
	.w2(32'hb8241df3),
	.w3(32'h37ace310),
	.w4(32'hb72a7c43),
	.w5(32'hb7f62cc2),
	.w6(32'hb7a945a9),
	.w7(32'hb7f6804c),
	.w8(32'hb79cdc37),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bebf7b),
	.w1(32'h378daaa1),
	.w2(32'h37885c35),
	.w3(32'h34d146d8),
	.w4(32'h372e69e2),
	.w5(32'h3738e039),
	.w6(32'h373716f1),
	.w7(32'h378dee01),
	.w8(32'hb72db399),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e4c7d),
	.w1(32'h384798c1),
	.w2(32'hb8388104),
	.w3(32'hb82b70d0),
	.w4(32'h38ca0219),
	.w5(32'hb81ab384),
	.w6(32'h3900c3e3),
	.w7(32'hb6962ae2),
	.w8(32'hb8d95902),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d68018),
	.w1(32'h3956032b),
	.w2(32'h399b589d),
	.w3(32'h3738d9b1),
	.w4(32'h3984323c),
	.w5(32'h392f5d7f),
	.w6(32'h38d7808f),
	.w7(32'h39a55d39),
	.w8(32'h38a440a0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bf977),
	.w1(32'hb9c08d40),
	.w2(32'hb99be68f),
	.w3(32'hb8b91bd7),
	.w4(32'hb996e63b),
	.w5(32'hb948f633),
	.w6(32'hb8b41558),
	.w7(32'hb96e85e8),
	.w8(32'hb92df75e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7688df9),
	.w1(32'hb7030eff),
	.w2(32'hb67b18d7),
	.w3(32'hb6bb9eac),
	.w4(32'h35afa506),
	.w5(32'h3710b58f),
	.w6(32'h369ed816),
	.w7(32'hb612296e),
	.w8(32'h36d542f9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85ec800),
	.w1(32'hb9ad7d1d),
	.w2(32'hb98b646c),
	.w3(32'h37bddefc),
	.w4(32'hb995a10d),
	.w5(32'hb9afd57e),
	.w6(32'h3930d8b1),
	.w7(32'hb908ab2f),
	.w8(32'hb9575815),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c34f08),
	.w1(32'hb7ad7574),
	.w2(32'h38ca53e8),
	.w3(32'hb9c595e6),
	.w4(32'h38dd60fe),
	.w5(32'h392d59c6),
	.w6(32'hb8742d54),
	.w7(32'h38745518),
	.w8(32'h38e9687b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39948b25),
	.w1(32'h36512aae),
	.w2(32'hb9e13f68),
	.w3(32'h38a599ea),
	.w4(32'hb987b057),
	.w5(32'hb9a51bcb),
	.w6(32'h39ae1743),
	.w7(32'hb8ea4748),
	.w8(32'hb99de8d5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977350c),
	.w1(32'hba328c0d),
	.w2(32'h38028ad2),
	.w3(32'h395f714c),
	.w4(32'hb985b69e),
	.w5(32'hb7efed6b),
	.w6(32'hb7981abd),
	.w7(32'h3722039b),
	.w8(32'h3939b818),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953ec0c),
	.w1(32'h35b5f114),
	.w2(32'h392972ff),
	.w3(32'hb9a91698),
	.w4(32'hb86f6bd4),
	.w5(32'h396a0d7d),
	.w6(32'hb84ec679),
	.w7(32'h399423b0),
	.w8(32'h39047e9c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9303ed8),
	.w1(32'hb933d2be),
	.w2(32'h391995f5),
	.w3(32'hb9e7efde),
	.w4(32'hba2121c7),
	.w5(32'hb9874874),
	.w6(32'hb998e460),
	.w7(32'hb9db6825),
	.w8(32'hb89cef73),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1018e8),
	.w1(32'hb56261f7),
	.w2(32'hb75a6d05),
	.w3(32'h39d87d03),
	.w4(32'h391c5eca),
	.w5(32'h38916e6e),
	.w6(32'h3807be07),
	.w7(32'h388ed2f1),
	.w8(32'h38fb5b70),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3838acf5),
	.w1(32'h3836ea31),
	.w2(32'h38f5d3a9),
	.w3(32'h38c58265),
	.w4(32'h38e3c97a),
	.w5(32'h38a47a67),
	.w6(32'h38be6241),
	.w7(32'h391f74bd),
	.w8(32'h36bd98f4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fce917),
	.w1(32'hb70368db),
	.w2(32'hb6e94bae),
	.w3(32'hb889dd32),
	.w4(32'h36920f61),
	.w5(32'hb84bd8b9),
	.w6(32'h378333cc),
	.w7(32'h38458098),
	.w8(32'hb88a72e1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8363394),
	.w1(32'hb8642b7d),
	.w2(32'hb92aabcc),
	.w3(32'hb8122450),
	.w4(32'hb89dedda),
	.w5(32'hb92f7e11),
	.w6(32'h3811365c),
	.w7(32'hb8b51fe1),
	.w8(32'hb91a4ed6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a2dafa),
	.w1(32'h37b6d988),
	.w2(32'h3855d3aa),
	.w3(32'hb78a00a9),
	.w4(32'h37a8077e),
	.w5(32'h37f4b3b4),
	.w6(32'hb78223fb),
	.w7(32'hb6bdd571),
	.w8(32'hb6eb0a65),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6298d),
	.w1(32'hb94c962e),
	.w2(32'hb980472f),
	.w3(32'hb8246ecc),
	.w4(32'hb88728d7),
	.w5(32'hb826ddb6),
	.w6(32'h3799cb96),
	.w7(32'hb9a103fa),
	.w8(32'hb9b20e6a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38894f98),
	.w1(32'h38944771),
	.w2(32'hb903ca85),
	.w3(32'h36ec85d8),
	.w4(32'h37a726dd),
	.w5(32'hb92220a2),
	.w6(32'h3864525b),
	.w7(32'hb812d76d),
	.w8(32'hb9079f5d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39289dbd),
	.w1(32'hb73ac0bc),
	.w2(32'h380df396),
	.w3(32'h3980a399),
	.w4(32'hb8058c43),
	.w5(32'h38f84b80),
	.w6(32'h3905391c),
	.w7(32'h38a03bac),
	.w8(32'h3916c560),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e6e9c2),
	.w1(32'hb9143cb0),
	.w2(32'hb8a3a1b0),
	.w3(32'hb74ef2d3),
	.w4(32'hb819c65e),
	.w5(32'hb888d35c),
	.w6(32'hb87c5aef),
	.w7(32'hb8ba28c4),
	.w8(32'hb9120983),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84f09d2),
	.w1(32'hb7effbc7),
	.w2(32'hb94f3d56),
	.w3(32'hb89fda86),
	.w4(32'hb8addcbe),
	.w5(32'hb8ecb595),
	.w6(32'hb7f57126),
	.w7(32'hb97ae8ea),
	.w8(32'hb9803726),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378239cf),
	.w1(32'hb7a69142),
	.w2(32'h3889ac5e),
	.w3(32'h37f7fbe0),
	.w4(32'hb82c522d),
	.w5(32'h37e3da29),
	.w6(32'hb6be8a74),
	.w7(32'hb790b298),
	.w8(32'h373730a5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a93c06),
	.w1(32'hb866ea6a),
	.w2(32'hb89378f7),
	.w3(32'h34b9b8f6),
	.w4(32'h37228705),
	.w5(32'hb86374f6),
	.w6(32'hb8995585),
	.w7(32'hb8cfe350),
	.w8(32'hb84d6f91),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b52d2e),
	.w1(32'h3981188a),
	.w2(32'h391a0f88),
	.w3(32'h39905fdc),
	.w4(32'h38b5ef66),
	.w5(32'h37a6905b),
	.w6(32'h3651deba),
	.w7(32'h3881b4d6),
	.w8(32'h3920c893),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993b99d),
	.w1(32'h379d97a9),
	.w2(32'hb9b0dca7),
	.w3(32'h3a2b9c8d),
	.w4(32'h3979f4ac),
	.w5(32'hb99b3e1d),
	.w6(32'h3985d97f),
	.w7(32'hb9548835),
	.w8(32'hb99383c4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4565c),
	.w1(32'hb9879297),
	.w2(32'hb9187d4c),
	.w3(32'hb9a18d3a),
	.w4(32'hb95cabef),
	.w5(32'hb8ecb1d4),
	.w6(32'hb8b5594c),
	.w7(32'hb95563e3),
	.w8(32'hb950c3ba),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb867bfbe),
	.w1(32'hb7c82879),
	.w2(32'h3908460d),
	.w3(32'h379c388e),
	.w4(32'h37114742),
	.w5(32'h38aac5dc),
	.w6(32'hb85c4f35),
	.w7(32'hb8e2129c),
	.w8(32'h38f63d21),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90026f6),
	.w1(32'hb984c676),
	.w2(32'hb84a5541),
	.w3(32'hb897a077),
	.w4(32'hb990e0b4),
	.w5(32'hb82b3436),
	.w6(32'hb8d48786),
	.w7(32'hb923545b),
	.w8(32'hb8bbfc51),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b3c83),
	.w1(32'hba51010f),
	.w2(32'hba0e1e3f),
	.w3(32'h38aa65e6),
	.w4(32'hba66c1ff),
	.w5(32'hb99041eb),
	.w6(32'hb8da7b23),
	.w7(32'hba35ce79),
	.w8(32'hba3c1d5e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c877ed),
	.w1(32'h38849c5f),
	.w2(32'h38eefc86),
	.w3(32'hb89b8aab),
	.w4(32'hb88fd3e9),
	.w5(32'h378ae6b8),
	.w6(32'hb8a3af5e),
	.w7(32'hb964d2dc),
	.w8(32'hb714bfa0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d821c),
	.w1(32'hb9e1af0d),
	.w2(32'hb9d18cd8),
	.w3(32'h3807a5fd),
	.w4(32'hb9ebac47),
	.w5(32'hb9d3c378),
	.w6(32'hb8d01137),
	.w7(32'hba11e2c9),
	.w8(32'hba07d12c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807242c),
	.w1(32'hb8b8408c),
	.w2(32'hb6c517c7),
	.w3(32'h3886572a),
	.w4(32'hb934137a),
	.w5(32'hb9231c84),
	.w6(32'hb6cce1e3),
	.w7(32'hb8d0ef5a),
	.w8(32'hb991f18f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39780e36),
	.w1(32'h38d1b037),
	.w2(32'h39441db6),
	.w3(32'h3918356c),
	.w4(32'h34ad43fd),
	.w5(32'h38ec52e2),
	.w6(32'h3914b3f3),
	.w7(32'hb88f6066),
	.w8(32'hb8a81793),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77dccec),
	.w1(32'hb675f9af),
	.w2(32'hb5b43077),
	.w3(32'hb75b4218),
	.w4(32'hb6e76517),
	.w5(32'hb5edc7db),
	.w6(32'h36d4fc9f),
	.w7(32'h36bfbe0c),
	.w8(32'h370d67e9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84caf8a),
	.w1(32'hb889db2f),
	.w2(32'hb84c14cf),
	.w3(32'hb87788c1),
	.w4(32'hb8b8b3c7),
	.w5(32'hb89b2e03),
	.w6(32'hb8010a3c),
	.w7(32'hb80e321c),
	.w8(32'hb7fe44b3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3766f91a),
	.w1(32'h384ca3c3),
	.w2(32'hb7b4e5c5),
	.w3(32'hb81170c2),
	.w4(32'hb6c01cc1),
	.w5(32'hb7bb2bc0),
	.w6(32'h37e8f377),
	.w7(32'h37b2020a),
	.w8(32'hb6c4d654),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89645df),
	.w1(32'hb96c975d),
	.w2(32'hb7ac47ab),
	.w3(32'hb95652f3),
	.w4(32'hb9ac9e58),
	.w5(32'hb75678ba),
	.w6(32'hb910d9a1),
	.w7(32'hb993e057),
	.w8(32'hb983dbb5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb636d418),
	.w1(32'hb6b8c6a8),
	.w2(32'h37057130),
	.w3(32'hb7042c6f),
	.w4(32'h36bb5b1c),
	.w5(32'h372a9ffb),
	.w6(32'hb75cf367),
	.w7(32'hb5c05726),
	.w8(32'h34a6c4b0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d359cc),
	.w1(32'hb7644904),
	.w2(32'hb7f766ae),
	.w3(32'hb708a055),
	.w4(32'hb7c7e365),
	.w5(32'hb73affdf),
	.w6(32'hb7693842),
	.w7(32'hb7253f0a),
	.w8(32'hb8048d7b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa98bd),
	.w1(32'hb8b652e8),
	.w2(32'hb746b095),
	.w3(32'h37a2884c),
	.w4(32'h37a29d56),
	.w5(32'h35e686ef),
	.w6(32'hb82ec9cc),
	.w7(32'h370b7143),
	.w8(32'h3882a06b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ec7fe2),
	.w1(32'h395c2624),
	.w2(32'hb8bc60a1),
	.w3(32'hb9b4a572),
	.w4(32'hb93f8281),
	.w5(32'hb812e423),
	.w6(32'h3790a8e1),
	.w7(32'hb837fd8d),
	.w8(32'hb9c506e7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994f8a6),
	.w1(32'h39433242),
	.w2(32'hb8891ad6),
	.w3(32'h37a68734),
	.w4(32'h38d52f42),
	.w5(32'hb972bddd),
	.w6(32'h39a2f5cc),
	.w7(32'h3915f58c),
	.w8(32'hb98875b9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36baa4a3),
	.w1(32'hb783ffd3),
	.w2(32'hb78dfc78),
	.w3(32'hb7f9db88),
	.w4(32'hb7d0ad05),
	.w5(32'hb7a70307),
	.w6(32'hb72eaec6),
	.w7(32'hb7c2082d),
	.w8(32'hb8086fbe),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3581fc68),
	.w1(32'hbaa73eea),
	.w2(32'hba984a4b),
	.w3(32'h3909db72),
	.w4(32'hba43263e),
	.w5(32'hb9ef885d),
	.w6(32'hb9bdfa4a),
	.w7(32'hba2241e2),
	.w8(32'hba207d7e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39556bc7),
	.w1(32'hb9e09d39),
	.w2(32'h39470194),
	.w3(32'h39939e6e),
	.w4(32'hba0879e2),
	.w5(32'h394a0a80),
	.w6(32'h399d1661),
	.w7(32'h398a933f),
	.w8(32'h3978e306),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38433f5d),
	.w1(32'h37250a70),
	.w2(32'hb8dde65e),
	.w3(32'h369b5b6a),
	.w4(32'hb8dfd8d4),
	.w5(32'hb9937257),
	.w6(32'h38e8a84f),
	.w7(32'hb92646e0),
	.w8(32'hb9271c12),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h341007bc),
	.w1(32'h37fc5b37),
	.w2(32'h37de5f6c),
	.w3(32'hb6327775),
	.w4(32'h36787539),
	.w5(32'h36383ef1),
	.w6(32'h37e9ff49),
	.w7(32'h379fc6f2),
	.w8(32'hb7a4b900),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373486d7),
	.w1(32'hb6ad705c),
	.w2(32'hb8c0fe27),
	.w3(32'hb7eebabb),
	.w4(32'h37976ec1),
	.w5(32'hb87100e0),
	.w6(32'hb889519a),
	.w7(32'hb8e3b34b),
	.w8(32'hb8c0780f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dcb37d),
	.w1(32'hb70b54af),
	.w2(32'hb725d146),
	.w3(32'hb72308da),
	.w4(32'h359b3f0b),
	.w5(32'hb659b6d5),
	.w6(32'hb6c6d7ee),
	.w7(32'hb6a9e072),
	.w8(32'hb6c5c308),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393610b3),
	.w1(32'h38ace7b5),
	.w2(32'hb98d2ccd),
	.w3(32'h38c206f2),
	.w4(32'h3866e066),
	.w5(32'hb9149562),
	.w6(32'h378f8e87),
	.w7(32'hb88570ba),
	.w8(32'hb9921744),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7269d),
	.w1(32'hb7d6da0f),
	.w2(32'h37d49fb0),
	.w3(32'h37307302),
	.w4(32'hb849c0eb),
	.w5(32'hb951d22e),
	.w6(32'h36c90497),
	.w7(32'hb95c6da2),
	.w8(32'hb9616c90),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c20536),
	.w1(32'h37ea1c4b),
	.w2(32'h399c8387),
	.w3(32'hb92ac2f9),
	.w4(32'h3896c290),
	.w5(32'h3951cc83),
	.w6(32'hb916b6fb),
	.w7(32'h38f41081),
	.w8(32'h384e33a0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3869dc9d),
	.w1(32'h383abfd8),
	.w2(32'h38447cfb),
	.w3(32'h382c0556),
	.w4(32'hb778ad09),
	.w5(32'h37f89bec),
	.w6(32'h381a6511),
	.w7(32'h380aaa3c),
	.w8(32'h38242fec),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fae673),
	.w1(32'hb976337a),
	.w2(32'hb9182201),
	.w3(32'h3700ab76),
	.w4(32'hb8f57de4),
	.w5(32'hb8841c59),
	.w6(32'hb8b060f8),
	.w7(32'hb93e0615),
	.w8(32'hb9298076),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78ba6f4),
	.w1(32'h383c6821),
	.w2(32'hb8c5d07f),
	.w3(32'hb8a5ac18),
	.w4(32'hb88a84b2),
	.w5(32'hb9513bc2),
	.w6(32'hb8aedca8),
	.w7(32'hb8f6260b),
	.w8(32'hb960b989),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67c957e),
	.w1(32'hb61cdf6f),
	.w2(32'hb6af433f),
	.w3(32'hb5be2d4a),
	.w4(32'hb6087e42),
	.w5(32'hb6ca5aba),
	.w6(32'h3702b32f),
	.w7(32'h36451ce4),
	.w8(32'h36904b27),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379d279d),
	.w1(32'hb8af86ae),
	.w2(32'h388d29e6),
	.w3(32'hb98c4c46),
	.w4(32'hb92f50fa),
	.w5(32'h35b4164a),
	.w6(32'hb803f7c4),
	.w7(32'hb9a44758),
	.w8(32'hb97a1224),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68ca302),
	.w1(32'hb6c9ce3e),
	.w2(32'hb6fe047d),
	.w3(32'hb63ff162),
	.w4(32'hb51e81cc),
	.w5(32'hb6604f21),
	.w6(32'h36fd3318),
	.w7(32'h372b359f),
	.w8(32'h37224f83),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8afe7ff),
	.w1(32'hb965194c),
	.w2(32'hb970969f),
	.w3(32'hb7aba15d),
	.w4(32'hb904d34e),
	.w5(32'hb90162b7),
	.w6(32'hb88f8b3c),
	.w7(32'hb95d0df0),
	.w8(32'hb950c86e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387c6114),
	.w1(32'h3969450d),
	.w2(32'h39ae94af),
	.w3(32'h390f5675),
	.w4(32'h39bf1ef1),
	.w5(32'h39ace08e),
	.w6(32'h390a64e9),
	.w7(32'h39a803b1),
	.w8(32'h394ea484),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387a80c5),
	.w1(32'h385c7bed),
	.w2(32'h39055ce7),
	.w3(32'h38820cf4),
	.w4(32'h387e70d9),
	.w5(32'h38905779),
	.w6(32'h36e1aac2),
	.w7(32'h3809bdd7),
	.w8(32'h364f0f46),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73736aa),
	.w1(32'hb6b9580c),
	.w2(32'h353d221d),
	.w3(32'h368af9ac),
	.w4(32'h374141db),
	.w5(32'hb6e0eb25),
	.w6(32'h3792b3ac),
	.w7(32'hb711ac6f),
	.w8(32'hb79db314),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ee779),
	.w1(32'hb88aa8d3),
	.w2(32'h3919f615),
	.w3(32'h37d3193b),
	.w4(32'hb85ebfd8),
	.w5(32'h38f7bfe2),
	.w6(32'hb84e44d2),
	.w7(32'h389b6609),
	.w8(32'h38ae3899),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df5c5c),
	.w1(32'hb975ccdb),
	.w2(32'hb8dd7cfc),
	.w3(32'hb9497617),
	.w4(32'hb95c7163),
	.w5(32'hb84316d7),
	.w6(32'hb91595ec),
	.w7(32'hb972c7a2),
	.w8(32'hb92bd144),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e9418),
	.w1(32'hb944fcbc),
	.w2(32'hb9310b71),
	.w3(32'h395a3e54),
	.w4(32'hb8792c4c),
	.w5(32'hb8f109d8),
	.w6(32'h3916c498),
	.w7(32'hb8b99e76),
	.w8(32'hb92e4d47),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84677ea),
	.w1(32'h378bf7e9),
	.w2(32'h37cefe59),
	.w3(32'hb7fa5baf),
	.w4(32'h378f16a2),
	.w5(32'h36cb0642),
	.w6(32'h373b4a0c),
	.w7(32'h366b9d7e),
	.w8(32'hb6bad3dc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb56c9371),
	.w1(32'h369edecc),
	.w2(32'h36f4a9a2),
	.w3(32'hb6954df8),
	.w4(32'h367fcb1c),
	.w5(32'h36d94f53),
	.w6(32'hb3502672),
	.w7(32'h3657c791),
	.w8(32'hb6d8d54c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ba0dc),
	.w1(32'hb91cca85),
	.w2(32'hb9d45cab),
	.w3(32'h396ef4fd),
	.w4(32'h397b4013),
	.w5(32'hb9523e02),
	.w6(32'hb90deba6),
	.w7(32'hb9fbd0ac),
	.w8(32'hb949d488),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912d47b),
	.w1(32'hb7ac33ae),
	.w2(32'hb98c7c0e),
	.w3(32'h39c276a4),
	.w4(32'hb81f46c1),
	.w5(32'hb905a2cd),
	.w6(32'h385fedbc),
	.w7(32'hb9d61220),
	.w8(32'hb9b68328),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886190c),
	.w1(32'h3906332a),
	.w2(32'h395b9781),
	.w3(32'h39472584),
	.w4(32'h399c99a2),
	.w5(32'h396a58ca),
	.w6(32'h3834d63d),
	.w7(32'h390af5ef),
	.w8(32'h39389b4e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942c50e),
	.w1(32'hb86ae14f),
	.w2(32'hba0220bb),
	.w3(32'hb9873e21),
	.w4(32'hba0659b8),
	.w5(32'hb9eecdb3),
	.w6(32'h39d01034),
	.w7(32'hb9fa9232),
	.w8(32'hba3950b8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb713d11d),
	.w1(32'hb8bbef40),
	.w2(32'hb84ca677),
	.w3(32'hb807c447),
	.w4(32'hb8b6a91a),
	.w5(32'hb70464d5),
	.w6(32'hb7600315),
	.w7(32'hb8d4df63),
	.w8(32'hb8d2be42),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b9cb45),
	.w1(32'hb8286815),
	.w2(32'h384cb4b4),
	.w3(32'hb794331a),
	.w4(32'hb7948ede),
	.w5(32'h38529677),
	.w6(32'hb847a722),
	.w7(32'hb87aa397),
	.w8(32'hb7d04f2e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d53a11),
	.w1(32'h39a64f1a),
	.w2(32'hba2e3451),
	.w3(32'h3968c48f),
	.w4(32'hb8189905),
	.w5(32'hba5b5591),
	.w6(32'h39ec8ab6),
	.w7(32'hb9481bee),
	.w8(32'hb9935632),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9565b06),
	.w1(32'hba237f50),
	.w2(32'hba1dcf7a),
	.w3(32'h3878eca9),
	.w4(32'hb9dc44ad),
	.w5(32'hb99dc7e6),
	.w6(32'hb8fae17e),
	.w7(32'hba2056a9),
	.w8(32'hba10a437),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39680aca),
	.w1(32'hb8526f35),
	.w2(32'hb9d37f43),
	.w3(32'h37ff3aeb),
	.w4(32'hb8139a11),
	.w5(32'hb9ce5900),
	.w6(32'h391d9e8c),
	.w7(32'hb981212a),
	.w8(32'hba0bb555),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a88d34),
	.w1(32'h3975c246),
	.w2(32'h391cb06d),
	.w3(32'h392aa10d),
	.w4(32'h397d41da),
	.w5(32'h38a0d991),
	.w6(32'h39713f55),
	.w7(32'h3993197a),
	.w8(32'h38d33612),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3cff4),
	.w1(32'h3901f77e),
	.w2(32'h3960e9af),
	.w3(32'h391264c9),
	.w4(32'h3957ed71),
	.w5(32'h394f3e0e),
	.w6(32'h3932fa31),
	.w7(32'h39bc7555),
	.w8(32'h39911c6d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816bece),
	.w1(32'h366bfd8c),
	.w2(32'h3607eb9c),
	.w3(32'hb8155d41),
	.w4(32'h36c2c1ed),
	.w5(32'h36814a9d),
	.w6(32'h360b76fd),
	.w7(32'h35012146),
	.w8(32'hb5bd58ba),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e53495),
	.w1(32'hb75986f3),
	.w2(32'h341f3148),
	.w3(32'h365490e9),
	.w4(32'h3615f779),
	.w5(32'h370fa6f7),
	.w6(32'hb65d63de),
	.w7(32'h36e94936),
	.w8(32'h372de7ba),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a85fbe),
	.w1(32'h37478895),
	.w2(32'hb8c79318),
	.w3(32'hb512f27d),
	.w4(32'hb800efc1),
	.w5(32'hb7d6af41),
	.w6(32'hb819a328),
	.w7(32'hb8fd3e6b),
	.w8(32'hb941eb88),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84d62ed),
	.w1(32'h36a368e8),
	.w2(32'h36a27cff),
	.w3(32'hb83dd342),
	.w4(32'hb72fa23c),
	.w5(32'h361183e7),
	.w6(32'h37286955),
	.w7(32'h37399990),
	.w8(32'hb7863034),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb659e32c),
	.w1(32'h37136747),
	.w2(32'hb91fb302),
	.w3(32'hb8de33bf),
	.w4(32'hb8d06b24),
	.w5(32'hb96fda4e),
	.w6(32'hb8a2a0d3),
	.w7(32'hb9338705),
	.w8(32'hb9362a16),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915e6eb),
	.w1(32'h38e338d3),
	.w2(32'hb5e8da11),
	.w3(32'h399e1475),
	.w4(32'h3905e14c),
	.w5(32'h399b2a8a),
	.w6(32'h394389c0),
	.w7(32'hb8c1a58b),
	.w8(32'hb8c3b9ce),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac8912),
	.w1(32'h37fd4382),
	.w2(32'h37adc6e4),
	.w3(32'h38994371),
	.w4(32'h38adfa5e),
	.w5(32'h3763ca00),
	.w6(32'h386615fd),
	.w7(32'h384c2d2f),
	.w8(32'h3833a587),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fce420),
	.w1(32'hb74e9b41),
	.w2(32'h3791151b),
	.w3(32'hb64a74ad),
	.w4(32'h36afef6d),
	.w5(32'h37a944b0),
	.w6(32'hb625ddaa),
	.w7(32'h3699b0b5),
	.w8(32'h37f4a9ce),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39887cd3),
	.w1(32'hb88dc70d),
	.w2(32'hba43a255),
	.w3(32'h398dd311),
	.w4(32'h391516ca),
	.w5(32'hb9bf3da2),
	.w6(32'h38cbbd16),
	.w7(32'hb9da4cdc),
	.w8(32'hba71a89e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380bc807),
	.w1(32'hb95582fd),
	.w2(32'hb980c7e3),
	.w3(32'h38d24687),
	.w4(32'hb8bdc7ca),
	.w5(32'hb921bd2c),
	.w6(32'h3762fcbe),
	.w7(32'hb9559224),
	.w8(32'hb9a7e64d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36830fde),
	.w1(32'h3672acc2),
	.w2(32'hb601e623),
	.w3(32'hb69e058d),
	.w4(32'hb6e9634e),
	.w5(32'hb6b189c8),
	.w6(32'h36628b49),
	.w7(32'hb60f4830),
	.w8(32'h3593df8c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e2f72f),
	.w1(32'hb9863182),
	.w2(32'hb9e773b0),
	.w3(32'hb7052a7a),
	.w4(32'hb9885a30),
	.w5(32'hb9a00e44),
	.w6(32'h389d36e3),
	.w7(32'hb96d26ef),
	.w8(32'hb9afab30),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885c050),
	.w1(32'hb8d781f2),
	.w2(32'hb8edf631),
	.w3(32'hb8905881),
	.w4(32'hb899149a),
	.w5(32'hb86600f1),
	.w6(32'hb886406b),
	.w7(32'hb89d8a82),
	.w8(32'hb8638ba6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72913dc),
	.w1(32'hb7250b87),
	.w2(32'h37dba001),
	.w3(32'h34f4ec2b),
	.w4(32'hb7faa42c),
	.w5(32'h35ccf6e4),
	.w6(32'hb84a8b6d),
	.w7(32'hb8306ec5),
	.w8(32'hb79f6506),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h346ac000),
	.w1(32'h3699ddbd),
	.w2(32'h368e37b2),
	.w3(32'h35da4bbd),
	.w4(32'hb6f81c38),
	.w5(32'hb688103b),
	.w6(32'h35335d25),
	.w7(32'hb6b600ae),
	.w8(32'h3238fe35),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7292784),
	.w1(32'h3433a055),
	.w2(32'hb7a7c8c4),
	.w3(32'hb79dbca1),
	.w4(32'hb597dd45),
	.w5(32'hb70a0c80),
	.w6(32'h36988c71),
	.w7(32'hb7456e15),
	.w8(32'hb7393eac),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68128e4),
	.w1(32'h38b525cd),
	.w2(32'h363d78e7),
	.w3(32'h38432900),
	.w4(32'h38d6b014),
	.w5(32'h37dc36fe),
	.w6(32'h38e44f5d),
	.w7(32'h3900f7fd),
	.w8(32'h388e1dca),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389382f9),
	.w1(32'hb98bef77),
	.w2(32'hb9c45ebd),
	.w3(32'hb8b018c8),
	.w4(32'hba1f3b2f),
	.w5(32'hb9e7cb9a),
	.w6(32'h3899be03),
	.w7(32'hb9a22a7a),
	.w8(32'hba0056cb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a6bc02),
	.w1(32'hb9a41b5a),
	.w2(32'hb9add0c7),
	.w3(32'h38971d6f),
	.w4(32'hb98e684d),
	.w5(32'hb9602955),
	.w6(32'h3883e65e),
	.w7(32'hb9788ff3),
	.w8(32'hb9940b0c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f95f9),
	.w1(32'hb9bd13ab),
	.w2(32'hb9c5bf36),
	.w3(32'h38c9f606),
	.w4(32'hb9c363ca),
	.w5(32'hb9837d05),
	.w6(32'h39282ef8),
	.w7(32'hb9eb38c5),
	.w8(32'hb9aeb90d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d3bb58),
	.w1(32'hb824ada1),
	.w2(32'hb833e0d2),
	.w3(32'hb7b112b5),
	.w4(32'hb842f8cf),
	.w5(32'hb82a45e7),
	.w6(32'hb7d72d6a),
	.w7(32'hb8093716),
	.w8(32'hb827a0ac),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d9bce8),
	.w1(32'hb84c4624),
	.w2(32'h380a0f3d),
	.w3(32'hb81142a0),
	.w4(32'hb85b864a),
	.w5(32'h36b21a26),
	.w6(32'hb7f2c76d),
	.w7(32'hb83e9c73),
	.w8(32'hb761653c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76c5dc3),
	.w1(32'h37b62c26),
	.w2(32'h37a849ec),
	.w3(32'h3759abd0),
	.w4(32'h37d04ee6),
	.w5(32'h37dda8e7),
	.w6(32'h379097c3),
	.w7(32'h36db5386),
	.w8(32'h35d470fb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb498c12c),
	.w1(32'hb5f529e8),
	.w2(32'h35d5a6ee),
	.w3(32'hb6bc0497),
	.w4(32'hb6cfdd06),
	.w5(32'hb60c5877),
	.w6(32'h35983207),
	.w7(32'h36781a70),
	.w8(32'h36bc2406),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ff8f46),
	.w1(32'hb9a2acc0),
	.w2(32'h386b7f20),
	.w3(32'hb81ce061),
	.w4(32'hb9b17125),
	.w5(32'hb89eb959),
	.w6(32'hb948b10b),
	.w7(32'hb9b7836c),
	.w8(32'hb99418b4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f0b4a),
	.w1(32'h38bee58a),
	.w2(32'h38fa21a1),
	.w3(32'h38c688be),
	.w4(32'h38fb264e),
	.w5(32'h38ab1370),
	.w6(32'h36350709),
	.w7(32'h3830932c),
	.w8(32'h37c6afea),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cbced2),
	.w1(32'hb8c25db0),
	.w2(32'hb8c015e3),
	.w3(32'hb8ee6dcc),
	.w4(32'hb9083ffd),
	.w5(32'hb9034f53),
	.w6(32'hb8a13eea),
	.w7(32'hb8ccf962),
	.w8(32'hb8b102d0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78c8584),
	.w1(32'hb932b4fe),
	.w2(32'hb890cfd5),
	.w3(32'hb925c92d),
	.w4(32'hb972b212),
	.w5(32'hb8c69a78),
	.w6(32'hb96148fb),
	.w7(32'hb952a991),
	.w8(32'hb90c73e4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fb4094),
	.w1(32'hb811ec64),
	.w2(32'hb7aa01a9),
	.w3(32'h37797d1f),
	.w4(32'hb6b8ea5c),
	.w5(32'hb4b0d258),
	.w6(32'h37368ae8),
	.w7(32'h3722dbe3),
	.w8(32'h37998382),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb760920f),
	.w1(32'hb916b810),
	.w2(32'hb8a87457),
	.w3(32'h37109e79),
	.w4(32'hb8e61a35),
	.w5(32'hb7fb69eb),
	.w6(32'hb75a2cc5),
	.w7(32'hb8b9528d),
	.w8(32'hb89f8629),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377bd734),
	.w1(32'hb710334e),
	.w2(32'h384e635c),
	.w3(32'hb7c0f5d5),
	.w4(32'hb80a577c),
	.w5(32'h37d3044d),
	.w6(32'hb84538d1),
	.w7(32'hb80d0aad),
	.w8(32'hb7f92433),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b0f2c),
	.w1(32'hba1d81f2),
	.w2(32'hb8472292),
	.w3(32'hb924c855),
	.w4(32'hba82c356),
	.w5(32'hb9f4bfcd),
	.w6(32'hb9e20a3b),
	.w7(32'hba84eace),
	.w8(32'hba802a9f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80537c0),
	.w1(32'hbaa48879),
	.w2(32'hbb05c2f0),
	.w3(32'hb56d0006),
	.w4(32'hba2bfbb9),
	.w5(32'hbac8edc0),
	.w6(32'hba751114),
	.w7(32'hba8f3d76),
	.w8(32'hba8baa1f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabda56a),
	.w1(32'hb9ab99c8),
	.w2(32'hba7f50a8),
	.w3(32'hba8a46c9),
	.w4(32'h399b0cb9),
	.w5(32'hba36343e),
	.w6(32'hb97df94c),
	.w7(32'hba00a16d),
	.w8(32'hb844bb9e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule