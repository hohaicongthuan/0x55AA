module layer_10_featuremap_370(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c077c36),
	.w1(32'hbb288c8a),
	.w2(32'h3be4ff0a),
	.w3(32'h3bf003b2),
	.w4(32'h3b39e58f),
	.w5(32'hbc2c8e4f),
	.w6(32'h3bb56f0b),
	.w7(32'hbb188a0a),
	.w8(32'h3c5fb684),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4fa8db),
	.w1(32'h3b9b9121),
	.w2(32'hbb71c5f4),
	.w3(32'hbb74892e),
	.w4(32'h399e211d),
	.w5(32'hbb1a7057),
	.w6(32'h3be9ead9),
	.w7(32'h3c3ad8ba),
	.w8(32'hbb18ea7b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c736b35),
	.w1(32'hbb8fbdd3),
	.w2(32'h3c0ed351),
	.w3(32'hbbcbd69d),
	.w4(32'h3c2d7fa0),
	.w5(32'h3b6acf9b),
	.w6(32'hbc9e0c34),
	.w7(32'h3bb16c1f),
	.w8(32'hbad8755f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c6e0d),
	.w1(32'hbcac0bc3),
	.w2(32'h3bd5e216),
	.w3(32'hbcb7ce12),
	.w4(32'h3ac3bc3f),
	.w5(32'hbc9ab908),
	.w6(32'h3adb1b95),
	.w7(32'h3bc40dd2),
	.w8(32'h3b81ff5b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10b9f3),
	.w1(32'hbc5016c2),
	.w2(32'h3b9eeef7),
	.w3(32'h3b46278f),
	.w4(32'h3a95063a),
	.w5(32'hb7ccf3e8),
	.w6(32'hbb268fa7),
	.w7(32'hbbf30ccc),
	.w8(32'h3c5d48c6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12278a),
	.w1(32'hbb5d55ef),
	.w2(32'h39a96768),
	.w3(32'h3b4b6c4d),
	.w4(32'h3b9fec17),
	.w5(32'h3bd5287a),
	.w6(32'hb98c6f8b),
	.w7(32'h3aa567dc),
	.w8(32'h3b937eb2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80805),
	.w1(32'hbb8c4321),
	.w2(32'hbbcdc7b9),
	.w3(32'h3c24e8b3),
	.w4(32'hbd18e1a6),
	.w5(32'hbc363d4e),
	.w6(32'hbc06244a),
	.w7(32'hbbaf60df),
	.w8(32'hbbbc106c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37739),
	.w1(32'hbb2438a6),
	.w2(32'hba11ed8c),
	.w3(32'hbcd840f8),
	.w4(32'h3bacb9cb),
	.w5(32'hbbe992a8),
	.w6(32'hbc8c47e3),
	.w7(32'h3b005f6d),
	.w8(32'h3a9e225f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cc441),
	.w1(32'hbbc6b76a),
	.w2(32'hbccf2efa),
	.w3(32'hbb783093),
	.w4(32'hbb887fc9),
	.w5(32'h3b8b922d),
	.w6(32'h3c1cc9a5),
	.w7(32'h3b9301c6),
	.w8(32'hba95e6b0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d6778),
	.w1(32'hbbf91980),
	.w2(32'hbbea70aa),
	.w3(32'h3c8efaa2),
	.w4(32'h3bae3848),
	.w5(32'hb9b91585),
	.w6(32'hbb8a00aa),
	.w7(32'hbc96aa3c),
	.w8(32'h384fde80),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0edfe3),
	.w1(32'hbbf1e680),
	.w2(32'hbb089b2f),
	.w3(32'h3bacd971),
	.w4(32'h3b10f207),
	.w5(32'h3c887c5c),
	.w6(32'hbb369688),
	.w7(32'hbb56caf9),
	.w8(32'hbb7bc8d9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9d75),
	.w1(32'h3c01e7c9),
	.w2(32'h3ca13d68),
	.w3(32'h3b83a0b8),
	.w4(32'h3c972a09),
	.w5(32'hb958cc6e),
	.w6(32'h3b798b64),
	.w7(32'hbb1cbc00),
	.w8(32'h3c41317b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c8b0f),
	.w1(32'h3c098dda),
	.w2(32'h3a5a93f0),
	.w3(32'h3c5660df),
	.w4(32'hbbceb354),
	.w5(32'h3b0094c4),
	.w6(32'hba1318a4),
	.w7(32'hbc1300a7),
	.w8(32'hbca54552),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa7d73),
	.w1(32'h3beb2152),
	.w2(32'hbba06aa6),
	.w3(32'h3be8674c),
	.w4(32'hbd8aafaa),
	.w5(32'hbcd40e76),
	.w6(32'hbd4b1c44),
	.w7(32'h3ca1778f),
	.w8(32'hbbd8d7ed),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6fb58),
	.w1(32'h3a617251),
	.w2(32'h3b3a691a),
	.w3(32'hbb9138d3),
	.w4(32'hbb6ca079),
	.w5(32'h3b96d1e4),
	.w6(32'hbb2d58c7),
	.w7(32'h3b826513),
	.w8(32'h3a94c83e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52178f),
	.w1(32'h3bba68ad),
	.w2(32'hbc296e38),
	.w3(32'hbc35bdc4),
	.w4(32'h3bbafa90),
	.w5(32'h3b9f892b),
	.w6(32'hbac55db6),
	.w7(32'hbb39f20c),
	.w8(32'h3d0f3c6b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb196d91),
	.w1(32'hbbaf989a),
	.w2(32'h3ba96eae),
	.w3(32'h3beee1c5),
	.w4(32'hb7a973d9),
	.w5(32'hbc77ed83),
	.w6(32'hbb1cd703),
	.w7(32'hbadc4761),
	.w8(32'h3b37e011),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75f776),
	.w1(32'hbd6ed792),
	.w2(32'hba1305f0),
	.w3(32'hbae20628),
	.w4(32'hbbfdee17),
	.w5(32'hbb0d1e4c),
	.w6(32'hbc3db07d),
	.w7(32'h3cd92a75),
	.w8(32'hbbd866bd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c877e36),
	.w1(32'h3cab7150),
	.w2(32'h3b982afb),
	.w3(32'h3ad718c3),
	.w4(32'hba0cc2dc),
	.w5(32'h3c56b5a9),
	.w6(32'h3c234ac7),
	.w7(32'h3bafd891),
	.w8(32'hba821552),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd3220a),
	.w1(32'hbbfb0dd6),
	.w2(32'h3c6aa87d),
	.w3(32'h3b649e7e),
	.w4(32'hbc9e366a),
	.w5(32'h3badbe95),
	.w6(32'hbc45e38c),
	.w7(32'h3a7eeef8),
	.w8(32'hbb919aed),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc6557),
	.w1(32'hbb52a4b8),
	.w2(32'hbc792745),
	.w3(32'hbb968e37),
	.w4(32'hbc05356c),
	.w5(32'h3be5adec),
	.w6(32'h3b6b2712),
	.w7(32'h3b0b8b07),
	.w8(32'hbbb81b64),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b0ea5),
	.w1(32'hbbf36a73),
	.w2(32'hbabe5565),
	.w3(32'h3b31554f),
	.w4(32'h3a4c2e8c),
	.w5(32'hbc479966),
	.w6(32'hbc3b0f44),
	.w7(32'h3a44252a),
	.w8(32'h3b41801c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12e67c),
	.w1(32'hba6022cc),
	.w2(32'h3c41ca06),
	.w3(32'h3bdd9949),
	.w4(32'h3b46f50b),
	.w5(32'hbbbc2009),
	.w6(32'hba053d38),
	.w7(32'h3b91a265),
	.w8(32'hbcb4d20f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6be98),
	.w1(32'h3be72d83),
	.w2(32'h3c32157d),
	.w3(32'hbb6ab509),
	.w4(32'h394d79d6),
	.w5(32'hbb97a8eb),
	.w6(32'hbbdbad7a),
	.w7(32'h3bf05ba5),
	.w8(32'h3b979ce7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8016f),
	.w1(32'hbc5c215a),
	.w2(32'hbb65037b),
	.w3(32'hb909483e),
	.w4(32'hb90a49e9),
	.w5(32'hbb6ec7de),
	.w6(32'h3c6c47fc),
	.w7(32'h3b1f17e4),
	.w8(32'h3b761b7b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca11840),
	.w1(32'hbc574f19),
	.w2(32'hbc2d9987),
	.w3(32'hbc14dcc0),
	.w4(32'hbc9473ce),
	.w5(32'hbb25f8fd),
	.w6(32'h3c1fae12),
	.w7(32'h3b1ccfcf),
	.w8(32'hba93256c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e895f),
	.w1(32'hbcdc1ed4),
	.w2(32'h3b6f213d),
	.w3(32'hbab2e167),
	.w4(32'hbbbf4e6b),
	.w5(32'hbbb49acb),
	.w6(32'h3bfa296e),
	.w7(32'h3aa557f2),
	.w8(32'h3a57fb32),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6056e6),
	.w1(32'h3ad4223e),
	.w2(32'h3cc6a449),
	.w3(32'hbab078e6),
	.w4(32'h3ba704c2),
	.w5(32'hbb242b65),
	.w6(32'h3bb42745),
	.w7(32'h3c883894),
	.w8(32'h3baf0d4f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba745cb6),
	.w1(32'h3aba481b),
	.w2(32'hbd067d88),
	.w3(32'h3c862d98),
	.w4(32'h3b9957b4),
	.w5(32'h3adb7ed8),
	.w6(32'hbc2273cb),
	.w7(32'hbbffe3b6),
	.w8(32'hbb0c1688),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5119b),
	.w1(32'h3bc12fbe),
	.w2(32'h3bafd150),
	.w3(32'h3b4ccef4),
	.w4(32'h3bcb6c71),
	.w5(32'hbc8878ed),
	.w6(32'h3c5e496a),
	.w7(32'hbbc9e180),
	.w8(32'h3b61fa74),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f31ed),
	.w1(32'hba7bc559),
	.w2(32'h3c4bc0bc),
	.w3(32'hbc71d7a2),
	.w4(32'hbc54aeb7),
	.w5(32'hbbe0072b),
	.w6(32'hbc31691d),
	.w7(32'h3a221816),
	.w8(32'h3bd0d05e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab517db),
	.w1(32'hbbbf1c22),
	.w2(32'h3c07ea85),
	.w3(32'h3c315e60),
	.w4(32'hbbe29209),
	.w5(32'hbd4dbcce),
	.w6(32'hbb830832),
	.w7(32'h3bb19636),
	.w8(32'h3b05c789),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c866a0f),
	.w1(32'h3b922756),
	.w2(32'hbc218186),
	.w3(32'hbb83b42d),
	.w4(32'hbacfbbd5),
	.w5(32'hbc4a96b0),
	.w6(32'hbc0f3278),
	.w7(32'hba95ba7d),
	.w8(32'hbb8fa8f1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c5987),
	.w1(32'h3d52bed3),
	.w2(32'hba975271),
	.w3(32'h3b68adae),
	.w4(32'h3bd8112b),
	.w5(32'h3bb2b974),
	.w6(32'h3aa19337),
	.w7(32'hbb436ae9),
	.w8(32'hbc02cefc),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd32935),
	.w1(32'hbb089969),
	.w2(32'hbb8ed878),
	.w3(32'h3b24f88a),
	.w4(32'h3bfca91f),
	.w5(32'hbbe000f1),
	.w6(32'h3bcca661),
	.w7(32'h3c470d2a),
	.w8(32'hbd85e3d7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4926ad),
	.w1(32'h3b66e553),
	.w2(32'h3c6175a5),
	.w3(32'hbc422187),
	.w4(32'h3c0eab9d),
	.w5(32'h3bcf7b8c),
	.w6(32'hbbbea61c),
	.w7(32'h39a32ddd),
	.w8(32'hbbefc521),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9c91d),
	.w1(32'hbc0f97ae),
	.w2(32'hbb9b243a),
	.w3(32'hbb14005c),
	.w4(32'hbb8b8ae7),
	.w5(32'hb9c6f011),
	.w6(32'hbb7f99b8),
	.w7(32'h3a11d6fe),
	.w8(32'hbc370327),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72cf96),
	.w1(32'h3ab69a0e),
	.w2(32'hbcf6ba31),
	.w3(32'h3c8cd2b9),
	.w4(32'hbc41cdff),
	.w5(32'hbb6896cb),
	.w6(32'h3ab05636),
	.w7(32'h3c1ba096),
	.w8(32'hbc3ab7f1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9a013),
	.w1(32'hbbbd08b2),
	.w2(32'hbb48497f),
	.w3(32'h3c94573c),
	.w4(32'hbbb0ff21),
	.w5(32'hbcb59cc4),
	.w6(32'h3b82a8f4),
	.w7(32'h3b8ab7b9),
	.w8(32'hbb9555e5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f57cd),
	.w1(32'hb7813cd9),
	.w2(32'h3896f65b),
	.w3(32'hba085147),
	.w4(32'hbb587fdc),
	.w5(32'h3c369d30),
	.w6(32'h3c36f32d),
	.w7(32'h3bfca73b),
	.w8(32'hbc994b9e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b7c9f),
	.w1(32'h3c000b08),
	.w2(32'h3c309992),
	.w3(32'h3ca9e2e3),
	.w4(32'h3ad18d01),
	.w5(32'h3b8869aa),
	.w6(32'h3ab095bc),
	.w7(32'h3c368242),
	.w8(32'hbaab8b0e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf958b8),
	.w1(32'hbb3bd5c0),
	.w2(32'hbad6f351),
	.w3(32'hbc3591e1),
	.w4(32'hbb3e948a),
	.w5(32'h3bd567cc),
	.w6(32'h3c5175d9),
	.w7(32'h3c5eb435),
	.w8(32'h3babf45a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedc85d),
	.w1(32'h3b98c116),
	.w2(32'h39ef56a6),
	.w3(32'hbb8f6aad),
	.w4(32'hb9d1ba87),
	.w5(32'hb9c37cf2),
	.w6(32'hbd187465),
	.w7(32'h3c0f950f),
	.w8(32'h3b32fe52),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35adb4),
	.w1(32'h3ae97cdb),
	.w2(32'hbbc5fdfe),
	.w3(32'h3b956eb7),
	.w4(32'h3af1e618),
	.w5(32'hbb275b89),
	.w6(32'hbc45077d),
	.w7(32'h3bf3130b),
	.w8(32'h3a89229c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0ed89),
	.w1(32'h3c7b41cf),
	.w2(32'h3b9e2e5a),
	.w3(32'h3b0b6998),
	.w4(32'hb79e2354),
	.w5(32'h3b355f35),
	.w6(32'h3af96c89),
	.w7(32'hbb46bf62),
	.w8(32'hba2048c9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3d2bd),
	.w1(32'hbb9a99b1),
	.w2(32'hba3cb007),
	.w3(32'hbbfa4977),
	.w4(32'h3bcec353),
	.w5(32'hbc918112),
	.w6(32'hbbfdd305),
	.w7(32'hbc180090),
	.w8(32'h3bd71c1d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d8335),
	.w1(32'hbaa4f5d8),
	.w2(32'h3bd74866),
	.w3(32'hbc610c23),
	.w4(32'hba641462),
	.w5(32'hbb69e605),
	.w6(32'hb8b16927),
	.w7(32'hbc7dd49c),
	.w8(32'h3c3cc0e1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97242d),
	.w1(32'hbb8dcea6),
	.w2(32'h3b530104),
	.w3(32'h3c6842f5),
	.w4(32'h3ba66be3),
	.w5(32'h3b8e2ce2),
	.w6(32'h3a3d92c6),
	.w7(32'hbcb4b3d8),
	.w8(32'hbcdc3367),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0cb5c),
	.w1(32'h39c6c633),
	.w2(32'hbc4f7b55),
	.w3(32'h3bb6dae3),
	.w4(32'h3b5fe440),
	.w5(32'h3ba46142),
	.w6(32'h3c2549f0),
	.w7(32'h3c0305c8),
	.w8(32'h3be5d92a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba5c58),
	.w1(32'h3c57e42d),
	.w2(32'hbd70d609),
	.w3(32'hbd1015e7),
	.w4(32'hbca3a8c8),
	.w5(32'h3ba68f58),
	.w6(32'h3b05756f),
	.w7(32'h3b2d0b0a),
	.w8(32'h3bc59780),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dd000),
	.w1(32'h3b39de18),
	.w2(32'h3b15fe2b),
	.w3(32'h3b923276),
	.w4(32'hbb69107e),
	.w5(32'hb9cc60fd),
	.w6(32'hbb1183d9),
	.w7(32'hbb90aed3),
	.w8(32'h3bcb8745),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9507de),
	.w1(32'h3b23834b),
	.w2(32'h3bcb996f),
	.w3(32'h3ce189e8),
	.w4(32'hbb941297),
	.w5(32'h3b1ddd03),
	.w6(32'h3bb92222),
	.w7(32'hb97618f2),
	.w8(32'hbb0dd3f0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95cda3),
	.w1(32'hbba2776a),
	.w2(32'hbc15d524),
	.w3(32'hbc0f42a8),
	.w4(32'h3b981634),
	.w5(32'h3b96a86b),
	.w6(32'hbbb17bcb),
	.w7(32'h3af9ba0d),
	.w8(32'h3c97db50),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1732c7),
	.w1(32'hbd56bacc),
	.w2(32'h3bfbf88f),
	.w3(32'h3bba8e95),
	.w4(32'hbc2f57c0),
	.w5(32'hbb9cb95f),
	.w6(32'h3b0659db),
	.w7(32'hbc1c99a8),
	.w8(32'h3be49625),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058eb5),
	.w1(32'hbc04f997),
	.w2(32'h3bcf939e),
	.w3(32'h3bfe290a),
	.w4(32'h3c277cf5),
	.w5(32'hbc022623),
	.w6(32'h3a0ca469),
	.w7(32'hbb99172d),
	.w8(32'h3b1811c9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa888a),
	.w1(32'h3b61b93c),
	.w2(32'hbc21ff64),
	.w3(32'hbcddb313),
	.w4(32'h3c390a11),
	.w5(32'h3bb7b9ee),
	.w6(32'hba4da650),
	.w7(32'hbbc5f4cc),
	.w8(32'hbb8eb0f0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5785e4),
	.w1(32'h38a71e31),
	.w2(32'hbc0ba29e),
	.w3(32'h3ccca85e),
	.w4(32'hbbb6c337),
	.w5(32'h3bfb569f),
	.w6(32'hba59aeca),
	.w7(32'hba126545),
	.w8(32'hbc613d36),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbf78f),
	.w1(32'hbaf1ea22),
	.w2(32'h3c91b199),
	.w3(32'hb918bad4),
	.w4(32'hba80a59b),
	.w5(32'h3bc3e765),
	.w6(32'h3b99f6ae),
	.w7(32'hbb5781f2),
	.w8(32'h3cbab3d8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b14ed),
	.w1(32'hb926eab3),
	.w2(32'hbba37123),
	.w3(32'h3b5546cd),
	.w4(32'h3b1e3a09),
	.w5(32'hbb50b817),
	.w6(32'hbc1af575),
	.w7(32'hbd62399f),
	.w8(32'hb69e37c0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841936),
	.w1(32'h3c236f5b),
	.w2(32'h3af282bf),
	.w3(32'h3d49b24a),
	.w4(32'h3a2e18a7),
	.w5(32'h3c3c328d),
	.w6(32'hba96029b),
	.w7(32'h3bededf0),
	.w8(32'h3c736dc6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981fd6f),
	.w1(32'h3bca1111),
	.w2(32'h3bb60dcf),
	.w3(32'hba92fd25),
	.w4(32'hbad49274),
	.w5(32'hbb851047),
	.w6(32'hbc8a2c60),
	.w7(32'hbbb0955e),
	.w8(32'hbaef2fb2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc398c46),
	.w1(32'h3b8fc602),
	.w2(32'hbab8de73),
	.w3(32'hbb7a143a),
	.w4(32'hbbbd0793),
	.w5(32'h3d04edde),
	.w6(32'h3b2cdc12),
	.w7(32'hbc241a35),
	.w8(32'h3be97263),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7566d3c),
	.w1(32'h3a9769d0),
	.w2(32'h3c0760ba),
	.w3(32'hbc1635fa),
	.w4(32'hbc5a8f1c),
	.w5(32'h3b99ba79),
	.w6(32'hbacec20a),
	.w7(32'hbb8fe0a2),
	.w8(32'hbb4822d1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c128c92),
	.w1(32'hbcc36042),
	.w2(32'h3c854b8c),
	.w3(32'h3a3e1ad0),
	.w4(32'hbaca841c),
	.w5(32'h3b9a444d),
	.w6(32'h3ba49843),
	.w7(32'h3bb83aa3),
	.w8(32'h3b0ccbf1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3b395),
	.w1(32'h3bf42db9),
	.w2(32'h3bb353f0),
	.w3(32'hbc5ec24b),
	.w4(32'hbc1affb1),
	.w5(32'h3bacb8ff),
	.w6(32'hbadda756),
	.w7(32'hbb62eda0),
	.w8(32'hbb8e3e03),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac22d40),
	.w1(32'h3be310fb),
	.w2(32'hbb933d9e),
	.w3(32'h3bb6676e),
	.w4(32'h3c2fe77d),
	.w5(32'hbba57418),
	.w6(32'hbceb292e),
	.w7(32'hbbeb0258),
	.w8(32'hbd8cdb03),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfde55b),
	.w1(32'hb96ecb9f),
	.w2(32'h3b8cab80),
	.w3(32'h3ba589bf),
	.w4(32'hbb008d31),
	.w5(32'h3cbafe0e),
	.w6(32'hbc1ec84e),
	.w7(32'h3b81493d),
	.w8(32'hbbe1b3d1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0d4ea),
	.w1(32'h3c36add6),
	.w2(32'hbcf2c3c8),
	.w3(32'h3b9dbef3),
	.w4(32'hbbab7c39),
	.w5(32'h3b9504cc),
	.w6(32'hbc8a0d49),
	.w7(32'hba070c3c),
	.w8(32'h3c1e975f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92e35a),
	.w1(32'hbdb167bf),
	.w2(32'h3abc896f),
	.w3(32'hbbae3aaa),
	.w4(32'hbb015d11),
	.w5(32'h3bb280b4),
	.w6(32'hbc2de8e9),
	.w7(32'hbd19cccb),
	.w8(32'h3a840d40),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3f615),
	.w1(32'h3bc073fd),
	.w2(32'hbc1a7dd4),
	.w3(32'h3c1ff41f),
	.w4(32'hbc25ec4c),
	.w5(32'hbc4adcb1),
	.w6(32'h3bae1c9f),
	.w7(32'hba0c126a),
	.w8(32'hbc69b667),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83ee26),
	.w1(32'h3d697237),
	.w2(32'h3b3969bc),
	.w3(32'h3ca6424a),
	.w4(32'h3a3deb33),
	.w5(32'h3bc25e69),
	.w6(32'hbcc5e4a4),
	.w7(32'hbaed74e1),
	.w8(32'hbc1ddbe3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f41262),
	.w1(32'hba0afd43),
	.w2(32'h39e047f5),
	.w3(32'hbbd21a4f),
	.w4(32'h3b0a7405),
	.w5(32'hbb3277d6),
	.w6(32'hbbfe184d),
	.w7(32'hba253b4f),
	.w8(32'hbb3c5d0c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca17d5),
	.w1(32'hb9f7fd07),
	.w2(32'h3b0705c1),
	.w3(32'hbbf59209),
	.w4(32'hbb192c31),
	.w5(32'h3c9bbcc7),
	.w6(32'h3b2365a7),
	.w7(32'hbc053c06),
	.w8(32'h3be38a5f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0503ad),
	.w1(32'h3a827503),
	.w2(32'h39bb6549),
	.w3(32'h381a3347),
	.w4(32'hbbcb42cd),
	.w5(32'h3b4393cb),
	.w6(32'hbacbd556),
	.w7(32'h391696ff),
	.w8(32'h3c737ce4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82ef53),
	.w1(32'hbac5b3ac),
	.w2(32'h3ab40c4b),
	.w3(32'hbb3f5b18),
	.w4(32'hbce2841a),
	.w5(32'h3b9902c7),
	.w6(32'h3bde4d98),
	.w7(32'h3bd3ec65),
	.w8(32'h3cb85b59),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba3a25),
	.w1(32'hbb71d0bb),
	.w2(32'hbd6ea7e0),
	.w3(32'h3c3e8408),
	.w4(32'h3c380827),
	.w5(32'h3a981a2b),
	.w6(32'hbc0590d2),
	.w7(32'h3b62dda2),
	.w8(32'hbb33adf2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a4a31),
	.w1(32'hbc198769),
	.w2(32'h3bd72ef3),
	.w3(32'h3b0cad51),
	.w4(32'hbb0aa9ae),
	.w5(32'h3bd80f10),
	.w6(32'h3ac86d16),
	.w7(32'h389bcbc6),
	.w8(32'hbb4a2d23),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcbc8d),
	.w1(32'h3a1350a8),
	.w2(32'hba8eeca5),
	.w3(32'hbba780b6),
	.w4(32'hbc76f854),
	.w5(32'h3a8e2c12),
	.w6(32'h3bbff80c),
	.w7(32'hbc9c7bd0),
	.w8(32'hbc7f0c0e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e8393),
	.w1(32'h3b90c35d),
	.w2(32'hbb0fc9fe),
	.w3(32'hbc871830),
	.w4(32'h3acc2df8),
	.w5(32'hbb06f24c),
	.w6(32'h3b2ac430),
	.w7(32'hbbca234c),
	.w8(32'hba6299be),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c523b14),
	.w1(32'hbabbd0a7),
	.w2(32'h3c4c395a),
	.w3(32'h3b3d5d96),
	.w4(32'hbbb07d49),
	.w5(32'h3c1c9684),
	.w6(32'h396edd78),
	.w7(32'h3d25051a),
	.w8(32'hbc31feff),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67c4a2),
	.w1(32'h3a835107),
	.w2(32'h3838fc0b),
	.w3(32'h3af46e60),
	.w4(32'hbcbd3fde),
	.w5(32'hbb67c323),
	.w6(32'hbb73c246),
	.w7(32'h3c147505),
	.w8(32'hbb209a3b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef9351),
	.w1(32'hbc13d7f0),
	.w2(32'hba478521),
	.w3(32'h3bad138d),
	.w4(32'h3b1ebaf8),
	.w5(32'h3b78327d),
	.w6(32'h3c25db06),
	.w7(32'h3c5a1ab0),
	.w8(32'h3c80a956),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c1c23),
	.w1(32'h3b829284),
	.w2(32'h3b84ecae),
	.w3(32'h3b0064ea),
	.w4(32'hba9cfbd6),
	.w5(32'h3a62f45c),
	.w6(32'h3be6ea16),
	.w7(32'h3b19b8a1),
	.w8(32'h3b8eedca),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7011dc),
	.w1(32'h3bcd1ebd),
	.w2(32'hbbddd67e),
	.w3(32'hbbad9718),
	.w4(32'hbbd54a2c),
	.w5(32'hbb842e1a),
	.w6(32'h3c32860a),
	.w7(32'h3b987efe),
	.w8(32'hbc1265d6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852450),
	.w1(32'h3ba78778),
	.w2(32'h3c5f556e),
	.w3(32'h3c03a5c6),
	.w4(32'h3c31ac52),
	.w5(32'hbb72d038),
	.w6(32'hbbde8338),
	.w7(32'hbb18bf41),
	.w8(32'hbbd8e361),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f5a4e),
	.w1(32'hbbcc50a0),
	.w2(32'h3ab0bb24),
	.w3(32'hba9ca382),
	.w4(32'hbbd4b0e1),
	.w5(32'h3b849e28),
	.w6(32'hbbd9e61c),
	.w7(32'hbc8274e4),
	.w8(32'h3c13cbf5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcea29c),
	.w1(32'h3d16b99e),
	.w2(32'h3b9bca12),
	.w3(32'h3bdb1cb7),
	.w4(32'h3be6bbe6),
	.w5(32'hbb0fc7d4),
	.w6(32'h3bfe91a2),
	.w7(32'h3be34c6d),
	.w8(32'h3ba2f64b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51d835),
	.w1(32'h3bcc5bca),
	.w2(32'hb79f4302),
	.w3(32'hbb505a53),
	.w4(32'hbb5eccf6),
	.w5(32'h3c72597c),
	.w6(32'hbb89ba98),
	.w7(32'h3cdb6884),
	.w8(32'hbb8d6fba),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1104c6),
	.w1(32'h3b9c1ca6),
	.w2(32'h3b5840b1),
	.w3(32'hba4280ae),
	.w4(32'hbc1094d3),
	.w5(32'h3c8562b7),
	.w6(32'hbbe66cea),
	.w7(32'hbc3afbe2),
	.w8(32'h3addfb8e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04e1e7),
	.w1(32'h39ce16f4),
	.w2(32'hbba58faf),
	.w3(32'hbc2fcdf3),
	.w4(32'hbcf4a78e),
	.w5(32'hbb4bfe79),
	.w6(32'hbb6ef2a7),
	.w7(32'h3bc68637),
	.w8(32'h3a9b8d27),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe65d2),
	.w1(32'h3c067fc6),
	.w2(32'hbba23163),
	.w3(32'h3bad1a14),
	.w4(32'h3b8c93da),
	.w5(32'h3ae650ff),
	.w6(32'hbceb578d),
	.w7(32'h3ad91e8e),
	.w8(32'hb91d3fa3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b348),
	.w1(32'hbb4cfa42),
	.w2(32'hbabd4b07),
	.w3(32'h389a5474),
	.w4(32'h3c8ae0ec),
	.w5(32'h3d069eef),
	.w6(32'h3bf1978a),
	.w7(32'h3b33e5ee),
	.w8(32'hbb2c80de),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdbfef),
	.w1(32'hbb07f3cc),
	.w2(32'h3b9e8b64),
	.w3(32'hbb84e677),
	.w4(32'hbbe236a4),
	.w5(32'hbba144ae),
	.w6(32'hbc2551c7),
	.w7(32'hbc1daefc),
	.w8(32'hbc0cba30),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac638d5),
	.w1(32'h3d0994c7),
	.w2(32'hbcd31370),
	.w3(32'hbb0406df),
	.w4(32'h3c59342a),
	.w5(32'hbb50a98c),
	.w6(32'hbb0bc77f),
	.w7(32'hbacdcbe2),
	.w8(32'h3b37b73e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd7dfb),
	.w1(32'hbd3eb4c5),
	.w2(32'hbb25fbfc),
	.w3(32'hbb8b44bb),
	.w4(32'h3bc9a1b6),
	.w5(32'h3bb7f9fb),
	.w6(32'hbaa58ae1),
	.w7(32'h3a9c0d26),
	.w8(32'h3c160dc4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30e326),
	.w1(32'h3a56cc95),
	.w2(32'h3b474ada),
	.w3(32'hbbf851c7),
	.w4(32'h3bac32be),
	.w5(32'hbc4d8a0d),
	.w6(32'h3c0521cf),
	.w7(32'hbaf30efd),
	.w8(32'h3a4559a6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb812b8e1),
	.w1(32'hbbffa138),
	.w2(32'h3b2e32bd),
	.w3(32'hbd2a16c2),
	.w4(32'h3bffbdb3),
	.w5(32'hbcfb9243),
	.w6(32'hbb89ebd3),
	.w7(32'hbae31669),
	.w8(32'hba506de7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd067e5b),
	.w1(32'hbc1ae40a),
	.w2(32'h3b82a3d7),
	.w3(32'hba7a72ad),
	.w4(32'hbad7d730),
	.w5(32'h3b51cdfc),
	.w6(32'h3ba1f132),
	.w7(32'h3ba5ce1b),
	.w8(32'h3b77cdd9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5627e3),
	.w1(32'hbd2626f7),
	.w2(32'hbc9ef8c6),
	.w3(32'hbad458e7),
	.w4(32'hbbda03a1),
	.w5(32'h3d96b57e),
	.w6(32'hbb8f091c),
	.w7(32'hbc7f8b3c),
	.w8(32'h39162471),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45ce2f),
	.w1(32'h3c17c2ae),
	.w2(32'h3bff8e76),
	.w3(32'hbc1e792c),
	.w4(32'h3b902cbd),
	.w5(32'h3b7f53a3),
	.w6(32'hbc44b6b8),
	.w7(32'hbb91ee23),
	.w8(32'h3b66190c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba02848),
	.w1(32'hbba31851),
	.w2(32'h3a958db0),
	.w3(32'h3c17f61c),
	.w4(32'h3c7e476f),
	.w5(32'hba0c9151),
	.w6(32'h3b83d4ff),
	.w7(32'h3bd17897),
	.w8(32'h3a0ea57d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c2304),
	.w1(32'h3a889423),
	.w2(32'h39b0b540),
	.w3(32'h3a91d34b),
	.w4(32'h3b3ab827),
	.w5(32'h3b0aedb1),
	.w6(32'hbd32a7a7),
	.w7(32'h3bd31a50),
	.w8(32'hbad193f1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7abc20),
	.w1(32'hbb38fea8),
	.w2(32'h3b86327c),
	.w3(32'hbc1435ec),
	.w4(32'h3bc35b06),
	.w5(32'h36c2213a),
	.w6(32'hbb521eb7),
	.w7(32'hbc130533),
	.w8(32'hbd4436fd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95192f9),
	.w1(32'h3c6a58c5),
	.w2(32'h3ba8ec4c),
	.w3(32'hbb88b554),
	.w4(32'h3abcca38),
	.w5(32'h3afd4d04),
	.w6(32'h3ac0fa93),
	.w7(32'hbb9afb55),
	.w8(32'hbb85430b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16df9c),
	.w1(32'hbcb6158e),
	.w2(32'hbc085d43),
	.w3(32'h3bc266a8),
	.w4(32'hbc331509),
	.w5(32'h3d250eee),
	.w6(32'hbb1b2308),
	.w7(32'hbc3483cb),
	.w8(32'h3b458002),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe7bd2),
	.w1(32'hbadc4d4d),
	.w2(32'hbc06e97a),
	.w3(32'h3bc17bad),
	.w4(32'hbbda4258),
	.w5(32'hbbcbf807),
	.w6(32'hbc08de5d),
	.w7(32'h3a8de04e),
	.w8(32'hbb88d47e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1c215),
	.w1(32'hbb8f581a),
	.w2(32'hbc0aa5cf),
	.w3(32'h3b31208e),
	.w4(32'hb97e8ca5),
	.w5(32'h3a9e5f89),
	.w6(32'hbb93651c),
	.w7(32'hbbde3df2),
	.w8(32'h3b443b15),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae42011),
	.w1(32'hb998b523),
	.w2(32'hb898ae86),
	.w3(32'h39e8358d),
	.w4(32'hba743c82),
	.w5(32'h3b8e3958),
	.w6(32'h3b4ed8c6),
	.w7(32'h3b4d282d),
	.w8(32'h3c11361f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39191f),
	.w1(32'h3c387ea6),
	.w2(32'h3bd670b0),
	.w3(32'h3bb81e4f),
	.w4(32'h3b66ba61),
	.w5(32'h3b2b0263),
	.w6(32'hbce7a348),
	.w7(32'hba8e76a5),
	.w8(32'h3c49c8e4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9cce),
	.w1(32'hbc0f8953),
	.w2(32'hbc210061),
	.w3(32'hbada671a),
	.w4(32'h3ae304f6),
	.w5(32'hbc0f5a37),
	.w6(32'hbb704f33),
	.w7(32'hbb952e48),
	.w8(32'h3bf67b40),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7382fb),
	.w1(32'h3ae242d4),
	.w2(32'hbae1e090),
	.w3(32'h3bf8f10b),
	.w4(32'h398f83ee),
	.w5(32'h3a76061a),
	.w6(32'h3c439dac),
	.w7(32'hbc3e3435),
	.w8(32'hb920b8bb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfde81),
	.w1(32'h3a7d5a00),
	.w2(32'h3bae4e70),
	.w3(32'h3a82ab52),
	.w4(32'h3b14baa8),
	.w5(32'hbbb835e3),
	.w6(32'hbb0400bf),
	.w7(32'h3bb61809),
	.w8(32'h3b9a142f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d389d),
	.w1(32'hbc43f031),
	.w2(32'hbbe9c384),
	.w3(32'hbb055356),
	.w4(32'h3c841e70),
	.w5(32'hbb611765),
	.w6(32'h3c021b69),
	.w7(32'hbbe6b3be),
	.w8(32'hbc45930d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc842bda),
	.w1(32'hbbde4380),
	.w2(32'h3a87a1b6),
	.w3(32'hbbbbf5e7),
	.w4(32'h3bd75287),
	.w5(32'hbbe615f0),
	.w6(32'h3b9c59e2),
	.w7(32'hbc076d34),
	.w8(32'h3c9723bf),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d9706),
	.w1(32'hbbe2af5d),
	.w2(32'hbb66ddbe),
	.w3(32'hbbef4514),
	.w4(32'h3b28322f),
	.w5(32'hbb4fead8),
	.w6(32'h3bbedfa4),
	.w7(32'hbcdbec2f),
	.w8(32'h3b8285a7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3808bd),
	.w1(32'hbca45591),
	.w2(32'hbba4e5ad),
	.w3(32'h3cb2d45e),
	.w4(32'h3c099e80),
	.w5(32'h3b90e620),
	.w6(32'h3c8d27b5),
	.w7(32'hbb9d8a47),
	.w8(32'hbade184a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85560e),
	.w1(32'hbc4e7de3),
	.w2(32'hba2211cd),
	.w3(32'hbbf55843),
	.w4(32'hba84a891),
	.w5(32'hbbc3fe6d),
	.w6(32'h3c6c38ef),
	.w7(32'hbba1851d),
	.w8(32'h3cb36d4d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba93eab),
	.w1(32'hbb9c870e),
	.w2(32'h3ca8730f),
	.w3(32'h3c6c905b),
	.w4(32'h3b2cc553),
	.w5(32'h3bdd3bb3),
	.w6(32'h3c6f2f9e),
	.w7(32'h3c405f1a),
	.w8(32'h3c94d4a7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09b929),
	.w1(32'h3b54cece),
	.w2(32'hbc04c4f1),
	.w3(32'h3b88e910),
	.w4(32'hbbbfa166),
	.w5(32'hbc2c1fe9),
	.w6(32'h3a55d66a),
	.w7(32'hb8946a81),
	.w8(32'hbc5c8421),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1d195f),
	.w1(32'h3c50d238),
	.w2(32'hbb176e19),
	.w3(32'hbc26db5a),
	.w4(32'hbbd7bd25),
	.w5(32'h3c5c1549),
	.w6(32'h3ba63d96),
	.w7(32'hbcf040a1),
	.w8(32'h3c1a445e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b652944),
	.w1(32'hbba51d35),
	.w2(32'h3c81bc5d),
	.w3(32'hbc9c4159),
	.w4(32'hbcbd86dd),
	.w5(32'h3c8864af),
	.w6(32'hbbbb012c),
	.w7(32'h3c8ecbf3),
	.w8(32'hbbe48221),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda9605),
	.w1(32'hbcade048),
	.w2(32'h3c223774),
	.w3(32'h3a06de47),
	.w4(32'h3d0afc40),
	.w5(32'h3bbecf74),
	.w6(32'hba9a70b3),
	.w7(32'hbc12daef),
	.w8(32'h3c02991e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90dbab),
	.w1(32'hbbecfda0),
	.w2(32'hbbad3df0),
	.w3(32'h3cec4c6d),
	.w4(32'h3d2dbd49),
	.w5(32'hbb789652),
	.w6(32'h3c07feb3),
	.w7(32'h3be17446),
	.w8(32'hbb07e865),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4a002),
	.w1(32'hbc0f963e),
	.w2(32'h3ca7cfb8),
	.w3(32'h3c021c5e),
	.w4(32'h3c6e83dd),
	.w5(32'h3c075bfb),
	.w6(32'h3babed16),
	.w7(32'hbc79b908),
	.w8(32'h3b9ef7a5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87d9ce),
	.w1(32'hbae5cfe3),
	.w2(32'h3b70cd78),
	.w3(32'h3c1374c5),
	.w4(32'h39adca9c),
	.w5(32'h39191a30),
	.w6(32'h3cbe131a),
	.w7(32'hbbac786a),
	.w8(32'hbbe1adb5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966ca4),
	.w1(32'h3a7182aa),
	.w2(32'hbcc2e215),
	.w3(32'h3ac6589c),
	.w4(32'hbc59e4f3),
	.w5(32'h3b10bf98),
	.w6(32'h3c6f00bf),
	.w7(32'hbc071a3a),
	.w8(32'h3c302dac),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd304a21),
	.w1(32'h3c411c9b),
	.w2(32'h3c778601),
	.w3(32'hbba4807f),
	.w4(32'h3a0ac4aa),
	.w5(32'h3bbf0338),
	.w6(32'h3b99c9f1),
	.w7(32'h3ccd472a),
	.w8(32'h3bbc6f2a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf63d14),
	.w1(32'h3b7648b9),
	.w2(32'hbbd36d76),
	.w3(32'hbc78e956),
	.w4(32'h3b326166),
	.w5(32'h3bb75402),
	.w6(32'h3a8620aa),
	.w7(32'h3c2b12c6),
	.w8(32'hb7877d7e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6da9fa),
	.w1(32'h3c428e18),
	.w2(32'h3bb15c31),
	.w3(32'hb97d3192),
	.w4(32'hbc8460b8),
	.w5(32'hbc1afecc),
	.w6(32'hbc401d4a),
	.w7(32'h3cced414),
	.w8(32'h3c31dc48),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30b910),
	.w1(32'hbb00c080),
	.w2(32'hbba7d885),
	.w3(32'hbc40508a),
	.w4(32'hba3502d2),
	.w5(32'hbac1db66),
	.w6(32'h3bbf6e64),
	.w7(32'hbabaae74),
	.w8(32'h3c2e6d48),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a1288),
	.w1(32'h3ac49270),
	.w2(32'h3c1f2c6b),
	.w3(32'h3bc949c8),
	.w4(32'h3c13d303),
	.w5(32'hbc48776f),
	.w6(32'h3a77aad0),
	.w7(32'h3c1f887b),
	.w8(32'hbc5728ad),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda8216),
	.w1(32'h39659a4a),
	.w2(32'hbbf47612),
	.w3(32'h3c970af1),
	.w4(32'h3c423a4d),
	.w5(32'h3c373a23),
	.w6(32'h3b3703bc),
	.w7(32'hbb40d518),
	.w8(32'hbcb1f34f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9dab86),
	.w1(32'h3a259625),
	.w2(32'hbc25d341),
	.w3(32'hbb3cb6fc),
	.w4(32'hbc9b757c),
	.w5(32'h3bd0943c),
	.w6(32'h3b7e3787),
	.w7(32'hbbc2d331),
	.w8(32'h3c90709f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b34d9),
	.w1(32'h3b5459e8),
	.w2(32'h3c0d2b17),
	.w3(32'h3c3346e9),
	.w4(32'hbb6554a8),
	.w5(32'hbac0f4bc),
	.w6(32'hbc687a1f),
	.w7(32'h3bbe0e07),
	.w8(32'h3c2816eb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf6ecb5),
	.w1(32'h3b0ef013),
	.w2(32'h3c10d422),
	.w3(32'h3a166017),
	.w4(32'h3a05a1d8),
	.w5(32'h3bcdcfb6),
	.w6(32'h3c008291),
	.w7(32'hbc82c66e),
	.w8(32'hba73a3e8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1e2f2),
	.w1(32'h3a6e7b6a),
	.w2(32'h3c116481),
	.w3(32'hbbb51e1a),
	.w4(32'hb994925c),
	.w5(32'hbbcbff3d),
	.w6(32'h3ba353d5),
	.w7(32'hbc9aa9fb),
	.w8(32'h3b8c3128),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8afc87),
	.w1(32'h3c42a690),
	.w2(32'h3c98fbf4),
	.w3(32'h3b0397be),
	.w4(32'hbbce9c4b),
	.w5(32'h3bb5bb1c),
	.w6(32'hba0ad155),
	.w7(32'hbd8d53c7),
	.w8(32'hbb94ec88),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93593c),
	.w1(32'h3c00418a),
	.w2(32'hbc01f625),
	.w3(32'h3c872e5d),
	.w4(32'h3b4dd510),
	.w5(32'h3c550c48),
	.w6(32'h3b9008c6),
	.w7(32'hbc068d84),
	.w8(32'h3b1bfb47),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5d833),
	.w1(32'hbc242008),
	.w2(32'h3c1875af),
	.w3(32'h3bfb46c9),
	.w4(32'h3ad798ec),
	.w5(32'h3cc1ff8e),
	.w6(32'h3c4d44a9),
	.w7(32'h3bf730b0),
	.w8(32'h3c4bd702),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8d36b),
	.w1(32'hba12ab5b),
	.w2(32'hbbe8d2a3),
	.w3(32'h3bd4adad),
	.w4(32'hbc94821d),
	.w5(32'h3ccf3499),
	.w6(32'h3c7c51e3),
	.w7(32'hbb94fa78),
	.w8(32'hbc652f37),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4dc2d7),
	.w1(32'hbadd163e),
	.w2(32'h3c06100a),
	.w3(32'hbac5d0cf),
	.w4(32'h3a153889),
	.w5(32'h3b36236f),
	.w6(32'h3b5b8066),
	.w7(32'h39d0ce36),
	.w8(32'hbbdf2d23),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87cbef),
	.w1(32'hbcd09811),
	.w2(32'hb99cb208),
	.w3(32'h3d759164),
	.w4(32'h3c0d6c6d),
	.w5(32'h3b028a91),
	.w6(32'hbc4bdea8),
	.w7(32'hbb052ecd),
	.w8(32'h3bd1d6af),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc18f78),
	.w1(32'h3c83b850),
	.w2(32'hbc36cf1e),
	.w3(32'h3b86adc8),
	.w4(32'h3ce01bae),
	.w5(32'hbc04f32e),
	.w6(32'hbba987f5),
	.w7(32'hbbeeece9),
	.w8(32'h3b6a8884),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbbc47),
	.w1(32'h39fe5db4),
	.w2(32'hba58debf),
	.w3(32'h3b77a8a4),
	.w4(32'hbb99f095),
	.w5(32'h3bf56d16),
	.w6(32'hbc21e94a),
	.w7(32'hbb1bdd67),
	.w8(32'h3b428bd7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8103d4),
	.w1(32'h3cb8f92f),
	.w2(32'hbcc10500),
	.w3(32'hbba00c73),
	.w4(32'h3bccfe73),
	.w5(32'hbc458fe0),
	.w6(32'h39494a9f),
	.w7(32'h391681af),
	.w8(32'h3c230137),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20985c),
	.w1(32'hbc7e4f28),
	.w2(32'hbb5ae000),
	.w3(32'h3a87affe),
	.w4(32'hbacb4eb2),
	.w5(32'hbc08da78),
	.w6(32'hbc195ee8),
	.w7(32'hbc43cdce),
	.w8(32'hbbf171eb),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f8663),
	.w1(32'h3c18e397),
	.w2(32'h3bd85543),
	.w3(32'hbb662fbf),
	.w4(32'hbb746355),
	.w5(32'hbc6d9f35),
	.w6(32'h3b7fb7d0),
	.w7(32'h3a2288e7),
	.w8(32'hbc0cc0f8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa460b5),
	.w1(32'hbbb6e4cc),
	.w2(32'h3b22ef22),
	.w3(32'hbbb709e1),
	.w4(32'hbb0f056f),
	.w5(32'hbbbffbeb),
	.w6(32'hbb240ed4),
	.w7(32'h3d375aa4),
	.w8(32'h3c19de34),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b1ed),
	.w1(32'h3a6f8471),
	.w2(32'hbb3d6c34),
	.w3(32'hbba5ca9b),
	.w4(32'h3a4bdc80),
	.w5(32'h3b3abc84),
	.w6(32'h3c27cd7a),
	.w7(32'h3be65e20),
	.w8(32'hbb999b54),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c639348),
	.w1(32'h3ba6e5f0),
	.w2(32'h3b9d4258),
	.w3(32'hbbb6546a),
	.w4(32'h3ba03dc3),
	.w5(32'hbb5a4211),
	.w6(32'hbc88c9f5),
	.w7(32'hbbe6b357),
	.w8(32'hba888154),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b890a8a),
	.w1(32'hbc687137),
	.w2(32'hba920e76),
	.w3(32'hbbd289fb),
	.w4(32'h3c31d616),
	.w5(32'hbb33bcae),
	.w6(32'h3c5e562b),
	.w7(32'h3bb50fc7),
	.w8(32'h3b25846e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc495f76),
	.w1(32'h3a3f25e6),
	.w2(32'h3c5a1172),
	.w3(32'hba6d3bcf),
	.w4(32'h3b3bf7aa),
	.w5(32'hbc7742c9),
	.w6(32'hbbaf9abb),
	.w7(32'hbb4d5a3e),
	.w8(32'h3a73a4cd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc359e01),
	.w1(32'h3c02a159),
	.w2(32'hbbacd051),
	.w3(32'h3b21cc43),
	.w4(32'hbc66fc6e),
	.w5(32'hbb2067c8),
	.w6(32'hbc3cd4c8),
	.w7(32'hbc8c14f7),
	.w8(32'hbbedda1c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c02b9),
	.w1(32'hbaf6a342),
	.w2(32'hbc492a37),
	.w3(32'hbb5dab47),
	.w4(32'hbb6202f9),
	.w5(32'hba3a0019),
	.w6(32'hbab1f40e),
	.w7(32'hbb1cc4e9),
	.w8(32'h3b8d55fa),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa863d0),
	.w1(32'h3bed4b1c),
	.w2(32'hbbb60f5f),
	.w3(32'hbc6a0172),
	.w4(32'hbb8b9738),
	.w5(32'hbc8ac3c4),
	.w6(32'hba04557f),
	.w7(32'h3b62706d),
	.w8(32'hbadda2d7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2866a2),
	.w1(32'h3b705525),
	.w2(32'h3af7ff16),
	.w3(32'h3a907a88),
	.w4(32'hbc16626c),
	.w5(32'hbc005404),
	.w6(32'h3cb18a48),
	.w7(32'hb9d98cc2),
	.w8(32'hbc07ef74),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a365b),
	.w1(32'hbbe1a5f2),
	.w2(32'h3bf363f3),
	.w3(32'hbb8916d6),
	.w4(32'hbc4dc765),
	.w5(32'h3c2ae37d),
	.w6(32'h3bec450c),
	.w7(32'hbba1e95e),
	.w8(32'hbb35f6a0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97c237),
	.w1(32'h3bc43590),
	.w2(32'hbaacf80e),
	.w3(32'h3ba357a1),
	.w4(32'hbb392264),
	.w5(32'h3b4a2ace),
	.w6(32'h3b847662),
	.w7(32'h3b7bdf0b),
	.w8(32'hbc0a597a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d7c30),
	.w1(32'hbba6654b),
	.w2(32'h3a57e62b),
	.w3(32'h3a664bc9),
	.w4(32'hbba6908c),
	.w5(32'hb9cda0bb),
	.w6(32'hbbfc8ba9),
	.w7(32'h3bb1f5ed),
	.w8(32'h3bd44f88),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ed37),
	.w1(32'hbb9d7a69),
	.w2(32'hbbdd92b6),
	.w3(32'hbb509324),
	.w4(32'hbbf327b5),
	.w5(32'h3c1080fd),
	.w6(32'h3c2fc030),
	.w7(32'h3b65234f),
	.w8(32'hbb13962e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b3eaa),
	.w1(32'h3bf90853),
	.w2(32'hbba3c1bb),
	.w3(32'h3b21930e),
	.w4(32'h3bc17108),
	.w5(32'h3b78b867),
	.w6(32'h3aaeed88),
	.w7(32'h3bb0ed3b),
	.w8(32'hbc3b3bae),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ff771),
	.w1(32'h3c285ef2),
	.w2(32'hbbb4a0c0),
	.w3(32'h3aeeda88),
	.w4(32'h3b493f73),
	.w5(32'hb9946392),
	.w6(32'h3b99087c),
	.w7(32'h3be34735),
	.w8(32'hba4a2c83),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5ec49),
	.w1(32'h3ab1ae0f),
	.w2(32'hbc02d044),
	.w3(32'h3b62295d),
	.w4(32'h3bd9ffda),
	.w5(32'hb9fc9a10),
	.w6(32'hbb626699),
	.w7(32'h3c8f65d2),
	.w8(32'hbb984de9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03eac0),
	.w1(32'h3b74acba),
	.w2(32'h3a1eb0d7),
	.w3(32'h3cc6a1ac),
	.w4(32'h3a87e35b),
	.w5(32'h3b07a18f),
	.w6(32'hbbf35a7b),
	.w7(32'hbc122498),
	.w8(32'hbb162f5d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fd5cb),
	.w1(32'hbb97fd50),
	.w2(32'h3c562ea1),
	.w3(32'hbbf7bd70),
	.w4(32'h3acbfff1),
	.w5(32'h3b91bced),
	.w6(32'hbb1848af),
	.w7(32'hb88d480a),
	.w8(32'h398db4b5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab7f0d),
	.w1(32'hba1cabd3),
	.w2(32'hbb977838),
	.w3(32'hbb50341a),
	.w4(32'hbb485875),
	.w5(32'hbc341d0e),
	.w6(32'hbca22e96),
	.w7(32'h39ce4555),
	.w8(32'hbb690e84),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bd294),
	.w1(32'h3bb085ee),
	.w2(32'h3c36aaea),
	.w3(32'hbbce5015),
	.w4(32'hbbd71fa2),
	.w5(32'hbbcbad57),
	.w6(32'hbb5ad0cf),
	.w7(32'h3a80ed3c),
	.w8(32'hbacf571b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe3ec0),
	.w1(32'h3bbb8571),
	.w2(32'hbbd4cc5a),
	.w3(32'h3bcc6cbf),
	.w4(32'hbbc9978e),
	.w5(32'hbc86408a),
	.w6(32'hbba019cd),
	.w7(32'hbc6e1c1c),
	.w8(32'hbc80b8ae),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1688b0),
	.w1(32'hb909088e),
	.w2(32'h3aecb7bb),
	.w3(32'hba6628ee),
	.w4(32'hbb8009c8),
	.w5(32'h3bbc4fb9),
	.w6(32'h3c65c57c),
	.w7(32'h3d3d6203),
	.w8(32'hb918f554),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53d364),
	.w1(32'hbb815f8e),
	.w2(32'hbb1fae14),
	.w3(32'h3c0975bc),
	.w4(32'hbb138f79),
	.w5(32'hbc15d842),
	.w6(32'hbc08255f),
	.w7(32'hbad79ee6),
	.w8(32'hbcc72aba),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad36e47),
	.w1(32'h3b974238),
	.w2(32'h3a4ec994),
	.w3(32'h3bec6f91),
	.w4(32'hb9dfa589),
	.w5(32'h3a7a0a8f),
	.w6(32'hbb9ad397),
	.w7(32'h3c911976),
	.w8(32'h3b88ea44),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c005e98),
	.w1(32'hbb4b6357),
	.w2(32'hbbae9bc9),
	.w3(32'hbb00f143),
	.w4(32'h3d17fc29),
	.w5(32'h3ba4da82),
	.w6(32'h3b573045),
	.w7(32'h3bf1f385),
	.w8(32'hbc6d5bd5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be06267),
	.w1(32'h3b18439b),
	.w2(32'hbb912825),
	.w3(32'hbc823849),
	.w4(32'hbb64b732),
	.w5(32'hb9bc5397),
	.w6(32'hbb7d9fc6),
	.w7(32'hbc2c9b67),
	.w8(32'h3b67141b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9e89a),
	.w1(32'hbc67fb8b),
	.w2(32'hbc90fd03),
	.w3(32'h3c3b4086),
	.w4(32'hbbb31eb3),
	.w5(32'hbbf87636),
	.w6(32'hbc245f07),
	.w7(32'hbc549929),
	.w8(32'h3b8372c4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d169e83),
	.w1(32'hbc3ed22f),
	.w2(32'h3c0ef5a2),
	.w3(32'hbcd16c89),
	.w4(32'h3b8b5d62),
	.w5(32'hbc8e0f7e),
	.w6(32'h3ab85370),
	.w7(32'h3b9b8654),
	.w8(32'h3c2350d3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4cb2a),
	.w1(32'hbb4ca878),
	.w2(32'hb93a047f),
	.w3(32'hbb15ae49),
	.w4(32'h3bb93e2b),
	.w5(32'hbb856d52),
	.w6(32'h3b2c6f68),
	.w7(32'hbac6e238),
	.w8(32'h3bef09a1),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af97e95),
	.w1(32'h3c3f57a7),
	.w2(32'h3c20b944),
	.w3(32'hbb9daabc),
	.w4(32'h3c5eb5a2),
	.w5(32'hbc6fc42b),
	.w6(32'hbc0bd3ac),
	.w7(32'hba40d934),
	.w8(32'hbc795ea9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce377),
	.w1(32'hbbde5d03),
	.w2(32'h3b979ec1),
	.w3(32'hbc033f62),
	.w4(32'hbb7b7040),
	.w5(32'hbb1ecdc6),
	.w6(32'h3b4cd735),
	.w7(32'h3bd0e5de),
	.w8(32'hbbdfd58c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a990c),
	.w1(32'hbba4211b),
	.w2(32'hb9ac9dba),
	.w3(32'hbc2a571e),
	.w4(32'hbb3f4af8),
	.w5(32'h3c6a11d6),
	.w6(32'h3bc2a440),
	.w7(32'h3cb5fe9d),
	.w8(32'hbb2372ad),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf47ec8),
	.w1(32'h3b689130),
	.w2(32'h3b8e52f8),
	.w3(32'h3c9b180f),
	.w4(32'h3b73f664),
	.w5(32'h3c4b507d),
	.w6(32'hbbfd3613),
	.w7(32'h3b1bccc0),
	.w8(32'h3c561d6a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93ecbc),
	.w1(32'hbb26b7b6),
	.w2(32'hbc475197),
	.w3(32'hbc06da69),
	.w4(32'hbb08a15a),
	.w5(32'h3caae094),
	.w6(32'hbb3d6d48),
	.w7(32'hbc9a5c16),
	.w8(32'h3be3c824),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6b823),
	.w1(32'h3affd90d),
	.w2(32'hb8c7521a),
	.w3(32'hb8b8dc4f),
	.w4(32'hbb124547),
	.w5(32'h3bf639af),
	.w6(32'h3a418dbd),
	.w7(32'hbca8d235),
	.w8(32'h3bc75226),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff3b37),
	.w1(32'hbbb153bc),
	.w2(32'hbbc77ad8),
	.w3(32'hba3e6b0d),
	.w4(32'h3a98a358),
	.w5(32'h3af93aed),
	.w6(32'hb89c0312),
	.w7(32'h3b77b100),
	.w8(32'h3c9a443e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a54aa),
	.w1(32'hbc1181ce),
	.w2(32'h3b5ba278),
	.w3(32'hbc190399),
	.w4(32'hbc649906),
	.w5(32'hbb5c3247),
	.w6(32'h3c5fa6ec),
	.w7(32'hbb1b71c8),
	.w8(32'hbb1f5d00),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb382cd),
	.w1(32'h3b8c8693),
	.w2(32'h3b68a02a),
	.w3(32'hbc0c2190),
	.w4(32'hbc38d994),
	.w5(32'hbc5b583b),
	.w6(32'hbc194ab5),
	.w7(32'h3b3ff891),
	.w8(32'hbca3f5f8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcbf94),
	.w1(32'hb81e8ce6),
	.w2(32'hbbb0d479),
	.w3(32'h3c00000f),
	.w4(32'h3be75047),
	.w5(32'h3b3007c2),
	.w6(32'hba891e66),
	.w7(32'h3acc5b8f),
	.w8(32'hbb807193),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0f00d),
	.w1(32'hbc21f70b),
	.w2(32'hbb3ed631),
	.w3(32'h3b43f328),
	.w4(32'hbac38f34),
	.w5(32'h3c01896b),
	.w6(32'h3a7ede6d),
	.w7(32'h3baadc48),
	.w8(32'h3ab1fa44),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b1a5e),
	.w1(32'hbbec5109),
	.w2(32'hbb0f65dd),
	.w3(32'hbb3f63ce),
	.w4(32'hbc2811a5),
	.w5(32'hbbe4bd3d),
	.w6(32'hbb7fd20c),
	.w7(32'hbbf6105b),
	.w8(32'h3c55f1d6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f0720),
	.w1(32'h3c4f323c),
	.w2(32'h3b1df3f9),
	.w3(32'hbca5435f),
	.w4(32'h3bd28ba1),
	.w5(32'h3c7f31ca),
	.w6(32'hbc0d464c),
	.w7(32'hbb1c509a),
	.w8(32'hbc89e90c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e89ac),
	.w1(32'hbc26b3fd),
	.w2(32'hbc4b94ac),
	.w3(32'hbc2cdceb),
	.w4(32'h3b84d7a1),
	.w5(32'hbb71e01a),
	.w6(32'hbc3fbd98),
	.w7(32'h3b518303),
	.w8(32'hbb782b77),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005172),
	.w1(32'hbc9a292e),
	.w2(32'hbb44afdc),
	.w3(32'h3b90f56e),
	.w4(32'hbb665a0f),
	.w5(32'hbc074ca3),
	.w6(32'hbb98c960),
	.w7(32'hbc12c33c),
	.w8(32'hbb394091),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd938e5),
	.w1(32'h3c7730e5),
	.w2(32'h3ba1bde7),
	.w3(32'hbbbba1ff),
	.w4(32'hbbb1bfd5),
	.w5(32'h3b486a2c),
	.w6(32'h3bf06a84),
	.w7(32'hbb936aaa),
	.w8(32'hbc120fca),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbb8d2),
	.w1(32'h3abefa4f),
	.w2(32'h3bd1b8db),
	.w3(32'h3badee74),
	.w4(32'hbb299538),
	.w5(32'hbb3913ef),
	.w6(32'h3b5cedef),
	.w7(32'h394ac512),
	.w8(32'h3a729e78),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed919),
	.w1(32'hb9b620fb),
	.w2(32'hbc1beab6),
	.w3(32'h39cf02ef),
	.w4(32'hbbdbf473),
	.w5(32'hba9cfe59),
	.w6(32'h3beb7352),
	.w7(32'h3bf3dec7),
	.w8(32'h3b0f0b7f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccc8d8),
	.w1(32'hbc9d2692),
	.w2(32'hbc330f1f),
	.w3(32'hbb641683),
	.w4(32'h3b8b83d9),
	.w5(32'h3c100b0d),
	.w6(32'h3bbd4f91),
	.w7(32'hba8f206d),
	.w8(32'hbaf5ca7e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb1b85),
	.w1(32'hb9322dc1),
	.w2(32'hbb57ba02),
	.w3(32'hbc94167d),
	.w4(32'hbb3b42cc),
	.w5(32'h3b5acc72),
	.w6(32'hbbe058db),
	.w7(32'hbcb5e776),
	.w8(32'hbae84fa7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1de4b7),
	.w1(32'h3c85833c),
	.w2(32'h3c04d909),
	.w3(32'h39e9c07e),
	.w4(32'h3bb6420f),
	.w5(32'hbc06ae00),
	.w6(32'h3ae05964),
	.w7(32'h37aa5572),
	.w8(32'h38b46cce),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ee674),
	.w1(32'h3b26e9cf),
	.w2(32'hbaf06d46),
	.w3(32'hbb905fa1),
	.w4(32'hbb7956dc),
	.w5(32'h3c453d4d),
	.w6(32'h3c10d853),
	.w7(32'h3a972f8a),
	.w8(32'hbb9116ff),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc04a95),
	.w1(32'h3c1ed360),
	.w2(32'hbb937f1b),
	.w3(32'h3a9c739c),
	.w4(32'h3b934d00),
	.w5(32'h3bb9d74a),
	.w6(32'h3d527bff),
	.w7(32'hbb523959),
	.w8(32'hb9fb11e0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08e9c8),
	.w1(32'hbc7cf6c2),
	.w2(32'hba173961),
	.w3(32'hbbd8fcc4),
	.w4(32'hbb9bdacd),
	.w5(32'h3bbd4b10),
	.w6(32'h3a0a5a66),
	.w7(32'hba833cd8),
	.w8(32'hbc791479),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc403ba9),
	.w1(32'h3bb29887),
	.w2(32'hbc16658d),
	.w3(32'hbc1e7466),
	.w4(32'hbbe01f8a),
	.w5(32'h3bad6e8e),
	.w6(32'h3a9778da),
	.w7(32'h3b8cba37),
	.w8(32'h38961dd9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41c5fc),
	.w1(32'h3909804c),
	.w2(32'hba34080a),
	.w3(32'h3bf34bfb),
	.w4(32'hbb56f9bf),
	.w5(32'hbb0d3682),
	.w6(32'hbb45560d),
	.w7(32'h3c2bb310),
	.w8(32'hbb455e5d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90790f),
	.w1(32'h3c00ec99),
	.w2(32'h3b64e672),
	.w3(32'h3c1cea20),
	.w4(32'hbd0d6f2e),
	.w5(32'h3c0c1a9e),
	.w6(32'hbbf896ef),
	.w7(32'h3c019b15),
	.w8(32'hbc0323bb),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc275b53),
	.w1(32'hbb104713),
	.w2(32'hba66b4ab),
	.w3(32'h397fa335),
	.w4(32'hbbf4fcc2),
	.w5(32'h3974b1dc),
	.w6(32'hbaab7fff),
	.w7(32'h3b20ec0e),
	.w8(32'hbb6fa25d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4bbef),
	.w1(32'hbbf45aa2),
	.w2(32'h3af216b7),
	.w3(32'h3c26fce2),
	.w4(32'h3b893793),
	.w5(32'h3a1ced3e),
	.w6(32'hbb03994d),
	.w7(32'h3b94ddbe),
	.w8(32'hbb82aafe),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b036520),
	.w1(32'h3c549ac5),
	.w2(32'hbab8634c),
	.w3(32'h3c226558),
	.w4(32'hbb0110fb),
	.w5(32'hbb8f6ebd),
	.w6(32'hbcb085e9),
	.w7(32'h3cab95e0),
	.w8(32'h3c1d913e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e80b),
	.w1(32'h3beb3820),
	.w2(32'hbbc35d07),
	.w3(32'hbc09267f),
	.w4(32'hbb136e53),
	.w5(32'h39231ebe),
	.w6(32'h3c24e7af),
	.w7(32'hbbfb4e91),
	.w8(32'hba9a4d9f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1b382),
	.w1(32'hbc0165d6),
	.w2(32'hbb0766db),
	.w3(32'hbb3049a6),
	.w4(32'hbc88c4e5),
	.w5(32'h3b94bbaf),
	.w6(32'h3b10fbce),
	.w7(32'h3b564479),
	.w8(32'h3a1d64c5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3a352),
	.w1(32'hbc95e46a),
	.w2(32'h3b80fce2),
	.w3(32'h3c35e94e),
	.w4(32'hba778e56),
	.w5(32'h3c9d6562),
	.w6(32'hbbc31eb1),
	.w7(32'h3b8c4ede),
	.w8(32'h397761af),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb842e7b),
	.w1(32'hbaaae7e9),
	.w2(32'h3af04e30),
	.w3(32'hbb331503),
	.w4(32'h3caf3a28),
	.w5(32'h3aaa4cb7),
	.w6(32'hbb1d9b49),
	.w7(32'h3c8e970f),
	.w8(32'h3c069e0c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca996a0),
	.w1(32'h39edb32a),
	.w2(32'h37fa93d4),
	.w3(32'h3af5cc18),
	.w4(32'hbad11733),
	.w5(32'hbb8df0f1),
	.w6(32'hbb7fe0ba),
	.w7(32'hbbc5999f),
	.w8(32'hbae8f399),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c205428),
	.w1(32'hbb7ea65f),
	.w2(32'hbbea236c),
	.w3(32'hbcc4444b),
	.w4(32'hbae5ca84),
	.w5(32'hbb5764f1),
	.w6(32'hbc276ec9),
	.w7(32'hba17bb8c),
	.w8(32'h3c7d3077),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99d8d5),
	.w1(32'h3c5d71ba),
	.w2(32'hb9213db7),
	.w3(32'hbc8203a9),
	.w4(32'hbb9489bd),
	.w5(32'hbc5c863e),
	.w6(32'hbbc42915),
	.w7(32'hba839f0c),
	.w8(32'h3c0b3f29),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02b37e),
	.w1(32'h3c021ab3),
	.w2(32'h3bd928ad),
	.w3(32'hbb85cdae),
	.w4(32'h3b274648),
	.w5(32'h3a37585a),
	.w6(32'h3a709918),
	.w7(32'hba76a429),
	.w8(32'hbc1ff77f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cecab),
	.w1(32'hbbda007e),
	.w2(32'hbb51fb97),
	.w3(32'hbbae551a),
	.w4(32'h391b6555),
	.w5(32'h3bfeb19d),
	.w6(32'h3b869e80),
	.w7(32'hbb2030db),
	.w8(32'hbbbcfea6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85787c),
	.w1(32'hbb021096),
	.w2(32'hbbee896e),
	.w3(32'hbbf944b2),
	.w4(32'hbca62759),
	.w5(32'hbb2053f9),
	.w6(32'h3b725058),
	.w7(32'hb9816703),
	.w8(32'h3c4c6ff7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de32c6),
	.w1(32'h3c7e197b),
	.w2(32'hbcff154f),
	.w3(32'h3bfeaca5),
	.w4(32'h3c23d864),
	.w5(32'h3cd71a9b),
	.w6(32'h3bfed474),
	.w7(32'hbbd1ca14),
	.w8(32'h3b7e54a9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba900144),
	.w1(32'hbbadb330),
	.w2(32'hbb88e399),
	.w3(32'h3a440e63),
	.w4(32'hbc5d82f1),
	.w5(32'hbbb52542),
	.w6(32'h370e7085),
	.w7(32'hbb6e3dcc),
	.w8(32'hb82d018c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f87ce),
	.w1(32'h3ba777ab),
	.w2(32'h3a0d0031),
	.w3(32'hbb428bbe),
	.w4(32'h3a0c58d4),
	.w5(32'hbb0e1dec),
	.w6(32'h3be9fccc),
	.w7(32'h3d329eff),
	.w8(32'hbbaa59d6),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb556db0),
	.w1(32'hbc07db30),
	.w2(32'hbb796d37),
	.w3(32'hbb457fdf),
	.w4(32'hbaed4b87),
	.w5(32'h3ce5e885),
	.w6(32'h3adc3373),
	.w7(32'h39d1f791),
	.w8(32'h3c6367ec),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6721d0),
	.w1(32'h3ca90097),
	.w2(32'hba6257e6),
	.w3(32'h3c235f07),
	.w4(32'hbc00f1f4),
	.w5(32'hbaf088dc),
	.w6(32'h39e68b3e),
	.w7(32'hbb72bbf9),
	.w8(32'hbc6c472c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2615ac),
	.w1(32'hbb09b92e),
	.w2(32'h3bee7965),
	.w3(32'hbb08d7a6),
	.w4(32'h3a91da41),
	.w5(32'hbc259dae),
	.w6(32'h3b01e816),
	.w7(32'hbbe7a48c),
	.w8(32'hbbadb1b4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc313f71),
	.w1(32'h3a95a2cf),
	.w2(32'h3ba604e4),
	.w3(32'h3cb3877f),
	.w4(32'hbbba29bd),
	.w5(32'h3bdd2038),
	.w6(32'h3ae46b8c),
	.w7(32'h3c3421a2),
	.w8(32'hb91a104b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2ef85),
	.w1(32'hba83f026),
	.w2(32'h39488dc1),
	.w3(32'h3a72dcd3),
	.w4(32'hbc589b6f),
	.w5(32'h39f53eb2),
	.w6(32'hb76579e2),
	.w7(32'hbaa76860),
	.w8(32'h3a606ccd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf17f25),
	.w1(32'h3c0f6f50),
	.w2(32'h3adc8ca6),
	.w3(32'h3c0a7559),
	.w4(32'h3bcc2050),
	.w5(32'h3a28a651),
	.w6(32'h3c63e371),
	.w7(32'hbae7f4db),
	.w8(32'hbb995ae3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dc781),
	.w1(32'hbb41674d),
	.w2(32'h3ac34a0f),
	.w3(32'hbbe802af),
	.w4(32'h3b4baafb),
	.w5(32'h3aebd1be),
	.w6(32'h3b251459),
	.w7(32'h3bd63b57),
	.w8(32'hbb65a804),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c6086),
	.w1(32'hbba67780),
	.w2(32'h3c2b9777),
	.w3(32'hbbfe88df),
	.w4(32'hbb59af3f),
	.w5(32'hbb80ad47),
	.w6(32'h3ad97156),
	.w7(32'hbc5ac3a1),
	.w8(32'hbdc22ff7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6f3ce),
	.w1(32'hba38fe41),
	.w2(32'hbbb4489d),
	.w3(32'hbb30aa8f),
	.w4(32'h3b71c949),
	.w5(32'h3d538a13),
	.w6(32'hbb44b4c3),
	.w7(32'hbcc48de0),
	.w8(32'h380e86dc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b4d2b),
	.w1(32'h3c42be7b),
	.w2(32'hbadf7024),
	.w3(32'hbacf1720),
	.w4(32'h3ba9e9a7),
	.w5(32'hbb84e9c8),
	.w6(32'hb8822ae6),
	.w7(32'h3de28581),
	.w8(32'hbb831d03),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04c311),
	.w1(32'hba82d6fa),
	.w2(32'hbac45b09),
	.w3(32'hbb519c09),
	.w4(32'hbb058ebd),
	.w5(32'hbc350c27),
	.w6(32'hbd97eeed),
	.w7(32'h3c0b0f0e),
	.w8(32'h3afd05bb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e11c4),
	.w1(32'hbb58c476),
	.w2(32'hbd04078f),
	.w3(32'hbb6518bf),
	.w4(32'h3b9986d4),
	.w5(32'hbb485b39),
	.w6(32'hbc132138),
	.w7(32'h3b606756),
	.w8(32'h3cb986dd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88f8ed),
	.w1(32'hbb953848),
	.w2(32'hbab2c7c6),
	.w3(32'hbb2bd5a7),
	.w4(32'hbbcce6bb),
	.w5(32'h3b14066a),
	.w6(32'hb9a10023),
	.w7(32'h3bac75bb),
	.w8(32'h3b093c84),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdf969),
	.w1(32'h3adaa353),
	.w2(32'hbb15e8f5),
	.w3(32'h39ee3291),
	.w4(32'hbce9dd7c),
	.w5(32'hbb8a71d7),
	.w6(32'hb8073737),
	.w7(32'h3bc9381c),
	.w8(32'h3cb17056),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bd730),
	.w1(32'h3b9e1676),
	.w2(32'hbc2efd4b),
	.w3(32'h3c59df28),
	.w4(32'hbb0f3118),
	.w5(32'hbb554489),
	.w6(32'hbac4aab9),
	.w7(32'h3c08e54f),
	.w8(32'h3b0ab02d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e26d4),
	.w1(32'hbb7d8c86),
	.w2(32'hbb09300b),
	.w3(32'hbc3d58ea),
	.w4(32'h3cc133a8),
	.w5(32'hbc1976f9),
	.w6(32'hbbeeb33b),
	.w7(32'h3b418c5f),
	.w8(32'h3c6d82c6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987cf60),
	.w1(32'h3b80967c),
	.w2(32'h3b82f7f4),
	.w3(32'hbc06bda6),
	.w4(32'hbb39a1f0),
	.w5(32'h3a87a0aa),
	.w6(32'h3b821e17),
	.w7(32'h3acb561e),
	.w8(32'hbd702c93),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0529),
	.w1(32'h3a20d95b),
	.w2(32'hbaac3a44),
	.w3(32'h3a89769b),
	.w4(32'hbb36ee01),
	.w5(32'h3b8d3cef),
	.w6(32'hbb81ac73),
	.w7(32'h3c1df8fc),
	.w8(32'hbb038226),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16a6dc),
	.w1(32'hbb956c2d),
	.w2(32'hbc3cf040),
	.w3(32'h3c571195),
	.w4(32'h3b8d707e),
	.w5(32'hb8bd8fc2),
	.w6(32'hbae8b700),
	.w7(32'h3bc27cdd),
	.w8(32'hbc1d8a6a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e6fd0),
	.w1(32'hbc2cf820),
	.w2(32'hbbce3036),
	.w3(32'hbb2cd009),
	.w4(32'hba557db3),
	.w5(32'hbb10319f),
	.w6(32'hbb582252),
	.w7(32'h3beed95e),
	.w8(32'h3a031c8d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c7b11),
	.w1(32'hba3d5581),
	.w2(32'hbbcd3dd3),
	.w3(32'hbaede718),
	.w4(32'h3b9af0e7),
	.w5(32'h3c933c76),
	.w6(32'hbb39d2d6),
	.w7(32'hbb5c1f52),
	.w8(32'h3b233d29),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803f19),
	.w1(32'hb9e67d6e),
	.w2(32'hbbd8e100),
	.w3(32'hbbb95cfb),
	.w4(32'hbc3a4962),
	.w5(32'h3c798fec),
	.w6(32'hbc02f996),
	.w7(32'hbdede318),
	.w8(32'hbbaba4e8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b761a),
	.w1(32'h3c264905),
	.w2(32'h3b59ad8f),
	.w3(32'hbc679ec5),
	.w4(32'hbc5564b2),
	.w5(32'h3b08972c),
	.w6(32'hb997c888),
	.w7(32'hbc7d4fff),
	.w8(32'h3ae8f3b8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcbb16),
	.w1(32'hba75aefe),
	.w2(32'h3c909a8a),
	.w3(32'hbb71ee36),
	.w4(32'hbbc6a625),
	.w5(32'h3a14e95d),
	.w6(32'h3bdf3803),
	.w7(32'h37b9c11d),
	.w8(32'h3b7b5dac),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b02e6),
	.w1(32'hbb0557fb),
	.w2(32'hbc18ac2d),
	.w3(32'hbbe7f438),
	.w4(32'h3c454ca5),
	.w5(32'hbba9ca3f),
	.w6(32'h3b8876f5),
	.w7(32'hbb6c36dd),
	.w8(32'hbb9932a0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad99161),
	.w1(32'hb9547f71),
	.w2(32'hbaacf23e),
	.w3(32'h3b954001),
	.w4(32'hba3fdc5f),
	.w5(32'h3c1623d9),
	.w6(32'hbbb50a40),
	.w7(32'h3b4552d5),
	.w8(32'hbd23d777),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b71dc),
	.w1(32'hbb13c5af),
	.w2(32'hbb77cd34),
	.w3(32'hb9ecf186),
	.w4(32'hbb66a10a),
	.w5(32'hbb941136),
	.w6(32'h3c8a9042),
	.w7(32'h3c9563b2),
	.w8(32'hbc084525),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1498ea),
	.w1(32'hbd19a35c),
	.w2(32'h3acd9e3d),
	.w3(32'h3b6f6373),
	.w4(32'hbb6801d9),
	.w5(32'hbbe44bf1),
	.w6(32'hbb6c8489),
	.w7(32'hbcee4234),
	.w8(32'hbbe0e912),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f4b2a),
	.w1(32'hbb06f58a),
	.w2(32'hbb4290e8),
	.w3(32'hbc17475b),
	.w4(32'h3c076b32),
	.w5(32'hbbb008ca),
	.w6(32'hbc49c18c),
	.w7(32'hbae7cb43),
	.w8(32'h3ad5e5fb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4606e),
	.w1(32'h3bd69114),
	.w2(32'hbb97f393),
	.w3(32'hbc46455a),
	.w4(32'h3c4e8e74),
	.w5(32'h3b57d4f8),
	.w6(32'hbb7671db),
	.w7(32'hbbfaca47),
	.w8(32'hbc581390),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdbcb3),
	.w1(32'hbc070257),
	.w2(32'h3a289950),
	.w3(32'h3bd0fe84),
	.w4(32'hbb8d847a),
	.w5(32'h3b6eef68),
	.w6(32'h3a142871),
	.w7(32'hbabdc70f),
	.w8(32'h3af382e9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc2d28),
	.w1(32'h3c91cb79),
	.w2(32'h3aab3ff0),
	.w3(32'hba16521e),
	.w4(32'h3bbc3318),
	.w5(32'h3beb188f),
	.w6(32'h3d54c4e9),
	.w7(32'hbcf0dd95),
	.w8(32'hba0f496c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cfe33),
	.w1(32'hbbf93434),
	.w2(32'h3ba266b6),
	.w3(32'hbccee5e5),
	.w4(32'hbb16cf81),
	.w5(32'hbb7e5b6f),
	.w6(32'hba4f983f),
	.w7(32'hbc25f751),
	.w8(32'hbb7535fc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb11fe6),
	.w1(32'h3bb26fb3),
	.w2(32'hbca712f4),
	.w3(32'h3a38cf54),
	.w4(32'h3c2e54d7),
	.w5(32'hbc0426c5),
	.w6(32'h3c0a0c56),
	.w7(32'h3ba1621a),
	.w8(32'h38d545b0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e209c),
	.w1(32'hbad06d14),
	.w2(32'hbbeeb737),
	.w3(32'h3ba160cd),
	.w4(32'hbbb49452),
	.w5(32'h3baf5c20),
	.w6(32'h3c2da0f0),
	.w7(32'hbb533a1f),
	.w8(32'h3be28837),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab67835),
	.w1(32'hba92dff3),
	.w2(32'hbb93d1db),
	.w3(32'h3aa84575),
	.w4(32'h3a8777f2),
	.w5(32'h3b8aff0c),
	.w6(32'hbb996aab),
	.w7(32'hbbc3ee1b),
	.w8(32'hbb23e073),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c272796),
	.w1(32'h3cb3582b),
	.w2(32'hbc984a66),
	.w3(32'hbc3016de),
	.w4(32'h3a0d3b38),
	.w5(32'hbc8d60a6),
	.w6(32'hbc7f552f),
	.w7(32'hbad330cd),
	.w8(32'hbc379970),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule