module layer_10_featuremap_503(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fdc59c),
	.w1(32'hb6efdf3d),
	.w2(32'h349bb6c9),
	.w3(32'hb81299dd),
	.w4(32'hb72032f2),
	.w5(32'h36243a5b),
	.w6(32'hb832e044),
	.w7(32'hb788eff3),
	.w8(32'hb6a5eb3b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c0997),
	.w1(32'hbba07dbf),
	.w2(32'hbba1d9ae),
	.w3(32'hbaf5fc21),
	.w4(32'hbb85e82e),
	.w5(32'hbb33cc84),
	.w6(32'hbac84137),
	.w7(32'hbaa7b499),
	.w8(32'hbaf8d570),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7942d3b),
	.w1(32'hb787b92d),
	.w2(32'hb730f857),
	.w3(32'hb78297f2),
	.w4(32'hb71cb7ab),
	.w5(32'hb61f0add),
	.w6(32'hb7432abd),
	.w7(32'hb6cf43d5),
	.w8(32'hb6c0b642),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ef29b),
	.w1(32'hb9e95e75),
	.w2(32'h3a163552),
	.w3(32'hb99441bd),
	.w4(32'hba32e776),
	.w5(32'hb9f77175),
	.w6(32'h37fd8926),
	.w7(32'hba16fe53),
	.w8(32'hb9298d66),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa2aa2),
	.w1(32'hb9f0bc7a),
	.w2(32'hb885b63a),
	.w3(32'hba1ac1f4),
	.w4(32'hba13b266),
	.w5(32'hb99a925b),
	.w6(32'hba20ece6),
	.w7(32'hba147feb),
	.w8(32'hb9e05e0b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5dc1957),
	.w1(32'h37ae4c6a),
	.w2(32'h370c2b3b),
	.w3(32'hb7cc6597),
	.w4(32'h353cd3a1),
	.w5(32'hb6a88977),
	.w6(32'hb7bd6041),
	.w7(32'hb6aa4e42),
	.w8(32'hb7b9e2ba),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69a6f0),
	.w1(32'hbaab274f),
	.w2(32'hba1b4f3e),
	.w3(32'hbb61e2f7),
	.w4(32'hbaeaaedd),
	.w5(32'h3a8315d5),
	.w6(32'hbb6e47f6),
	.w7(32'h39e60a92),
	.w8(32'h3bbce162),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcaf0d),
	.w1(32'h3ba35559),
	.w2(32'h3c00b1f3),
	.w3(32'h3bffde0e),
	.w4(32'h3c64c5fe),
	.w5(32'h3bed68e6),
	.w6(32'h3bc98f4e),
	.w7(32'h3b8b0b85),
	.w8(32'h3b736a45),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba822f),
	.w1(32'h3ac19144),
	.w2(32'h3a4b8a8c),
	.w3(32'h3aa21d72),
	.w4(32'h3a8a7209),
	.w5(32'h39fd1e32),
	.w6(32'h39f2de19),
	.w7(32'h394c2dbc),
	.w8(32'h396fb000),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b245f4c),
	.w1(32'h39ac479c),
	.w2(32'hbbac515e),
	.w3(32'h3b5527e9),
	.w4(32'hb9b49659),
	.w5(32'hbb702942),
	.w6(32'h3ac789b6),
	.w7(32'hba073510),
	.w8(32'hbae53ae5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ba4d9),
	.w1(32'hb84919b3),
	.w2(32'h3a37b7bf),
	.w3(32'hb98d4511),
	.w4(32'hb9dc878c),
	.w5(32'h39e7ceb6),
	.w6(32'hba2f5f46),
	.w7(32'hba0f0763),
	.w8(32'h36bd7af4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb461b78),
	.w1(32'hbada1984),
	.w2(32'h3a5d82e5),
	.w3(32'hbb47763c),
	.w4(32'hbb86999d),
	.w5(32'hba80d914),
	.w6(32'hbb3db3ee),
	.w7(32'hbb3735c7),
	.w8(32'h3b6db204),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b199f60),
	.w1(32'h3ab9ba6e),
	.w2(32'hb9be1053),
	.w3(32'h3aa8ea51),
	.w4(32'h3aae0964),
	.w5(32'h3a86e04c),
	.w6(32'hbae1265a),
	.w7(32'h3a30615e),
	.w8(32'h3a9b8d73),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a63ca),
	.w1(32'h38839f24),
	.w2(32'h3a50b4fd),
	.w3(32'hb88eb1ec),
	.w4(32'hb9ab1ac0),
	.w5(32'hb9b2fef1),
	.w6(32'hba14874f),
	.w7(32'h39d56c6f),
	.w8(32'hb95ed67d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83bf75),
	.w1(32'hbb2bbf2d),
	.w2(32'hbb24b328),
	.w3(32'hb9b03498),
	.w4(32'hbb00ae51),
	.w5(32'hbb06c7e2),
	.w6(32'hba8fb6d3),
	.w7(32'hbb177926),
	.w8(32'hbb0c52ad),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfa1f9),
	.w1(32'h38035eb4),
	.w2(32'hba6a91e6),
	.w3(32'h3b0b8612),
	.w4(32'hb8f368c8),
	.w5(32'hba28e963),
	.w6(32'h3b665b0e),
	.w7(32'h3b8d8262),
	.w8(32'h3a094f73),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba301b63),
	.w1(32'hba18bf18),
	.w2(32'hba386cee),
	.w3(32'h39b5d719),
	.w4(32'h3929c4f5),
	.w5(32'hb7a31e75),
	.w6(32'h39ebdbc3),
	.w7(32'h3929a28f),
	.w8(32'hb97bfa9b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6dac8),
	.w1(32'h3c7a685e),
	.w2(32'h3c86f457),
	.w3(32'h3c1218a2),
	.w4(32'h3c7b68c9),
	.w5(32'h3c4558a8),
	.w6(32'h3c04c23c),
	.w7(32'h3c3b78c8),
	.w8(32'h3c20cdf3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebb87e),
	.w1(32'h3bc8db20),
	.w2(32'h3bb94972),
	.w3(32'h3b81d8f7),
	.w4(32'h3bd6c9b2),
	.w5(32'h3b8beeff),
	.w6(32'h3b5292f3),
	.w7(32'h3b99fa69),
	.w8(32'h3b7cd39b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ace03),
	.w1(32'hb87a735f),
	.w2(32'hb85baaec),
	.w3(32'hb895fb08),
	.w4(32'hb8963265),
	.w5(32'hb8408125),
	.w6(32'hb8089bef),
	.w7(32'hb7baf257),
	.w8(32'h36ead0d5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b84f5),
	.w1(32'h38397805),
	.w2(32'h360a1d98),
	.w3(32'hb79f70a2),
	.w4(32'h38b8cc2b),
	.w5(32'h378608e3),
	.w6(32'hb7a47f20),
	.w7(32'h382cb721),
	.w8(32'hb8e34377),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba757fe9),
	.w1(32'hbabd6908),
	.w2(32'hba6ec845),
	.w3(32'hbaee76b0),
	.w4(32'hbb0d5952),
	.w5(32'hba93e88a),
	.w6(32'hbac39349),
	.w7(32'hbac755b5),
	.w8(32'hba369098),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d216d),
	.w1(32'h3c9c5f2e),
	.w2(32'h3c78247b),
	.w3(32'h3c48f375),
	.w4(32'h3c4c2422),
	.w5(32'h3c44f5fa),
	.w6(32'h3c867dc5),
	.w7(32'h3c45bf29),
	.w8(32'h3c5cb498),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a2ddf),
	.w1(32'hba888579),
	.w2(32'hbc087cc5),
	.w3(32'h3a103642),
	.w4(32'hbb72c838),
	.w5(32'hbbd63040),
	.w6(32'hb9ba491f),
	.w7(32'hbb4d0e5c),
	.w8(32'hbba3b850),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8dab),
	.w1(32'hbb4bc1c0),
	.w2(32'hbc0e4ba8),
	.w3(32'hba02c168),
	.w4(32'hbc09824d),
	.w5(32'hbc05a3d6),
	.w6(32'h3aba58e7),
	.w7(32'hbb272da1),
	.w8(32'hbb948527),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995a4e0),
	.w1(32'hb9b01931),
	.w2(32'hb9c27b14),
	.w3(32'h39835b33),
	.w4(32'h38bb3e2f),
	.w5(32'h38ec3832),
	.w6(32'h3946c88f),
	.w7(32'hb926d19f),
	.w8(32'hb96aeddf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9377b10),
	.w1(32'hb8fb5d23),
	.w2(32'hb90d151a),
	.w3(32'hb981a298),
	.w4(32'hb939f7da),
	.w5(32'hb911362e),
	.w6(32'hb9488495),
	.w7(32'hb8bdf94e),
	.w8(32'hb9033db3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1cdb9),
	.w1(32'hbb10f6b9),
	.w2(32'hbb870a9c),
	.w3(32'hba967369),
	.w4(32'hbbbb130e),
	.w5(32'hbb803913),
	.w6(32'hbae9c7ed),
	.w7(32'h3ac326a1),
	.w8(32'h39bc5038),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69b5c8),
	.w1(32'hba5d695a),
	.w2(32'hb896e919),
	.w3(32'hbb12e950),
	.w4(32'hbb1c6837),
	.w5(32'hbab64352),
	.w6(32'hbb0c0e6f),
	.w7(32'hbac8f698),
	.w8(32'hbaaadc35),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b000d03),
	.w1(32'hbbb27e9d),
	.w2(32'hbc19e4f6),
	.w3(32'h395da48b),
	.w4(32'hbbcc9edf),
	.w5(32'hbbee9754),
	.w6(32'hbb113528),
	.w7(32'hbb5eeb1c),
	.w8(32'hbb95f3a1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f7526),
	.w1(32'hb80f3e65),
	.w2(32'hb8745134),
	.w3(32'hb83014df),
	.w4(32'hb7d86181),
	.w5(32'hb86e35ca),
	.w6(32'hb89c9d07),
	.w7(32'hb887221b),
	.w8(32'hb89a4c48),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb738fe24),
	.w1(32'hb6833c87),
	.w2(32'hb92674c3),
	.w3(32'h37348217),
	.w4(32'hb8afcca6),
	.w5(32'hb987a865),
	.w6(32'hb871bac0),
	.w7(32'hb96b9b85),
	.w8(32'hb9afecff),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f20fc),
	.w1(32'h398eee72),
	.w2(32'hba8cc0b1),
	.w3(32'h3aacc862),
	.w4(32'h38b5c150),
	.w5(32'hbac5bd8c),
	.w6(32'h39c153ed),
	.w7(32'hba1f1beb),
	.w8(32'hba99b60a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1db8d9),
	.w1(32'hba8b9c44),
	.w2(32'hbae75cbe),
	.w3(32'h398e9f41),
	.w4(32'hba3b16c9),
	.w5(32'hbaa61eb7),
	.w6(32'h3a1b9ead),
	.w7(32'h37beaf55),
	.w8(32'hba95c056),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0953ae),
	.w1(32'hb8e907c1),
	.w2(32'hb87ea4ea),
	.w3(32'h38aecfb2),
	.w4(32'hb982924e),
	.w5(32'hb9c8e21f),
	.w6(32'hb8b09232),
	.w7(32'h3a34fc21),
	.w8(32'h3a07cddc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e7fa9),
	.w1(32'hba74378b),
	.w2(32'hba69ec32),
	.w3(32'hb9cc70af),
	.w4(32'hb9f43d57),
	.w5(32'h39b2c592),
	.w6(32'hb98853ee),
	.w7(32'hbacdb0a6),
	.w8(32'h3a461333),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba790ee),
	.w1(32'h3ab3bbb6),
	.w2(32'h3bcb1e2c),
	.w3(32'hbb28fc51),
	.w4(32'h37e6e531),
	.w5(32'hbb3daf43),
	.w6(32'hb97cad7a),
	.w7(32'hbb39cec4),
	.w8(32'h3b10df99),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba78e31),
	.w1(32'hbc395f8e),
	.w2(32'hbc676ab1),
	.w3(32'hbbc954fb),
	.w4(32'hbc83ce22),
	.w5(32'hbc58768a),
	.w6(32'hbb89bde6),
	.w7(32'hbbf21c86),
	.w8(32'hbc0c98c7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a6cb9),
	.w1(32'hbc396c3a),
	.w2(32'hbc37a72b),
	.w3(32'hbbc2cde7),
	.w4(32'hbc533506),
	.w5(32'hbc04f493),
	.w6(32'hbc044d19),
	.w7(32'hbba80b99),
	.w8(32'hbb7e4a7a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92942c7),
	.w1(32'hbaf54643),
	.w2(32'hbb1d18a5),
	.w3(32'hbac10274),
	.w4(32'hbb096f19),
	.w5(32'hbb06a83f),
	.w6(32'hba383077),
	.w7(32'hba983880),
	.w8(32'hba9c94cd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f83ab3),
	.w1(32'h393584dc),
	.w2(32'h38f10bbb),
	.w3(32'h39ab526b),
	.w4(32'h38a27a5e),
	.w5(32'hb8440942),
	.w6(32'h399a2ce5),
	.w7(32'h390e4cf6),
	.w8(32'hb8ae3c50),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9341499),
	.w1(32'hb92d2318),
	.w2(32'hb9244826),
	.w3(32'hb9a1391c),
	.w4(32'hb94a2a6a),
	.w5(32'hb911cd9e),
	.w6(32'hb990bb39),
	.w7(32'hb907a6d6),
	.w8(32'hb89dc20c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d99af),
	.w1(32'hbaa24325),
	.w2(32'hba846fac),
	.w3(32'hb81c2a59),
	.w4(32'hbaae69ff),
	.w5(32'hb9c59784),
	.w6(32'h399eabf8),
	.w7(32'hba3cb833),
	.w8(32'hb96baf0d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9b592),
	.w1(32'h3b15f41c),
	.w2(32'hbb36bfaa),
	.w3(32'h3c028ee7),
	.w4(32'h3b1606a3),
	.w5(32'hb97bc809),
	.w6(32'h3b2e31c8),
	.w7(32'h3b3655e6),
	.w8(32'hba509b17),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ae1e6),
	.w1(32'hbaf03cdb),
	.w2(32'hbbb1972b),
	.w3(32'h3afca027),
	.w4(32'hbb71e4bc),
	.w5(32'hbb93175d),
	.w6(32'hb82d3c92),
	.w7(32'hbb6290c0),
	.w8(32'hbb90f201),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae2ef7),
	.w1(32'hba35ad96),
	.w2(32'hbc0ca241),
	.w3(32'h3a635789),
	.w4(32'hbb0d6079),
	.w5(32'hbb8d2b16),
	.w6(32'h3abecde5),
	.w7(32'hbb412e46),
	.w8(32'hbbb3dfea),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91a367),
	.w1(32'h3b039b64),
	.w2(32'hbad54be2),
	.w3(32'h3b807ad7),
	.w4(32'h3b0408ef),
	.w5(32'hbb0b0293),
	.w6(32'h3bf8eca8),
	.w7(32'h3b6a86cc),
	.w8(32'hbaa1a38b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d32e7),
	.w1(32'h3c781ea7),
	.w2(32'h3c93b9b0),
	.w3(32'h3bf9867f),
	.w4(32'h3c842b14),
	.w5(32'h3c5a3de0),
	.w6(32'h3c0dedb9),
	.w7(32'h3c220c6e),
	.w8(32'h3c290706),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371f82e4),
	.w1(32'hb9ac60ec),
	.w2(32'hb9abeb73),
	.w3(32'h38e2a081),
	.w4(32'hb9b45215),
	.w5(32'hb9cb32ba),
	.w6(32'hb962da41),
	.w7(32'hb999df08),
	.w8(32'hb9817ba6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6638f),
	.w1(32'h3ac998e3),
	.w2(32'h3aba2838),
	.w3(32'h3af91695),
	.w4(32'h3b211554),
	.w5(32'h3b0dc0f2),
	.w6(32'h3b0c0827),
	.w7(32'h3b27f6dc),
	.w8(32'h3b19d3be),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942f0c7),
	.w1(32'hb9e90eca),
	.w2(32'hb95a602b),
	.w3(32'hba09beb3),
	.w4(32'hb91af333),
	.w5(32'hb941eeda),
	.w6(32'hba3f3fbc),
	.w7(32'h3500670f),
	.w8(32'h3953a882),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae35b2d),
	.w1(32'h3aaa4837),
	.w2(32'hb9fe78ac),
	.w3(32'h3a9499e5),
	.w4(32'hbadb98db),
	.w5(32'hb910acb0),
	.w6(32'h3a28c559),
	.w7(32'h39869211),
	.w8(32'h3acd7560),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e5b59),
	.w1(32'h3abd480a),
	.w2(32'h3ad33299),
	.w3(32'h3a5a633b),
	.w4(32'h3afbccdc),
	.w5(32'h3ac358e2),
	.w6(32'h3ada0f2b),
	.w7(32'h3aab4084),
	.w8(32'h3a8ee445),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10611f),
	.w1(32'h3c2a3217),
	.w2(32'h3c1ce8b6),
	.w3(32'h3bedc433),
	.w4(32'h3c3da9d0),
	.w5(32'h3b8077d3),
	.w6(32'h3ba198dc),
	.w7(32'h3bf5bd90),
	.w8(32'h3bb58721),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01bc1b),
	.w1(32'h3aaa7d45),
	.w2(32'h3ad64762),
	.w3(32'h39a66bf3),
	.w4(32'h3a573ca7),
	.w5(32'h3a89caef),
	.w6(32'h38a1e0a2),
	.w7(32'h395208a5),
	.w8(32'h39a20763),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9717856),
	.w1(32'hb95433c6),
	.w2(32'hb5ddd42b),
	.w3(32'hb94b5e37),
	.w4(32'hb94e6546),
	.w5(32'hb895ee4b),
	.w6(32'hb833fccc),
	.w7(32'hb890b50a),
	.w8(32'hb828b4e6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34f61072),
	.w1(32'hb746d111),
	.w2(32'hb7cfcd65),
	.w3(32'hb84e8b8f),
	.w4(32'hb831acfe),
	.w5(32'hb80aa6f8),
	.w6(32'hb7e1d816),
	.w7(32'hb82a3f64),
	.w8(32'hb80ff725),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388977a9),
	.w1(32'h39871c86),
	.w2(32'hb92dd3fc),
	.w3(32'hb9160105),
	.w4(32'hb89a954a),
	.w5(32'hb930d452),
	.w6(32'hb92c8f3a),
	.w7(32'h38b13c00),
	.w8(32'hb892e303),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9895c2e),
	.w1(32'hba3ca98d),
	.w2(32'hba1ff4f0),
	.w3(32'hba1f4c28),
	.w4(32'hba8c6a8b),
	.w5(32'hba36a6fc),
	.w6(32'hb9f76f70),
	.w7(32'hba4a947c),
	.w8(32'hb9e025dd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dbf87f),
	.w1(32'hb9b54e78),
	.w2(32'hba153ed7),
	.w3(32'hb9260151),
	.w4(32'hba2b04a1),
	.w5(32'hb9bcfa3d),
	.w6(32'hba9b734c),
	.w7(32'hba620544),
	.w8(32'hb9c81af1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85f405),
	.w1(32'h3b8d6ebe),
	.w2(32'h3b86bdf1),
	.w3(32'h3b2f5c7a),
	.w4(32'h3b787874),
	.w5(32'h3b624313),
	.w6(32'h3af8b87e),
	.w7(32'h3b3de9cf),
	.w8(32'h3b5aa558),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5a2a),
	.w1(32'h3bae6f69),
	.w2(32'h3b115922),
	.w3(32'h3bf73d9a),
	.w4(32'h3b253c20),
	.w5(32'h3b9e67b2),
	.w6(32'h3bb5ffe2),
	.w7(32'h3b838bd0),
	.w8(32'h3b9fee7e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3854532e),
	.w1(32'h3801791f),
	.w2(32'hb88088a0),
	.w3(32'h38cbf392),
	.w4(32'h37b44e52),
	.w5(32'hb89c911b),
	.w6(32'h38868617),
	.w7(32'h37db6b45),
	.w8(32'hb881fbe7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361978d1),
	.w1(32'h374e2caa),
	.w2(32'hb79d8885),
	.w3(32'h37b775bf),
	.w4(32'h37e685b7),
	.w5(32'hb69a67f6),
	.w6(32'h377abaa5),
	.w7(32'h37702b1b),
	.w8(32'hb756be8e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a0b24),
	.w1(32'hb949561a),
	.w2(32'hb814b29e),
	.w3(32'hb9b9633d),
	.w4(32'hb9589c44),
	.w5(32'hb90ddf68),
	.w6(32'hb9a0d5bd),
	.w7(32'hb95f800b),
	.w8(32'hb8e00322),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e16422),
	.w1(32'h37534263),
	.w2(32'hb85da0d6),
	.w3(32'hb89715fa),
	.w4(32'hb847fc3f),
	.w5(32'hb8899bd6),
	.w6(32'hb886273e),
	.w7(32'hb8367e24),
	.w8(32'hb8b463a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb330c66),
	.w1(32'h3b10c40f),
	.w2(32'h3aa73ffd),
	.w3(32'h39a96e75),
	.w4(32'hb871074d),
	.w5(32'hbb9d90d1),
	.w6(32'h3a4f1aa3),
	.w7(32'h3bb58053),
	.w8(32'h3b7b5523),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514f59),
	.w1(32'hbb3e5982),
	.w2(32'hbbc556d9),
	.w3(32'hbb07df48),
	.w4(32'hbab8e145),
	.w5(32'h379b7dd2),
	.w6(32'h3a8e4f45),
	.w7(32'hbb751f6e),
	.w8(32'hbb3911f5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5513c),
	.w1(32'h3c149483),
	.w2(32'h3bb186b3),
	.w3(32'h3ba55ba4),
	.w4(32'h3b552a60),
	.w5(32'h3bb108e5),
	.w6(32'h3be92c5f),
	.w7(32'h3bc14c4e),
	.w8(32'h3be44875),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb22d2),
	.w1(32'hbbde973e),
	.w2(32'hbc7b4557),
	.w3(32'hbad59c26),
	.w4(32'hbc6d205d),
	.w5(32'hbc5734df),
	.w6(32'h39c17e57),
	.w7(32'hbbf39266),
	.w8(32'hbc113571),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2069cf),
	.w1(32'h3a2ab2e5),
	.w2(32'hbbab4941),
	.w3(32'hbb9f3a27),
	.w4(32'hbb045dc6),
	.w5(32'hbb9770f6),
	.w6(32'hbb98df47),
	.w7(32'hbaa79250),
	.w8(32'hbb931d20),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5eab8),
	.w1(32'h395672d8),
	.w2(32'hbb9ed00f),
	.w3(32'hbb489fea),
	.w4(32'h3b7561ac),
	.w5(32'hbc26975c),
	.w6(32'hbb4cf4d7),
	.w7(32'hba452895),
	.w8(32'hba0b7aa1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b32b1),
	.w1(32'hbb2f0800),
	.w2(32'h3ab918a6),
	.w3(32'h3b8a3cab),
	.w4(32'hbb4823ff),
	.w5(32'h3c1d7e27),
	.w6(32'h3b4fc5ee),
	.w7(32'hbb25abac),
	.w8(32'h3b5cfdc6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386b244a),
	.w1(32'h3b264d57),
	.w2(32'h3befc597),
	.w3(32'hbb391d82),
	.w4(32'h3b5bb7f8),
	.w5(32'h3b00795a),
	.w6(32'hba4766da),
	.w7(32'h3ba4cbae),
	.w8(32'h3a491c3c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9523fe),
	.w1(32'hb960f506),
	.w2(32'hbb045842),
	.w3(32'hbae9462e),
	.w4(32'hb8deea72),
	.w5(32'hb999f0d9),
	.w6(32'h3b9adb27),
	.w7(32'h3a6de9de),
	.w8(32'hbb96a8d2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd9099),
	.w1(32'h3c104f2e),
	.w2(32'h3c36f8a8),
	.w3(32'h3b46c265),
	.w4(32'h3c3433fb),
	.w5(32'h3a067f8f),
	.w6(32'h3acbb104),
	.w7(32'h3bc7e737),
	.w8(32'h3b074235),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb821c4f7),
	.w1(32'h3bd276a4),
	.w2(32'h3bbd9b6f),
	.w3(32'h3b7ad769),
	.w4(32'h3c859016),
	.w5(32'h3a83983d),
	.w6(32'h3bfc16ef),
	.w7(32'h3c4ea14d),
	.w8(32'h3c14021d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fda63),
	.w1(32'hbbf6496a),
	.w2(32'h3b272542),
	.w3(32'hb9428b03),
	.w4(32'hbc806685),
	.w5(32'h3c2a456f),
	.w6(32'hba6b4027),
	.w7(32'hbab1d641),
	.w8(32'hbac8285d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac45aaf),
	.w1(32'h3b47d32d),
	.w2(32'h3add9f05),
	.w3(32'hbba12f5e),
	.w4(32'hba99ae43),
	.w5(32'h3c21568f),
	.w6(32'h3c36b51a),
	.w7(32'h3ab504c7),
	.w8(32'h3a5abbd8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98434b),
	.w1(32'hbb66c278),
	.w2(32'hbb9ecfe9),
	.w3(32'h3b25bd72),
	.w4(32'hbb714c73),
	.w5(32'hbbd497a3),
	.w6(32'h3c0fe1f4),
	.w7(32'h3b43bc7d),
	.w8(32'h3b6c4b1f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9964),
	.w1(32'hbae079eb),
	.w2(32'h3aa11d5b),
	.w3(32'hbb8d85bf),
	.w4(32'h3b2c6a38),
	.w5(32'hbb83111d),
	.w6(32'hba4307e2),
	.w7(32'h3b7f47bf),
	.w8(32'hbb3ff2c7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b3870),
	.w1(32'h3b6dc8cd),
	.w2(32'h3bdecd29),
	.w3(32'h3c29f4cc),
	.w4(32'h3b480b12),
	.w5(32'h3b7b166c),
	.w6(32'h3bcc6a75),
	.w7(32'h3b2d1db2),
	.w8(32'h3b74e531),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37a55b),
	.w1(32'hbac13314),
	.w2(32'h391ba942),
	.w3(32'h3b321211),
	.w4(32'h3b3b07d6),
	.w5(32'hbb4675e1),
	.w6(32'h3955d1a3),
	.w7(32'h3ae437c2),
	.w8(32'hbba1bb3c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33cfad),
	.w1(32'hbb2572e5),
	.w2(32'h3bd35d25),
	.w3(32'h3b0109ee),
	.w4(32'hba8567b9),
	.w5(32'h3b1d32da),
	.w6(32'h3ae86e3b),
	.w7(32'h3b76c873),
	.w8(32'hbaf84a7e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39024403),
	.w1(32'hbb563c75),
	.w2(32'hbb5711b5),
	.w3(32'hbb881edd),
	.w4(32'hbb7ffd91),
	.w5(32'h3b9672e1),
	.w6(32'hbb11b535),
	.w7(32'hbbc44f9e),
	.w8(32'h3b34c8f8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277d8a),
	.w1(32'hbbc920cf),
	.w2(32'hbb0129ee),
	.w3(32'hbbdb2d46),
	.w4(32'hba198dad),
	.w5(32'hbbae056d),
	.w6(32'hbb1b0e9e),
	.w7(32'hb9879d0e),
	.w8(32'hbb8829e1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4ca7c),
	.w1(32'hbbd2e665),
	.w2(32'h3ba05169),
	.w3(32'hbac078c5),
	.w4(32'hbc823bee),
	.w5(32'h3caf2ab0),
	.w6(32'h386f532d),
	.w7(32'hbb12aeb6),
	.w8(32'hbbc82e29),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba033e9e),
	.w1(32'hbafc8c3b),
	.w2(32'h3b53b56d),
	.w3(32'hbba5ba3d),
	.w4(32'hbc05633e),
	.w5(32'h3c69e1c5),
	.w6(32'h3b8f52e8),
	.w7(32'hb990a91f),
	.w8(32'h3b3a854d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86645d),
	.w1(32'h3bade299),
	.w2(32'hbb13e4d2),
	.w3(32'hbc17b2c9),
	.w4(32'h3b8866fe),
	.w5(32'hbad940c8),
	.w6(32'h3bc274c0),
	.w7(32'h3b78a79c),
	.w8(32'h3bc06767),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a1587),
	.w1(32'h3c940d49),
	.w2(32'h3c87b9cd),
	.w3(32'h3c5cdf52),
	.w4(32'h3c8838fe),
	.w5(32'h3cc26eea),
	.w6(32'h3c5fc3ec),
	.w7(32'h3c6f5b6b),
	.w8(32'h3c82e328),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8155f),
	.w1(32'hbbb493da),
	.w2(32'hbb9b6af7),
	.w3(32'hbb5d3a6f),
	.w4(32'hbbd02a6a),
	.w5(32'hbbb1cbe5),
	.w6(32'hbb126d04),
	.w7(32'hbbb1f046),
	.w8(32'hbb53ab23),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8167),
	.w1(32'h3acf4695),
	.w2(32'h3a031d19),
	.w3(32'hbb216971),
	.w4(32'h3abbd90f),
	.w5(32'h38e60147),
	.w6(32'hbb431f6c),
	.w7(32'h3b766b44),
	.w8(32'h3b9fa438),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3950d),
	.w1(32'hbbac6bf1),
	.w2(32'hbc2898ae),
	.w3(32'hbb903333),
	.w4(32'hbab623cb),
	.w5(32'hbc4a76fb),
	.w6(32'hbb16ddf0),
	.w7(32'hbc13f973),
	.w8(32'hbc05e628),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4c010),
	.w1(32'h3ba4a7bd),
	.w2(32'h3a7b6a09),
	.w3(32'h3c222e32),
	.w4(32'h3c0200ca),
	.w5(32'hbac70a7d),
	.w6(32'h3a69b70b),
	.w7(32'h3c0b9de7),
	.w8(32'h3b1172c6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09b5cc),
	.w1(32'hbb8aa5d5),
	.w2(32'hbb2297ca),
	.w3(32'h3b23c97e),
	.w4(32'hbb9a093f),
	.w5(32'hbb926ebc),
	.w6(32'hbac096ef),
	.w7(32'hb998eef5),
	.w8(32'h3ac2ce0f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9c2cf),
	.w1(32'hbbaa297f),
	.w2(32'hbbd201c5),
	.w3(32'hbbc07a64),
	.w4(32'hba92496a),
	.w5(32'hbc0b3dfa),
	.w6(32'hbbe71e3b),
	.w7(32'hbb44504c),
	.w8(32'hbba8e426),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a21cd1),
	.w1(32'hbbceaf6b),
	.w2(32'hbbbd0397),
	.w3(32'hbaecdc48),
	.w4(32'hbbcc2960),
	.w5(32'hbb89a47b),
	.w6(32'hbb6b9d1a),
	.w7(32'hbba5949c),
	.w8(32'hba59f12c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9f750),
	.w1(32'h3bc0c1ef),
	.w2(32'h3c03ed6d),
	.w3(32'h3a228450),
	.w4(32'h3c1181cc),
	.w5(32'h3c4d88fe),
	.w6(32'h3b85eef5),
	.w7(32'h3be457dd),
	.w8(32'h3bd3bfab),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b548b15),
	.w1(32'h3b77520f),
	.w2(32'hba360f97),
	.w3(32'h3b065524),
	.w4(32'hbb52207e),
	.w5(32'hbae05202),
	.w6(32'h39adcd5e),
	.w7(32'h390a34a4),
	.w8(32'h3c0e314b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a450d),
	.w1(32'h3c877f39),
	.w2(32'h3c1a6da5),
	.w3(32'h3b2e5408),
	.w4(32'h3bf89cd6),
	.w5(32'h3bbdb44d),
	.w6(32'h3c0c1d82),
	.w7(32'h3b3e481f),
	.w8(32'hba4ac4d5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3747c),
	.w1(32'hbc2e38da),
	.w2(32'hbbcdf168),
	.w3(32'hbc067afc),
	.w4(32'hbc4bbcbf),
	.w5(32'hbc38b2d1),
	.w6(32'h3a49aead),
	.w7(32'hbba5d78e),
	.w8(32'hbb3815a9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0117f2),
	.w1(32'hbb691e8f),
	.w2(32'hbc2c3da1),
	.w3(32'hbacfe429),
	.w4(32'hbb9bb1c0),
	.w5(32'hbb82d6b9),
	.w6(32'hbac78982),
	.w7(32'hbbb33ba4),
	.w8(32'hbbb8ea0f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab232d4),
	.w1(32'hbbefea0a),
	.w2(32'hbb951d8c),
	.w3(32'h3a1f0302),
	.w4(32'hbc048b44),
	.w5(32'hbc20ea94),
	.w6(32'hba34ba41),
	.w7(32'hbbe9ebbe),
	.w8(32'h3c04b2ee),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d98be),
	.w1(32'h3b883683),
	.w2(32'h3bef5e50),
	.w3(32'hbc003f3f),
	.w4(32'hbc24df0a),
	.w5(32'h3c84600b),
	.w6(32'hbbe6ba75),
	.w7(32'hbc61147f),
	.w8(32'h3b6bf9f7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4df949),
	.w1(32'h3cb94738),
	.w2(32'h3ca4314d),
	.w3(32'h3b146f81),
	.w4(32'h3cb643e1),
	.w5(32'h3aa46536),
	.w6(32'h3c625964),
	.w7(32'h3c4534ab),
	.w8(32'h3b74122e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b088984),
	.w1(32'hbbd21cf8),
	.w2(32'hbbe28c25),
	.w3(32'h3b680f6c),
	.w4(32'hbb9efafa),
	.w5(32'hbb25ce26),
	.w6(32'hbb981b76),
	.w7(32'hbbabaf2c),
	.w8(32'hbb5de043),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9d51e),
	.w1(32'h3b1cb17b),
	.w2(32'hba0a1f06),
	.w3(32'h3ac5f7fc),
	.w4(32'h3b869f86),
	.w5(32'h3b221863),
	.w6(32'h3a40427c),
	.w7(32'h3af06215),
	.w8(32'hbafc41ff),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ddd1e8),
	.w1(32'hbad4f809),
	.w2(32'hbae57ff5),
	.w3(32'h39f8cb78),
	.w4(32'h3a13d2d5),
	.w5(32'hba62dc84),
	.w6(32'h3bbb7734),
	.w7(32'h3adcd167),
	.w8(32'h3a974528),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf6904),
	.w1(32'hbaf32b1e),
	.w2(32'hbb7f539f),
	.w3(32'hbbf1020f),
	.w4(32'h3b19ebb5),
	.w5(32'hbbe1778f),
	.w6(32'hbb403664),
	.w7(32'hbb4aa195),
	.w8(32'hbb370f2b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06730f),
	.w1(32'h3abfffbd),
	.w2(32'hbbecb430),
	.w3(32'h3a7e57b3),
	.w4(32'h3b8f50fd),
	.w5(32'hbb430589),
	.w6(32'hbbff104b),
	.w7(32'hbb3b6032),
	.w8(32'hba9a4e69),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c049188),
	.w1(32'h39b50306),
	.w2(32'h3a9f1a4d),
	.w3(32'h3c44d0f9),
	.w4(32'h3be2388e),
	.w5(32'h3b0bb840),
	.w6(32'h3b85cbae),
	.w7(32'h3b8e54ff),
	.w8(32'h3a6a1583),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e4354),
	.w1(32'hbbe0c8ba),
	.w2(32'hbaff1721),
	.w3(32'h3b5c4ab0),
	.w4(32'hbc28d4ee),
	.w5(32'hbc107818),
	.w6(32'hbaec018e),
	.w7(32'hba817f8a),
	.w8(32'hbb448650),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b520f42),
	.w1(32'hbb87c48d),
	.w2(32'hbbaba495),
	.w3(32'hb993b579),
	.w4(32'hbba5e9ba),
	.w5(32'hbb53fcf6),
	.w6(32'hb8b7dc47),
	.w7(32'hbc04458d),
	.w8(32'hbbf8a307),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa90612),
	.w1(32'h3b91177c),
	.w2(32'h3bab302d),
	.w3(32'hba15724f),
	.w4(32'hba83f16f),
	.w5(32'hbb5093ad),
	.w6(32'h38b0b98c),
	.w7(32'h3bddeaeb),
	.w8(32'h3aabaa3e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13f124),
	.w1(32'hbb90cacc),
	.w2(32'hbc1582e5),
	.w3(32'h3c13b9d3),
	.w4(32'hbbbd5a63),
	.w5(32'hba9af024),
	.w6(32'h3c5afc51),
	.w7(32'hbb24984e),
	.w8(32'hbbe31b09),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a9ef1),
	.w1(32'hbb388e8a),
	.w2(32'hba42fdc8),
	.w3(32'h3b718d4e),
	.w4(32'hbb92c2b0),
	.w5(32'hbb333ad8),
	.w6(32'h3b53ec45),
	.w7(32'hbb2760a2),
	.w8(32'hbb6e4fd1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba746d6e),
	.w1(32'hb96a6191),
	.w2(32'hba9ae3fb),
	.w3(32'hbb741f99),
	.w4(32'h3c041d2e),
	.w5(32'hba5f0f38),
	.w6(32'hbab8680a),
	.w7(32'h3a0f98ad),
	.w8(32'hbab8f7cb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb4fc0),
	.w1(32'h3af763ec),
	.w2(32'hb98dd257),
	.w3(32'h3c1d7f55),
	.w4(32'hbb0b6bc6),
	.w5(32'hbbe29573),
	.w6(32'h3b3ddb6d),
	.w7(32'hbaf36f78),
	.w8(32'hbbf46526),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b545489),
	.w1(32'hbbf5c4b8),
	.w2(32'h3b36fff8),
	.w3(32'h3b665ca9),
	.w4(32'hbc047716),
	.w5(32'hbae2b97d),
	.w6(32'hbaf5eda7),
	.w7(32'hba0df361),
	.w8(32'hbb11318d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f6597),
	.w1(32'hbc039059),
	.w2(32'hbc10830d),
	.w3(32'hbbe870b3),
	.w4(32'h3b0f158d),
	.w5(32'hbbd191dc),
	.w6(32'hbb43081b),
	.w7(32'h3b97b90c),
	.w8(32'hbbe0bd39),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09f1d1),
	.w1(32'h3bdcdb91),
	.w2(32'h3a0d8d02),
	.w3(32'h3b4b9e30),
	.w4(32'h3c017c7f),
	.w5(32'hbaa1b328),
	.w6(32'hbaa1bbf0),
	.w7(32'h3a88539f),
	.w8(32'h3a92b723),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace9a00),
	.w1(32'h3bc9cd87),
	.w2(32'h3a6eb398),
	.w3(32'h3be609d6),
	.w4(32'h3ad378f2),
	.w5(32'hba8fac0e),
	.w6(32'h3bded213),
	.w7(32'hbab0e7d5),
	.w8(32'h3b1261b7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf5315),
	.w1(32'hbc1569e2),
	.w2(32'hbc320e49),
	.w3(32'h38ee041b),
	.w4(32'hbc12b0e6),
	.w5(32'hbc2ffff5),
	.w6(32'hbbce1bc6),
	.w7(32'hbb3fd03f),
	.w8(32'hba9bb86c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b0b44),
	.w1(32'hbb89f36e),
	.w2(32'hbc12afab),
	.w3(32'hbbb44697),
	.w4(32'h3ba09a69),
	.w5(32'hbc0a1c75),
	.w6(32'hbb0d0f11),
	.w7(32'h3b6f0809),
	.w8(32'hbae13307),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfba49),
	.w1(32'h3b887773),
	.w2(32'hba4f34f8),
	.w3(32'h3b9317a3),
	.w4(32'h3c0c382a),
	.w5(32'hbb293291),
	.w6(32'hbba9101f),
	.w7(32'hbad61d9f),
	.w8(32'h3ac62a1a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1244e),
	.w1(32'h3b038cdb),
	.w2(32'hbb8c893b),
	.w3(32'h3bcd6278),
	.w4(32'h397f41c4),
	.w5(32'hbc1798fb),
	.w6(32'h3a7b28a6),
	.w7(32'hbb890f8b),
	.w8(32'hbb48dad5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5e755),
	.w1(32'h3b8f4ba7),
	.w2(32'hbbbd3388),
	.w3(32'h3b8b194f),
	.w4(32'hbb336b95),
	.w5(32'hbb6ff67e),
	.w6(32'hb8e978b5),
	.w7(32'h3b2f3c20),
	.w8(32'h3b11f1cb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb288015),
	.w1(32'hbb848610),
	.w2(32'hbb5a4650),
	.w3(32'hbc3e0a96),
	.w4(32'h3b56b8df),
	.w5(32'h39bb8676),
	.w6(32'hbbc725a8),
	.w7(32'h3a09a046),
	.w8(32'h38b0e42f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d90b9),
	.w1(32'hb948d9f1),
	.w2(32'hbb14a108),
	.w3(32'hba07d801),
	.w4(32'h3b44281f),
	.w5(32'hbaf773a2),
	.w6(32'hbb86ea65),
	.w7(32'h3a5436c8),
	.w8(32'h39d9527f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa111fc),
	.w1(32'hbad3a949),
	.w2(32'h3b2f187c),
	.w3(32'hb994e4e9),
	.w4(32'hbb443fe1),
	.w5(32'h3bb9b427),
	.w6(32'hbb01f71c),
	.w7(32'hbaad3f74),
	.w8(32'hbb4c45eb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86635a),
	.w1(32'hbb541dba),
	.w2(32'hba0bc319),
	.w3(32'h3b9e86aa),
	.w4(32'h3b653360),
	.w5(32'h3ac58089),
	.w6(32'h3c3ae73f),
	.w7(32'h3aa2838b),
	.w8(32'h3b035fab),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6fa60),
	.w1(32'hb9fcc115),
	.w2(32'h39fbfd18),
	.w3(32'h3aae495e),
	.w4(32'hb87fcf3a),
	.w5(32'hb98da06c),
	.w6(32'hb9c58a60),
	.w7(32'hbbaca178),
	.w8(32'hbb226991),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f726f),
	.w1(32'h3aec48ab),
	.w2(32'hbb85f131),
	.w3(32'h3bdf759b),
	.w4(32'h3b391b27),
	.w5(32'hbb53e794),
	.w6(32'h3c2246ce),
	.w7(32'h3aad0093),
	.w8(32'hba854b23),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4905cb),
	.w1(32'h3b1537bd),
	.w2(32'hbc2228bc),
	.w3(32'hba74823b),
	.w4(32'hbb7274fc),
	.w5(32'hbc593ed6),
	.w6(32'hbb5d6074),
	.w7(32'h3bbd351f),
	.w8(32'hbc0ed3c0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41918e),
	.w1(32'h3bfcfa42),
	.w2(32'h3c2cf285),
	.w3(32'h39d0a377),
	.w4(32'h3b71366c),
	.w5(32'h3b14c4b6),
	.w6(32'h3b86cb7f),
	.w7(32'h3bffb13f),
	.w8(32'h3bcfc5c6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f7172),
	.w1(32'hba9b963c),
	.w2(32'hb9044c60),
	.w3(32'hbbca423c),
	.w4(32'hbb06c58c),
	.w5(32'hbbf83623),
	.w6(32'hbb774f54),
	.w7(32'h3b9809d0),
	.w8(32'hbb12ceab),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940ab04),
	.w1(32'h3b8d18e6),
	.w2(32'h3b7078df),
	.w3(32'h3ae7c9e6),
	.w4(32'hbbb5efa9),
	.w5(32'h3bb56517),
	.w6(32'h3b24e41e),
	.w7(32'hbb94f923),
	.w8(32'h3b02b2eb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3dda0),
	.w1(32'h3be4f666),
	.w2(32'h3b6d5c73),
	.w3(32'h3b58879c),
	.w4(32'h3bd2e703),
	.w5(32'hbc08a29d),
	.w6(32'h3c17f790),
	.w7(32'h3a6cc1bf),
	.w8(32'hbabb1bfc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b5ecc),
	.w1(32'hbbbdc385),
	.w2(32'hbb9f2d2b),
	.w3(32'h3aa2794a),
	.w4(32'hbbb58fe5),
	.w5(32'hbb4ed565),
	.w6(32'hba163482),
	.w7(32'hbb47b9ea),
	.w8(32'hbb87a219),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cd4a6),
	.w1(32'hbb031be2),
	.w2(32'hbba840e2),
	.w3(32'h3b016dc9),
	.w4(32'h3b4a0db3),
	.w5(32'hbafad019),
	.w6(32'h3b584656),
	.w7(32'h3b401c8e),
	.w8(32'hb98cd6f2),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac939ef),
	.w1(32'h3b974021),
	.w2(32'hba793fad),
	.w3(32'h3bcffc6d),
	.w4(32'h3a81d5e8),
	.w5(32'hbaf9ee97),
	.w6(32'h3a93d25a),
	.w7(32'h3a325f4d),
	.w8(32'hbc5bd203),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27da5c),
	.w1(32'hbb1e5f77),
	.w2(32'hbbcebd15),
	.w3(32'h3b9e3596),
	.w4(32'hbbcb09b9),
	.w5(32'h3b04a7a4),
	.w6(32'h3ba5a73f),
	.w7(32'hbbd287b9),
	.w8(32'h3b3616c9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8555c0),
	.w1(32'hbb01c391),
	.w2(32'hba908173),
	.w3(32'hbbd01d16),
	.w4(32'h3b13e555),
	.w5(32'h3af0fc1c),
	.w6(32'hba91afef),
	.w7(32'hbb0e5625),
	.w8(32'hba089c86),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99d8ee),
	.w1(32'hbaed363b),
	.w2(32'hbb8e7843),
	.w3(32'h3b416835),
	.w4(32'h3a80d220),
	.w5(32'h3a8f21a3),
	.w6(32'hbb33c86e),
	.w7(32'h39f7d893),
	.w8(32'h3a0bc9ae),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d997e),
	.w1(32'h3aad5ffd),
	.w2(32'hb94210d3),
	.w3(32'hbbd3d699),
	.w4(32'h3b848933),
	.w5(32'h3b8084d4),
	.w6(32'hbb98fe16),
	.w7(32'hba492f01),
	.w8(32'h3ac070d0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafea2fb),
	.w1(32'h3a87f372),
	.w2(32'hbb9104d0),
	.w3(32'h3a3893fd),
	.w4(32'h3b578c96),
	.w5(32'hba5eaf65),
	.w6(32'hba7a8a57),
	.w7(32'hbb05e9b0),
	.w8(32'h3bb48469),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80b208),
	.w1(32'hbaec8a52),
	.w2(32'h3b66350b),
	.w3(32'hbbd5e3dc),
	.w4(32'hbb65cdd1),
	.w5(32'h3b194222),
	.w6(32'hbbabf87a),
	.w7(32'h39b21145),
	.w8(32'h3b99fb35),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83bb3c),
	.w1(32'h3b267ef6),
	.w2(32'hbaff0b5f),
	.w3(32'h3b8c7649),
	.w4(32'h3ac4ec86),
	.w5(32'h3add7f53),
	.w6(32'h3ae4f01d),
	.w7(32'hbb98eba6),
	.w8(32'hbbd95c69),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb167859),
	.w1(32'h3a8d1e1c),
	.w2(32'hbb135af7),
	.w3(32'hbc1aa7b7),
	.w4(32'h3b144a69),
	.w5(32'hbb1203e9),
	.w6(32'h3b976cf7),
	.w7(32'h3baab090),
	.w8(32'hb901e73c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e74cc),
	.w1(32'hba0e4419),
	.w2(32'hbac4c153),
	.w3(32'h3b80441c),
	.w4(32'hbb7921d8),
	.w5(32'hbb931e95),
	.w6(32'h3b755f83),
	.w7(32'h3a94d289),
	.w8(32'hb9f252fa),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc932f),
	.w1(32'h3a328261),
	.w2(32'h3b3c64a9),
	.w3(32'h3aa43e3d),
	.w4(32'h3b57b4e6),
	.w5(32'hbb41ad00),
	.w6(32'hbb01004e),
	.w7(32'h3ba11d41),
	.w8(32'h3b28ffd6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c125d4c),
	.w1(32'hba500d60),
	.w2(32'h3befb6b8),
	.w3(32'h3b8932bc),
	.w4(32'hbb15b1dd),
	.w5(32'h3b4c6eeb),
	.w6(32'h3aefb284),
	.w7(32'h3a16b59c),
	.w8(32'h3c3c7a8c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21aafc),
	.w1(32'hbb08571c),
	.w2(32'hbbd7a2b9),
	.w3(32'hbb03cd57),
	.w4(32'hbc47e267),
	.w5(32'h3bbb1214),
	.w6(32'hbbe8c7f7),
	.w7(32'hbb698796),
	.w8(32'h3b9f0427),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39beeddd),
	.w1(32'h3aaeb240),
	.w2(32'hbb179e4a),
	.w3(32'hbc09c054),
	.w4(32'h3b29d1ad),
	.w5(32'hbb4f6a68),
	.w6(32'hbb4329b9),
	.w7(32'h3b9c0ab5),
	.w8(32'hbb570afe),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2239c9),
	.w1(32'hbb710a3d),
	.w2(32'hbb3330a3),
	.w3(32'hbb23afc0),
	.w4(32'hbba707b5),
	.w5(32'hbc083dee),
	.w6(32'hbae381e0),
	.w7(32'hbb5ebba2),
	.w8(32'hbb5b86f6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5658bb),
	.w1(32'h3ae2d3de),
	.w2(32'hbb01b4f3),
	.w3(32'h3a79d030),
	.w4(32'h3af6130d),
	.w5(32'hbb6f53b6),
	.w6(32'hbaf41913),
	.w7(32'hb8d1d4b6),
	.w8(32'hbb32aa58),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34eb16),
	.w1(32'hba95042c),
	.w2(32'hbb69d46c),
	.w3(32'hbaf33385),
	.w4(32'hbb2235df),
	.w5(32'hbbe1d2f2),
	.w6(32'hbb8874b6),
	.w7(32'h3b6fb835),
	.w8(32'hbb25165f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195d01),
	.w1(32'hbbaef60f),
	.w2(32'hbc0d9751),
	.w3(32'hbb6ae460),
	.w4(32'hbb6a47b3),
	.w5(32'hbc20a830),
	.w6(32'hba227f17),
	.w7(32'hba7dca2e),
	.w8(32'hbb60a726),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba898ea3),
	.w1(32'h3bd1fe93),
	.w2(32'hbaa3ff03),
	.w3(32'h3a8dd3d2),
	.w4(32'h3c161db9),
	.w5(32'h3a6ae66b),
	.w6(32'hbb2f1efe),
	.w7(32'h3bbfc093),
	.w8(32'h3b3b46ed),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb642ac0),
	.w1(32'hb9c48937),
	.w2(32'hbac00bea),
	.w3(32'hbb874f3d),
	.w4(32'h3a62c8ec),
	.w5(32'hb9357cf8),
	.w6(32'hb9ededd7),
	.w7(32'h3bb7cf30),
	.w8(32'hbbbbf2b3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8c68e),
	.w1(32'hbb183cf3),
	.w2(32'h3c20344e),
	.w3(32'h3bca6d0a),
	.w4(32'hbb05eb32),
	.w5(32'h3c50630c),
	.w6(32'h3a82dfef),
	.w7(32'h3a9c47b0),
	.w8(32'h3b938585),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9054584),
	.w1(32'hba020f8f),
	.w2(32'hb8d2cd60),
	.w3(32'hbbd83974),
	.w4(32'hbb5447b2),
	.w5(32'hbb36c1e4),
	.w6(32'h39b49763),
	.w7(32'hb893bebb),
	.w8(32'hbaa1af71),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0b796),
	.w1(32'h3b900230),
	.w2(32'h3b5789db),
	.w3(32'hb94aa4ae),
	.w4(32'hbaa43371),
	.w5(32'h3b8ba969),
	.w6(32'hbabf88d0),
	.w7(32'hba73a106),
	.w8(32'h3b9a5051),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f41f59),
	.w1(32'hba4e8732),
	.w2(32'h3ac58b50),
	.w3(32'hbb9681da),
	.w4(32'hba5d2518),
	.w5(32'h3bdacd1f),
	.w6(32'hbb04317e),
	.w7(32'hba04edb2),
	.w8(32'h39fcdaba),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb34e81),
	.w1(32'hbbbc3097),
	.w2(32'hb9c4187b),
	.w3(32'hb9844ce1),
	.w4(32'hbbf75df0),
	.w5(32'h3bf7cce0),
	.w6(32'h3a917f81),
	.w7(32'hbb1a99b1),
	.w8(32'h3aa35073),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab69ce1),
	.w1(32'hba604625),
	.w2(32'h3bdfdbf7),
	.w3(32'h3b0f1c07),
	.w4(32'hbc180ee9),
	.w5(32'h3c7a6f1b),
	.w6(32'h3ba567e9),
	.w7(32'hbb5927d4),
	.w8(32'hbba07b36),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e01b6),
	.w1(32'hba9821fb),
	.w2(32'hbba1322e),
	.w3(32'h3a55f872),
	.w4(32'h3b1272a0),
	.w5(32'hbbd77d16),
	.w6(32'h3c3a5c99),
	.w7(32'hb9e7c701),
	.w8(32'hbb35f7a1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95a87c),
	.w1(32'hba895758),
	.w2(32'h3be83f1e),
	.w3(32'h3b776827),
	.w4(32'hbba24d53),
	.w5(32'h3c4053cc),
	.w6(32'hbb317b0a),
	.w7(32'hbb678965),
	.w8(32'hbba46775),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bc3bb),
	.w1(32'h3b90aab9),
	.w2(32'hbba82037),
	.w3(32'h3bc6f7cf),
	.w4(32'h3c8f4e1f),
	.w5(32'hbc1721a9),
	.w6(32'h3c9cc485),
	.w7(32'h3bc6d113),
	.w8(32'h3b9525b5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8a84),
	.w1(32'hbb13457b),
	.w2(32'hbb151eee),
	.w3(32'hbb0561d0),
	.w4(32'hba2e2edc),
	.w5(32'hba8bdfa8),
	.w6(32'hba954497),
	.w7(32'hbb064290),
	.w8(32'h397cc8e1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b488083),
	.w1(32'hbb13b2a4),
	.w2(32'h39f66220),
	.w3(32'hb91aa7e7),
	.w4(32'hbbec177a),
	.w5(32'h3c65bc17),
	.w6(32'hbb44f494),
	.w7(32'hbbfdb2e6),
	.w8(32'hba4c2c19),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf84776),
	.w1(32'hbaaf756f),
	.w2(32'hbb8c1adb),
	.w3(32'hbad936dc),
	.w4(32'hba978332),
	.w5(32'hbbe830e2),
	.w6(32'h3b682bad),
	.w7(32'hbb007f02),
	.w8(32'hbb019202),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c7bee),
	.w1(32'h3b45d8a1),
	.w2(32'h3b20aed7),
	.w3(32'h3aca638a),
	.w4(32'hba7e6c73),
	.w5(32'h3a78b38a),
	.w6(32'hb636ea64),
	.w7(32'h3ab65a48),
	.w8(32'h3b44c94d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b633ae),
	.w1(32'h3abb68f6),
	.w2(32'hbbc1d74c),
	.w3(32'hbabda179),
	.w4(32'hba9f60e3),
	.w5(32'hbb847d9c),
	.w6(32'h3abc3502),
	.w7(32'hbac11dae),
	.w8(32'h390bcf50),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1440c5),
	.w1(32'h3b4d36fa),
	.w2(32'hbb8916d3),
	.w3(32'hbaa6e8af),
	.w4(32'h3c3ca94b),
	.w5(32'hbb4ba460),
	.w6(32'hba3c497f),
	.w7(32'h3b7aa427),
	.w8(32'h3a132043),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b9b9a),
	.w1(32'hbb01187f),
	.w2(32'h3b6ec571),
	.w3(32'h3b94fe16),
	.w4(32'hbacd674c),
	.w5(32'h39c93970),
	.w6(32'h3aacd3dc),
	.w7(32'hba939b32),
	.w8(32'hbb0f0c93),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18ea35),
	.w1(32'h3b962efe),
	.w2(32'hbbdced77),
	.w3(32'h3a24ed2e),
	.w4(32'h3bf5eb31),
	.w5(32'hbbc71541),
	.w6(32'h39d3880c),
	.w7(32'h3aa349dc),
	.w8(32'h3ad98053),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1edb98),
	.w1(32'hbb32fd33),
	.w2(32'hbc2d8652),
	.w3(32'h3afc6750),
	.w4(32'h3c22d4f5),
	.w5(32'hbbef1492),
	.w6(32'h3aea7e51),
	.w7(32'h3c0334fe),
	.w8(32'hbb5b7f7c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb61344),
	.w1(32'h3b98118a),
	.w2(32'h39c630b1),
	.w3(32'h3c061032),
	.w4(32'h3b2b02c9),
	.w5(32'hb91ee0d6),
	.w6(32'hbb1c4a5d),
	.w7(32'h3b82eba4),
	.w8(32'h3be02454),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917831),
	.w1(32'hbbbac740),
	.w2(32'h3beb580f),
	.w3(32'h3b9571bf),
	.w4(32'hbbba1396),
	.w5(32'h3a94a1cd),
	.w6(32'h3a1fb789),
	.w7(32'hbb761fbe),
	.w8(32'hbb121e74),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add19a1),
	.w1(32'hb855e5c8),
	.w2(32'hbabdc5b4),
	.w3(32'h3a7c5b7c),
	.w4(32'hbb3c82a2),
	.w5(32'hbac560b0),
	.w6(32'h3b7e07e2),
	.w7(32'h3b7cb64b),
	.w8(32'h3afda916),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb103c3e),
	.w1(32'hbb462989),
	.w2(32'h3bfa50fa),
	.w3(32'hbbb41f7f),
	.w4(32'hbbbc33a9),
	.w5(32'h3c8ddc8e),
	.w6(32'hbb4a3efb),
	.w7(32'h3a91f524),
	.w8(32'h3b205eeb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb744d12),
	.w1(32'h3a44ff56),
	.w2(32'h3b952039),
	.w3(32'hbc0876d1),
	.w4(32'hbbaad455),
	.w5(32'h3c752635),
	.w6(32'h3af94cd0),
	.w7(32'hbaab0a5a),
	.w8(32'hbbc5c1e7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850d4b),
	.w1(32'h39042a0b),
	.w2(32'h3b6cf5a2),
	.w3(32'hbb8eb740),
	.w4(32'hbc402f15),
	.w5(32'h3cc475e9),
	.w6(32'h3bad9196),
	.w7(32'hbb171a15),
	.w8(32'hbb6848b2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf763e6),
	.w1(32'h3b87a364),
	.w2(32'hb9ee83a7),
	.w3(32'hbc3e4a66),
	.w4(32'hbaae8b78),
	.w5(32'hbbd9f06d),
	.w6(32'h3b2a6f66),
	.w7(32'h3b882e1f),
	.w8(32'h3ade70ac),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62bb31),
	.w1(32'h3a01367a),
	.w2(32'h3ad106fd),
	.w3(32'h39ce1f94),
	.w4(32'hbb834f65),
	.w5(32'hbab229c0),
	.w6(32'h3b8d08c4),
	.w7(32'hbb47b962),
	.w8(32'hbab39579),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c6e24),
	.w1(32'h3b831494),
	.w2(32'h3bd9ea4c),
	.w3(32'hbb82be48),
	.w4(32'hbb0311ca),
	.w5(32'h3bdf439c),
	.w6(32'h3ad95b55),
	.w7(32'hbbd06142),
	.w8(32'hb8d042f5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba131ea5),
	.w1(32'h3c0ae762),
	.w2(32'h3bc19283),
	.w3(32'h3b77be54),
	.w4(32'h3b430abc),
	.w5(32'h3ca58667),
	.w6(32'h3b0d09c3),
	.w7(32'h3be98a7c),
	.w8(32'h3b894317),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a616966),
	.w1(32'hbbda491f),
	.w2(32'hbc51dd61),
	.w3(32'hbbe906c1),
	.w4(32'hbc0957b6),
	.w5(32'hbc26a1e8),
	.w6(32'hbaf68b36),
	.w7(32'h3b02661e),
	.w8(32'h3b05b263),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f9ed3),
	.w1(32'hbb6752e8),
	.w2(32'hbb03a7bf),
	.w3(32'hbba63289),
	.w4(32'h3b0eb19c),
	.w5(32'hbb78fadb),
	.w6(32'hba932304),
	.w7(32'hbbad46dd),
	.w8(32'hbaa80621),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a010f68),
	.w1(32'hbab07288),
	.w2(32'h3acc0c1c),
	.w3(32'h3b936f49),
	.w4(32'h390a38d7),
	.w5(32'h3c391cfa),
	.w6(32'hb935323f),
	.w7(32'hb98bcea1),
	.w8(32'h3bfb5eb0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab23eb1),
	.w1(32'h3b90a232),
	.w2(32'h3aebba36),
	.w3(32'hb93dc1db),
	.w4(32'h3bb42a02),
	.w5(32'hbae7d448),
	.w6(32'h3b88305c),
	.w7(32'h3bc2c25a),
	.w8(32'h3b934d03),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394556a6),
	.w1(32'h3b2918bf),
	.w2(32'h3b21d8a7),
	.w3(32'h3a95e8da),
	.w4(32'h3b945110),
	.w5(32'h3b16224a),
	.w6(32'hba12c1a0),
	.w7(32'h3b5e033c),
	.w8(32'h3a05400f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6563b1),
	.w1(32'hbb2b919b),
	.w2(32'hbbca6f74),
	.w3(32'h3a96dffd),
	.w4(32'h3b82f3a7),
	.w5(32'hbb3c4ef8),
	.w6(32'h3b3bfdbc),
	.w7(32'hb957daf5),
	.w8(32'hbad82b89),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc25d8),
	.w1(32'hba5637fc),
	.w2(32'h3b5dcbde),
	.w3(32'h39a0f989),
	.w4(32'h3b0352c1),
	.w5(32'h3ab2054a),
	.w6(32'hbb82c7ad),
	.w7(32'h3b24b614),
	.w8(32'h3b053f7b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd73189),
	.w1(32'hbb91a94e),
	.w2(32'hbc0929fc),
	.w3(32'h3ae81b59),
	.w4(32'hbbff0ca3),
	.w5(32'hbc0b8313),
	.w6(32'hbb0d5ae1),
	.w7(32'hbbaa6643),
	.w8(32'hbbd0afc8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affe5cd),
	.w1(32'hbc143621),
	.w2(32'hbaee8756),
	.w3(32'h39696aee),
	.w4(32'hbc03cf6b),
	.w5(32'h3a00510a),
	.w6(32'hbb6ac65c),
	.w7(32'hbb64e8b6),
	.w8(32'hbbdd7b05),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73a6a8),
	.w1(32'h3a05ad54),
	.w2(32'hba126972),
	.w3(32'hb9a3c285),
	.w4(32'h3a56fc50),
	.w5(32'h3b66ab71),
	.w6(32'hbba797f9),
	.w7(32'h3b1bf090),
	.w8(32'h3b74205a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b4557),
	.w1(32'hbb083aea),
	.w2(32'hbae95224),
	.w3(32'hbb29bceb),
	.w4(32'hbb067c0a),
	.w5(32'hbac8d69c),
	.w6(32'hba205ec4),
	.w7(32'hbb7bf364),
	.w8(32'hbb3ad5d9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba901e78),
	.w1(32'hb9f9f56c),
	.w2(32'hbae4f553),
	.w3(32'hb927933f),
	.w4(32'h39eccad3),
	.w5(32'h3a2fc6c3),
	.w6(32'hbab02c70),
	.w7(32'hb9c1c30a),
	.w8(32'hba488412),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0811ea),
	.w1(32'h3afb9218),
	.w2(32'h3b48e3e9),
	.w3(32'h3a5b858b),
	.w4(32'h3b584017),
	.w5(32'h398acaf9),
	.w6(32'h3a30b4e6),
	.w7(32'hbafb3dd0),
	.w8(32'h398b5410),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2469fd),
	.w1(32'h39bcf847),
	.w2(32'hb905e5a1),
	.w3(32'hbb2d7f43),
	.w4(32'hb9915022),
	.w5(32'h39c504c5),
	.w6(32'hbb011a2e),
	.w7(32'h3aa3b778),
	.w8(32'h3a85e081),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efb8ed),
	.w1(32'h3b33a851),
	.w2(32'h3b26345a),
	.w3(32'h3b0fdb25),
	.w4(32'h3afdd882),
	.w5(32'h3af15112),
	.w6(32'h3a7b885d),
	.w7(32'h3962f312),
	.w8(32'h3b1702a6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba01abf),
	.w1(32'hbbaa772b),
	.w2(32'hbbe7a913),
	.w3(32'h39e5bfef),
	.w4(32'hbbd387db),
	.w5(32'hbbc9b060),
	.w6(32'h3adb4072),
	.w7(32'hbaa83422),
	.w8(32'hbb0f90d9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1aec3c),
	.w1(32'hbb3286c1),
	.w2(32'hbb8f82f6),
	.w3(32'hba52c9b6),
	.w4(32'hbb81b093),
	.w5(32'hbb206c71),
	.w6(32'hba9d282c),
	.w7(32'hbb72760c),
	.w8(32'hbacbc8b3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a181b8),
	.w1(32'hba5e6c7d),
	.w2(32'hb98afb24),
	.w3(32'hba935b1d),
	.w4(32'hbb2b3842),
	.w5(32'hbb4d978a),
	.w6(32'h3aa290d2),
	.w7(32'hba9c13b0),
	.w8(32'hbadd48c5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073470),
	.w1(32'hbb700c9d),
	.w2(32'hbbacbd0c),
	.w3(32'hbabde458),
	.w4(32'hbb56ee69),
	.w5(32'hbb3f59b9),
	.w6(32'hbbba0658),
	.w7(32'hbaf8b326),
	.w8(32'hbb72f23f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e9e7f),
	.w1(32'h3a0edc90),
	.w2(32'h3aac8522),
	.w3(32'h3b9f80ea),
	.w4(32'h3ac0df7e),
	.w5(32'h3ba28688),
	.w6(32'h3b3fabb7),
	.w7(32'h3b00804b),
	.w8(32'h3a3f3102),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfe3b6),
	.w1(32'h3b88acf1),
	.w2(32'hba8f1c07),
	.w3(32'hba4e08d0),
	.w4(32'h3b024863),
	.w5(32'hbaf10822),
	.w6(32'hbb819882),
	.w7(32'h3b3e91ee),
	.w8(32'h3af87389),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819127),
	.w1(32'h3a0c7d38),
	.w2(32'h3a0a66ef),
	.w3(32'h3b57a01b),
	.w4(32'h398e5149),
	.w5(32'h3a2175a1),
	.w6(32'h3bb214b5),
	.w7(32'hb7ada0d1),
	.w8(32'hb8c4f1e7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6a21d),
	.w1(32'h39cbaa95),
	.w2(32'hb95802e2),
	.w3(32'hb9b13bcb),
	.w4(32'hba3bdf9b),
	.w5(32'h3937a892),
	.w6(32'hba226358),
	.w7(32'hbac7c0e4),
	.w8(32'hbabca59b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84393b2),
	.w1(32'hbb87445c),
	.w2(32'hbbe74f57),
	.w3(32'hbb9f67ef),
	.w4(32'hbb17771b),
	.w5(32'hbb6f7032),
	.w6(32'hba8ae7d3),
	.w7(32'hbb417130),
	.w8(32'hbbb0faac),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dbcf0),
	.w1(32'h3bca9378),
	.w2(32'h3b254c69),
	.w3(32'hb88e29e3),
	.w4(32'h3b8d81f4),
	.w5(32'h391491ea),
	.w6(32'h3bd15f8a),
	.w7(32'h3b6f199c),
	.w8(32'h3b20d883),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b630d64),
	.w1(32'hbb72a042),
	.w2(32'hbbcc33df),
	.w3(32'h3a751307),
	.w4(32'hbb5f5f0a),
	.w5(32'hbb8ecae0),
	.w6(32'h39eb92ea),
	.w7(32'hbb2c233a),
	.w8(32'hbb78dd08),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f5294),
	.w1(32'hb9dc8ea1),
	.w2(32'hba6b9400),
	.w3(32'hbab553b6),
	.w4(32'hbbde34ca),
	.w5(32'hbc1526c2),
	.w6(32'hbad4a909),
	.w7(32'hb98ee344),
	.w8(32'h3b4041ff),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55fb54),
	.w1(32'hba292892),
	.w2(32'hb980cc1b),
	.w3(32'hba5fe25a),
	.w4(32'hb7d6cb62),
	.w5(32'h39171413),
	.w6(32'hba12e49a),
	.w7(32'h39e25858),
	.w8(32'h3b1691a9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d8e98),
	.w1(32'h39f82686),
	.w2(32'hba86ac4a),
	.w3(32'h3a256689),
	.w4(32'hba4b61f0),
	.w5(32'h38e50d93),
	.w6(32'h3a20afb2),
	.w7(32'hb9e5893f),
	.w8(32'hbaa28e14),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55e84c),
	.w1(32'hbb6afc9b),
	.w2(32'h3ab1d32b),
	.w3(32'hbb8393ed),
	.w4(32'hbad5c4ea),
	.w5(32'h3b4bff48),
	.w6(32'h3a681060),
	.w7(32'hbb567d56),
	.w8(32'h3a015e51),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b530f02),
	.w1(32'h3c3c21f3),
	.w2(32'h3bceb480),
	.w3(32'h3bdc724e),
	.w4(32'h3bf94d54),
	.w5(32'h3bdab327),
	.w6(32'h3b6ee29a),
	.w7(32'h3b9848cc),
	.w8(32'h3be86a09),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba05b9b),
	.w1(32'h3a8e5d8c),
	.w2(32'h3b74e682),
	.w3(32'hba6b9246),
	.w4(32'h3bd170ca),
	.w5(32'h3b3520f7),
	.w6(32'h3baa25d0),
	.w7(32'h3b723b23),
	.w8(32'h3b3b6c74),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdd98d),
	.w1(32'hbac1fd06),
	.w2(32'hbb24dbc0),
	.w3(32'hbaafc0df),
	.w4(32'hbb475006),
	.w5(32'hbb367911),
	.w6(32'hba690e6a),
	.w7(32'hb9738bd9),
	.w8(32'hbb1145b3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b970177),
	.w1(32'hbb589e53),
	.w2(32'hbb9a1eef),
	.w3(32'h3b6682e3),
	.w4(32'hbb544d05),
	.w5(32'hbb80a54c),
	.w6(32'h3b1cddbb),
	.w7(32'h3ac813f3),
	.w8(32'hba3622e4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e8175),
	.w1(32'h3916ed1d),
	.w2(32'hba942a29),
	.w3(32'hbaff0436),
	.w4(32'hb9c1e6b7),
	.w5(32'hb9c7cbdc),
	.w6(32'hba8c14c7),
	.w7(32'h3737a69b),
	.w8(32'hbadbe2fc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfacbb),
	.w1(32'hb9ea4efc),
	.w2(32'hba66acdc),
	.w3(32'hbabb2f9c),
	.w4(32'hb961110a),
	.w5(32'h39c53fa0),
	.w6(32'hbab387e4),
	.w7(32'h3809cf86),
	.w8(32'h3b0ad9ba),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa70c84),
	.w1(32'hba0ce722),
	.w2(32'h3986db6f),
	.w3(32'h3a11b518),
	.w4(32'h3986c6ee),
	.w5(32'h3aaaab9a),
	.w6(32'h38c7564f),
	.w7(32'h39bef690),
	.w8(32'h39a945b7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b1099),
	.w1(32'h3abb2a7d),
	.w2(32'h3a21672d),
	.w3(32'h3813c343),
	.w4(32'hba189996),
	.w5(32'h39f85ed4),
	.w6(32'hbadfa8f3),
	.w7(32'h394cdddb),
	.w8(32'h37ae914c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015a27),
	.w1(32'hba5edafe),
	.w2(32'h3a773a9e),
	.w3(32'h3a3d5dd1),
	.w4(32'h3a00d74f),
	.w5(32'h3b460cb8),
	.w6(32'hbaab86f9),
	.w7(32'h3a0658e2),
	.w8(32'h3aae7b4a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93bce7f),
	.w1(32'h3aaca74d),
	.w2(32'h3a08c6a9),
	.w3(32'h3b38c135),
	.w4(32'hbb17c999),
	.w5(32'h3b41922e),
	.w6(32'h3b7bc673),
	.w7(32'hbada8cd4),
	.w8(32'hbab68a9a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2c8df),
	.w1(32'hba7cbd07),
	.w2(32'hbb068945),
	.w3(32'h3ade58b2),
	.w4(32'hbacaef3c),
	.w5(32'hbab20b15),
	.w6(32'hbafc2251),
	.w7(32'hb9b503ce),
	.w8(32'hb9dd9545),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987ce1f),
	.w1(32'hba2bd43f),
	.w2(32'hb8df5c8e),
	.w3(32'hb9223013),
	.w4(32'hb9ec13ae),
	.w5(32'hba1c3db9),
	.w6(32'h3a816d1a),
	.w7(32'hb9049ac8),
	.w8(32'hba8cf47b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc6464),
	.w1(32'h3bdfb712),
	.w2(32'h3c17191c),
	.w3(32'h3b83f736),
	.w4(32'h3bdd0b03),
	.w5(32'h3bcd7f66),
	.w6(32'h3b91f986),
	.w7(32'h3b8c1e9a),
	.w8(32'h3bc7cb06),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2ed99),
	.w1(32'h3b2a02fb),
	.w2(32'h3b74a393),
	.w3(32'h3b419ca7),
	.w4(32'h3b17f8f8),
	.w5(32'h3a029830),
	.w6(32'hb8eefc00),
	.w7(32'h3b5b59fe),
	.w8(32'h39af0187),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94a48b),
	.w1(32'h3919adc7),
	.w2(32'h391d5d3d),
	.w3(32'h3a8eb934),
	.w4(32'hba57c878),
	.w5(32'hbae2e875),
	.w6(32'hba60258f),
	.w7(32'hbad96623),
	.w8(32'hbb131336),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7939f),
	.w1(32'h3ba825a1),
	.w2(32'h3b70efe4),
	.w3(32'h3b65a904),
	.w4(32'h3b76b861),
	.w5(32'h3abeac18),
	.w6(32'h3addb1d1),
	.w7(32'h3ac41027),
	.w8(32'h3aea2eb2),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939b06a),
	.w1(32'h3ab31134),
	.w2(32'h3a803881),
	.w3(32'hba15a2d3),
	.w4(32'h3acbae55),
	.w5(32'h3a810f32),
	.w6(32'hba15a49d),
	.w7(32'h3aac38f3),
	.w8(32'h3a8cd058),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaac197),
	.w1(32'h3a9c5739),
	.w2(32'hb7fc1ed5),
	.w3(32'h3ac08768),
	.w4(32'h3ac5f0ca),
	.w5(32'h3a4707eb),
	.w6(32'h3a9ff4ce),
	.w7(32'hb9fc5c33),
	.w8(32'h39fbffdc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a174b88),
	.w1(32'h3a96d29a),
	.w2(32'h3b12c756),
	.w3(32'h3aba9c78),
	.w4(32'h3a178e4a),
	.w5(32'hba38baa6),
	.w6(32'h3b0180ba),
	.w7(32'h3a931c25),
	.w8(32'h3a139d9b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac278db),
	.w1(32'hbaf8ecb3),
	.w2(32'hba2fdbec),
	.w3(32'h3afed96a),
	.w4(32'hba06aa6f),
	.w5(32'hbb2028b4),
	.w6(32'h3b091126),
	.w7(32'hba47b138),
	.w8(32'hbab0aa32),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace5761),
	.w1(32'h39ae5964),
	.w2(32'h3a247aa6),
	.w3(32'h3925161b),
	.w4(32'h39d340c3),
	.w5(32'hba2592a7),
	.w6(32'hba8cb16e),
	.w7(32'hb9cdefee),
	.w8(32'hbb4ef988),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fdd2e),
	.w1(32'h3a56cd63),
	.w2(32'h399d878b),
	.w3(32'h3b7115ec),
	.w4(32'hbae33c49),
	.w5(32'hbb4ddedf),
	.w6(32'h38a82047),
	.w7(32'h3b49c89b),
	.w8(32'h39f18a4f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae61a5a),
	.w1(32'h3bb4cfd6),
	.w2(32'h3b6cd004),
	.w3(32'h3abd4d49),
	.w4(32'h3b46a378),
	.w5(32'h3b07af00),
	.w6(32'hbabc234f),
	.w7(32'h3a9325c7),
	.w8(32'h3b15a3f1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba62af0),
	.w1(32'h3bbf6a95),
	.w2(32'h3b316208),
	.w3(32'h3bf040a7),
	.w4(32'h3b948083),
	.w5(32'h3b6ea765),
	.w6(32'h3b84d5be),
	.w7(32'h3bbe4130),
	.w8(32'h3b7b6e81),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b8c7f),
	.w1(32'hbabe3ccb),
	.w2(32'hbaa1459e),
	.w3(32'h3960443e),
	.w4(32'hba461c0f),
	.w5(32'hba02e886),
	.w6(32'h3a1184fb),
	.w7(32'hba1b1a83),
	.w8(32'hbb1ae7ae),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f95876),
	.w1(32'hbb14c57a),
	.w2(32'hbaf1e27d),
	.w3(32'hba7d829b),
	.w4(32'hbacb7fad),
	.w5(32'hb79bd0d5),
	.w6(32'hb9d9ace9),
	.w7(32'hbb01ad5e),
	.w8(32'hba811fa1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac57785),
	.w1(32'hba52de94),
	.w2(32'h36b0f8fe),
	.w3(32'hbb031a4c),
	.w4(32'h3a8125f2),
	.w5(32'hbb019455),
	.w6(32'hbad43996),
	.w7(32'h3a872b69),
	.w8(32'h39f460d0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abce5f4),
	.w1(32'hb9217b18),
	.w2(32'h390fd04c),
	.w3(32'h3aa287e7),
	.w4(32'h399d6d0d),
	.w5(32'hb9f70380),
	.w6(32'h3a5f2c5e),
	.w7(32'h3a63c78b),
	.w8(32'hba04cb65),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38906f6c),
	.w1(32'h3b5aa197),
	.w2(32'h3b8e69d7),
	.w3(32'hb937f383),
	.w4(32'h3b543256),
	.w5(32'h3b7c86a9),
	.w6(32'h38277f5b),
	.w7(32'h3b881f89),
	.w8(32'h3b9ed66e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae31cfc),
	.w1(32'h3a0b9ecd),
	.w2(32'h3b07d597),
	.w3(32'h3b19f2bb),
	.w4(32'h3ac69d5e),
	.w5(32'hb836ecba),
	.w6(32'h3aef4684),
	.w7(32'h3af198f1),
	.w8(32'h3a85951b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4052c),
	.w1(32'hb9afd15e),
	.w2(32'hbaaf6700),
	.w3(32'hbabf4f93),
	.w4(32'hb9a6a340),
	.w5(32'h3a2386d6),
	.w6(32'hb95e32e4),
	.w7(32'hb961aae4),
	.w8(32'h39fb0c61),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b78c6),
	.w1(32'hbb082403),
	.w2(32'hbb057e24),
	.w3(32'hbacfb735),
	.w4(32'hba6bddf8),
	.w5(32'hba94e488),
	.w6(32'h3a3da166),
	.w7(32'hbb0807f4),
	.w8(32'hba825a5a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3dad6),
	.w1(32'hb95c2a21),
	.w2(32'hb9335a05),
	.w3(32'hb8908f45),
	.w4(32'hb99b20d9),
	.w5(32'hb9805969),
	.w6(32'h39aafeb1),
	.w7(32'hbab1d4d3),
	.w8(32'hba450a55),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5ebff),
	.w1(32'hb95a4b26),
	.w2(32'h39b748a1),
	.w3(32'hbace0a52),
	.w4(32'h3a4ba524),
	.w5(32'hba155aae),
	.w6(32'hbb2c265e),
	.w7(32'hb9aabd08),
	.w8(32'hb9a0819f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae12a6e),
	.w1(32'hba3b2b68),
	.w2(32'hb99225ab),
	.w3(32'h3b4eab37),
	.w4(32'hb86e23ae),
	.w5(32'hbb2ebba3),
	.w6(32'h3a91b602),
	.w7(32'h3a9c9537),
	.w8(32'h3a8c040b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59b3ed),
	.w1(32'h3b888955),
	.w2(32'h3bab8dcf),
	.w3(32'h3b66dbcf),
	.w4(32'h3b164bcb),
	.w5(32'h3bfe2682),
	.w6(32'h3bf6402a),
	.w7(32'h3c2588a2),
	.w8(32'h3babec08),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392420de),
	.w1(32'hbb85e0ae),
	.w2(32'hbb413b5b),
	.w3(32'h3974ecd8),
	.w4(32'hbb69f6b3),
	.w5(32'hbb2b10cc),
	.w6(32'hba02c1c7),
	.w7(32'h3a1325b9),
	.w8(32'hbab27d4b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b9da3),
	.w1(32'h3b5c7f74),
	.w2(32'hbb1e1c8c),
	.w3(32'hba89c6e7),
	.w4(32'h3a8dbafe),
	.w5(32'hbae94f54),
	.w6(32'h3b8ab3f4),
	.w7(32'hbab7a5fd),
	.w8(32'hbb3af11c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule