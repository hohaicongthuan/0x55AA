module layer_10_featuremap_61(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3763e),
	.w1(32'hbc0884cc),
	.w2(32'hba9ec5a8),
	.w3(32'hbc1823ed),
	.w4(32'hbbf0770e),
	.w5(32'hb94d1699),
	.w6(32'hbb7db3b9),
	.w7(32'hbc6d13da),
	.w8(32'h3b709e6f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade020d),
	.w1(32'hbacbf239),
	.w2(32'hbbfada05),
	.w3(32'h3ba8a7eb),
	.w4(32'hbb9430f9),
	.w5(32'hbbbc6325),
	.w6(32'h3baf5ceb),
	.w7(32'h39982647),
	.w8(32'hba05bae1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b112b),
	.w1(32'hbbf1bad3),
	.w2(32'h3b186eed),
	.w3(32'h394fcdac),
	.w4(32'hbbe48e5a),
	.w5(32'h3ac1d26d),
	.w6(32'hb97b5951),
	.w7(32'hbc7cbac7),
	.w8(32'hbb3c64af),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f4bc1),
	.w1(32'h3ba4b2d8),
	.w2(32'h3c005149),
	.w3(32'h3b756642),
	.w4(32'hb8e0a5c2),
	.w5(32'h3b45c73c),
	.w6(32'hbb913758),
	.w7(32'h3b47d823),
	.w8(32'h3b31004e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e24d5),
	.w1(32'hba2ed2ec),
	.w2(32'h3c1e57da),
	.w3(32'h3b035f5b),
	.w4(32'h3a497fce),
	.w5(32'h3be1d6bd),
	.w6(32'h3c0e3d10),
	.w7(32'h3b9173b9),
	.w8(32'h3c06f305),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1359a2),
	.w1(32'h3acc81c3),
	.w2(32'h3c32fae0),
	.w3(32'h3bfa7932),
	.w4(32'h3c0fecf9),
	.w5(32'h3c2c0301),
	.w6(32'h3bb4de60),
	.w7(32'h3c04290f),
	.w8(32'hba3582cc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c664559),
	.w1(32'hba32ec8a),
	.w2(32'hbc43b6ea),
	.w3(32'hbaf95ea1),
	.w4(32'hbc49f7b3),
	.w5(32'hbc5a4054),
	.w6(32'hbc4ee40f),
	.w7(32'hbc931b1c),
	.w8(32'h3a462711),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79579f),
	.w1(32'h3a05a5a6),
	.w2(32'h39d9a882),
	.w3(32'hbc35358a),
	.w4(32'hbc54bdbe),
	.w5(32'h3c382de1),
	.w6(32'hbbbca7ed),
	.w7(32'hbb47e882),
	.w8(32'hbbb1d6c7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b2a89),
	.w1(32'hbb6774ae),
	.w2(32'hbbae1299),
	.w3(32'hbbf249d2),
	.w4(32'hbbdb2a4d),
	.w5(32'hbb6cb688),
	.w6(32'hba2b6c22),
	.w7(32'hbb888b50),
	.w8(32'hb9c46fe3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0adae9),
	.w1(32'hbb282c87),
	.w2(32'h3c5fb348),
	.w3(32'hbc0162f9),
	.w4(32'h3b0c88fc),
	.w5(32'h3b9c98f0),
	.w6(32'hba3b5d12),
	.w7(32'h3c2efaf8),
	.w8(32'h3bdabf5e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf242e7),
	.w1(32'h3c2a2be7),
	.w2(32'h3be0fafd),
	.w3(32'hbc2c68ec),
	.w4(32'hbb565103),
	.w5(32'h3bd1a228),
	.w6(32'hbc0713cd),
	.w7(32'hbb3869c4),
	.w8(32'h3c178ab6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec7db2),
	.w1(32'h3ba28931),
	.w2(32'hbd21259f),
	.w3(32'h3b99ec2e),
	.w4(32'h3b82591b),
	.w5(32'hbd102cef),
	.w6(32'h3bfc21bd),
	.w7(32'h3c59ba0d),
	.w8(32'hbcf928ec),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd027268),
	.w1(32'hbce3c7a8),
	.w2(32'hbb701d25),
	.w3(32'hbcdadea8),
	.w4(32'hbca17742),
	.w5(32'hbc0b7e92),
	.w6(32'hbccc9c36),
	.w7(32'hbc9e8a7d),
	.w8(32'hba8cc493),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb349b),
	.w1(32'hbaebb4dc),
	.w2(32'h3c1f04d4),
	.w3(32'hbb934de2),
	.w4(32'h3b93e21b),
	.w5(32'h3bd9c326),
	.w6(32'hbb8137fb),
	.w7(32'hbb331cd7),
	.w8(32'h3c15414f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b043d8a),
	.w1(32'hbb2df098),
	.w2(32'hbb9990b4),
	.w3(32'h3ad6be61),
	.w4(32'hb9f07956),
	.w5(32'hbb831f59),
	.w6(32'h3b860c74),
	.w7(32'h3b58584b),
	.w8(32'hbb9ad6b6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac25239),
	.w1(32'hba8df97d),
	.w2(32'h3c8a5394),
	.w3(32'hbb96bf68),
	.w4(32'h3ab0d7aa),
	.w5(32'h3b8bfcd2),
	.w6(32'hbc147b0d),
	.w7(32'hbb11591e),
	.w8(32'h3ab2420e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b444907),
	.w1(32'h3acaf57b),
	.w2(32'hbb8a5210),
	.w3(32'hbca4627e),
	.w4(32'hbc8c5730),
	.w5(32'hbbac5868),
	.w6(32'hbcb5953d),
	.w7(32'hbc9479d3),
	.w8(32'h3c0d5610),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb29971),
	.w1(32'h3beb8f79),
	.w2(32'h3c2eb86c),
	.w3(32'hbc319a30),
	.w4(32'h3bc68701),
	.w5(32'h3b201690),
	.w6(32'hb90426bc),
	.w7(32'h3c8487d4),
	.w8(32'h3b125e2c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ac91c),
	.w1(32'hba354ad0),
	.w2(32'hba76be3d),
	.w3(32'hbb5e56f7),
	.w4(32'hbc0955cb),
	.w5(32'h39877007),
	.w6(32'hbb4a155b),
	.w7(32'hb8d99027),
	.w8(32'h3abf558d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75a1b8),
	.w1(32'hbb5faadb),
	.w2(32'hbb8c4baa),
	.w3(32'hbae53ab6),
	.w4(32'hbbd96b47),
	.w5(32'hbb91f57a),
	.w6(32'hbb8cd344),
	.w7(32'hba584de1),
	.w8(32'hbab64d69),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b9564),
	.w1(32'h345cfe90),
	.w2(32'hbb815d21),
	.w3(32'hbaac81a7),
	.w4(32'hba4607ba),
	.w5(32'hbb3ffaed),
	.w6(32'h3a411d99),
	.w7(32'h3aff57c1),
	.w8(32'hbbceb21d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a249287),
	.w1(32'h3afa84d2),
	.w2(32'hbbab3b99),
	.w3(32'hbb4aa40d),
	.w4(32'h39c7e21f),
	.w5(32'hbb87f851),
	.w6(32'h3ab4b206),
	.w7(32'h381826c2),
	.w8(32'hbc199de3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97702c),
	.w1(32'h3ab718bd),
	.w2(32'hbbf57f41),
	.w3(32'hbba31f6d),
	.w4(32'hbb907bd1),
	.w5(32'hbc3f0522),
	.w6(32'hbc7eb0e5),
	.w7(32'hbb7e7552),
	.w8(32'hbc52b473),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd69be0),
	.w1(32'hbccde7ea),
	.w2(32'hbb8f57b6),
	.w3(32'hbcdccfe7),
	.w4(32'hbce3d3c0),
	.w5(32'hbb95744a),
	.w6(32'hbcb35f63),
	.w7(32'hbca50358),
	.w8(32'hbb626827),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c5fbc),
	.w1(32'hbc83623f),
	.w2(32'hbbecadb6),
	.w3(32'hbb872802),
	.w4(32'hbc54b99b),
	.w5(32'hbb866381),
	.w6(32'hba9f2946),
	.w7(32'hbb5474ec),
	.w8(32'h3a3559fc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c025800),
	.w1(32'h3b41b58e),
	.w2(32'hbb6eb5c5),
	.w3(32'h3b8318b4),
	.w4(32'hba1453a1),
	.w5(32'hbb8dfbc6),
	.w6(32'hb8c90fe1),
	.w7(32'hbc29de2f),
	.w8(32'hbb319cf7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560820),
	.w1(32'h3b4ea361),
	.w2(32'h3974f381),
	.w3(32'hbbb13ff5),
	.w4(32'hbc02e5bd),
	.w5(32'hba6bd333),
	.w6(32'h3a5bde45),
	.w7(32'hb801a593),
	.w8(32'h39645bf6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c079344),
	.w1(32'h3b7ce819),
	.w2(32'hbc2d15ee),
	.w3(32'h3a20cd6f),
	.w4(32'h3c001eb0),
	.w5(32'hbc59db97),
	.w6(32'h3c5339da),
	.w7(32'h3c62cb44),
	.w8(32'hbbaa6ff3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a1716),
	.w1(32'hbbd8d41e),
	.w2(32'h3b2a3bb2),
	.w3(32'hbc5c97f3),
	.w4(32'hbc150dd4),
	.w5(32'h3b66d1a6),
	.w6(32'hbc839d01),
	.w7(32'hbc2987f8),
	.w8(32'h3c074aec),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35ab6a),
	.w1(32'hbb420383),
	.w2(32'hbb33c9f6),
	.w3(32'h3b51c5e9),
	.w4(32'hbbcfce79),
	.w5(32'hbb0ecc1f),
	.w6(32'h3c460844),
	.w7(32'hbbd5f06f),
	.w8(32'h3c06641c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998003d),
	.w1(32'h3b3795b9),
	.w2(32'hbc42c9c9),
	.w3(32'hbb46272c),
	.w4(32'hbb400250),
	.w5(32'hbb95b937),
	.w6(32'hbb57246f),
	.w7(32'hbb3fc0f2),
	.w8(32'hbbee91ea),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dfe77),
	.w1(32'hbc56c05b),
	.w2(32'hbc5148f4),
	.w3(32'h3b71a072),
	.w4(32'h3a5fc823),
	.w5(32'hbc6e7d5e),
	.w6(32'hbb0da69e),
	.w7(32'hbb76df29),
	.w8(32'hbc37790d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91e73f),
	.w1(32'hbc35ff98),
	.w2(32'hbb2d3767),
	.w3(32'hbcb0a430),
	.w4(32'hbc97b9cc),
	.w5(32'hbaa98e2c),
	.w6(32'h3af65d16),
	.w7(32'h3c076d42),
	.w8(32'h3be25a3f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d4da0),
	.w1(32'h3a1ab1b0),
	.w2(32'h3a97eeda),
	.w3(32'hba321bc6),
	.w4(32'h3b31ccf7),
	.w5(32'h3b8e39bb),
	.w6(32'h3c132814),
	.w7(32'h3bc16d60),
	.w8(32'hbb29fd70),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1caa9c),
	.w1(32'hbb855ef4),
	.w2(32'hbba56d4a),
	.w3(32'h3b841461),
	.w4(32'hbbb57a19),
	.w5(32'hbbd60065),
	.w6(32'hbb6d682a),
	.w7(32'h3aa5e916),
	.w8(32'hbb034393),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c4c2b),
	.w1(32'hbb779268),
	.w2(32'h3c06d258),
	.w3(32'hbbeba05f),
	.w4(32'hba9a5af0),
	.w5(32'h3b8cbd8c),
	.w6(32'hbadd3088),
	.w7(32'h3a7de39e),
	.w8(32'h3bdf1594),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac392b1),
	.w1(32'hba92bce6),
	.w2(32'hbc970328),
	.w3(32'hbc8ad52d),
	.w4(32'hbc59eb43),
	.w5(32'hbc509fa3),
	.w6(32'hbc7f3d74),
	.w7(32'hbc0895e4),
	.w8(32'hbc185965),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc851737),
	.w1(32'hbc7ff6cf),
	.w2(32'hbcee4444),
	.w3(32'hbb61a43d),
	.w4(32'hbc0b3d07),
	.w5(32'hbc8b2188),
	.w6(32'h3c1f124f),
	.w7(32'hba811d6d),
	.w8(32'hbbde5240),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a4847),
	.w1(32'hbc971e59),
	.w2(32'hbbc908a5),
	.w3(32'hbb343e5f),
	.w4(32'hbc51f243),
	.w5(32'h3a43b3c5),
	.w6(32'h3c6cc7a9),
	.w7(32'h3c52d757),
	.w8(32'h3c667979),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73beb9),
	.w1(32'h3aa7d5c6),
	.w2(32'hbb3b09b9),
	.w3(32'hbb31f7a5),
	.w4(32'hbad6e26b),
	.w5(32'h39225847),
	.w6(32'h3bd1c822),
	.w7(32'h3b43e2d3),
	.w8(32'h3b95f293),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bef4a1),
	.w1(32'h3b093342),
	.w2(32'h3ba182b0),
	.w3(32'h3a08d93d),
	.w4(32'h3b3a1d05),
	.w5(32'hbc26607a),
	.w6(32'h3aff2def),
	.w7(32'h3b582f48),
	.w8(32'hbc701ed9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14f7f2),
	.w1(32'hbb535487),
	.w2(32'hbc08069c),
	.w3(32'hbcce5f8f),
	.w4(32'hbc6daeb5),
	.w5(32'hbbee19e4),
	.w6(32'hbc0d1e31),
	.w7(32'hbbc44580),
	.w8(32'hbba6517d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c233d),
	.w1(32'hbc0e7405),
	.w2(32'hbc3528ec),
	.w3(32'hbbee2f1c),
	.w4(32'hbbbad200),
	.w5(32'hbc0d9390),
	.w6(32'hbc73b66d),
	.w7(32'hbc059809),
	.w8(32'hbb3a5d7c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8788de),
	.w1(32'h3a43e6ac),
	.w2(32'h3ba75711),
	.w3(32'hba1f481c),
	.w4(32'h3c554cab),
	.w5(32'hba58e8c7),
	.w6(32'h3c0243b5),
	.w7(32'h3c81442d),
	.w8(32'hbb4e00b6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a38e),
	.w1(32'hbbe41b70),
	.w2(32'hbbb82abf),
	.w3(32'h3b1db6bd),
	.w4(32'hbbb5486a),
	.w5(32'hbc184ed5),
	.w6(32'hbac39a7a),
	.w7(32'hbb6eca2e),
	.w8(32'hbab8a390),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfc71f),
	.w1(32'hbbf0178b),
	.w2(32'h3a7fe210),
	.w3(32'h395fa466),
	.w4(32'hbbca6a6f),
	.w5(32'hbbcba75a),
	.w6(32'hbc009b72),
	.w7(32'hbbfd4dce),
	.w8(32'hbba47530),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f77dc),
	.w1(32'hbc03e1ee),
	.w2(32'h3c091d3f),
	.w3(32'hbc17892b),
	.w4(32'hbc24bff7),
	.w5(32'h3c187181),
	.w6(32'hbc0e91d4),
	.w7(32'hbbdd58c3),
	.w8(32'h3bd0d8a9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7987e),
	.w1(32'h3c95d786),
	.w2(32'h3beb936a),
	.w3(32'h3bd09d1f),
	.w4(32'h3c40e963),
	.w5(32'h3be07f76),
	.w6(32'hbba5b2c1),
	.w7(32'h3c0169ee),
	.w8(32'h3c0ee6e9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d5882),
	.w1(32'hbb2fcf5a),
	.w2(32'hbab66396),
	.w3(32'h3b32800a),
	.w4(32'h3b931989),
	.w5(32'hbb83414d),
	.w6(32'h3b83000a),
	.w7(32'h3be7daa8),
	.w8(32'h3bc40cce),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4cddc),
	.w1(32'hbb30e53a),
	.w2(32'hb9dd5542),
	.w3(32'hbbed20c8),
	.w4(32'hbbfe5d22),
	.w5(32'hbc212c2c),
	.w6(32'hbb8fa0ca),
	.w7(32'hbb85acd4),
	.w8(32'hbb4d9b7d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc542040),
	.w1(32'hbc0db639),
	.w2(32'h3bb4ffe7),
	.w3(32'hbc3e0dd7),
	.w4(32'hbc25ac92),
	.w5(32'h3c23085b),
	.w6(32'hbb695b7f),
	.w7(32'hbb927cf6),
	.w8(32'hbc144dac),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4bfa8),
	.w1(32'hbc83ca94),
	.w2(32'h3a065dac),
	.w3(32'hba44297e),
	.w4(32'hbc8a00e1),
	.w5(32'hbbaaa8d5),
	.w6(32'hbcc01a3d),
	.w7(32'hbca9975e),
	.w8(32'h3b136d81),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba66af2),
	.w1(32'hbb5b35f8),
	.w2(32'h3b1323e0),
	.w3(32'hbb9997f5),
	.w4(32'hbb98ad4e),
	.w5(32'h3be7a6ab),
	.w6(32'h3a6970d9),
	.w7(32'h3bb0c6eb),
	.w8(32'h3b7e522f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12c99f),
	.w1(32'h3c75ddb8),
	.w2(32'h3be12b17),
	.w3(32'h3c74f167),
	.w4(32'h3c476085),
	.w5(32'h3bd12ea2),
	.w6(32'h3b83e332),
	.w7(32'h3b859415),
	.w8(32'h3c0b1161),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6235e4),
	.w1(32'h3c71ecb5),
	.w2(32'hbb28eb6d),
	.w3(32'h3b850626),
	.w4(32'h3be6a440),
	.w5(32'h3afd8867),
	.w6(32'h39a35155),
	.w7(32'h38dd534f),
	.w8(32'hbb3c7caf),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991f025),
	.w1(32'h3ac47b19),
	.w2(32'h3b1e0b96),
	.w3(32'h3adbc430),
	.w4(32'hbaa1e232),
	.w5(32'h3c0825ec),
	.w6(32'h3c3eaef9),
	.w7(32'h3c6f165f),
	.w8(32'h3b34f8e3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c4208),
	.w1(32'hbb57f61a),
	.w2(32'hbbdfdbab),
	.w3(32'hba05614b),
	.w4(32'h39291293),
	.w5(32'hbc6294ed),
	.w6(32'h3a984447),
	.w7(32'h3bf5ead1),
	.w8(32'hbc50a797),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a6abe),
	.w1(32'hbc8654e0),
	.w2(32'hbb1cac37),
	.w3(32'hbca76cd0),
	.w4(32'hbc2751bd),
	.w5(32'hbb047ea2),
	.w6(32'hbc45e8d3),
	.w7(32'h3bfbd809),
	.w8(32'h3b918c60),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba217a),
	.w1(32'h3b836dec),
	.w2(32'hbbd55d9e),
	.w3(32'hbbb72509),
	.w4(32'h3b1eb570),
	.w5(32'hbcabbb35),
	.w6(32'h3ae92f33),
	.w7(32'h3c138fc3),
	.w8(32'hbc7e42af),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39a046),
	.w1(32'hbc1686e2),
	.w2(32'h3c47d889),
	.w3(32'hbcb77f18),
	.w4(32'hbc5d0f4f),
	.w5(32'h3bd619f4),
	.w6(32'hbbc056fe),
	.w7(32'h3b894657),
	.w8(32'hbc1258a6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92c6bf),
	.w1(32'h3c4aaf9c),
	.w2(32'hbc28ddfc),
	.w3(32'h3b9d6d00),
	.w4(32'hbb34fb6f),
	.w5(32'hbc220552),
	.w6(32'hbc8c2ce2),
	.w7(32'hbc9db070),
	.w8(32'h3bd1c37d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43e7a1),
	.w1(32'h3a009632),
	.w2(32'h3bc72eb8),
	.w3(32'h3931f03a),
	.w4(32'h3c3b927d),
	.w5(32'h3a15d92a),
	.w6(32'h3c65b8a4),
	.w7(32'h3c58478a),
	.w8(32'hba828769),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47b05b),
	.w1(32'h3a1bd6bc),
	.w2(32'hbaf49199),
	.w3(32'h3bca1737),
	.w4(32'hbbd5f39c),
	.w5(32'hbbba2636),
	.w6(32'h3b207c57),
	.w7(32'h3b3a627e),
	.w8(32'h3b8f1a00),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20f5b3),
	.w1(32'h3b8d02d0),
	.w2(32'hba30e95d),
	.w3(32'hbb940686),
	.w4(32'hb8cf1551),
	.w5(32'hbb7d1888),
	.w6(32'h3bed419d),
	.w7(32'h3be0f612),
	.w8(32'hba378bf8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba6a6d),
	.w1(32'h3a1b0858),
	.w2(32'hbb155dff),
	.w3(32'hbb61898e),
	.w4(32'hbbfdf66b),
	.w5(32'hb965a267),
	.w6(32'hbc053e95),
	.w7(32'hba99ebb3),
	.w8(32'h3b0e19b0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace267e),
	.w1(32'hb94e45d7),
	.w2(32'hbc2b8adb),
	.w3(32'h3a99166e),
	.w4(32'h3b2b3386),
	.w5(32'hbb9ae468),
	.w6(32'h3b57968b),
	.w7(32'h3b0ed060),
	.w8(32'h3a2c353b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7fbb0),
	.w1(32'h3b9e7350),
	.w2(32'h3b82287a),
	.w3(32'h3bd90738),
	.w4(32'h3c518050),
	.w5(32'hbc114fa0),
	.w6(32'h3cb342f5),
	.w7(32'h3cb2b1f5),
	.w8(32'hba7e6e32),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc063c70),
	.w1(32'hbb018ec0),
	.w2(32'h3be82763),
	.w3(32'hbbdf278d),
	.w4(32'hbb8eb6b7),
	.w5(32'h3c540950),
	.w6(32'hbc6a2d7e),
	.w7(32'h3a705c0e),
	.w8(32'h3aab62fb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7201ad),
	.w1(32'h3c12eb91),
	.w2(32'h3c9820a4),
	.w3(32'h3b7f5fd3),
	.w4(32'h3b19dd20),
	.w5(32'h3c6a564e),
	.w6(32'hbb9cea56),
	.w7(32'hb9f1edd7),
	.w8(32'h3c615dc2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a32e8),
	.w1(32'hbb01884c),
	.w2(32'hbbe34098),
	.w3(32'h3c5602ff),
	.w4(32'hbb29547f),
	.w5(32'h3bcf0ddc),
	.w6(32'h3c7a3491),
	.w7(32'h3b9896fd),
	.w8(32'h3c8b2f68),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50a248),
	.w1(32'h3c67fbf7),
	.w2(32'hbbc4ddcb),
	.w3(32'h3c870198),
	.w4(32'h3c4bf235),
	.w5(32'hbb1421e6),
	.w6(32'h3ba60547),
	.w7(32'hb97c12bb),
	.w8(32'hbb4c7bda),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96a905),
	.w1(32'hbb11baa8),
	.w2(32'hbba96ca8),
	.w3(32'h38e62d01),
	.w4(32'hbb338985),
	.w5(32'hbbb63999),
	.w6(32'hba1e4deb),
	.w7(32'hbb93e2e6),
	.w8(32'hbc1e82d1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd746a4),
	.w1(32'hbb8eb61e),
	.w2(32'hbc2889b7),
	.w3(32'hbc31e0d5),
	.w4(32'h3b546178),
	.w5(32'hbc1b9199),
	.w6(32'hbc0ce0ef),
	.w7(32'h3ab5a9e4),
	.w8(32'h3afa7587),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b7133),
	.w1(32'hbbf8b501),
	.w2(32'h3c2567a1),
	.w3(32'hbc0508c9),
	.w4(32'h3a81d980),
	.w5(32'h3bcbde9f),
	.w6(32'hbac0589b),
	.w7(32'h3b9aec86),
	.w8(32'h3c37c2fa),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb809c31),
	.w1(32'h3b94b67d),
	.w2(32'hbc4db875),
	.w3(32'hbbdbc96e),
	.w4(32'h3b03eda6),
	.w5(32'hbc83cf3f),
	.w6(32'hbb21a8fe),
	.w7(32'h3b751a31),
	.w8(32'hbc250f53),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99c046),
	.w1(32'hbc0e598b),
	.w2(32'h3c36eb76),
	.w3(32'hbc915ebe),
	.w4(32'hbc62558d),
	.w5(32'hbab8f487),
	.w6(32'hbc545fb0),
	.w7(32'hbc1e66cd),
	.w8(32'h38bd398b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37b58c),
	.w1(32'hbb9fc536),
	.w2(32'hbba8358b),
	.w3(32'hbc7f2c54),
	.w4(32'hbb6dd506),
	.w5(32'hbb5f9f60),
	.w6(32'hbc866969),
	.w7(32'h3bb63aa3),
	.w8(32'hbb3e88f8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bad56),
	.w1(32'hbc6e186b),
	.w2(32'h3aa524bc),
	.w3(32'hbc590f5e),
	.w4(32'hbc8aaaad),
	.w5(32'hbb2a1ea1),
	.w6(32'hbc9256b6),
	.w7(32'hbc80c4d8),
	.w8(32'h3b90871a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf39612),
	.w1(32'hbb5f9fca),
	.w2(32'hb9533710),
	.w3(32'h3b0c92e5),
	.w4(32'h3bc0ac18),
	.w5(32'h3b16b61b),
	.w6(32'hbb4e59eb),
	.w7(32'hbb13acea),
	.w8(32'hb97512ad),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0598),
	.w1(32'hbaf70b4a),
	.w2(32'h3c2fc28c),
	.w3(32'h3b91218b),
	.w4(32'hba613f1b),
	.w5(32'h3c829df7),
	.w6(32'h3bb5e921),
	.w7(32'h3b8ae809),
	.w8(32'h3cb38014),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e7dfc),
	.w1(32'h3c56c96e),
	.w2(32'hbab72709),
	.w3(32'h3c8a1aeb),
	.w4(32'h3c6f1d0c),
	.w5(32'hbb81d76e),
	.w6(32'h3c632bca),
	.w7(32'h3c47904a),
	.w8(32'h3a0adcb6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4d98a),
	.w1(32'h3b23acb1),
	.w2(32'h3c512dcf),
	.w3(32'hbc034d27),
	.w4(32'h3a7d19db),
	.w5(32'h3c3f113b),
	.w6(32'hbbe363c1),
	.w7(32'h3b0fcf49),
	.w8(32'h3b30f66d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c38ec),
	.w1(32'hba93ce0a),
	.w2(32'hbba1c7af),
	.w3(32'hbb2f9308),
	.w4(32'hbb84dd92),
	.w5(32'hbbe3a917),
	.w6(32'hbb6529ba),
	.w7(32'h3b963dd6),
	.w8(32'h3b3af5b3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1211c),
	.w1(32'h3a88753e),
	.w2(32'h376c8754),
	.w3(32'hb9ba94d5),
	.w4(32'hbc0c72d9),
	.w5(32'h3b89ad36),
	.w6(32'h3a8d19ab),
	.w7(32'h3b7fb4be),
	.w8(32'hbbce4ef0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc3de),
	.w1(32'h3b00d32d),
	.w2(32'hbc794265),
	.w3(32'hbbf23438),
	.w4(32'hbbacb8fd),
	.w5(32'hbc5e0a76),
	.w6(32'hbbf00b64),
	.w7(32'hbb919f81),
	.w8(32'hbc158c62),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb739940),
	.w1(32'h3b00b466),
	.w2(32'hbbb05a42),
	.w3(32'hbbd7aa66),
	.w4(32'hbb7805d6),
	.w5(32'hbc1f352f),
	.w6(32'hbadb1afb),
	.w7(32'h3c10f787),
	.w8(32'hbbd0d57d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85bc4b),
	.w1(32'hbc23ea59),
	.w2(32'hbbfc3223),
	.w3(32'hbc88bd58),
	.w4(32'hbc03177e),
	.w5(32'hbbfed296),
	.w6(32'hbbea829b),
	.w7(32'hbb6871da),
	.w8(32'hbb90c1e8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8b9d4),
	.w1(32'h3a5ca9d8),
	.w2(32'h3b1b93f5),
	.w3(32'hbb16e0cf),
	.w4(32'hba013b35),
	.w5(32'hba802159),
	.w6(32'h385b2571),
	.w7(32'h3b0a9e4c),
	.w8(32'hbaeb45f4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cdadfc),
	.w1(32'hbb710373),
	.w2(32'hbba93db4),
	.w3(32'hbc2170f6),
	.w4(32'hbc7b8f2e),
	.w5(32'h3bd756ee),
	.w6(32'hbbfd27a6),
	.w7(32'hb7ee425f),
	.w8(32'h3bcfb0f1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b530387),
	.w1(32'h3c6e9083),
	.w2(32'h3c86688e),
	.w3(32'h3ce45c2a),
	.w4(32'h3c78b5a0),
	.w5(32'h3c709cc7),
	.w6(32'h3bccb9f6),
	.w7(32'h3b99bcbb),
	.w8(32'h3c83f3a3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca56685),
	.w1(32'h3c64eb58),
	.w2(32'hbc3eb587),
	.w3(32'h3cb476c0),
	.w4(32'h3c6b7453),
	.w5(32'hbba5eef5),
	.w6(32'h3caf7bbb),
	.w7(32'h3c0e923e),
	.w8(32'hbc8ee577),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21cdae),
	.w1(32'hbbd01767),
	.w2(32'h3bd6e52e),
	.w3(32'hbc1bfb88),
	.w4(32'hbb815e46),
	.w5(32'h3b8bd483),
	.w6(32'hbc684360),
	.w7(32'hbc4b0f33),
	.w8(32'h3c2ca385),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc42d30),
	.w1(32'h3ab2cc77),
	.w2(32'hbb420561),
	.w3(32'h3bf22cf8),
	.w4(32'h3a8e999a),
	.w5(32'hbb36e456),
	.w6(32'h3c4fca42),
	.w7(32'h3bb13edd),
	.w8(32'hbbd36ad8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba111ab),
	.w1(32'h3b77d5ae),
	.w2(32'h3c61bb83),
	.w3(32'h3ab84cc0),
	.w4(32'h3a8f222f),
	.w5(32'h3bc1c478),
	.w6(32'hbb935ce2),
	.w7(32'hbb792982),
	.w8(32'h3ba1d8d1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd92a2e),
	.w1(32'hbbae24e8),
	.w2(32'h3b91a5ad),
	.w3(32'h3aea1a26),
	.w4(32'hbb29c523),
	.w5(32'hbad6d41b),
	.w6(32'h3af88622),
	.w7(32'h3aaa3bb8),
	.w8(32'hbc1568f2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab40dbb),
	.w1(32'hbc14c966),
	.w2(32'h3a593e35),
	.w3(32'h3b7497fb),
	.w4(32'h39ea8e2c),
	.w5(32'hb90e9922),
	.w6(32'h3ba8e4fb),
	.w7(32'h3c316876),
	.w8(32'h3caa8835),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b33c5f),
	.w1(32'h3b2ee09b),
	.w2(32'hbad51e5a),
	.w3(32'hb7573172),
	.w4(32'h3bb5c531),
	.w5(32'hba6e8165),
	.w6(32'h3bee8470),
	.w7(32'h3b5b002b),
	.w8(32'h3ba33ca4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7487e),
	.w1(32'h3b41e92f),
	.w2(32'h3c2dd78f),
	.w3(32'hbbf7eb4a),
	.w4(32'h3af25dd4),
	.w5(32'h3bb115f5),
	.w6(32'h37800f67),
	.w7(32'hba5d4e4f),
	.w8(32'h3c5dcae9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be00724),
	.w1(32'h3ba889d1),
	.w2(32'h3b8d84fe),
	.w3(32'h3c807c7a),
	.w4(32'h3c2cabb4),
	.w5(32'h3c46f69b),
	.w6(32'h3cfb302c),
	.w7(32'h3a2df003),
	.w8(32'h3c5fe665),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f538c),
	.w1(32'h3cab0428),
	.w2(32'h3af1f15e),
	.w3(32'h3b7d1406),
	.w4(32'h3cbef5b2),
	.w5(32'hbbf5d089),
	.w6(32'h3a99d0f9),
	.w7(32'h3c948417),
	.w8(32'hbbe30047),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32f00a),
	.w1(32'hbc839a9c),
	.w2(32'hbc5a1ce0),
	.w3(32'hbb8ff8e3),
	.w4(32'hbb8a3b67),
	.w5(32'hbc5398ae),
	.w6(32'h3b800838),
	.w7(32'h39402a9e),
	.w8(32'hbbdce6fa),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02c4e3),
	.w1(32'hbc706725),
	.w2(32'hbc54dbdd),
	.w3(32'hbc3bc62d),
	.w4(32'hbc8eb5f8),
	.w5(32'hbc858454),
	.w6(32'hbbf9362e),
	.w7(32'hbc80c689),
	.w8(32'hbb7e78bb),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae2add),
	.w1(32'h3ad6e0df),
	.w2(32'h3c61a541),
	.w3(32'hbc8400ac),
	.w4(32'h3b7e40b8),
	.w5(32'h3c7ad5b9),
	.w6(32'hbb25d622),
	.w7(32'h3c03d978),
	.w8(32'h3c83f4f7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8232e0),
	.w1(32'h3c65477d),
	.w2(32'h3a8e3328),
	.w3(32'h3c80bdb6),
	.w4(32'h3c71868e),
	.w5(32'h3c098aa0),
	.w6(32'h3c5e70a9),
	.w7(32'h3b974dce),
	.w8(32'h38a03333),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005204),
	.w1(32'h3bcae010),
	.w2(32'hbc0445e0),
	.w3(32'hbacf9e46),
	.w4(32'hbb829317),
	.w5(32'hbbf155c4),
	.w6(32'hbc033f7f),
	.w7(32'hbc143ca6),
	.w8(32'hbbe60803),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc628108),
	.w1(32'hbbad3c8c),
	.w2(32'hbc77c3a5),
	.w3(32'hbc44b426),
	.w4(32'hbc1c96f9),
	.w5(32'hbc6a6c1d),
	.w6(32'hbadc9d5b),
	.w7(32'hbad2c84a),
	.w8(32'hbb996536),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd4c6d),
	.w1(32'h39644393),
	.w2(32'hbbc5f0cd),
	.w3(32'hbbf5b368),
	.w4(32'h3a556e4d),
	.w5(32'hbb7a147d),
	.w6(32'hbb8e4760),
	.w7(32'h37c89e4b),
	.w8(32'h3a6e31ed),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc970194),
	.w1(32'hbbd15f9c),
	.w2(32'h3b843476),
	.w3(32'hbc82ba14),
	.w4(32'hbb898c8c),
	.w5(32'h3b2eebcb),
	.w6(32'hbba32c8a),
	.w7(32'h3aa65173),
	.w8(32'h3c1eee95),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc168b43),
	.w1(32'hbb5fb489),
	.w2(32'hba81baa0),
	.w3(32'hbb59b816),
	.w4(32'hbc32b331),
	.w5(32'hbbdfdf79),
	.w6(32'hba829d9e),
	.w7(32'h3b3b2647),
	.w8(32'h3b64554d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfef5dd),
	.w1(32'hbc18e11c),
	.w2(32'hbb08fad7),
	.w3(32'hbb9b1508),
	.w4(32'hba820bd7),
	.w5(32'h3a04a2f3),
	.w6(32'h3bb899a8),
	.w7(32'h3ad8f97f),
	.w8(32'h3b8c769c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c144f3d),
	.w1(32'h3bb34e81),
	.w2(32'hb98811a1),
	.w3(32'hbb703bd0),
	.w4(32'hbb28ac23),
	.w5(32'h3b8fd3c1),
	.w6(32'h3a9bb246),
	.w7(32'h3becf085),
	.w8(32'h3be25e4e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978b45b),
	.w1(32'hbbb5d274),
	.w2(32'hbb1577ca),
	.w3(32'h3c4e0508),
	.w4(32'hbb8f8bc9),
	.w5(32'hbc27fb9b),
	.w6(32'h3bc89b03),
	.w7(32'hbb6df51c),
	.w8(32'hbb1ac465),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ebf1d),
	.w1(32'hbbe83e68),
	.w2(32'hbbff5b9d),
	.w3(32'hbc8a00db),
	.w4(32'hbc956ef3),
	.w5(32'hbc202054),
	.w6(32'hbc1f5a36),
	.w7(32'h3b3eab87),
	.w8(32'hbc0f946e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21f97b),
	.w1(32'hbb59e922),
	.w2(32'h3c91e90b),
	.w3(32'hbb25377f),
	.w4(32'h3b7231d2),
	.w5(32'hbb71fffa),
	.w6(32'h3aa97c40),
	.w7(32'hbaf50526),
	.w8(32'hbbbcdf6f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6202a7),
	.w1(32'hbc59f8b3),
	.w2(32'hbc0f98f2),
	.w3(32'hbcd11907),
	.w4(32'hbcefd0e2),
	.w5(32'hbc498893),
	.w6(32'hbce0081b),
	.w7(32'hbcd73041),
	.w8(32'hbc40a261),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83e699),
	.w1(32'hbc4e0c9e),
	.w2(32'h3c3223fb),
	.w3(32'hbc9ed620),
	.w4(32'hbc861b71),
	.w5(32'h3ccb5e6b),
	.w6(32'hbc81231f),
	.w7(32'hbc3aefdc),
	.w8(32'h3c44c3dc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd0bafe),
	.w1(32'h3caefd44),
	.w2(32'hbc50f564),
	.w3(32'h3cffefd2),
	.w4(32'h3c98ee79),
	.w5(32'hbcc48395),
	.w6(32'h3c13bafe),
	.w7(32'hbbc2b8f4),
	.w8(32'hbc3fd3f5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88784d),
	.w1(32'hbc6fa5f2),
	.w2(32'hbc0a911b),
	.w3(32'hbcf3c741),
	.w4(32'hbcc8443f),
	.w5(32'hb9a7364b),
	.w6(32'hbc48cc3c),
	.w7(32'hbbe395e5),
	.w8(32'hbb7d76d5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe48179),
	.w1(32'hbb94858c),
	.w2(32'hbb72a533),
	.w3(32'h3b710f3b),
	.w4(32'h3bad3f4a),
	.w5(32'hbbfa50a8),
	.w6(32'h3c0b151e),
	.w7(32'h3c5d93aa),
	.w8(32'hbb819d1e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee848),
	.w1(32'hbc209699),
	.w2(32'hb9d5c237),
	.w3(32'hbc0448d1),
	.w4(32'hbbcf9015),
	.w5(32'hbbe01fe5),
	.w6(32'hbc2ea957),
	.w7(32'hbc04c534),
	.w8(32'hbbc55a90),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32b78d),
	.w1(32'hbb35b280),
	.w2(32'h3bf9d5ef),
	.w3(32'hbb674b41),
	.w4(32'hb981736f),
	.w5(32'h3bac1fd5),
	.w6(32'hbbdc402d),
	.w7(32'hbba8b477),
	.w8(32'h3af335ce),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13176c),
	.w1(32'h3b231d0d),
	.w2(32'h3b602b66),
	.w3(32'hbb96ab97),
	.w4(32'hbb4397fb),
	.w5(32'hba39f533),
	.w6(32'hbbb32831),
	.w7(32'hbba13bcc),
	.w8(32'h3abf32d3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3937872a),
	.w1(32'hbbc7f330),
	.w2(32'hbc4c7051),
	.w3(32'hbb2808ab),
	.w4(32'hbc181581),
	.w5(32'hbc2e6470),
	.w6(32'hba872d12),
	.w7(32'hbbaa25a5),
	.w8(32'hbb5ba926),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca38e45),
	.w1(32'hbc28c3f2),
	.w2(32'hbc8beff4),
	.w3(32'hbcd56645),
	.w4(32'hbc30f0a1),
	.w5(32'hbcb6adcb),
	.w6(32'hbc0899a9),
	.w7(32'h3adc5160),
	.w8(32'hbc892050),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a528c),
	.w1(32'hbc7871c8),
	.w2(32'hbbf4cbec),
	.w3(32'hbccd61ed),
	.w4(32'hbc8b70a7),
	.w5(32'hbc2d38da),
	.w6(32'hbc7a58d5),
	.w7(32'hbbf09f20),
	.w8(32'hbbab0e12),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1e908),
	.w1(32'hbc51d407),
	.w2(32'hbb9be99e),
	.w3(32'hbc9113e3),
	.w4(32'hbc418700),
	.w5(32'hbc376743),
	.w6(32'hbb25e8bf),
	.w7(32'h3c274540),
	.w8(32'hbc6f5da1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc437730),
	.w1(32'hbb8303ac),
	.w2(32'hbbb1212f),
	.w3(32'hbc777a23),
	.w4(32'hbb3ceec1),
	.w5(32'hbabe4215),
	.w6(32'hbc2c8590),
	.w7(32'h3b423c74),
	.w8(32'hbb92e813),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab5d57),
	.w1(32'hbb8c5965),
	.w2(32'h3c7c573a),
	.w3(32'hbb8d7a8c),
	.w4(32'hbba83e69),
	.w5(32'h3c744ef9),
	.w6(32'hbbaa0068),
	.w7(32'h3b947bbe),
	.w8(32'h3c050289),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa6879),
	.w1(32'h3b714330),
	.w2(32'h3a21a2bd),
	.w3(32'h3ac8c903),
	.w4(32'hba6d5c6b),
	.w5(32'h3b926b5f),
	.w6(32'hbc08824f),
	.w7(32'hbb5d3518),
	.w8(32'h3bcd757e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f33a12),
	.w1(32'h3bac3a23),
	.w2(32'h3b1e0453),
	.w3(32'hbacc0dcb),
	.w4(32'h3ac5fa81),
	.w5(32'hbae270b3),
	.w6(32'h3b95f24b),
	.w7(32'h3bbfd302),
	.w8(32'hbb57eb47),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b76bc),
	.w1(32'h3ac281e2),
	.w2(32'hbbdabcc0),
	.w3(32'h3aff67e9),
	.w4(32'h3bbaa67c),
	.w5(32'hbbc5d48e),
	.w6(32'h3b104045),
	.w7(32'h3c8b6e62),
	.w8(32'hbb893300),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcf801),
	.w1(32'h3ae84f84),
	.w2(32'hbc852721),
	.w3(32'hbc513d6b),
	.w4(32'hbb1cf368),
	.w5(32'hbb0bf9bc),
	.w6(32'hbc183999),
	.w7(32'hbbc4b42d),
	.w8(32'hbb474e66),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb661c41),
	.w1(32'h39c596a3),
	.w2(32'hba640e76),
	.w3(32'h3c382095),
	.w4(32'h3c48effa),
	.w5(32'h3b6d1cd5),
	.w6(32'h3be9d919),
	.w7(32'h3bfe29e7),
	.w8(32'h3b815faa),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96c1b6),
	.w1(32'h3b3aab2f),
	.w2(32'h3bb312c8),
	.w3(32'h3b18eecc),
	.w4(32'h3ad8b208),
	.w5(32'hb8a5832a),
	.w6(32'h3af09dd3),
	.w7(32'h3b3b9ba6),
	.w8(32'h3b0d84bc),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d029f),
	.w1(32'h3b761ac8),
	.w2(32'hbc1f7ca1),
	.w3(32'hbc9330e0),
	.w4(32'hbb2e2154),
	.w5(32'hbbc62651),
	.w6(32'hbc804d55),
	.w7(32'hba7f14b6),
	.w8(32'h3bd7914c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e302a),
	.w1(32'hbc45b836),
	.w2(32'hbb5c625b),
	.w3(32'hbbac155d),
	.w4(32'hbbc6b5e5),
	.w5(32'hba976892),
	.w6(32'h3c16bf42),
	.w7(32'hba17ebea),
	.w8(32'h3bc004ab),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e1505),
	.w1(32'h3c338121),
	.w2(32'h3bdaa919),
	.w3(32'h3c5585ae),
	.w4(32'h3b9bfc65),
	.w5(32'h3c26bba3),
	.w6(32'h3c6d4a68),
	.w7(32'h3c176641),
	.w8(32'h3b0681cd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc53642),
	.w1(32'h3c73e892),
	.w2(32'h3b1c2ef9),
	.w3(32'h3c0d42c5),
	.w4(32'h3c1753b6),
	.w5(32'h3ab73a8c),
	.w6(32'hbc02130d),
	.w7(32'hbbfb06aa),
	.w8(32'hba4e4701),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982b6a5),
	.w1(32'hbae6af45),
	.w2(32'h3aeca5ee),
	.w3(32'hbba6394b),
	.w4(32'hbc0f27fb),
	.w5(32'hbc0c074c),
	.w6(32'hbc215562),
	.w7(32'hbc3f07f8),
	.w8(32'hbb9f168b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d7be8),
	.w1(32'h3985ba01),
	.w2(32'h3c0ce82b),
	.w3(32'hbbd5e9ce),
	.w4(32'h3aa6f11c),
	.w5(32'h3c055eec),
	.w6(32'hbb9b6708),
	.w7(32'h3a978a81),
	.w8(32'h3bab5731),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9887f6),
	.w1(32'h3b75b14c),
	.w2(32'h3ba97894),
	.w3(32'h3b03b38a),
	.w4(32'h3a701ccd),
	.w5(32'h3c2aff64),
	.w6(32'hbb2aa69b),
	.w7(32'hbbb1b1b1),
	.w8(32'hba363477),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30ba3e),
	.w1(32'h3ad4f687),
	.w2(32'hbb13b36f),
	.w3(32'h3c868781),
	.w4(32'h3baff2ea),
	.w5(32'hbc0911e6),
	.w6(32'h3c8e5e59),
	.w7(32'hba3bab3e),
	.w8(32'hbb904a63),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acde8b),
	.w1(32'hba984626),
	.w2(32'hb9ac5ebb),
	.w3(32'hbb8e20f2),
	.w4(32'hbbc7281c),
	.w5(32'hbc17d269),
	.w6(32'hbbf68acf),
	.w7(32'hbc24d4fb),
	.w8(32'hba832702),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb754),
	.w1(32'hbbb443a5),
	.w2(32'hbab857f5),
	.w3(32'hbc779ef2),
	.w4(32'hbc5036a3),
	.w5(32'hbab1380e),
	.w6(32'hbbbcf50d),
	.w7(32'hba58bbe3),
	.w8(32'hbb94d26e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef5d97),
	.w1(32'hbb60d7ce),
	.w2(32'h3c7129b1),
	.w3(32'hbb4252f5),
	.w4(32'hbbcbc710),
	.w5(32'h3cc3744c),
	.w6(32'hbbbb3035),
	.w7(32'hbbe7a28e),
	.w8(32'h3c5ffd5e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5f4a8),
	.w1(32'h3c8c0b87),
	.w2(32'h3ba1d1ac),
	.w3(32'h3d0cb474),
	.w4(32'h3cd5d0ab),
	.w5(32'h3b744995),
	.w6(32'h3cc49262),
	.w7(32'h3c155072),
	.w8(32'h3b6afe2a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbf02f),
	.w1(32'h3b6b9d24),
	.w2(32'hbc7691df),
	.w3(32'h3c03f396),
	.w4(32'hba9a6ee5),
	.w5(32'hbc48fd4b),
	.w6(32'h3b771a7a),
	.w7(32'hbbd045e2),
	.w8(32'hbb8fef24),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc885b89),
	.w1(32'hbbd377ba),
	.w2(32'h3b6d8d54),
	.w3(32'hbc5247ef),
	.w4(32'h3b227759),
	.w5(32'h3c057d40),
	.w6(32'hb9dcf53c),
	.w7(32'h3bba3bc6),
	.w8(32'h3c216903),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf502de),
	.w1(32'h3bc505b3),
	.w2(32'h3b28e96f),
	.w3(32'h3c39c1eb),
	.w4(32'h3bb25c8a),
	.w5(32'h3a841bdc),
	.w6(32'h3bf54973),
	.w7(32'h3b8ed719),
	.w8(32'h3bb04003),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd4405),
	.w1(32'hbaa4e648),
	.w2(32'hbc2ad4cf),
	.w3(32'hbab6971b),
	.w4(32'hbb4d35b9),
	.w5(32'hbc493440),
	.w6(32'h3b06645e),
	.w7(32'h39a2bf1c),
	.w8(32'h3bafae0d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eaeb7),
	.w1(32'hbb9f1e5e),
	.w2(32'h39d2d493),
	.w3(32'hbb4791d8),
	.w4(32'h3967bba3),
	.w5(32'hbac4e49d),
	.w6(32'h3b72c8ee),
	.w7(32'hbb817fdf),
	.w8(32'hba9180a5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b8718),
	.w1(32'h3b84430a),
	.w2(32'h3ba7e404),
	.w3(32'hbc34e84a),
	.w4(32'hb9aef650),
	.w5(32'h3c3833b6),
	.w6(32'hbc1a60b6),
	.w7(32'hbbecdce5),
	.w8(32'h3bbfd567),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9add9a),
	.w1(32'h3bae8d73),
	.w2(32'hbc097c16),
	.w3(32'h3c57bc81),
	.w4(32'h3a336acd),
	.w5(32'hbb25f985),
	.w6(32'h3c8f22e7),
	.w7(32'h3b44d13b),
	.w8(32'hbb6107e5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc3a9b),
	.w1(32'h3a90d1b2),
	.w2(32'h3bbcdcde),
	.w3(32'h3bf04b8e),
	.w4(32'h3bfb7e99),
	.w5(32'hbb431827),
	.w6(32'h39c22b74),
	.w7(32'hbb69cced),
	.w8(32'hbc04d9ee),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94544a),
	.w1(32'hbbdbb22a),
	.w2(32'hb91300a2),
	.w3(32'hbc1d5e44),
	.w4(32'hbc108d24),
	.w5(32'hb9682d87),
	.w6(32'hbbe0c3f6),
	.w7(32'hb9f2ecb2),
	.w8(32'hb9ae20a1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f4ade),
	.w1(32'hba5b2e23),
	.w2(32'h3c1c135c),
	.w3(32'h3a8e3450),
	.w4(32'hba4198e5),
	.w5(32'h3c582e4f),
	.w6(32'h3abc1661),
	.w7(32'hbaa31628),
	.w8(32'h3c462e0a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9975bf),
	.w1(32'h3bb0d0b2),
	.w2(32'h3c293422),
	.w3(32'h3cc00542),
	.w4(32'h3c69fa9e),
	.w5(32'h3bd8439e),
	.w6(32'h3c75310b),
	.w7(32'h3c0eeabc),
	.w8(32'h3a412c83),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510d69),
	.w1(32'hbaec3d46),
	.w2(32'hba8db90e),
	.w3(32'h3c2539ad),
	.w4(32'h3b1d7c9f),
	.w5(32'hbb1cac5a),
	.w6(32'hb900d058),
	.w7(32'h3bab47f5),
	.w8(32'hbb8e9546),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac25374),
	.w1(32'hba24255d),
	.w2(32'hba3fc869),
	.w3(32'hbac6f4c2),
	.w4(32'hbae6e5ae),
	.w5(32'h3a3bf8c1),
	.w6(32'hbb26b79e),
	.w7(32'hbaced29c),
	.w8(32'hbb976041),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd13143),
	.w1(32'hbc1b9f96),
	.w2(32'h3b354c79),
	.w3(32'hbacb05c9),
	.w4(32'hbbd47eb5),
	.w5(32'h3b41107b),
	.w6(32'h3b3cc8b8),
	.w7(32'h3b8aa682),
	.w8(32'hba4440a1),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5408fd),
	.w1(32'hbc3b5b75),
	.w2(32'h3b3e43ca),
	.w3(32'h3b173696),
	.w4(32'hbbbb6e9e),
	.w5(32'h3af45821),
	.w6(32'hba96671e),
	.w7(32'h3c0ea2e2),
	.w8(32'h3b23e141),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe64b9d),
	.w1(32'hbc68533b),
	.w2(32'hbae64787),
	.w3(32'hbb6d8b02),
	.w4(32'hbc37d80e),
	.w5(32'hbbc06e73),
	.w6(32'h3a80002e),
	.w7(32'hbb3e7d64),
	.w8(32'h3a9de3a5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c14e1),
	.w1(32'hb8c5a901),
	.w2(32'hbb807c2f),
	.w3(32'hbb188d7c),
	.w4(32'hbc6f0ee7),
	.w5(32'hbae2ee99),
	.w6(32'hbb854bd4),
	.w7(32'hbb9d019d),
	.w8(32'hba875aed),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddebb1),
	.w1(32'hbb82815c),
	.w2(32'hbc27e9cb),
	.w3(32'hba8cee6f),
	.w4(32'hbb160c94),
	.w5(32'h3afea271),
	.w6(32'hba1f9098),
	.w7(32'hb9c9d60e),
	.w8(32'h3b8ac614),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c7fb6),
	.w1(32'hbc97724f),
	.w2(32'hbb2f558a),
	.w3(32'h3b0073a5),
	.w4(32'hbc3b0350),
	.w5(32'hbac3af3a),
	.w6(32'h3be25e8f),
	.w7(32'h3c2e219d),
	.w8(32'h3b6ddc7e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d65e),
	.w1(32'hbc96daef),
	.w2(32'hbb1fb4c8),
	.w3(32'hbb6a8fdc),
	.w4(32'hbc243cc0),
	.w5(32'hbbdaeda5),
	.w6(32'h38e7bcd1),
	.w7(32'hbb56ecfd),
	.w8(32'hbbaa7280),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a133119),
	.w1(32'hbbdac2e5),
	.w2(32'hbbdc802a),
	.w3(32'hbc172841),
	.w4(32'hbb83219c),
	.w5(32'hbbe5b229),
	.w6(32'hbc05846b),
	.w7(32'hbbf814f7),
	.w8(32'hbc1958a7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b553e47),
	.w1(32'h3bb8f4f3),
	.w2(32'hba5db1c4),
	.w3(32'hbb8a05a6),
	.w4(32'h3b14a7ab),
	.w5(32'hba2b7cea),
	.w6(32'hba98a01e),
	.w7(32'hb97d7781),
	.w8(32'hbb5cecdd),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8f770),
	.w1(32'h38e24392),
	.w2(32'h3baa2a0b),
	.w3(32'hbab97a11),
	.w4(32'hbb3b2bcd),
	.w5(32'h3b949f19),
	.w6(32'hbc2a1be0),
	.w7(32'h3a8a7d15),
	.w8(32'h3aa84d04),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbd01c),
	.w1(32'hbbc8e282),
	.w2(32'hbbec4e73),
	.w3(32'h3b5442a1),
	.w4(32'hbbc7b1ab),
	.w5(32'hbb8ca8c9),
	.w6(32'h38c8e7a9),
	.w7(32'h3b84d76a),
	.w8(32'hbb5aae2c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc029ad3),
	.w1(32'hbbe6db1c),
	.w2(32'hbbe23de2),
	.w3(32'hbad7bab0),
	.w4(32'hbb8c525c),
	.w5(32'hbb7b57e7),
	.w6(32'hbb851d58),
	.w7(32'hba3b1832),
	.w8(32'hb97665d9),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91c533),
	.w1(32'hbaa9d73f),
	.w2(32'h3ac58888),
	.w3(32'hbaad469c),
	.w4(32'h3b3c6247),
	.w5(32'hbb43354f),
	.w6(32'h3a4802f0),
	.w7(32'h3aef6d6b),
	.w8(32'hbb2c32de),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be217c8),
	.w1(32'h3b3357b8),
	.w2(32'h3c4ff33f),
	.w3(32'hbbc4b51f),
	.w4(32'h3bd5f93b),
	.w5(32'h39c57306),
	.w6(32'hb8fc6aa8),
	.w7(32'h3b7bd40d),
	.w8(32'h3b39c973),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe51d6b),
	.w1(32'hba384d87),
	.w2(32'h3bf8bebf),
	.w3(32'hba9d5d9e),
	.w4(32'hb940dc36),
	.w5(32'h3aac0048),
	.w6(32'hbadda73f),
	.w7(32'hba891029),
	.w8(32'h3a5d1b14),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dbf68),
	.w1(32'h3c0a240e),
	.w2(32'hbb1916d9),
	.w3(32'h3b17bbda),
	.w4(32'h3b908f61),
	.w5(32'hbb1a7497),
	.w6(32'h3b517f9c),
	.w7(32'h3ad8357a),
	.w8(32'hbb3c9b97),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb621f6e),
	.w1(32'hbbd07cfc),
	.w2(32'hbaaa49e8),
	.w3(32'hbb5e17d4),
	.w4(32'hbaf1f769),
	.w5(32'h39df2a0c),
	.w6(32'h3971b199),
	.w7(32'h3b329d0e),
	.w8(32'h3ac35cfc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a476819),
	.w1(32'hbae37aca),
	.w2(32'h3a817c2b),
	.w3(32'h3ae60af3),
	.w4(32'h3b20159a),
	.w5(32'hbaefefda),
	.w6(32'h3b8020fb),
	.w7(32'h3ae213ba),
	.w8(32'h3ac23f44),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9f5a1),
	.w1(32'hba861630),
	.w2(32'h3aab27e9),
	.w3(32'hbb367284),
	.w4(32'h3ae8ad90),
	.w5(32'h3a87ec34),
	.w6(32'h39149762),
	.w7(32'hbb998fc1),
	.w8(32'hbb696fe5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1695d5),
	.w1(32'hbb896b25),
	.w2(32'hb9f5e0b7),
	.w3(32'hb9de3ad7),
	.w4(32'hbbff59de),
	.w5(32'h3a200806),
	.w6(32'hbb9eaecb),
	.w7(32'h3aa532f6),
	.w8(32'hbb4089d3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038102),
	.w1(32'hbc27bd41),
	.w2(32'h3924a08c),
	.w3(32'h39f07191),
	.w4(32'hbad327f9),
	.w5(32'hbb93209c),
	.w6(32'h3a3f420a),
	.w7(32'hb9e27ed5),
	.w8(32'h390db141),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de07f3),
	.w1(32'hbc50d08f),
	.w2(32'h3c9be2b0),
	.w3(32'hbbc49fbf),
	.w4(32'hbb54a6b6),
	.w5(32'h3c13eb79),
	.w6(32'hbbcfaae6),
	.w7(32'hba763838),
	.w8(32'hbb467eca),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6bc24),
	.w1(32'hbbd3ba3d),
	.w2(32'hbc08df96),
	.w3(32'h3c224adf),
	.w4(32'h3bed2b0a),
	.w5(32'hbbaefd48),
	.w6(32'h3b448357),
	.w7(32'h3bd97518),
	.w8(32'hbaff1cf0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3c63),
	.w1(32'hbb43ee7e),
	.w2(32'hbb134ddb),
	.w3(32'hbc4d30c8),
	.w4(32'h3a21a5c4),
	.w5(32'hbb305d5a),
	.w6(32'hbb808224),
	.w7(32'hbba85b0d),
	.w8(32'hba9b655b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877b69),
	.w1(32'hbabdec87),
	.w2(32'h3c8d522a),
	.w3(32'hbbd03240),
	.w4(32'hbbf72a9f),
	.w5(32'h3c2fcf70),
	.w6(32'hbb79ceb4),
	.w7(32'hbb061275),
	.w8(32'h3c08e3f0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55f9fb),
	.w1(32'hbc0bc346),
	.w2(32'h3c611b37),
	.w3(32'h3c4ac4e6),
	.w4(32'h3bc69b99),
	.w5(32'h3be764a6),
	.w6(32'h3c4d1ce8),
	.w7(32'h3c4be0dd),
	.w8(32'h3aec50df),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd632a7),
	.w1(32'h3c73d878),
	.w2(32'hba6bb9d0),
	.w3(32'h3c1ee91f),
	.w4(32'h3c6d1160),
	.w5(32'hb8ee8d79),
	.w6(32'h3b3aaef9),
	.w7(32'h3c2ab849),
	.w8(32'hbb8d57ff),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4716f),
	.w1(32'hbb127ece),
	.w2(32'hba63d2f1),
	.w3(32'h3b1939d8),
	.w4(32'hbaeda5c7),
	.w5(32'hbbc8eac3),
	.w6(32'hbb48fdcf),
	.w7(32'hbb893abd),
	.w8(32'hbc10ee7a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0ff68),
	.w1(32'hbb56bd45),
	.w2(32'h3b7527d8),
	.w3(32'hbc66d473),
	.w4(32'hbb5fcf10),
	.w5(32'h3b87df0d),
	.w6(32'hbc17e213),
	.w7(32'h3b73bfd7),
	.w8(32'h3c59ecc8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfba30),
	.w1(32'h3be9381b),
	.w2(32'h3ae66f13),
	.w3(32'h3ab310f4),
	.w4(32'h3b9fd6e8),
	.w5(32'hbb5597b7),
	.w6(32'h3c1a2b89),
	.w7(32'h3b8344ad),
	.w8(32'h3a3c33d5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a4de2),
	.w1(32'h3b287e5c),
	.w2(32'hbb65240b),
	.w3(32'hbac1706f),
	.w4(32'h3ba4fc24),
	.w5(32'hbbe0e4b0),
	.w6(32'hbbdb6892),
	.w7(32'h3bc163f2),
	.w8(32'hbb63d846),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca50d6),
	.w1(32'hbb708259),
	.w2(32'hbb9474fb),
	.w3(32'hbbf37ab3),
	.w4(32'hbc13f01a),
	.w5(32'hbb1fda1b),
	.w6(32'hbbf16e0d),
	.w7(32'hbbd834f3),
	.w8(32'hbbcaaaf9),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d6e6f),
	.w1(32'hbb8ae1a4),
	.w2(32'hb8524cbb),
	.w3(32'hbb4f111e),
	.w4(32'hbb8717cc),
	.w5(32'hba9bc0ae),
	.w6(32'hbad389cf),
	.w7(32'h3a946ce0),
	.w8(32'h37eebdad),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e62fa),
	.w1(32'h3af00545),
	.w2(32'h3bfc2781),
	.w3(32'hbbc9bf14),
	.w4(32'hbbdb6e66),
	.w5(32'h3c148b6d),
	.w6(32'h3a8f4a8c),
	.w7(32'h39c5da3d),
	.w8(32'h3bab7e37),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb624),
	.w1(32'h3a52c362),
	.w2(32'h3ad9ee2c),
	.w3(32'h3c0bb8f8),
	.w4(32'h3b95aba5),
	.w5(32'h3a58fccc),
	.w6(32'h3c0590f0),
	.w7(32'h3c26e06d),
	.w8(32'h3b6795a3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ad50e),
	.w1(32'h3a42e3a6),
	.w2(32'h3ba4003e),
	.w3(32'hb862ede3),
	.w4(32'h3bab3420),
	.w5(32'hbba6f821),
	.w6(32'hbb215bf2),
	.w7(32'h3b93037f),
	.w8(32'h3b121379),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd28903),
	.w1(32'hbc04baf4),
	.w2(32'hbc30e62b),
	.w3(32'hbba04421),
	.w4(32'hbc1f592c),
	.w5(32'hbb9a91e7),
	.w6(32'hbad19346),
	.w7(32'h3af7309c),
	.w8(32'hbbfd7194),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf70e8f),
	.w1(32'hbb997544),
	.w2(32'h3a96acf7),
	.w3(32'hbb732c74),
	.w4(32'hbb807064),
	.w5(32'h3ad2a236),
	.w6(32'hbbe43c98),
	.w7(32'h3a95156f),
	.w8(32'h399e6de6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4dac1),
	.w1(32'h3b02826a),
	.w2(32'hbb32a59b),
	.w3(32'h39e8f0aa),
	.w4(32'h3b2b3e43),
	.w5(32'hbbc11c00),
	.w6(32'hba3e8435),
	.w7(32'h3b5b24e0),
	.w8(32'hbbd19259),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc895c4),
	.w1(32'h3c254c33),
	.w2(32'h3adebed1),
	.w3(32'hbc20dfcc),
	.w4(32'h3b3015fb),
	.w5(32'h3ac0f71d),
	.w6(32'hbb88cf1b),
	.w7(32'h3bfcf613),
	.w8(32'hbb1668c9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be76652),
	.w1(32'h39da3133),
	.w2(32'hbb5f5df2),
	.w3(32'h3c08feb5),
	.w4(32'h3b9479fc),
	.w5(32'hbacada43),
	.w6(32'h3b13ff8a),
	.w7(32'h3b84b1fb),
	.w8(32'h3aea445d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39c488),
	.w1(32'hbbe6e140),
	.w2(32'h3b21ffdb),
	.w3(32'h3b8f9053),
	.w4(32'hbaf5f83a),
	.w5(32'h3b39102e),
	.w6(32'h3b076987),
	.w7(32'hba200bfc),
	.w8(32'h3aa4eb36),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954e9b3),
	.w1(32'h3bb021ac),
	.w2(32'hbae552f5),
	.w3(32'hba86559b),
	.w4(32'h3bc2b493),
	.w5(32'hbb812f0c),
	.w6(32'h3a3f18bc),
	.w7(32'h3bb7a983),
	.w8(32'hbbff5442),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade0da2),
	.w1(32'hb9bfeee3),
	.w2(32'h3a734e11),
	.w3(32'hba5418cf),
	.w4(32'hba46156f),
	.w5(32'hbaf795f6),
	.w6(32'hbbca1c97),
	.w7(32'hbab7866f),
	.w8(32'h39b78caf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c17d8d),
	.w1(32'hbb8af42e),
	.w2(32'hbb912c37),
	.w3(32'hba58ae77),
	.w4(32'hbab76854),
	.w5(32'hbac2a69a),
	.w6(32'h3ac067c3),
	.w7(32'h3ac5f099),
	.w8(32'hbb57c73e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91e55e),
	.w1(32'hbc1ea423),
	.w2(32'hbb0a5cef),
	.w3(32'h396c4d7b),
	.w4(32'hbb92cd42),
	.w5(32'hbb4a4828),
	.w6(32'hbba00c78),
	.w7(32'hbb0fd8c5),
	.w8(32'hbc123f43),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f5243),
	.w1(32'hbbd692f6),
	.w2(32'h3b340e45),
	.w3(32'hbb190a75),
	.w4(32'hbbe19924),
	.w5(32'hb95de78b),
	.w6(32'hbb4ce085),
	.w7(32'hbbcab2bf),
	.w8(32'h3ab977fa),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75c00d),
	.w1(32'h3a049536),
	.w2(32'hbb777517),
	.w3(32'h3c4906be),
	.w4(32'h3c044a98),
	.w5(32'hbb5c575b),
	.w6(32'h3ba533fc),
	.w7(32'h3b35dca7),
	.w8(32'hbb01df6e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ce5e9),
	.w1(32'hb970a778),
	.w2(32'hbb3dab51),
	.w3(32'hbb6ee3f1),
	.w4(32'h3a1f6246),
	.w5(32'hbbb5d991),
	.w6(32'hbb8652c8),
	.w7(32'hbaae6886),
	.w8(32'hbb97d16f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3ee89),
	.w1(32'hbbada3d9),
	.w2(32'hbb1cd26c),
	.w3(32'hbc56afa5),
	.w4(32'hbba9cdc9),
	.w5(32'hbb02a1ca),
	.w6(32'hbc0c670d),
	.w7(32'h3b0dcd9d),
	.w8(32'hbaca4cd1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32110b),
	.w1(32'hbbe6304d),
	.w2(32'hbaed5ee1),
	.w3(32'hbba1c55e),
	.w4(32'hbbeae10b),
	.w5(32'hb6cf7e07),
	.w6(32'hbb9da218),
	.w7(32'hbbcfdb1f),
	.w8(32'h3c0c9238),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f44e),
	.w1(32'hbbd0af48),
	.w2(32'hbc8e0814),
	.w3(32'h3c483002),
	.w4(32'h3aa70f9a),
	.w5(32'hbcb09b37),
	.w6(32'h3c363747),
	.w7(32'h3b8f3a49),
	.w8(32'hbc971f17),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31ed88),
	.w1(32'hbc55f7a3),
	.w2(32'h3ac6fc7f),
	.w3(32'hbc75e789),
	.w4(32'hbc7c922f),
	.w5(32'hba9cf2eb),
	.w6(32'hbcc92e1c),
	.w7(32'hbc1ca9d6),
	.w8(32'hbb688099),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6a49a),
	.w1(32'hbbf87117),
	.w2(32'hba4f89d8),
	.w3(32'hbb75df9a),
	.w4(32'hbb984641),
	.w5(32'hbbcd0273),
	.w6(32'hbb6d9af3),
	.w7(32'hbc1d5b27),
	.w8(32'hbb8ef176),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50798e),
	.w1(32'hbcb68276),
	.w2(32'h3bbba5e4),
	.w3(32'hbc4052df),
	.w4(32'hbcb7373e),
	.w5(32'h3ba7ca92),
	.w6(32'hbbdb95a4),
	.w7(32'hbc4b5caf),
	.w8(32'h3b5040ae),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce4328),
	.w1(32'h39d53e04),
	.w2(32'hbade8f94),
	.w3(32'h3c4f6dbb),
	.w4(32'h3b8d3756),
	.w5(32'hbb883ca0),
	.w6(32'h3ca2c609),
	.w7(32'h3c89b9a3),
	.w8(32'h3ab6fed6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c572b),
	.w1(32'h3b2473b8),
	.w2(32'h3b737bcb),
	.w3(32'h395e18ba),
	.w4(32'h3b3ef866),
	.w5(32'h3ac7f170),
	.w6(32'hbb41eb4c),
	.w7(32'h3ac0db28),
	.w8(32'h3aef7945),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ee9d1),
	.w1(32'hbaae1f58),
	.w2(32'h3b7faffb),
	.w3(32'hbba1e452),
	.w4(32'hbbd7cce8),
	.w5(32'hbaf4609e),
	.w6(32'hbb24f46c),
	.w7(32'hb9306223),
	.w8(32'hba961e0f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb001f1c),
	.w1(32'h376f483c),
	.w2(32'h3c3e0edc),
	.w3(32'hbb1ad791),
	.w4(32'hbb7fb9b9),
	.w5(32'h3ca9923b),
	.w6(32'hbb6ce986),
	.w7(32'h3a69bdea),
	.w8(32'h3cac7ba4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf91386),
	.w1(32'h3bfaf986),
	.w2(32'h3a639f42),
	.w3(32'h3c668db8),
	.w4(32'h3cc17ad0),
	.w5(32'h3bd6adc6),
	.w6(32'h3c839a99),
	.w7(32'h3cb7e115),
	.w8(32'h3c4369d9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f84a3),
	.w1(32'h3bde4028),
	.w2(32'h3b8e0420),
	.w3(32'hbb2d7e44),
	.w4(32'h3bdf6734),
	.w5(32'h3bc9f04d),
	.w6(32'hbb375c18),
	.w7(32'h3893f7f2),
	.w8(32'h3b46131a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad62f51),
	.w1(32'hbb5377d5),
	.w2(32'hbbd87e90),
	.w3(32'h3b424178),
	.w4(32'h397e59a9),
	.w5(32'hbbe6d921),
	.w6(32'h3b2f438f),
	.w7(32'h3b0e981a),
	.w8(32'hbbab2a90),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b477494),
	.w1(32'h3b34dd47),
	.w2(32'hbc1d89db),
	.w3(32'hba784024),
	.w4(32'h38cab284),
	.w5(32'hbc1ee277),
	.w6(32'hba883477),
	.w7(32'hbb09fecb),
	.w8(32'hbb385243),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadad9f1),
	.w1(32'hba2c5ebe),
	.w2(32'h3be9ea6c),
	.w3(32'hbb19313d),
	.w4(32'hba3725d5),
	.w5(32'hbb8e7133),
	.w6(32'hbb8dec54),
	.w7(32'hb91046fc),
	.w8(32'h3a52dad0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f0d91),
	.w1(32'hbbdbfda7),
	.w2(32'hbb507d9c),
	.w3(32'hbbe4cfdc),
	.w4(32'hbc273dfa),
	.w5(32'h392d708a),
	.w6(32'hb9da3b38),
	.w7(32'h3972663e),
	.w8(32'hba9f6a2d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992dd29),
	.w1(32'hbb592883),
	.w2(32'h3b7add5c),
	.w3(32'h3a04f2f4),
	.w4(32'hbaaab150),
	.w5(32'hbbad90cb),
	.w6(32'hb9f6bf0a),
	.w7(32'hba73b7d6),
	.w8(32'hbafa1034),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d7517),
	.w1(32'h3b501974),
	.w2(32'hbba30e53),
	.w3(32'h39b65032),
	.w4(32'hbad88f15),
	.w5(32'h3b644327),
	.w6(32'hbc2bd912),
	.w7(32'hba04dfc4),
	.w8(32'hba15b417),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb125ffa),
	.w1(32'hbc25adbd),
	.w2(32'hbbc373f8),
	.w3(32'h3b2a7483),
	.w4(32'hbbafb70f),
	.w5(32'hbb90dd59),
	.w6(32'h3b19cd52),
	.w7(32'h3b20d55d),
	.w8(32'h3735c1dc),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc652876),
	.w1(32'hbac5698c),
	.w2(32'h3bb7aefa),
	.w3(32'hbc7ed252),
	.w4(32'hbb88ac80),
	.w5(32'h3afdef0b),
	.w6(32'hbc89f89c),
	.w7(32'hbbd8e617),
	.w8(32'hb9ea43f2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc284f6f),
	.w1(32'hbc483a45),
	.w2(32'hbba873f7),
	.w3(32'hbb1dab40),
	.w4(32'hb9ffa980),
	.w5(32'hbb81e36c),
	.w6(32'hbb4d79e6),
	.w7(32'hbb8e1c5c),
	.w8(32'hbb8b9f08),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34ee89),
	.w1(32'hbc8093b8),
	.w2(32'hbb23f482),
	.w3(32'hbbeb0724),
	.w4(32'hbb6bcdfd),
	.w5(32'hbb39059a),
	.w6(32'hbab29907),
	.w7(32'hb7a87a62),
	.w8(32'hbb34475c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cbc29),
	.w1(32'h3acb027f),
	.w2(32'hba531836),
	.w3(32'hbbba1d59),
	.w4(32'h3ac41b52),
	.w5(32'hbb803d56),
	.w6(32'hbbf4cbc3),
	.w7(32'h3b9e3d8b),
	.w8(32'hbbbd2725),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56d9c8),
	.w1(32'hbc233e5d),
	.w2(32'hbb605002),
	.w3(32'hbc113e83),
	.w4(32'hbbb01a3d),
	.w5(32'hbb4a272e),
	.w6(32'hbc0c4e6c),
	.w7(32'hbb818210),
	.w8(32'h3b2e6117),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae504b3),
	.w1(32'hbb471905),
	.w2(32'hbac54669),
	.w3(32'hbbc0914f),
	.w4(32'hbbc46ea8),
	.w5(32'hbb9983e2),
	.w6(32'h3b40436e),
	.w7(32'hbb368db9),
	.w8(32'hbbc22dd7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bd7ed),
	.w1(32'h3b2452a6),
	.w2(32'h3c08d28e),
	.w3(32'h3b6616cf),
	.w4(32'h3bcf7d3f),
	.w5(32'h3bda4516),
	.w6(32'hbb21db32),
	.w7(32'h3b8d414c),
	.w8(32'h3a4735e2),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c601649),
	.w1(32'h3b9355db),
	.w2(32'h396c1b70),
	.w3(32'h3c500971),
	.w4(32'h3c2688b1),
	.w5(32'hbba15dce),
	.w6(32'h3bc2d7e6),
	.w7(32'h3c1e153a),
	.w8(32'hbbce45a5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2fb05),
	.w1(32'h3b97fb0b),
	.w2(32'hba01d974),
	.w3(32'hbbd80252),
	.w4(32'h3b02dd6b),
	.w5(32'hbb43999b),
	.w6(32'hbc124ab6),
	.w7(32'hba69f208),
	.w8(32'hbb96f481),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42779e),
	.w1(32'hbc05b6c0),
	.w2(32'h39d84bda),
	.w3(32'hbae13944),
	.w4(32'h374ef3ef),
	.w5(32'hbb0b6cd0),
	.w6(32'hba998274),
	.w7(32'hba9a367c),
	.w8(32'hbba935a5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa337f7),
	.w1(32'hbbb7e32e),
	.w2(32'h38d8495a),
	.w3(32'hbb8ad402),
	.w4(32'h3badac1d),
	.w5(32'hbbd325eb),
	.w6(32'hbba13986),
	.w7(32'hbb593b80),
	.w8(32'hbc122c4c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7bb58),
	.w1(32'hbbb42923),
	.w2(32'hbba8dc5c),
	.w3(32'hbbb1999b),
	.w4(32'hbbd47bd3),
	.w5(32'hbc36afa1),
	.w6(32'hbbfab0bf),
	.w7(32'h3ad4598b),
	.w8(32'hbbaa59a8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ff62c),
	.w1(32'hbc36f34f),
	.w2(32'h3b1312f9),
	.w3(32'hb883d582),
	.w4(32'hbb58f885),
	.w5(32'h3b327b95),
	.w6(32'h3c0ef55a),
	.w7(32'h3befa476),
	.w8(32'h3bfb5c77),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b635e9e),
	.w1(32'h3c10236f),
	.w2(32'h3bdc391e),
	.w3(32'hbab3475e),
	.w4(32'h3ac79b1b),
	.w5(32'hbb090512),
	.w6(32'hbbc0e186),
	.w7(32'hb8b8ac1c),
	.w8(32'hbc36121d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6d3bd),
	.w1(32'hbb0248cf),
	.w2(32'h3aea7e8d),
	.w3(32'hba7359a0),
	.w4(32'h39383b8e),
	.w5(32'h3a171c16),
	.w6(32'hbb92e9e2),
	.w7(32'h3bd5a102),
	.w8(32'h3bcf6984),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc032b9f),
	.w1(32'hbbebaa1d),
	.w2(32'hbba0ea8e),
	.w3(32'hbae6664f),
	.w4(32'hbc2da32d),
	.w5(32'hbbe35451),
	.w6(32'h38feb8a9),
	.w7(32'hbb5ac99e),
	.w8(32'hbbc6201a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe92ae0),
	.w1(32'hbb61cf17),
	.w2(32'h3c3048ff),
	.w3(32'hbc07c871),
	.w4(32'hbb8bb913),
	.w5(32'h3bcca4ef),
	.w6(32'hbbef7e0d),
	.w7(32'hbb085118),
	.w8(32'hbb9173f0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f72d1),
	.w1(32'h3c920d26),
	.w2(32'hbbecf5b9),
	.w3(32'h3c5f8c45),
	.w4(32'h3cbad9ca),
	.w5(32'hbc046f7d),
	.w6(32'h3bcceaae),
	.w7(32'h3c41886f),
	.w8(32'hbc5605af),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0513a2),
	.w1(32'hbc376f74),
	.w2(32'hbb8689d6),
	.w3(32'hbc1a97ef),
	.w4(32'hbc1a3950),
	.w5(32'hbb5b71ec),
	.w6(32'hbc32f74c),
	.w7(32'hbbdc1392),
	.w8(32'hbbc5e4d5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe614c4),
	.w1(32'h3aecc776),
	.w2(32'hba38ceb3),
	.w3(32'h3b524510),
	.w4(32'hbb8fef91),
	.w5(32'h3bf0c395),
	.w6(32'hb9787b0b),
	.w7(32'h3b902c04),
	.w8(32'h3b489679),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce8be4),
	.w1(32'hbbec0ea7),
	.w2(32'hbb84ac58),
	.w3(32'h3a851d6c),
	.w4(32'hbb925ff8),
	.w5(32'h39f981d6),
	.w6(32'h3b15cb61),
	.w7(32'h3b970f98),
	.w8(32'hbbd87212),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82928a),
	.w1(32'hbb8c8203),
	.w2(32'h3b39ed1d),
	.w3(32'hbb03e081),
	.w4(32'hbb85d1a4),
	.w5(32'h3b12dfed),
	.w6(32'hbbc805f2),
	.w7(32'hbc1ca15b),
	.w8(32'h39a86553),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70d3fd),
	.w1(32'h3aef61f9),
	.w2(32'h3ad75d3e),
	.w3(32'h3b8eb2a4),
	.w4(32'h3b402fe2),
	.w5(32'hb9ee77e6),
	.w6(32'h3b9a8e8c),
	.w7(32'h3b35a8f2),
	.w8(32'hbb8ca36b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b322615),
	.w1(32'h3b8ba75d),
	.w2(32'hbc147a55),
	.w3(32'h3b05714b),
	.w4(32'h3ac7f00a),
	.w5(32'hbc0396fa),
	.w6(32'hbb0820d0),
	.w7(32'h3b21e8a4),
	.w8(32'hbc2b3f57),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7c0ef),
	.w1(32'hba6a674c),
	.w2(32'h3b97a20a),
	.w3(32'hb9996265),
	.w4(32'h3bf3a01a),
	.w5(32'h3b8fa7c9),
	.w6(32'hbb70f590),
	.w7(32'h3bd670ee),
	.w8(32'h3ad2c23d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09ea61),
	.w1(32'hba377123),
	.w2(32'hbbd1ac88),
	.w3(32'h3b77efe1),
	.w4(32'h3b036099),
	.w5(32'hbbc8d28e),
	.w6(32'h3a3a6911),
	.w7(32'h3b35479e),
	.w8(32'hba998890),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea365),
	.w1(32'h3a89b44e),
	.w2(32'h3bd16f25),
	.w3(32'h3b1801e8),
	.w4(32'h3ba389a9),
	.w5(32'h3c034313),
	.w6(32'h3bc558d2),
	.w7(32'h3b11f494),
	.w8(32'h3c3758fd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5e84d),
	.w1(32'hbbfe39a7),
	.w2(32'hbb716e7f),
	.w3(32'hbba7b4bc),
	.w4(32'hbc17ef9a),
	.w5(32'h3b14719e),
	.w6(32'hbacc1b56),
	.w7(32'h38e26260),
	.w8(32'h3bbc946b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32f343),
	.w1(32'hbc48615d),
	.w2(32'h3b0edcd7),
	.w3(32'h39e3be44),
	.w4(32'hbc36009d),
	.w5(32'hbb427bb6),
	.w6(32'hbae65a8b),
	.w7(32'hbc74969e),
	.w8(32'hbc5572df),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule