module layer_10_featuremap_164(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff8de5),
	.w1(32'hbc991a18),
	.w2(32'hbc99ff32),
	.w3(32'h3b171670),
	.w4(32'h3c16ec79),
	.w5(32'hbb4aa20b),
	.w6(32'hbca8e9d4),
	.w7(32'hbceea067),
	.w8(32'hbbbe179c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc8660c),
	.w1(32'hbc02696a),
	.w2(32'hbb9900a5),
	.w3(32'hbbfbc756),
	.w4(32'hb983e942),
	.w5(32'h3ac74438),
	.w6(32'h3b45536e),
	.w7(32'h3aa9d005),
	.w8(32'h39d8cfcf),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a821a08),
	.w1(32'hbadc28b4),
	.w2(32'h39193462),
	.w3(32'h390abdc0),
	.w4(32'hba69c685),
	.w5(32'hbb97ff10),
	.w6(32'hba71b381),
	.w7(32'hba40df4c),
	.w8(32'h38ba567b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb001795),
	.w1(32'hbb2e0c9a),
	.w2(32'h3ae94162),
	.w3(32'hba95e915),
	.w4(32'hbbba55b6),
	.w5(32'hb9cdd7af),
	.w6(32'h3b921120),
	.w7(32'h3b1cd616),
	.w8(32'hbc1a7f40),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60ecdd),
	.w1(32'h3b2dfefc),
	.w2(32'hbbb5626a),
	.w3(32'hbb0db500),
	.w4(32'hbb982113),
	.w5(32'hbb73c5e9),
	.w6(32'h3c46fd16),
	.w7(32'h3b98bb43),
	.w8(32'hbc2c898d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd75d7),
	.w1(32'hbaf42bbc),
	.w2(32'hbab4d6a7),
	.w3(32'h3c4df6cd),
	.w4(32'h3b65dd8e),
	.w5(32'h3bf0d78e),
	.w6(32'hbbe708e2),
	.w7(32'hbc39d3fc),
	.w8(32'hbbffda44),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5e665),
	.w1(32'h3c46ce3d),
	.w2(32'h3b4eba20),
	.w3(32'h3a9678d8),
	.w4(32'h3bec154d),
	.w5(32'h3b966bc9),
	.w6(32'h3a907b60),
	.w7(32'h3bc1ed0d),
	.w8(32'hbaaa268a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0099fb),
	.w1(32'h3cea7207),
	.w2(32'h3c11aa29),
	.w3(32'hbc2ad644),
	.w4(32'h3b0b0fcb),
	.w5(32'hbab1d4c5),
	.w6(32'hbb6a7799),
	.w7(32'hbaee7e99),
	.w8(32'hbc374df8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dad47),
	.w1(32'h3a7e0f93),
	.w2(32'h3b3f5017),
	.w3(32'hb9359d80),
	.w4(32'h3a4b8fd6),
	.w5(32'h3b136645),
	.w6(32'hba84036e),
	.w7(32'h37bf9348),
	.w8(32'hba56c540),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c046f47),
	.w1(32'h3c054e0f),
	.w2(32'h3beea9ed),
	.w3(32'h3b35f190),
	.w4(32'h3c2461b2),
	.w5(32'h3c3928e0),
	.w6(32'hbbde0b9a),
	.w7(32'h3a6406dc),
	.w8(32'h3bc290a9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00bf24),
	.w1(32'hbcac6a72),
	.w2(32'hbca7a57a),
	.w3(32'h3be4a091),
	.w4(32'hbc6cd8ae),
	.w5(32'hbc845eab),
	.w6(32'hbc38b101),
	.w7(32'hbc4f886c),
	.w8(32'hbc6c90fa),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce09099),
	.w1(32'h3c9d49e6),
	.w2(32'h3c6281c3),
	.w3(32'hbcd2913d),
	.w4(32'h3c84b065),
	.w5(32'h3ca793d3),
	.w6(32'h3b469bc3),
	.w7(32'h3c41fb15),
	.w8(32'h3c11e90b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc964fc),
	.w1(32'h3bf8f2c9),
	.w2(32'h3aeb9f60),
	.w3(32'h3c37888c),
	.w4(32'hba613292),
	.w5(32'hbb9afebd),
	.w6(32'hbbd975e7),
	.w7(32'hbbd572fc),
	.w8(32'hbbab8359),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59bf87),
	.w1(32'h3bd27987),
	.w2(32'hbad02b0b),
	.w3(32'h3a7d8a4c),
	.w4(32'h3aaa3e2b),
	.w5(32'hbc7b70b5),
	.w6(32'h3c6d13e9),
	.w7(32'h3cac62e4),
	.w8(32'h3c71fb9a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc45e4),
	.w1(32'h3b29cfa9),
	.w2(32'h3c9f82f2),
	.w3(32'hbc5330d4),
	.w4(32'h39e1edc1),
	.w5(32'h3c9579e9),
	.w6(32'h3c395c29),
	.w7(32'h3c1f5036),
	.w8(32'hbbe30d2d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4cc4e),
	.w1(32'h3bc5c1c3),
	.w2(32'h3b173b2d),
	.w3(32'h3c8b8387),
	.w4(32'h3bd3bd54),
	.w5(32'h3b9287aa),
	.w6(32'h3a4b3fb3),
	.w7(32'h3b016aeb),
	.w8(32'hbacd53fc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad032f6),
	.w1(32'h3aa38eff),
	.w2(32'h3a871b40),
	.w3(32'hba99b81d),
	.w4(32'h3a5a8ff2),
	.w5(32'h3b1a7790),
	.w6(32'hbb8b11e2),
	.w7(32'hbb4a7da9),
	.w8(32'hbbde322e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7411e),
	.w1(32'h3c9f2594),
	.w2(32'hb89ffd9c),
	.w3(32'hba257c53),
	.w4(32'h3b94ae17),
	.w5(32'hbbbeec2f),
	.w6(32'hbc4826f7),
	.w7(32'hbc1aac71),
	.w8(32'hbc3104cd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8ebf6),
	.w1(32'h3c07a956),
	.w2(32'h3b34bc00),
	.w3(32'hbb43eb8b),
	.w4(32'h3afe0048),
	.w5(32'hbb901665),
	.w6(32'hbbd140c9),
	.w7(32'hbbde610b),
	.w8(32'hbbd9384f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefefc3),
	.w1(32'h39f1bdc1),
	.w2(32'hb8e1f18f),
	.w3(32'hbb1b0d20),
	.w4(32'hb97a7da1),
	.w5(32'h3a88fc02),
	.w6(32'hbb0019b1),
	.w7(32'hbb39b5dc),
	.w8(32'hbb715d4d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6e100),
	.w1(32'hbb234a52),
	.w2(32'hbb845bd1),
	.w3(32'hbb994116),
	.w4(32'h3aa119cb),
	.w5(32'h3b0cfb66),
	.w6(32'h39c843ef),
	.w7(32'h3b5558cb),
	.w8(32'h3a77b2c7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcba7e1),
	.w1(32'hbbf1a881),
	.w2(32'h39e47f5f),
	.w3(32'h3a627d5b),
	.w4(32'hbb23ab8d),
	.w5(32'hbc74054f),
	.w6(32'hbabc67fa),
	.w7(32'hbc105c3c),
	.w8(32'h37a4a1d7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c140009),
	.w1(32'h3c86e8a9),
	.w2(32'h3c4c8840),
	.w3(32'h3b445739),
	.w4(32'h3c82c733),
	.w5(32'h3bb8ce41),
	.w6(32'hba24afb7),
	.w7(32'hbbc8b336),
	.w8(32'hbc294572),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da2271),
	.w1(32'hb94742cf),
	.w2(32'hbaf46c32),
	.w3(32'h3b617e92),
	.w4(32'hbb87ed59),
	.w5(32'hbba971ff),
	.w6(32'hbb21ba60),
	.w7(32'hb91798ce),
	.w8(32'hba7c908b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3542ef),
	.w1(32'hbc844ccd),
	.w2(32'hbbdb0832),
	.w3(32'hbbf9bb02),
	.w4(32'hbc021d7a),
	.w5(32'hbabd178e),
	.w6(32'h3a5eb85e),
	.w7(32'hbbf49429),
	.w8(32'hba01a56e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2030bf),
	.w1(32'h3b9af4fe),
	.w2(32'h3cc810c5),
	.w3(32'h3adb5be1),
	.w4(32'h3c4ad82a),
	.w5(32'h3c75849b),
	.w6(32'h3b8c501b),
	.w7(32'h3c61ee26),
	.w8(32'h3c1de8fa),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0e852),
	.w1(32'hb9ceeb0b),
	.w2(32'h39cd1f25),
	.w3(32'h3bc26b52),
	.w4(32'hba10c2fd),
	.w5(32'h38c1039a),
	.w6(32'hba207245),
	.w7(32'hba444baa),
	.w8(32'hbb3dee6f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b7eb6),
	.w1(32'hbb5d1d54),
	.w2(32'h3c22f781),
	.w3(32'h3c7339ad),
	.w4(32'h3c7343f0),
	.w5(32'h3c4aaf44),
	.w6(32'hbc70d7d2),
	.w7(32'h3a24d634),
	.w8(32'h3c9db62f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf23b5d),
	.w1(32'h3aa3f58b),
	.w2(32'hbbc9a300),
	.w3(32'hbbaad6da),
	.w4(32'h3c16950a),
	.w5(32'h3bcb844b),
	.w6(32'h3aecf222),
	.w7(32'hbb541262),
	.w8(32'hbbb3b56a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73c8bc),
	.w1(32'hbc7ea4a4),
	.w2(32'hbbde387d),
	.w3(32'h3b864833),
	.w4(32'h3b3f5b32),
	.w5(32'h3be6a3ae),
	.w6(32'h3b25ff24),
	.w7(32'h3c263583),
	.w8(32'h3c08504f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c1b7e),
	.w1(32'hba0ff24b),
	.w2(32'hbb2c0547),
	.w3(32'h3b5622c7),
	.w4(32'hba394b47),
	.w5(32'hba8a9827),
	.w6(32'h398b7ba9),
	.w7(32'h3b0745dd),
	.w8(32'h3aa0364d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb2192),
	.w1(32'hb786b963),
	.w2(32'hb9c91504),
	.w3(32'hbad7e6d6),
	.w4(32'hb8404587),
	.w5(32'h39ee7558),
	.w6(32'hba9f8184),
	.w7(32'hbac77dfc),
	.w8(32'hbac7338c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d02920),
	.w1(32'h3af80af8),
	.w2(32'h3a9b7248),
	.w3(32'hb961b095),
	.w4(32'h3a922069),
	.w5(32'h3a3e02bc),
	.w6(32'hbc3252f8),
	.w7(32'hbc2a6838),
	.w8(32'hbb86286c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9a40),
	.w1(32'hba42e1af),
	.w2(32'h3c375caa),
	.w3(32'hbc591e0d),
	.w4(32'hbc445f32),
	.w5(32'h3bc5b264),
	.w6(32'h3bfdd173),
	.w7(32'hbb872bab),
	.w8(32'hbc51dc7e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16d32e),
	.w1(32'h3ab78306),
	.w2(32'h3b316848),
	.w3(32'h3bc7195b),
	.w4(32'h3bd27566),
	.w5(32'h3c390a86),
	.w6(32'hbb601eba),
	.w7(32'hbabf77de),
	.w8(32'h3a6d474c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a8a9e),
	.w1(32'h3bc8cf74),
	.w2(32'h3b9f591e),
	.w3(32'h3b7dacfc),
	.w4(32'hba7e49df),
	.w5(32'hb9dac6e5),
	.w6(32'hbc058e5d),
	.w7(32'hbbef1b36),
	.w8(32'hbbd0f3fa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfda097),
	.w1(32'h3c464cc7),
	.w2(32'h3c7bc303),
	.w3(32'hbcc3a00b),
	.w4(32'h3b9d31bc),
	.w5(32'h3c5891a1),
	.w6(32'h3a19a3a6),
	.w7(32'h3b6bf19d),
	.w8(32'hbab47f2e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90250a),
	.w1(32'hbc8a59af),
	.w2(32'hbc6d5de5),
	.w3(32'h3c16ecf8),
	.w4(32'hbb265d4b),
	.w5(32'hbc532914),
	.w6(32'h3c8c7080),
	.w7(32'h3caa1466),
	.w8(32'h3b8d39b8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c63bf),
	.w1(32'hbc597eea),
	.w2(32'hbbe264f5),
	.w3(32'h3b111435),
	.w4(32'h3b86b1ca),
	.w5(32'hbaf07eb2),
	.w6(32'h3c0780ba),
	.w7(32'h3c71e9aa),
	.w8(32'h3c490da2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ca925),
	.w1(32'h3b011851),
	.w2(32'h3b452558),
	.w3(32'h3a74a333),
	.w4(32'h3aaf51a1),
	.w5(32'h3aa80038),
	.w6(32'h3b94d72a),
	.w7(32'h3b88c36c),
	.w8(32'hba2bcadf),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af919e9),
	.w1(32'h3b62d321),
	.w2(32'hbb5f7768),
	.w3(32'hba84c076),
	.w4(32'h3bc061f7),
	.w5(32'h3b227ff8),
	.w6(32'hbae50841),
	.w7(32'hbb8bf509),
	.w8(32'hbbb7454d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e44b4),
	.w1(32'hbbe7d9af),
	.w2(32'hbc016f8c),
	.w3(32'h3b121931),
	.w4(32'hbc2641e9),
	.w5(32'hbc039cd0),
	.w6(32'hbaf5f6bb),
	.w7(32'hbb8a1b61),
	.w8(32'hbb9c2929),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe786c4),
	.w1(32'h3a3af85b),
	.w2(32'hb9d6de1b),
	.w3(32'hbc47fe85),
	.w4(32'hba1ebdb4),
	.w5(32'hbaf32649),
	.w6(32'hbb8db7f0),
	.w7(32'hbb439a2c),
	.w8(32'hbb8ee51a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9f7a0),
	.w1(32'h3c2921c4),
	.w2(32'h3bfa98cf),
	.w3(32'h3c31ad79),
	.w4(32'h3b5faa1a),
	.w5(32'h3bae184f),
	.w6(32'hbc2863a9),
	.w7(32'hbc1dbaff),
	.w8(32'hbbcedcb8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45b223),
	.w1(32'hbc9d8f06),
	.w2(32'hbc187c6f),
	.w3(32'h3a146157),
	.w4(32'hbcb9c808),
	.w5(32'hbcf1b93f),
	.w6(32'hbab06877),
	.w7(32'hbac43348),
	.w8(32'h3bc0e9f8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc725a28),
	.w1(32'hbc2c52a5),
	.w2(32'hbc49cfab),
	.w3(32'hbcfee51e),
	.w4(32'hbca39562),
	.w5(32'hbcd4dc3a),
	.w6(32'hba73fe83),
	.w7(32'hbc03e556),
	.w8(32'hbc4c2b53),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc269c0b),
	.w1(32'h3b549c92),
	.w2(32'h3bfbb1b2),
	.w3(32'hbc2a1bad),
	.w4(32'h3c3142ca),
	.w5(32'h3c7d86a7),
	.w6(32'h3be0a3d8),
	.w7(32'h3cb2b373),
	.w8(32'h3c5b3597),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd278ce),
	.w1(32'h3cbe8cf7),
	.w2(32'h3b8720ff),
	.w3(32'h3bdff991),
	.w4(32'h3b983b70),
	.w5(32'h38f10b6a),
	.w6(32'hbc8ca220),
	.w7(32'hbc8af6fb),
	.w8(32'hbc9bd5e3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fe94b),
	.w1(32'hba874ba1),
	.w2(32'hb9ff8d54),
	.w3(32'hba5117bb),
	.w4(32'h380a02e1),
	.w5(32'h39bed7f3),
	.w6(32'hbb9be150),
	.w7(32'hbbc1fb67),
	.w8(32'hbbb86c49),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46d617),
	.w1(32'h3b7c63f5),
	.w2(32'h3a999c9a),
	.w3(32'hbb1504a2),
	.w4(32'hbb1f1643),
	.w5(32'hbbda1e59),
	.w6(32'h3be21b94),
	.w7(32'h3c02f5d5),
	.w8(32'h3b604e8c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae653d),
	.w1(32'h3be08ebd),
	.w2(32'h3bd0b138),
	.w3(32'hbb537c05),
	.w4(32'hba94db15),
	.w5(32'hbbd67b0d),
	.w6(32'h3c1d2194),
	.w7(32'h3c85f1eb),
	.w8(32'h3bf7d7e6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcbb4e),
	.w1(32'h3bc30ef2),
	.w2(32'h3c202739),
	.w3(32'hbb14a19b),
	.w4(32'h3bf0fc26),
	.w5(32'h3cc8b577),
	.w6(32'hbc6cf3cf),
	.w7(32'hbc337134),
	.w8(32'h3c84b852),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca28d14),
	.w1(32'h3b4c9399),
	.w2(32'hba9c67a8),
	.w3(32'h3aa1ffb6),
	.w4(32'h3bc7b9ae),
	.w5(32'h3c00d0aa),
	.w6(32'hbbade3ac),
	.w7(32'hbc0a665a),
	.w8(32'hbb8769b8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca451a5),
	.w1(32'h3c873ac2),
	.w2(32'hbb6b5a49),
	.w3(32'h3c0f24dd),
	.w4(32'h3c1f90a3),
	.w5(32'hbb20b923),
	.w6(32'hbbc9e1bf),
	.w7(32'hbc97027d),
	.w8(32'hbcddcb59),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80d757),
	.w1(32'h3a8a5c32),
	.w2(32'hbb2bce4f),
	.w3(32'h3bf9bddc),
	.w4(32'h3a8e3b42),
	.w5(32'h3a04fc10),
	.w6(32'hbb3d28e0),
	.w7(32'hbbb259a6),
	.w8(32'hbaee48f4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2de79),
	.w1(32'hbb9e939a),
	.w2(32'hbc1d8fb6),
	.w3(32'hba9c46b4),
	.w4(32'h3b9e9330),
	.w5(32'hbbe77257),
	.w6(32'hbb5f7f0f),
	.w7(32'hbbdd1833),
	.w8(32'hbb80d686),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb280d),
	.w1(32'hbb119956),
	.w2(32'hbb48e49f),
	.w3(32'hbb0e9e48),
	.w4(32'hbb77349b),
	.w5(32'hbb882300),
	.w6(32'h3b9f822c),
	.w7(32'h3bc0cc2f),
	.w8(32'h3bb8dead),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b057ac8),
	.w1(32'h3a83db32),
	.w2(32'hbbc02b8f),
	.w3(32'h3a1e209f),
	.w4(32'hbc1f1de5),
	.w5(32'hbc34a052),
	.w6(32'h3c2dbf28),
	.w7(32'h3bfac189),
	.w8(32'hbc38b150),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb21826),
	.w1(32'h3a87f1e5),
	.w2(32'hb79f9e4f),
	.w3(32'h3c0b3e95),
	.w4(32'h398da3cb),
	.w5(32'h3ad424fb),
	.w6(32'hba3fbf49),
	.w7(32'hbb630772),
	.w8(32'hbaf385bb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b578f51),
	.w1(32'h3b874e35),
	.w2(32'h3b1b41f5),
	.w3(32'h3aadd751),
	.w4(32'h3b73bae2),
	.w5(32'hb8e4f9a0),
	.w6(32'h3af43715),
	.w7(32'h3b189a86),
	.w8(32'hba5a3695),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7d489),
	.w1(32'h3b94901e),
	.w2(32'h3a14603d),
	.w3(32'h3aad0c16),
	.w4(32'h3aa7609f),
	.w5(32'hbb006812),
	.w6(32'hbaa8806e),
	.w7(32'hbb6f2033),
	.w8(32'hbb08bece),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fd28e),
	.w1(32'hbb89a358),
	.w2(32'hbb7be150),
	.w3(32'h3bbaa6fd),
	.w4(32'hbaf840d0),
	.w5(32'hbbd5297c),
	.w6(32'hba880b4c),
	.w7(32'hbaac9953),
	.w8(32'h39a043d6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf74806),
	.w1(32'hbb0a2ada),
	.w2(32'h3a2e8007),
	.w3(32'hbc123e1c),
	.w4(32'hbb0e8d28),
	.w5(32'hbb91c6a8),
	.w6(32'h3abef2b3),
	.w7(32'hbbc253d0),
	.w8(32'hbb6073c5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82c4e4),
	.w1(32'hbaf388bc),
	.w2(32'h3a54910f),
	.w3(32'hbc1fb6eb),
	.w4(32'hbaf119c5),
	.w5(32'h3b5d3057),
	.w6(32'hbb853b1a),
	.w7(32'hbbb633ea),
	.w8(32'hbb39cefe),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24cfba),
	.w1(32'hbbd11b48),
	.w2(32'hb8b4d8a9),
	.w3(32'h3b215c61),
	.w4(32'hbbafc9db),
	.w5(32'hbb590419),
	.w6(32'hbbf6da13),
	.w7(32'hbbd6e418),
	.w8(32'hbbb5b9a1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1968c),
	.w1(32'hbb82799c),
	.w2(32'hbc00a078),
	.w3(32'hbb9c55d6),
	.w4(32'hbc4911a5),
	.w5(32'hbc536782),
	.w6(32'hba711fbc),
	.w7(32'h3a6173ac),
	.w8(32'hbc39c793),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca44623),
	.w1(32'h3c84a0f6),
	.w2(32'hbc4f3bdb),
	.w3(32'h3c794079),
	.w4(32'h3ce3fec2),
	.w5(32'h3b9c285b),
	.w6(32'hbba17317),
	.w7(32'h3be99c48),
	.w8(32'h3c077c92),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fdfac),
	.w1(32'h3c0afdeb),
	.w2(32'h3a4d2485),
	.w3(32'hba8f54ef),
	.w4(32'h3b190d6f),
	.w5(32'h3b6036b2),
	.w6(32'hbb13689a),
	.w7(32'hbc89c142),
	.w8(32'hbcc8823c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedfa9b),
	.w1(32'h3c0e18cf),
	.w2(32'h3b8cd508),
	.w3(32'h3bdc8ff2),
	.w4(32'h3a3b637d),
	.w5(32'h3ba8b6b3),
	.w6(32'hb9370f8b),
	.w7(32'hbb8a547d),
	.w8(32'hbb8c7263),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca552c),
	.w1(32'hbcc514ec),
	.w2(32'hbc4b0c9e),
	.w3(32'hbb4b3bb8),
	.w4(32'hbce80984),
	.w5(32'hbd00f743),
	.w6(32'h3cc4e76c),
	.w7(32'h3d019530),
	.w8(32'h3b378096),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3a519),
	.w1(32'hbb33c3ea),
	.w2(32'hbb1beb3a),
	.w3(32'hbb94bd3a),
	.w4(32'hbb8fcd1b),
	.w5(32'hbb1f10c9),
	.w6(32'hbb8f59b2),
	.w7(32'hbbaeb30d),
	.w8(32'hbb988b82),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb348198),
	.w1(32'hbb4720df),
	.w2(32'hbb1bfe51),
	.w3(32'hbb3bd7d5),
	.w4(32'hbbbcfa89),
	.w5(32'hbb4a1d3e),
	.w6(32'h39d4d716),
	.w7(32'h3ade8262),
	.w8(32'hbb6da306),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba414678),
	.w1(32'h3b78a9b9),
	.w2(32'h3b747e17),
	.w3(32'hba4cd7da),
	.w4(32'h3b242912),
	.w5(32'h3a7eb42a),
	.w6(32'h3a628346),
	.w7(32'h3adbae28),
	.w8(32'h3811c222),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd50c8b),
	.w1(32'h3b57b741),
	.w2(32'h3a50ad45),
	.w3(32'h3a67ba67),
	.w4(32'h3b026fcd),
	.w5(32'hba8aba38),
	.w6(32'hbbc1b59d),
	.w7(32'hbc05be61),
	.w8(32'hbc0776c4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4beb04),
	.w1(32'h3a6dbb76),
	.w2(32'h39e7ca9f),
	.w3(32'hbaf3da47),
	.w4(32'h3938cfe5),
	.w5(32'h3b75668c),
	.w6(32'hbbd72fc2),
	.w7(32'hbc1186d4),
	.w8(32'hbb08ce58),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32be76),
	.w1(32'h3c0ab053),
	.w2(32'h3c6290c5),
	.w3(32'hbab5f853),
	.w4(32'h3af81b1a),
	.w5(32'h3c78538d),
	.w6(32'hbc5ae5e0),
	.w7(32'hbb6afd3d),
	.w8(32'h3bb22852),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34ef37),
	.w1(32'h3c8b4fcf),
	.w2(32'h3bdc1c85),
	.w3(32'hbc8a7147),
	.w4(32'h3ad373e3),
	.w5(32'hbb93a42e),
	.w6(32'hbb5b6699),
	.w7(32'h3b5e10f2),
	.w8(32'hbb9084e8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f82dc),
	.w1(32'hbc21463a),
	.w2(32'hbb504733),
	.w3(32'hb99aa976),
	.w4(32'hbbc9cb4d),
	.w5(32'hbbf1fa96),
	.w6(32'h3ba567eb),
	.w7(32'h3b659f3f),
	.w8(32'h3b9d0052),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb141cf),
	.w1(32'h3b7283ca),
	.w2(32'h3c1ec98b),
	.w3(32'hbbd3eb9b),
	.w4(32'h3bb49156),
	.w5(32'h3be37486),
	.w6(32'hbc3d15ed),
	.w7(32'hbbaac37e),
	.w8(32'hba8a8bd4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbdc16),
	.w1(32'h3c383f7c),
	.w2(32'hbaa41936),
	.w3(32'hbbb76fa8),
	.w4(32'h3c3a8df5),
	.w5(32'h3b11d705),
	.w6(32'hb9b9185d),
	.w7(32'h3c0c13b0),
	.w8(32'h3b160a6e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf1cb8),
	.w1(32'hbb254110),
	.w2(32'hbc12a1fe),
	.w3(32'h3b9afc3a),
	.w4(32'h3bae209d),
	.w5(32'h3a30add4),
	.w6(32'h3b7b5863),
	.w7(32'hba2de9ad),
	.w8(32'h38bec84e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64b271),
	.w1(32'h3c41ea2a),
	.w2(32'h3bbbd1b2),
	.w3(32'hba576675),
	.w4(32'h3b5d8356),
	.w5(32'h3b875ad7),
	.w6(32'h3ac23628),
	.w7(32'h3a80dc81),
	.w8(32'h39a42c4d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee9c04),
	.w1(32'h3a7d6e4c),
	.w2(32'hba59e51c),
	.w3(32'h3b2b3a6f),
	.w4(32'h39b07ff4),
	.w5(32'h39c2db20),
	.w6(32'hbbbccf18),
	.w7(32'hbc1c943b),
	.w8(32'hbbb32aab),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1d5e1),
	.w1(32'hbae99e16),
	.w2(32'hbae31fc3),
	.w3(32'hbb982536),
	.w4(32'hbadfcead),
	.w5(32'hba49a31a),
	.w6(32'hbabc56a7),
	.w7(32'hbab78e4b),
	.w8(32'h3a309e92),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0274b6),
	.w1(32'hbc0341e9),
	.w2(32'hbba8b6df),
	.w3(32'hbaa88aa1),
	.w4(32'hbc806020),
	.w5(32'hbc3274c8),
	.w6(32'hbb481dd9),
	.w7(32'hbb747d7a),
	.w8(32'hbbdb8617),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0ab12),
	.w1(32'h3ab97254),
	.w2(32'hbb10e607),
	.w3(32'hbba6cefd),
	.w4(32'h3b5c7f62),
	.w5(32'h3b16e71e),
	.w6(32'h3bbd94a6),
	.w7(32'h3bf0b71c),
	.w8(32'h3c06fb7d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b1d8e),
	.w1(32'hbbc61d72),
	.w2(32'h3bbadd7a),
	.w3(32'h3ad2d6be),
	.w4(32'h3b06196d),
	.w5(32'h3b2ba4bc),
	.w6(32'h3c5fdc7d),
	.w7(32'h3c940228),
	.w8(32'h3c534f06),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f9019),
	.w1(32'hb9f244b7),
	.w2(32'hba722437),
	.w3(32'h3aa63cff),
	.w4(32'h3aa88f15),
	.w5(32'h3aa989d4),
	.w6(32'h3970fa67),
	.w7(32'h3adb225b),
	.w8(32'h3a934386),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b50a),
	.w1(32'hbb869a77),
	.w2(32'hbb8b45bf),
	.w3(32'hbb2919de),
	.w4(32'hbab9dd17),
	.w5(32'h3a26495d),
	.w6(32'hb9ccaff2),
	.w7(32'hbb8751a9),
	.w8(32'hbb2b0b5b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1784e1),
	.w1(32'h3c624d5e),
	.w2(32'h3ba1cf87),
	.w3(32'hbab464aa),
	.w4(32'h3b8f7da4),
	.w5(32'h3b769626),
	.w6(32'hbbd00104),
	.w7(32'hbae1c0d0),
	.w8(32'hba37b0a1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a435dae),
	.w1(32'hbbde3298),
	.w2(32'hbbaee74b),
	.w3(32'h3bea138f),
	.w4(32'h3a1466a2),
	.w5(32'hbac44403),
	.w6(32'h3b592e99),
	.w7(32'h3bee3bb2),
	.w8(32'h3b93d7ad),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0625d),
	.w1(32'h3c221c3d),
	.w2(32'hbb9a6a25),
	.w3(32'hba3cf535),
	.w4(32'h3bb86e09),
	.w5(32'hbc0321a9),
	.w6(32'h3bc3d213),
	.w7(32'h3bfc0ed4),
	.w8(32'h3b25bbab),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc22932),
	.w1(32'hbbb84b88),
	.w2(32'hbc43deb7),
	.w3(32'hbb7a8a81),
	.w4(32'h3af4c5bd),
	.w5(32'h3b31894d),
	.w6(32'hbbb2e5ec),
	.w7(32'hbbaa1c41),
	.w8(32'hbb644711),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c146dd5),
	.w1(32'h3c06d4f9),
	.w2(32'hbc85b687),
	.w3(32'h3b78b0ff),
	.w4(32'h3c7036e2),
	.w5(32'hbb34a48d),
	.w6(32'hba209828),
	.w7(32'hbc51e230),
	.w8(32'hbc68784c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4efc5),
	.w1(32'hbb0933ae),
	.w2(32'hbbb5bfa2),
	.w3(32'h3b475ebf),
	.w4(32'h3b8be28d),
	.w5(32'hbb48d2f6),
	.w6(32'h3b7f4dc9),
	.w7(32'h3bbd0639),
	.w8(32'h3b93d7c2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb469d4a),
	.w1(32'hbccbe0eb),
	.w2(32'hbcafed6d),
	.w3(32'h3bf69a80),
	.w4(32'hba2145d8),
	.w5(32'hbad0ea2c),
	.w6(32'hbc340e6e),
	.w7(32'hbc99d158),
	.w8(32'hbca5568c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59897c),
	.w1(32'h3b2d1cb5),
	.w2(32'h3ba73fbc),
	.w3(32'h3bbb3f1f),
	.w4(32'h39d1f05a),
	.w5(32'h3aba1de5),
	.w6(32'h3b57666f),
	.w7(32'h3bafdce7),
	.w8(32'hbb4527f9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c108736),
	.w1(32'h3b5c3627),
	.w2(32'hbb8d229b),
	.w3(32'h3beea8c2),
	.w4(32'h3bbe1142),
	.w5(32'h39c2f992),
	.w6(32'hbc8571f5),
	.w7(32'hbcaac6a7),
	.w8(32'hbbee9007),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0966c9),
	.w1(32'h3c7118af),
	.w2(32'hbba510f7),
	.w3(32'hbbe1021b),
	.w4(32'h3bcac767),
	.w5(32'hb8cf88bf),
	.w6(32'hbaefe72f),
	.w7(32'hbadf0c40),
	.w8(32'hbb8bc899),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc662449),
	.w1(32'h3ca0e5af),
	.w2(32'h3c777c5a),
	.w3(32'hbc2f9143),
	.w4(32'h39c2aab3),
	.w5(32'h3c266f4b),
	.w6(32'h3bd83419),
	.w7(32'hbc105db2),
	.w8(32'hbbe1fdab),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb452260),
	.w1(32'hbc99a466),
	.w2(32'hbc9cb5fb),
	.w3(32'h3c825e77),
	.w4(32'hbc72984b),
	.w5(32'hbc8740b8),
	.w6(32'h3c96da60),
	.w7(32'h3c2ffa97),
	.w8(32'hbc772c7e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ac854),
	.w1(32'hbca52830),
	.w2(32'hbcaccb1e),
	.w3(32'h3b9204d4),
	.w4(32'hbcbcd070),
	.w5(32'hbc8cc667),
	.w6(32'h3ba4db90),
	.w7(32'hbc2d3765),
	.w8(32'hbc67fe0f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf161a6),
	.w1(32'h3c82c2c1),
	.w2(32'hbb56b3a8),
	.w3(32'hbaa06eea),
	.w4(32'hbb485f92),
	.w5(32'hbc6b3f79),
	.w6(32'hbb421034),
	.w7(32'h3b86c6ca),
	.w8(32'h3a8e57b3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2534ab),
	.w1(32'h39b09d0d),
	.w2(32'h39ec065d),
	.w3(32'hbb148646),
	.w4(32'hbb966f6e),
	.w5(32'hba2fc507),
	.w6(32'hb9bdd291),
	.w7(32'h3b733da2),
	.w8(32'hbaffe7a9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b015c85),
	.w1(32'h3c86e7c2),
	.w2(32'h3c82bfc2),
	.w3(32'hbb980e57),
	.w4(32'hbb8c7af5),
	.w5(32'hbaacf8ec),
	.w6(32'hbbda5af8),
	.w7(32'hbb2d70c6),
	.w8(32'hbb07691e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906a086),
	.w1(32'h3ac49e28),
	.w2(32'h3b91aabf),
	.w3(32'hbb34116d),
	.w4(32'hba8850bb),
	.w5(32'h3a9a72f7),
	.w6(32'hbb2fcc21),
	.w7(32'hbaf80b87),
	.w8(32'hba988e5f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60503d),
	.w1(32'h3a1c5e58),
	.w2(32'h3a0d319d),
	.w3(32'hbb7a3bb5),
	.w4(32'hbb1cd3d0),
	.w5(32'hbb362444),
	.w6(32'h3b248bd6),
	.w7(32'h3b0292b6),
	.w8(32'h3afd17fb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb001270),
	.w1(32'hbbc0c860),
	.w2(32'hbbd9a365),
	.w3(32'h3a8097d6),
	.w4(32'h3a3a6c17),
	.w5(32'hba655800),
	.w6(32'h3ba77d5b),
	.w7(32'h3bc17df9),
	.w8(32'h3afffef5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f77590),
	.w1(32'h3bdb685a),
	.w2(32'h3b881c2f),
	.w3(32'hba1bccdf),
	.w4(32'hb9adc5dd),
	.w5(32'hbba04b01),
	.w6(32'hbadd8980),
	.w7(32'h3b5b547b),
	.w8(32'hba86bcbe),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812425),
	.w1(32'hbb86e7a7),
	.w2(32'h3b6eb0a3),
	.w3(32'hbae09268),
	.w4(32'hbc031186),
	.w5(32'hbc290bf8),
	.w6(32'h3c20254c),
	.w7(32'h3c5062d9),
	.w8(32'h3c6c83f2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6cc2a),
	.w1(32'h3ae9c505),
	.w2(32'h3b4dac6e),
	.w3(32'hbbd8eb7c),
	.w4(32'h3bebe74f),
	.w5(32'h3b16373b),
	.w6(32'hba0c8164),
	.w7(32'h39839bee),
	.w8(32'h3b970fcc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15ad29),
	.w1(32'hbc3a77f2),
	.w2(32'hbb990e3a),
	.w3(32'hba2a1b0c),
	.w4(32'hba8f0dd2),
	.w5(32'hbb8e0cdf),
	.w6(32'hbbb8f783),
	.w7(32'hbc79a16f),
	.w8(32'h3bb62283),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc035ddd),
	.w1(32'h3c3c8a12),
	.w2(32'h3b160116),
	.w3(32'hbcb196aa),
	.w4(32'hbb49ef8b),
	.w5(32'hbbae781a),
	.w6(32'hb8c7dad9),
	.w7(32'hbc2ad5d9),
	.w8(32'hbc3493be),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94d66c),
	.w1(32'h3c0f4b33),
	.w2(32'h3b078bb1),
	.w3(32'h3c63bce5),
	.w4(32'h3c629524),
	.w5(32'h3bd2f1ad),
	.w6(32'h3bf052b7),
	.w7(32'h3c0ccc66),
	.w8(32'h3b612437),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b095539),
	.w1(32'h3ae2cb85),
	.w2(32'hbb5f75b2),
	.w3(32'h391e08bb),
	.w4(32'h3a452641),
	.w5(32'hbbf980aa),
	.w6(32'h3ba8109c),
	.w7(32'h3af01518),
	.w8(32'h3c1cf3ee),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe4eae),
	.w1(32'hb954a656),
	.w2(32'h37f57914),
	.w3(32'hbba0b250),
	.w4(32'hbb7cab60),
	.w5(32'hbc08e5d8),
	.w6(32'h3b679bd5),
	.w7(32'h3c05d5ed),
	.w8(32'h3b4edf64),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae240e9),
	.w1(32'hbb672938),
	.w2(32'hbb2a8aee),
	.w3(32'hbaab7d32),
	.w4(32'hbb44d866),
	.w5(32'hbbb820c1),
	.w6(32'h39efd5f8),
	.w7(32'h3a8dab7f),
	.w8(32'hba6a4dc0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aefab),
	.w1(32'hbb26b502),
	.w2(32'hbb27a6e6),
	.w3(32'hbb5337c7),
	.w4(32'hbb247ad1),
	.w5(32'hbb721dde),
	.w6(32'hbabe60b4),
	.w7(32'hba3ad78e),
	.w8(32'hbb34532b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cae17),
	.w1(32'hbc828891),
	.w2(32'hbc945ea9),
	.w3(32'hbaaee82a),
	.w4(32'hbc7e42b6),
	.w5(32'hbcee4b34),
	.w6(32'hbc816a25),
	.w7(32'hbcc9c64c),
	.w8(32'hbc5c5b34),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccabb6c),
	.w1(32'hbbbee8dd),
	.w2(32'hbb85f5df),
	.w3(32'hbcbbfa37),
	.w4(32'hbc23e576),
	.w5(32'hbc3eccb6),
	.w6(32'hba244ca7),
	.w7(32'hba15c25e),
	.w8(32'hbc04ebef),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb95033),
	.w1(32'h3b175dcc),
	.w2(32'h3ab3211d),
	.w3(32'hbaf5d164),
	.w4(32'hbbcd7ffa),
	.w5(32'hbae62259),
	.w6(32'h3b40cff5),
	.w7(32'h3b1665e6),
	.w8(32'hbafed173),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd964c6),
	.w1(32'h3c03c477),
	.w2(32'hbacd4068),
	.w3(32'hbb019b49),
	.w4(32'h3b1169da),
	.w5(32'h39a49809),
	.w6(32'hbba632a5),
	.w7(32'hbbf15f9c),
	.w8(32'hbc24b28e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56f2c4),
	.w1(32'hbc55dcc5),
	.w2(32'hbbd462f4),
	.w3(32'hbb75a728),
	.w4(32'hbb98d6ed),
	.w5(32'hbbdd733d),
	.w6(32'h3c23f0fa),
	.w7(32'h3c49f44c),
	.w8(32'h3b9e6c34),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a181409),
	.w1(32'hbc9d9d11),
	.w2(32'hbc85c06c),
	.w3(32'hba5f01b6),
	.w4(32'hbc19935b),
	.w5(32'hbca1c513),
	.w6(32'hbc7c402d),
	.w7(32'hbcff1da6),
	.w8(32'hbcb18e64),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca16c0d),
	.w1(32'h3ae2bfe8),
	.w2(32'hbb81bcf3),
	.w3(32'hbc18fff0),
	.w4(32'h3c02115b),
	.w5(32'h3c5ab526),
	.w6(32'hbbf1867c),
	.w7(32'hbc76aff9),
	.w8(32'hbc2eac59),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ebf45),
	.w1(32'hbb5c6eb3),
	.w2(32'hbb1f3b0f),
	.w3(32'h3c4e48a9),
	.w4(32'hba739752),
	.w5(32'h3ad4e76c),
	.w6(32'hbadf2bda),
	.w7(32'h3959e1aa),
	.w8(32'hba82a57a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4d0bd),
	.w1(32'h391a0c8a),
	.w2(32'hb89dab03),
	.w3(32'hba85656d),
	.w4(32'hb8631a2f),
	.w5(32'hb98d2fcf),
	.w6(32'h39774484),
	.w7(32'h38e3e2e5),
	.w8(32'hb93a85cf),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96aed3),
	.w1(32'h3bf692b4),
	.w2(32'h3b983518),
	.w3(32'hbc6b3203),
	.w4(32'hbb3b2765),
	.w5(32'h35242000),
	.w6(32'h3b9e9c20),
	.w7(32'h3a473661),
	.w8(32'hbc318ee8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31f082),
	.w1(32'h3c0ddabd),
	.w2(32'h3997fea6),
	.w3(32'h3bb7a544),
	.w4(32'h3c0cf379),
	.w5(32'h3ad88353),
	.w6(32'hbba69259),
	.w7(32'hbb8e2892),
	.w8(32'hbbbc2cf0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac46d85),
	.w1(32'h3b0a8013),
	.w2(32'hb96a8cf8),
	.w3(32'h3a5b4c1a),
	.w4(32'h3adb3d28),
	.w5(32'hb8f2a6cc),
	.w6(32'hba01f305),
	.w7(32'h38b5beb5),
	.w8(32'hb58a02d4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d9fce),
	.w1(32'h3b0deced),
	.w2(32'hbac3c9a1),
	.w3(32'hbb39262f),
	.w4(32'h38cae02e),
	.w5(32'hbb1f48e0),
	.w6(32'hbab32466),
	.w7(32'hbae0a97e),
	.w8(32'hbadaedce),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58ae84),
	.w1(32'hbae9cc98),
	.w2(32'hbaaeb36d),
	.w3(32'hb9343d2f),
	.w4(32'hba0bb029),
	.w5(32'hba8119a9),
	.w6(32'hb9c55daa),
	.w7(32'h3a2ced27),
	.w8(32'hb8c7186b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0560e7),
	.w1(32'h3aa819c5),
	.w2(32'hba894d72),
	.w3(32'hb8fa9fa1),
	.w4(32'h3aa98e45),
	.w5(32'hbaafce99),
	.w6(32'hba485511),
	.w7(32'hba8ba395),
	.w8(32'hbaa2a6ff),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ca7e),
	.w1(32'hbbb40a42),
	.w2(32'h3ace844f),
	.w3(32'h3b9ff360),
	.w4(32'h3b799cba),
	.w5(32'h3b4c42ad),
	.w6(32'h3b812e89),
	.w7(32'h3bdd3b23),
	.w8(32'h3bcb2f6a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c997395),
	.w1(32'h3cab34ff),
	.w2(32'h3bcdc13d),
	.w3(32'h3b328aa1),
	.w4(32'h3c40759c),
	.w5(32'hba86408c),
	.w6(32'hbc0047d6),
	.w7(32'hbbfd713a),
	.w8(32'hbbea43cf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c4c4),
	.w1(32'hbbff3615),
	.w2(32'hbb4d2bbc),
	.w3(32'hb9dcc64a),
	.w4(32'hbb1d877c),
	.w5(32'hbb02060a),
	.w6(32'h3b4b4b57),
	.w7(32'h3b89cd47),
	.w8(32'h3a6e5aac),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7fbea),
	.w1(32'h3b834ff3),
	.w2(32'hb8858f17),
	.w3(32'h3ba98149),
	.w4(32'h3bba241d),
	.w5(32'h3aa38817),
	.w6(32'h3b48a2e4),
	.w7(32'h3a9dbc46),
	.w8(32'hbb23b281),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b89c7),
	.w1(32'h3c26a460),
	.w2(32'h3b235977),
	.w3(32'hbb190321),
	.w4(32'h39830fba),
	.w5(32'hba96bd11),
	.w6(32'hbbfba2de),
	.w7(32'hbbbf872c),
	.w8(32'hbb35d8ac),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa2d1),
	.w1(32'hbb9460c2),
	.w2(32'hbac68d58),
	.w3(32'hbb607b13),
	.w4(32'hbbe5a475),
	.w5(32'hbb9191a7),
	.w6(32'h3a9ac40e),
	.w7(32'hba22fb8a),
	.w8(32'hbb452405),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fc701),
	.w1(32'h3bc53be1),
	.w2(32'h39efbb41),
	.w3(32'h3aebff5d),
	.w4(32'h3b7d4786),
	.w5(32'h3a9421d2),
	.w6(32'hbb860de6),
	.w7(32'hbb060e94),
	.w8(32'hbb1a9e20),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9e240),
	.w1(32'hba2e13ca),
	.w2(32'hb9db51f5),
	.w3(32'hb94f42e7),
	.w4(32'hb9e58d78),
	.w5(32'hb9e67c84),
	.w6(32'hb9e8fe45),
	.w7(32'hb9a81c98),
	.w8(32'hb9e72026),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b167a),
	.w1(32'hbbf0f8d9),
	.w2(32'hbbca4662),
	.w3(32'h3b0d54bc),
	.w4(32'hbb7d2396),
	.w5(32'hbb42ca6f),
	.w6(32'h3bdf465b),
	.w7(32'h3c120e84),
	.w8(32'h3813874d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3035d),
	.w1(32'hbb31a6fc),
	.w2(32'hb8c75f29),
	.w3(32'h39051278),
	.w4(32'h37f8433e),
	.w5(32'hba625213),
	.w6(32'h3ae414b8),
	.w7(32'h38a87379),
	.w8(32'hbb1e3cf5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e2225),
	.w1(32'h3a0a9053),
	.w2(32'h394ab335),
	.w3(32'h39b53bc3),
	.w4(32'h398f5198),
	.w5(32'h396d25da),
	.w6(32'h3a411bb0),
	.w7(32'h39d608fe),
	.w8(32'hb8a542a2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969f2ba),
	.w1(32'h3788dbef),
	.w2(32'hb8dba70c),
	.w3(32'hb77714a6),
	.w4(32'h386918a6),
	.w5(32'hb8cf9031),
	.w6(32'hb8474d29),
	.w7(32'hb8aae8fa),
	.w8(32'hb8b0e00b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac192c0),
	.w1(32'hba93a9bf),
	.w2(32'hba25f14f),
	.w3(32'h3ab4fec2),
	.w4(32'h3a1e79e1),
	.w5(32'h3a62ce76),
	.w6(32'hbb0025aa),
	.w7(32'hbaf0e7f6),
	.w8(32'hbab7e4ca),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8d1a8),
	.w1(32'hbc1bfc03),
	.w2(32'h39941c92),
	.w3(32'h3a41c680),
	.w4(32'hb9f59ff4),
	.w5(32'h3b1440fc),
	.w6(32'h3b97cfad),
	.w7(32'h3bb81f7e),
	.w8(32'h39d2ecf9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3379f9),
	.w1(32'h3b0e3c87),
	.w2(32'h3aef2d61),
	.w3(32'hb98d5044),
	.w4(32'h39e6bfa3),
	.w5(32'h39cfec92),
	.w6(32'hbb34ecb6),
	.w7(32'hbb560ca7),
	.w8(32'hbb16c183),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857d414),
	.w1(32'h3893a92a),
	.w2(32'h37d334b8),
	.w3(32'h38777beb),
	.w4(32'h38741d72),
	.w5(32'h389282ba),
	.w6(32'hb66f89eb),
	.w7(32'h38522999),
	.w8(32'h38d43f79),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8d1db),
	.w1(32'h3bbe2c0c),
	.w2(32'h393baa65),
	.w3(32'h3b841f7d),
	.w4(32'h3bab6a90),
	.w5(32'h3a96e8fe),
	.w6(32'hbb70708f),
	.w7(32'hbad1d36a),
	.w8(32'hba9eb742),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c2e0a),
	.w1(32'hba9e3714),
	.w2(32'hba8cd0d1),
	.w3(32'hba664cc7),
	.w4(32'hbaec829d),
	.w5(32'hbaf06da2),
	.w6(32'hbac109ab),
	.w7(32'hbacb11a8),
	.w8(32'hbad8dc96),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3996e),
	.w1(32'h3c65e91c),
	.w2(32'h3b37c843),
	.w3(32'hbbdb2624),
	.w4(32'h3b0d9281),
	.w5(32'hbb967357),
	.w6(32'hbbb806ec),
	.w7(32'hbba58022),
	.w8(32'hbb98b080),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d36af),
	.w1(32'hbc4f9786),
	.w2(32'hbbedcd1e),
	.w3(32'h3beaf9de),
	.w4(32'h3be1e670),
	.w5(32'hbb96c163),
	.w6(32'h3c22583a),
	.w7(32'h3c821684),
	.w8(32'h3c270087),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb450f6c),
	.w1(32'hbb8d0788),
	.w2(32'h38b4fa88),
	.w3(32'h3a19b261),
	.w4(32'h399044f9),
	.w5(32'h39f88174),
	.w6(32'h3b88db3c),
	.w7(32'h3b72345d),
	.w8(32'h3b12a0a9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a104029),
	.w1(32'h3a4b54f8),
	.w2(32'h3a4ffafc),
	.w3(32'h3aa00254),
	.w4(32'h3ab46ca7),
	.w5(32'h3a3d6044),
	.w6(32'h3ad5a1b6),
	.w7(32'h3ad61e44),
	.w8(32'h3a3849f9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402563),
	.w1(32'hbbb89f3e),
	.w2(32'hbb83890d),
	.w3(32'hbafaddad),
	.w4(32'hbb916188),
	.w5(32'hbb4de2d5),
	.w6(32'hb983f4cc),
	.w7(32'hbaa248be),
	.w8(32'hbb040b58),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a087c47),
	.w1(32'hbb6979a1),
	.w2(32'hb9a31629),
	.w3(32'h3b334bd8),
	.w4(32'h3ab8da89),
	.w5(32'hb950d190),
	.w6(32'h3b0390f0),
	.w7(32'h3b4d18f6),
	.w8(32'h3ad1b8a4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb959886),
	.w1(32'hbbb91258),
	.w2(32'hbb613367),
	.w3(32'hbb06503d),
	.w4(32'hbaf6b637),
	.w5(32'hbb0fb0cb),
	.w6(32'h3aaf98d3),
	.w7(32'h3b5139b2),
	.w8(32'h3ad6d475),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae43a05),
	.w1(32'h3b844d19),
	.w2(32'h3af90e1b),
	.w3(32'hb7a04cfb),
	.w4(32'h3a54f4d4),
	.w5(32'h3a36a363),
	.w6(32'hbaf28a71),
	.w7(32'hbaaa10da),
	.w8(32'hb97dc350),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c7700),
	.w1(32'hba456cfb),
	.w2(32'hb95a2437),
	.w3(32'hb9dc897a),
	.w4(32'hb91e040b),
	.w5(32'hba6babfc),
	.w6(32'h3a41745c),
	.w7(32'h3921d782),
	.w8(32'h3703b196),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb6055),
	.w1(32'h3c070133),
	.w2(32'h38c290d3),
	.w3(32'h3b14cb82),
	.w4(32'h3b67deec),
	.w5(32'hba88510d),
	.w6(32'hbb1ebde3),
	.w7(32'hbaf03a02),
	.w8(32'hbb739298),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d097d),
	.w1(32'h3ad5768b),
	.w2(32'h3a1fe837),
	.w3(32'hba922a07),
	.w4(32'h3a0b5696),
	.w5(32'h39edd657),
	.w6(32'hb8738cd6),
	.w7(32'h39ab9cde),
	.w8(32'hb9c45cfe),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9694c),
	.w1(32'hbb76333d),
	.w2(32'hbb92d447),
	.w3(32'hb853cfa8),
	.w4(32'hbb772b22),
	.w5(32'hbb77009c),
	.w6(32'h3b1876d6),
	.w7(32'h3a4a494e),
	.w8(32'hbae22aaa),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886a217),
	.w1(32'h394fbc40),
	.w2(32'h38fe1d1a),
	.w3(32'hb7e9b6f5),
	.w4(32'h398473e3),
	.w5(32'h3959f88f),
	.w6(32'h37fa6a1f),
	.w7(32'h3985cb54),
	.w8(32'h38d68521),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06bc61),
	.w1(32'h3aaff058),
	.w2(32'h3a0bf003),
	.w3(32'hbb3645ad),
	.w4(32'h3b82d781),
	.w5(32'h3b87130b),
	.w6(32'h39659261),
	.w7(32'h3a3103a9),
	.w8(32'hbb586e61),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e5a5cd),
	.w1(32'h38250b85),
	.w2(32'h38dbb6c3),
	.w3(32'hb823ee71),
	.w4(32'h375688a7),
	.w5(32'h38ac6858),
	.w6(32'h3833560d),
	.w7(32'h38ae20a2),
	.w8(32'h3908e4f1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a470c53),
	.w1(32'h3a4a77a2),
	.w2(32'h3a037f65),
	.w3(32'h3a46243d),
	.w4(32'h3a1f1622),
	.w5(32'h39a73b44),
	.w6(32'h3a174c3f),
	.w7(32'h39bea8cc),
	.w8(32'h3989607f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4f04c),
	.w1(32'hbb8733d2),
	.w2(32'hbaef33a4),
	.w3(32'h3a5db0dd),
	.w4(32'hba11b9ea),
	.w5(32'hba433255),
	.w6(32'h3a91d0cf),
	.w7(32'h3b22b2b1),
	.w8(32'h39ac6183),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f56e5),
	.w1(32'h3c243176),
	.w2(32'h3b878e87),
	.w3(32'hbbf7e94d),
	.w4(32'hbac1bdb9),
	.w5(32'hba54125d),
	.w6(32'hbb83ab35),
	.w7(32'hbbfea9c7),
	.w8(32'hbc22466b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a1507),
	.w1(32'h397e3d43),
	.w2(32'h39a6422d),
	.w3(32'h39aab926),
	.w4(32'h3a373a88),
	.w5(32'h39cb32d9),
	.w6(32'h3a25d7c4),
	.w7(32'h3a5f2546),
	.w8(32'h389fff25),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e243d),
	.w1(32'hbbd88d81),
	.w2(32'hbb79dce3),
	.w3(32'hba3d71e2),
	.w4(32'hbb2da455),
	.w5(32'hbb058593),
	.w6(32'h3b21bc6e),
	.w7(32'h3b00032a),
	.w8(32'h3a5d36ad),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39640a),
	.w1(32'hba774a2a),
	.w2(32'h3b305194),
	.w3(32'h3b505eda),
	.w4(32'h3bf1b356),
	.w5(32'h3bcd1382),
	.w6(32'h385db5b4),
	.w7(32'h3b3b9010),
	.w8(32'h3b8ce7ec),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c92b4),
	.w1(32'h3bc9dfd5),
	.w2(32'h3b6ab7cf),
	.w3(32'h3c23e2f4),
	.w4(32'h3b750caa),
	.w5(32'h3b31460e),
	.w6(32'hbb112a9f),
	.w7(32'hbb37d121),
	.w8(32'h3a2a2e41),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cbefd),
	.w1(32'h3ba615ec),
	.w2(32'h3b2741e5),
	.w3(32'h37b208bc),
	.w4(32'h3b20c120),
	.w5(32'h3abd2314),
	.w6(32'hbae0cefc),
	.w7(32'hba944d41),
	.w8(32'h39cc23c2),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf67c8b),
	.w1(32'h3bddbbd7),
	.w2(32'h3acbdc03),
	.w3(32'h3a97425c),
	.w4(32'h3b58a9f2),
	.w5(32'h39736f2d),
	.w6(32'hbbbc3e02),
	.w7(32'hbbadc915),
	.w8(32'hbb99bea6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7192f10),
	.w1(32'h39b9c1aa),
	.w2(32'h39c970fe),
	.w3(32'hb8dabbef),
	.w4(32'h39bb621c),
	.w5(32'h39d46ca0),
	.w6(32'hb8a9a21b),
	.w7(32'h39e0735d),
	.w8(32'h3a0a1dcc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cae70),
	.w1(32'hb9b0c09a),
	.w2(32'hbb1ba2ba),
	.w3(32'h3b500a76),
	.w4(32'h3b464f9d),
	.w5(32'hb9bd7497),
	.w6(32'h39edfd44),
	.w7(32'h3a91aaec),
	.w8(32'h3a59d1e7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38454ff9),
	.w1(32'h379deb9b),
	.w2(32'h3797f0cb),
	.w3(32'h3732997b),
	.w4(32'h37d7d5ec),
	.w5(32'h37ff8a04),
	.w6(32'h3787e00d),
	.w7(32'h37fe4fbf),
	.w8(32'h3837ced7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affc0ad),
	.w1(32'h3a25fa24),
	.w2(32'h3a7cbe51),
	.w3(32'h39b1ae74),
	.w4(32'hb959df20),
	.w5(32'h3800ddd2),
	.w6(32'hb8cf1e55),
	.w7(32'hba506746),
	.w8(32'hb84aa49f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e6c7c),
	.w1(32'hbaacc63d),
	.w2(32'hba914e9a),
	.w3(32'hba462597),
	.w4(32'hb9a6f9c6),
	.w5(32'hb9857575),
	.w6(32'h3aab79e9),
	.w7(32'h3aef0454),
	.w8(32'h3aa95dd3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b827e),
	.w1(32'h3a9804ac),
	.w2(32'hbb536541),
	.w3(32'h3bcddbfb),
	.w4(32'h3b3f73ed),
	.w5(32'hba8ab3bd),
	.w6(32'h3ac539cf),
	.w7(32'h3aa900be),
	.w8(32'hb941124b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ef4032),
	.w1(32'hb84f11c6),
	.w2(32'hb506a814),
	.w3(32'hb760249b),
	.w4(32'hb80251b1),
	.w5(32'hb709344c),
	.w6(32'h3735bcf8),
	.w7(32'h37557ac6),
	.w8(32'h37c55eba),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37db9096),
	.w1(32'h37abdeaa),
	.w2(32'h37a78f62),
	.w3(32'h383920ae),
	.w4(32'h384087d2),
	.w5(32'h37978e3f),
	.w6(32'hb73ac941),
	.w7(32'hb669f8ee),
	.w8(32'hb866f94c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9cc16),
	.w1(32'hbb66b862),
	.w2(32'hbb85a5bb),
	.w3(32'hbaae90f7),
	.w4(32'hba88a5bc),
	.w5(32'hbac83ff3),
	.w6(32'h3b3e4439),
	.w7(32'h3a0e24b7),
	.w8(32'h39b24ef6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d97c),
	.w1(32'h3c1fce79),
	.w2(32'h3b547a93),
	.w3(32'h3b61e5f2),
	.w4(32'h3ac1a771),
	.w5(32'h3af398ee),
	.w6(32'h3ad76ed4),
	.w7(32'h3a649ad9),
	.w8(32'h3c1c60fc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb762919),
	.w1(32'h39daeede),
	.w2(32'h3b1234d4),
	.w3(32'hbaaf93fa),
	.w4(32'hbb0ebb35),
	.w5(32'h3b9eaf86),
	.w6(32'h38ddb5c6),
	.w7(32'hbabe4264),
	.w8(32'h3ad30d64),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0200c6),
	.w1(32'hb8a4f42f),
	.w2(32'h38a1bbbb),
	.w3(32'hb9d7e61b),
	.w4(32'hb9803f17),
	.w5(32'h38be919d),
	.w6(32'hb9f73b78),
	.w7(32'hb98c8737),
	.w8(32'hb827f734),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77f8a0),
	.w1(32'h3c46aa69),
	.w2(32'h3b82d094),
	.w3(32'h3b125d4d),
	.w4(32'h39fbf0d9),
	.w5(32'hbbb0a615),
	.w6(32'hbb8721e6),
	.w7(32'hbc167db5),
	.w8(32'hbc2daa3c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c647cb4),
	.w1(32'hbc274ba5),
	.w2(32'hbb90eba4),
	.w3(32'h3c5a0e58),
	.w4(32'h3c3098d1),
	.w5(32'h3b0e8383),
	.w6(32'h3bdbfaeb),
	.w7(32'h3c421e2b),
	.w8(32'h3c262ffc),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46e06b),
	.w1(32'h3bca54f8),
	.w2(32'h3ab52151),
	.w3(32'hbb34ac54),
	.w4(32'h3b1b66cd),
	.w5(32'h3b197fb9),
	.w6(32'hba99d718),
	.w7(32'h3aba322b),
	.w8(32'h3afc37f9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c6e96c),
	.w1(32'h37691750),
	.w2(32'h36656e77),
	.w3(32'h381fbe17),
	.w4(32'h3798e458),
	.w5(32'h378a4188),
	.w6(32'h38a4f0bf),
	.w7(32'h374cdfd1),
	.w8(32'h3816009b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f8c2af),
	.w1(32'hb6d7253d),
	.w2(32'h38a83b99),
	.w3(32'h3907a3e1),
	.w4(32'h3820c003),
	.w5(32'hb60ca4ef),
	.w6(32'h380bad42),
	.w7(32'hb8cfe65c),
	.w8(32'hb919c244),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381bd414),
	.w1(32'h37d870c1),
	.w2(32'h37549612),
	.w3(32'h37f40487),
	.w4(32'h37af015e),
	.w5(32'h378e63c1),
	.w6(32'h3700419e),
	.w7(32'hb62cc567),
	.w8(32'h3729f5f8),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6af998),
	.w1(32'h3beb5fe9),
	.w2(32'h3a884fda),
	.w3(32'hbbc6369f),
	.w4(32'h3adc909f),
	.w5(32'h3b0af571),
	.w6(32'hbb311037),
	.w7(32'h3a9425d2),
	.w8(32'h370d417e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bd9c0),
	.w1(32'h3b4b71f5),
	.w2(32'h3b12d8c7),
	.w3(32'h39d0b792),
	.w4(32'h3a3ecf67),
	.w5(32'h39dd1628),
	.w6(32'hba8981eb),
	.w7(32'hbab73779),
	.w8(32'hbaf4ff81),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104c47),
	.w1(32'hbc0f888c),
	.w2(32'hbb32cf67),
	.w3(32'hbb3b11cf),
	.w4(32'hbbb5bfe6),
	.w5(32'hba8bc470),
	.w6(32'h3b9c0083),
	.w7(32'h3b86ed29),
	.w8(32'h3b794045),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0acb29),
	.w1(32'hbb050cd8),
	.w2(32'hbaabcfb7),
	.w3(32'hbaa6f888),
	.w4(32'hbb1603b4),
	.w5(32'hbaff5c1e),
	.w6(32'h391dc086),
	.w7(32'hba0a81f3),
	.w8(32'hba80d600),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde9343),
	.w1(32'h3bfc1f92),
	.w2(32'h3b854062),
	.w3(32'h3a5f24ad),
	.w4(32'h3b2d1f78),
	.w5(32'h3ac8bb64),
	.w6(32'hbbadb64b),
	.w7(32'hbb92d74f),
	.w8(32'hbb6da61b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb2c5d),
	.w1(32'hba01a9ad),
	.w2(32'h3b2693ee),
	.w3(32'h3a9177b1),
	.w4(32'hbb1e6aa7),
	.w5(32'h3ab8b0a8),
	.w6(32'h3b3048a7),
	.w7(32'h3a8f81c5),
	.w8(32'h3af5f919),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79b2c8b),
	.w1(32'hb7f06506),
	.w2(32'h358b3184),
	.w3(32'hb611c27a),
	.w4(32'hb715482e),
	.w5(32'h36d4157d),
	.w6(32'h37a3b9b4),
	.w7(32'h37b37b47),
	.w8(32'h37e9bf3d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf361fb),
	.w1(32'h3b3ba217),
	.w2(32'hbaba7327),
	.w3(32'h3b3654ef),
	.w4(32'hba964674),
	.w5(32'hbb0734d3),
	.w6(32'hb9575992),
	.w7(32'hbb1d5079),
	.w8(32'hbb320673),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37639109),
	.w1(32'hb89fd02a),
	.w2(32'h37850c50),
	.w3(32'h37323fa1),
	.w4(32'hb796dad0),
	.w5(32'h37e41143),
	.w6(32'h3885c2c5),
	.w7(32'h38927335),
	.w8(32'h38ac3b76),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d36b3),
	.w1(32'h3b1cb410),
	.w2(32'h3a2d368a),
	.w3(32'hba9bb500),
	.w4(32'h3a832ec6),
	.w5(32'h393cb88c),
	.w6(32'hbb4277a6),
	.w7(32'hbac31b00),
	.w8(32'hbb04b5dd),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb26650),
	.w1(32'hbc200054),
	.w2(32'hbb4a7bb3),
	.w3(32'hba44c8ad),
	.w4(32'hba15aa07),
	.w5(32'hbb3aa4f2),
	.w6(32'h3c1364f3),
	.w7(32'h3c2903bc),
	.w8(32'h3b92236b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac151e8),
	.w1(32'hbb861863),
	.w2(32'hbb1a9c1d),
	.w3(32'hbabde5a6),
	.w4(32'hbb1b2fe0),
	.w5(32'hbb072040),
	.w6(32'hba627ba4),
	.w7(32'h3a1ffa4f),
	.w8(32'hb9374dce),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82f6164),
	.w1(32'h394a6b28),
	.w2(32'h39614014),
	.w3(32'hb83edd9c),
	.w4(32'h3990bb15),
	.w5(32'h393098ff),
	.w6(32'hb7277f37),
	.w7(32'h39380599),
	.w8(32'hb7d17fa4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa80071),
	.w1(32'hbc2c1652),
	.w2(32'hbb26cd27),
	.w3(32'hba0ab215),
	.w4(32'hbb599e55),
	.w5(32'hba8f1598),
	.w6(32'h3b47312d),
	.w7(32'h3b6e40df),
	.w8(32'h3b3ae991),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b670e77),
	.w1(32'h3b43f2b9),
	.w2(32'hbae5ff82),
	.w3(32'hb8478a5c),
	.w4(32'h3b3646c4),
	.w5(32'hbb177759),
	.w6(32'hbb1d38b7),
	.w7(32'hba875cc9),
	.w8(32'hbb27c50b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e7d9f),
	.w1(32'h3a94ac9e),
	.w2(32'h3a86114b),
	.w3(32'hba86d2a3),
	.w4(32'hba8cbc39),
	.w5(32'hb938433f),
	.w6(32'hbb40502b),
	.w7(32'hbb802360),
	.w8(32'hbb190da2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e233bd),
	.w1(32'hb91372b7),
	.w2(32'hb91fc8a1),
	.w3(32'hb74ed36d),
	.w4(32'hb7d6044c),
	.w5(32'hb8d2f005),
	.w6(32'hb6b37198),
	.w7(32'h36a28106),
	.w8(32'hb7f9c72c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9617483),
	.w1(32'hb901de14),
	.w2(32'hb955d951),
	.w3(32'hb8a75530),
	.w4(32'h3991b6fd),
	.w5(32'h38b5fe87),
	.w6(32'h38918d89),
	.w7(32'h386b6826),
	.w8(32'h391d5e02),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34199b),
	.w1(32'h3bb32938),
	.w2(32'h3affb7f5),
	.w3(32'hbc041bc0),
	.w4(32'hbb98d2c3),
	.w5(32'hbb50c3c4),
	.w6(32'h3ab2cb6c),
	.w7(32'hbb88363d),
	.w8(32'hbc2d958b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e58b91),
	.w1(32'h3b7dca8e),
	.w2(32'h3a44d629),
	.w3(32'hba99124f),
	.w4(32'hbb9a6c0e),
	.w5(32'hbb74e990),
	.w6(32'hb986cdf4),
	.w7(32'hbbb136d5),
	.w8(32'hbc1df519),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcedad3),
	.w1(32'hbbf053cb),
	.w2(32'hbbc94fea),
	.w3(32'hbba3f79e),
	.w4(32'hbbb82433),
	.w5(32'hbb85f626),
	.w6(32'hba413d9a),
	.w7(32'hbb006eea),
	.w8(32'hbab9cf3c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd7b22),
	.w1(32'h3c271927),
	.w2(32'hbc098ada),
	.w3(32'hbc19a971),
	.w4(32'h3c4e7c3a),
	.w5(32'h3b0e7c98),
	.w6(32'hbbd9a6d9),
	.w7(32'h3b972438),
	.w8(32'hba35f80d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcdc93),
	.w1(32'hb9cabc42),
	.w2(32'h39a6e453),
	.w3(32'h3b0947a8),
	.w4(32'hba14d0dc),
	.w5(32'h3a287fcf),
	.w6(32'h3ac7c499),
	.w7(32'h3a63ef2b),
	.w8(32'hba899991),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad63c7),
	.w1(32'h3aa87f82),
	.w2(32'hb9bca29b),
	.w3(32'hb98c4a5a),
	.w4(32'h3a9faa7d),
	.w5(32'hba3b5c40),
	.w6(32'hb9249828),
	.w7(32'h395d66bd),
	.w8(32'hba14ca89),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30920e),
	.w1(32'h3c60d105),
	.w2(32'h3c30a7fe),
	.w3(32'hbc40c566),
	.w4(32'h3b850399),
	.w5(32'h3bb4fc91),
	.w6(32'hba08f9df),
	.w7(32'h3bb0c6df),
	.w8(32'hbb37b775),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d91c3),
	.w1(32'h3c3842cf),
	.w2(32'h3abbfe94),
	.w3(32'hbb00394c),
	.w4(32'h3b0e7a31),
	.w5(32'hbb6f79b5),
	.w6(32'hbbeca2b9),
	.w7(32'hbbf51e6d),
	.w8(32'hbc188b1b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aec9d4),
	.w1(32'h3c18c6fc),
	.w2(32'h3b548f1e),
	.w3(32'hbb8fcc06),
	.w4(32'hb7746fd6),
	.w5(32'hb9581ddb),
	.w6(32'hbb963cc6),
	.w7(32'hbbc3dea7),
	.w8(32'hbbd0fb5a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801421),
	.w1(32'hbc0e9582),
	.w2(32'hbbe161d9),
	.w3(32'hbadd7664),
	.w4(32'hbb8eca1a),
	.w5(32'hbb982360),
	.w6(32'h3b96ba72),
	.w7(32'h3bd7981d),
	.w8(32'h3ae1a64d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937290),
	.w1(32'hbc4cac29),
	.w2(32'hbba7dad7),
	.w3(32'h3b0c2117),
	.w4(32'hba7eebab),
	.w5(32'hbb6547c4),
	.w6(32'h3bf665e9),
	.w7(32'h3c10d12a),
	.w8(32'h3b91251a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76d9fc4),
	.w1(32'hb77f88e7),
	.w2(32'h3570228a),
	.w3(32'hb69240c9),
	.w4(32'hb6194dfb),
	.w5(32'h3717f19a),
	.w6(32'h3724de24),
	.w7(32'h3794023b),
	.w8(32'h3778e93b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60485f8),
	.w1(32'hb5c231dd),
	.w2(32'h372c71dc),
	.w3(32'h369befb7),
	.w4(32'h3732bb4a),
	.w5(32'h375810b1),
	.w6(32'h378d7e59),
	.w7(32'h3745041e),
	.w8(32'h378c705f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab66aea),
	.w1(32'hba8afecb),
	.w2(32'hbb316f91),
	.w3(32'hba6ff80a),
	.w4(32'h3a5e57ae),
	.w5(32'hb9d6465e),
	.w6(32'hba9fc674),
	.w7(32'hbaf9c367),
	.w8(32'hbb9cf380),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a283f0),
	.w1(32'hb6833204),
	.w2(32'hb6b24179),
	.w3(32'h356a4d38),
	.w4(32'hb70d6ef2),
	.w5(32'hb6e0779f),
	.w6(32'h37a07299),
	.w7(32'h3751c5c4),
	.w8(32'h373bb866),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad69b66),
	.w1(32'h3b89cf25),
	.w2(32'h3b84c50c),
	.w3(32'hba14fb9d),
	.w4(32'h3b8c4913),
	.w5(32'h3b8215c6),
	.w6(32'hba095213),
	.w7(32'h3ae7a3dc),
	.w8(32'h3b02fe39),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb743af0),
	.w1(32'h3b4719c9),
	.w2(32'hba8f5c34),
	.w3(32'hbb45aa3c),
	.w4(32'hbb485063),
	.w5(32'hba31be54),
	.w6(32'hb9baf25c),
	.w7(32'hbaeb7d45),
	.w8(32'hbbe47ed2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a69f4),
	.w1(32'hba172f1b),
	.w2(32'hb9b82405),
	.w3(32'hb9a7bfa4),
	.w4(32'hbaa6f35f),
	.w5(32'hba20045b),
	.w6(32'hb94ec95c),
	.w7(32'hba0ef03a),
	.w8(32'hba899501),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb808819a),
	.w1(32'hb824b898),
	.w2(32'h369be897),
	.w3(32'hb52a499a),
	.w4(32'h3523a87e),
	.w5(32'h365a7f07),
	.w6(32'h3838a236),
	.w7(32'h383c74af),
	.w8(32'h3736f57c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e09e1),
	.w1(32'h3c8cfac8),
	.w2(32'h3b5031b8),
	.w3(32'hbc283f0f),
	.w4(32'h3a709982),
	.w5(32'hbb8692ed),
	.w6(32'hbc1f4683),
	.w7(32'hbc571cc3),
	.w8(32'hbc1dcb07),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7930af),
	.w1(32'h3ba275ea),
	.w2(32'h3abac876),
	.w3(32'hb97a3dff),
	.w4(32'h3b01b443),
	.w5(32'h3a13c583),
	.w6(32'hbb4b6659),
	.w7(32'hbb1e79e7),
	.w8(32'hbb2a65f8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f90c34),
	.w1(32'hb7669a13),
	.w2(32'hb80b4004),
	.w3(32'h38468e60),
	.w4(32'hb8cf9e04),
	.w5(32'hb7140e9f),
	.w6(32'h3840a85c),
	.w7(32'hb7e1e67a),
	.w8(32'hb77439a1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd771ec),
	.w1(32'h3c1f26e8),
	.w2(32'h3b56bd15),
	.w3(32'hba7e44f6),
	.w4(32'h3b1ce3cc),
	.w5(32'h38994f98),
	.w6(32'hbb95a5c0),
	.w7(32'hbb2535f5),
	.w8(32'hbb67f588),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c84bed),
	.w1(32'h38beef1a),
	.w2(32'h38d1ca42),
	.w3(32'h3906bc9f),
	.w4(32'h3905c950),
	.w5(32'h38a7930b),
	.w6(32'h38e8e3e1),
	.w7(32'h38ce14db),
	.w8(32'h383215f3),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10f173),
	.w1(32'hb9a68224),
	.w2(32'hb998ced2),
	.w3(32'hb9d0994f),
	.w4(32'hb813d549),
	.w5(32'h38953032),
	.w6(32'hb9c94e4e),
	.w7(32'hb930a380),
	.w8(32'hb9a2fe80),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b0e944),
	.w1(32'hb6e182f6),
	.w2(32'hb6f9320e),
	.w3(32'h3771e89c),
	.w4(32'hb7ff2b33),
	.w5(32'h36bf4034),
	.w6(32'hb68cc140),
	.w7(32'h34377eee),
	.w8(32'h3798570c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ed4e05),
	.w1(32'h371b089d),
	.w2(32'hb8b7bb5a),
	.w3(32'hb8b1e34c),
	.w4(32'hb9113c88),
	.w5(32'hb8c1d088),
	.w6(32'hb5bed0f1),
	.w7(32'hb8518ba3),
	.w8(32'hb80cc177),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65047f),
	.w1(32'hbbaf72a8),
	.w2(32'hbb542b44),
	.w3(32'hbadf7445),
	.w4(32'hbb775f54),
	.w5(32'hbae90307),
	.w6(32'h3a2013e8),
	.w7(32'h3a307f31),
	.w8(32'hb9d321a2),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c452e9f),
	.w1(32'h3b8e4448),
	.w2(32'hba45965b),
	.w3(32'h3c0b53d1),
	.w4(32'h3c0d966b),
	.w5(32'h3b58760d),
	.w6(32'hbb4b8432),
	.w7(32'h3adaeb84),
	.w8(32'h3b3c3812),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa99b2),
	.w1(32'h3c0f1623),
	.w2(32'h3aefb436),
	.w3(32'h3aef17f4),
	.w4(32'h3b49ffb7),
	.w5(32'hba971364),
	.w6(32'hbb9b4b2a),
	.w7(32'hbb9caa86),
	.w8(32'hbb9690e4),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e19df),
	.w1(32'h3c1a2aca),
	.w2(32'h3b31a563),
	.w3(32'h3bbfc693),
	.w4(32'h3c0db9fb),
	.w5(32'h3a9e1239),
	.w6(32'hbb9fe4ba),
	.w7(32'hbb21f87d),
	.w8(32'hbaf105d6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3863c944),
	.w1(32'h380a036d),
	.w2(32'h38aef1ab),
	.w3(32'h38bf327f),
	.w4(32'h38a41c67),
	.w5(32'h38bbc2a9),
	.w6(32'h390106fe),
	.w7(32'h390b3afa),
	.w8(32'h38de2f9b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8185f),
	.w1(32'hb98fa01f),
	.w2(32'hb8f66905),
	.w3(32'h391a0f2f),
	.w4(32'h3a704953),
	.w5(32'h3a3e36a6),
	.w6(32'hb990f12a),
	.w7(32'hb897492a),
	.w8(32'h398b43df),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a2313f),
	.w1(32'hb744bdfd),
	.w2(32'hb736a3d4),
	.w3(32'hb73e8234),
	.w4(32'hb790de6a),
	.w5(32'hb75d7967),
	.w6(32'h3607f0a0),
	.w7(32'hb61b824d),
	.w8(32'hb5f6c412),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3715d208),
	.w1(32'h3477c500),
	.w2(32'hb7d79413),
	.w3(32'hb746820a),
	.w4(32'hb70cea9b),
	.w5(32'hb7f4168f),
	.w6(32'h37b5be0b),
	.w7(32'h3788cd2a),
	.w8(32'hb7984654),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c004cf0),
	.w1(32'h3ade9be4),
	.w2(32'hbb5b0ff4),
	.w3(32'h3b207a0d),
	.w4(32'h3b1b6537),
	.w5(32'hb8c6591b),
	.w6(32'hbb0898d3),
	.w7(32'hbb61e685),
	.w8(32'hbb918dce),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f1cb2),
	.w1(32'hb97b0b70),
	.w2(32'hb94b4c87),
	.w3(32'hb9309025),
	.w4(32'hb988142a),
	.w5(32'hb97efd08),
	.w6(32'hb9925191),
	.w7(32'hb9b32f64),
	.w8(32'hb9a82f44),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d7812a),
	.w1(32'h39eec518),
	.w2(32'h39af8b62),
	.w3(32'h39b01b86),
	.w4(32'h3a29f891),
	.w5(32'h39ce0c5b),
	.w6(32'h3965a3fd),
	.w7(32'h39d3b96e),
	.w8(32'h391211f9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fda74),
	.w1(32'hb997cf24),
	.w2(32'h3ace83a0),
	.w3(32'h3b6779e7),
	.w4(32'hb9d339bc),
	.w5(32'h3ad7fa09),
	.w6(32'h3b0055a5),
	.w7(32'h3a9209f4),
	.w8(32'h3afded02),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e4329),
	.w1(32'h38226e60),
	.w2(32'hb6acba57),
	.w3(32'hb6c9a1e4),
	.w4(32'hb6e4b05a),
	.w5(32'hb8576219),
	.w6(32'hb582c4ef),
	.w7(32'hb7c3f233),
	.w8(32'hb8630379),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19c72f),
	.w1(32'h3b127af1),
	.w2(32'h3a920762),
	.w3(32'h39c18e47),
	.w4(32'h39f1e04a),
	.w5(32'hb8e4b739),
	.w6(32'hba8f6821),
	.w7(32'hbacb2bbd),
	.w8(32'hbac74638),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb2d5e),
	.w1(32'h39583900),
	.w2(32'hb936c870),
	.w3(32'h399b2d9f),
	.w4(32'h3a042ac8),
	.w5(32'h399263b9),
	.w6(32'h3999fd02),
	.w7(32'h3a26b340),
	.w8(32'h39879700),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3477f),
	.w1(32'h3bb9d5c4),
	.w2(32'hbb3c5085),
	.w3(32'h3c5d268b),
	.w4(32'h3c5e723f),
	.w5(32'h3ae6af8c),
	.w6(32'h3b383e97),
	.w7(32'h3ab5d65b),
	.w8(32'h3a08b80e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9834281),
	.w1(32'h394f100c),
	.w2(32'h39d1b78b),
	.w3(32'hb973a62a),
	.w4(32'h397ed482),
	.w5(32'h39f9b198),
	.w6(32'hb8fa8cc7),
	.w7(32'hb8b17304),
	.w8(32'h37116673),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ec730),
	.w1(32'hbb8b6d0e),
	.w2(32'hbb8b1e22),
	.w3(32'hbb9893ab),
	.w4(32'hbc003314),
	.w5(32'hbbdcb942),
	.w6(32'h3b347b96),
	.w7(32'hbbbf1184),
	.w8(32'hbba928d1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule