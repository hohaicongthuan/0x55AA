module layer_10_featuremap_105(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba839c1a),
	.w1(32'hba172dd8),
	.w2(32'hbab11781),
	.w3(32'hba89f720),
	.w4(32'h3a426e33),
	.w5(32'hb9c38ebc),
	.w6(32'h3a2ad7dd),
	.w7(32'hb7d496c3),
	.w8(32'hba11d04b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d224f),
	.w1(32'hb986fceb),
	.w2(32'hb92f89b3),
	.w3(32'hbb800674),
	.w4(32'h39e73e1c),
	.w5(32'hb95b6cfc),
	.w6(32'hbaa8e6d4),
	.w7(32'h39ddad41),
	.w8(32'hba8d5a47),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39886fd3),
	.w1(32'h3948a59f),
	.w2(32'h39c26b1e),
	.w3(32'h39216414),
	.w4(32'h3884a353),
	.w5(32'hb93eeade),
	.w6(32'hb84da5f5),
	.w7(32'hb91f3fb8),
	.w8(32'hba02dc4b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf937c),
	.w1(32'h39f25c02),
	.w2(32'h3a1fa072),
	.w3(32'hb9a69774),
	.w4(32'hb9d8dadd),
	.w5(32'hb9a251eb),
	.w6(32'hba572acf),
	.w7(32'hba6ddab3),
	.w8(32'hba063e22),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cf1c45),
	.w1(32'hb93c2784),
	.w2(32'hb888f0e7),
	.w3(32'hb9e1b8b1),
	.w4(32'h3907da62),
	.w5(32'hba18aed5),
	.w6(32'hb933eb9d),
	.w7(32'hb9a9100f),
	.w8(32'h3a2dd0b9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab41416),
	.w1(32'hb9c7404f),
	.w2(32'hba72dbd2),
	.w3(32'hb8406d90),
	.w4(32'hba0eb23c),
	.w5(32'hbabdb2e4),
	.w6(32'hb9862294),
	.w7(32'hba3695f0),
	.w8(32'hba49ca54),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09bd87),
	.w1(32'hba9b9489),
	.w2(32'hbb494545),
	.w3(32'hbb1f5f0b),
	.w4(32'hba7c4d60),
	.w5(32'hbb1085e7),
	.w6(32'h3b362cf4),
	.w7(32'h39a3e89d),
	.w8(32'hbab64e05),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2d393),
	.w1(32'hbb102702),
	.w2(32'hbb737be7),
	.w3(32'hbbf4a08d),
	.w4(32'hbba786bc),
	.w5(32'hbae96dfc),
	.w6(32'hbbe587be),
	.w7(32'hbb8d6831),
	.w8(32'hbb0a66a3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9f306),
	.w1(32'hba6d38e6),
	.w2(32'hba77850e),
	.w3(32'hba8bcb44),
	.w4(32'hba89d5bf),
	.w5(32'hba809d63),
	.w6(32'hbaa3f08d),
	.w7(32'hba8fc818),
	.w8(32'hba663ba2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08f20),
	.w1(32'hbaa36b8b),
	.w2(32'hbba14905),
	.w3(32'hbbaac5bf),
	.w4(32'h38ec961a),
	.w5(32'hbad1d838),
	.w6(32'hbbb9234b),
	.w7(32'hba64c87d),
	.w8(32'hbb32cc3a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a638d4d),
	.w1(32'hba471707),
	.w2(32'hba240d13),
	.w3(32'h3a8eb1f5),
	.w4(32'hb90543e3),
	.w5(32'h38ba4d1a),
	.w6(32'hba59f6ed),
	.w7(32'hba897cfb),
	.w8(32'hba4d5a66),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55542d),
	.w1(32'h3a68fc62),
	.w2(32'hbb1c3365),
	.w3(32'hbb350b3f),
	.w4(32'h389c79f2),
	.w5(32'hbb072794),
	.w6(32'h3b09c9d0),
	.w7(32'h3b379a87),
	.w8(32'hba9d2a18),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc707),
	.w1(32'hbaf85bb8),
	.w2(32'hbbb6eef6),
	.w3(32'hbbc08734),
	.w4(32'hbb13de8b),
	.w5(32'hbb1cf60a),
	.w6(32'hbbb96d2d),
	.w7(32'hbb36abaa),
	.w8(32'hbb65079f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da84e5),
	.w1(32'hba0695de),
	.w2(32'hb9ceb95d),
	.w3(32'hb90c5f7e),
	.w4(32'hb8cb6fe3),
	.w5(32'hb82245b5),
	.w6(32'hb9d65a11),
	.w7(32'hb9b81d50),
	.w8(32'h39a4f6df),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb013bdb),
	.w1(32'hba7740aa),
	.w2(32'hbac67e09),
	.w3(32'hba9d3870),
	.w4(32'h3a84f20a),
	.w5(32'hba3095ad),
	.w6(32'hbb618491),
	.w7(32'h39874db1),
	.w8(32'hbac581f1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5d3a8),
	.w1(32'hbb84e4c7),
	.w2(32'hbbfa5212),
	.w3(32'hbb892426),
	.w4(32'hb9bb9443),
	.w5(32'hbb6b4433),
	.w6(32'hbbccc64d),
	.w7(32'hbb244a66),
	.w8(32'hbb8818b6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba253946),
	.w1(32'hba21680c),
	.w2(32'hb9ecbbdc),
	.w3(32'hb9f8b7d3),
	.w4(32'h3998443c),
	.w5(32'hb8b9b3f5),
	.w6(32'h39a15caf),
	.w7(32'h38b4f31b),
	.w8(32'h3a115113),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b865),
	.w1(32'hbaf681f1),
	.w2(32'hbbd49e1a),
	.w3(32'hbbb21b62),
	.w4(32'h399c68f8),
	.w5(32'hb9d8b7e7),
	.w6(32'hbbbbe5e8),
	.w7(32'hbaa81d96),
	.w8(32'hba54f2a9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb068934),
	.w1(32'hbab00a61),
	.w2(32'hbb73fd74),
	.w3(32'hbb1ddf5a),
	.w4(32'hba9ea874),
	.w5(32'hbb22cf9b),
	.w6(32'hbb9422ce),
	.w7(32'hbb323b28),
	.w8(32'hbb2f473d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bae7c6),
	.w1(32'hb9ab020c),
	.w2(32'hb9e20356),
	.w3(32'hb8c443d4),
	.w4(32'hb9b07b48),
	.w5(32'hb9bab302),
	.w6(32'hb9b46e00),
	.w7(32'hb9bf6784),
	.w8(32'hb943dfd3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994d072),
	.w1(32'h3a50ab37),
	.w2(32'h3a43ecbb),
	.w3(32'hb94ba8a4),
	.w4(32'h3a56a6ff),
	.w5(32'h3a53b0d2),
	.w6(32'h3a61945c),
	.w7(32'h3a5a52ef),
	.w8(32'h3a844457),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8682ff),
	.w1(32'h3a5cb82f),
	.w2(32'h3970a566),
	.w3(32'h3a6c0121),
	.w4(32'h3ab21580),
	.w5(32'h39f45e6e),
	.w6(32'h3a011a2d),
	.w7(32'h3b0f071f),
	.w8(32'hba724e09),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a5073),
	.w1(32'hb8f1cfae),
	.w2(32'hbc0b26ce),
	.w3(32'hbb9ee1fd),
	.w4(32'h3b224056),
	.w5(32'hbb78ac18),
	.w6(32'hbb495a0c),
	.w7(32'h3b925cfe),
	.w8(32'h38010a80),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58a71a),
	.w1(32'hba6d9b6f),
	.w2(32'hbb7a980b),
	.w3(32'hba6ffafc),
	.w4(32'h3a7d7be6),
	.w5(32'hbae96693),
	.w6(32'hbb349ccc),
	.w7(32'h3abf34d2),
	.w8(32'hbaa90839),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba63bd5),
	.w1(32'h3b129a6d),
	.w2(32'h39205957),
	.w3(32'hbbb5a9ca),
	.w4(32'h3a830eb4),
	.w5(32'hba454ae7),
	.w6(32'hbbeda0e3),
	.w7(32'h3a89191b),
	.w8(32'hb99ffab4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a64b62),
	.w1(32'hbae69b6f),
	.w2(32'hbad24a45),
	.w3(32'hb91fe89e),
	.w4(32'hb93f6bb5),
	.w5(32'hba2306d9),
	.w6(32'hbac2f03d),
	.w7(32'hbb01e1c8),
	.w8(32'hbaf05b4f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab118f7),
	.w1(32'hb9dd2025),
	.w2(32'hb9f87895),
	.w3(32'hba07f1b8),
	.w4(32'hb9a5d18d),
	.w5(32'hb9a52e51),
	.w6(32'hb987d885),
	.w7(32'hb9b58e1b),
	.w8(32'hb95c2b3a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02bb93),
	.w1(32'hba27e382),
	.w2(32'hbad4cbd0),
	.w3(32'hbaf31a1d),
	.w4(32'hbb79c799),
	.w5(32'hbb691d68),
	.w6(32'hbbe8fc4d),
	.w7(32'hbb8db810),
	.w8(32'hbb47c179),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb204936),
	.w1(32'h398ae4db),
	.w2(32'hb9b89d90),
	.w3(32'hbb1f515c),
	.w4(32'hba09c579),
	.w5(32'hba636844),
	.w6(32'hb9d71951),
	.w7(32'h3aeae045),
	.w8(32'h3aa4f606),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bbf1a),
	.w1(32'h3b1241be),
	.w2(32'h3a97da6f),
	.w3(32'hbb3a88a2),
	.w4(32'hba74a133),
	.w5(32'hbb0c6216),
	.w6(32'hbbf8c9ef),
	.w7(32'hbb6132bb),
	.w8(32'hbb6b9659),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392548e3),
	.w1(32'h39bee4f3),
	.w2(32'h39294a2a),
	.w3(32'h390a1731),
	.w4(32'h39fef86a),
	.w5(32'h39aef908),
	.w6(32'h39f85cf8),
	.w7(32'h39ce2d97),
	.w8(32'h39e1db2b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377089d8),
	.w1(32'hb946d365),
	.w2(32'hb8a6a041),
	.w3(32'h39cbfb14),
	.w4(32'h384082b9),
	.w5(32'hb86a79b4),
	.w6(32'hb8e560ea),
	.w7(32'h381922ea),
	.w8(32'hb827f3a2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6752c),
	.w1(32'hbaa0445a),
	.w2(32'hbb5d1216),
	.w3(32'hba4703b6),
	.w4(32'hb88a2acb),
	.w5(32'hbad42a1c),
	.w6(32'hbaec35eb),
	.w7(32'hba16fc9f),
	.w8(32'h373604ad),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabea2d9),
	.w1(32'hb9a16c8b),
	.w2(32'hba692837),
	.w3(32'hba9ba965),
	.w4(32'hb9b51c84),
	.w5(32'hb9ab0f3d),
	.w6(32'hbb0d194f),
	.w7(32'hb8b9e8a7),
	.w8(32'hbaad1957),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba545ba3),
	.w1(32'hb808c32e),
	.w2(32'hb93bb8a8),
	.w3(32'hba7b56a7),
	.w4(32'hb8acb784),
	.w5(32'h370141c3),
	.w6(32'hb9b61fa8),
	.w7(32'h3a04caeb),
	.w8(32'h395c27f6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e5b43),
	.w1(32'hba826e27),
	.w2(32'hbb176480),
	.w3(32'hba962e43),
	.w4(32'hbac4c2d7),
	.w5(32'hbaed0b54),
	.w6(32'h3acc8584),
	.w7(32'h3998b127),
	.w8(32'hba7b9687),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13d870),
	.w1(32'h39d16d96),
	.w2(32'hbb98bdba),
	.w3(32'hbbf195ca),
	.w4(32'h3b11d4e4),
	.w5(32'hb7b727e1),
	.w6(32'hbb8e8e8f),
	.w7(32'h3b7587b9),
	.w8(32'hbb3c1d38),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd527c),
	.w1(32'h3b5153af),
	.w2(32'h3b5634ab),
	.w3(32'hbb854d03),
	.w4(32'h3ba327a3),
	.w5(32'h3a90c803),
	.w6(32'hbaefe7ab),
	.w7(32'h3c076a32),
	.w8(32'h3b1d221b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac5e69),
	.w1(32'h3bb68131),
	.w2(32'h3b9ba7f8),
	.w3(32'hbaea0d0a),
	.w4(32'h3b0be6ce),
	.w5(32'hbaaf6fe0),
	.w6(32'hbb0d358e),
	.w7(32'h3b449357),
	.w8(32'hb953760c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05653e),
	.w1(32'h3a80ac5f),
	.w2(32'h3aac787a),
	.w3(32'hbaf968b3),
	.w4(32'h3a3b7da0),
	.w5(32'h3a50a18c),
	.w6(32'hba7b07e0),
	.w7(32'h3a714829),
	.w8(32'h39ed00c1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f2ffb),
	.w1(32'h3685a2e7),
	.w2(32'hb956cdc2),
	.w3(32'h37b7ebb3),
	.w4(32'h39c34c5d),
	.w5(32'h398dac55),
	.w6(32'h396b7319),
	.w7(32'h370c7dab),
	.w8(32'h3a292a46),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39650195),
	.w1(32'h38bac6e7),
	.w2(32'h39fee175),
	.w3(32'h39aa4640),
	.w4(32'h3a09bb5d),
	.w5(32'h39edf7c3),
	.w6(32'h39b78c13),
	.w7(32'hb753db17),
	.w8(32'hb8aa4aa4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9cb3a),
	.w1(32'h3a25487a),
	.w2(32'hb9b60655),
	.w3(32'hbaf92338),
	.w4(32'h398fcaeb),
	.w5(32'hba82844c),
	.w6(32'hba5b4548),
	.w7(32'h3a92a685),
	.w8(32'hbab11828),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfc14d),
	.w1(32'hbb1e31d0),
	.w2(32'hbbdccbda),
	.w3(32'hbbdc3c92),
	.w4(32'h32e9c200),
	.w5(32'hbb069cb4),
	.w6(32'hbc0b43d1),
	.w7(32'hbb2043b8),
	.w8(32'hbb386c78),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7bd4d),
	.w1(32'h3abbba1f),
	.w2(32'hb9ae6a05),
	.w3(32'hb947e42f),
	.w4(32'h3b0a7829),
	.w5(32'hba066b48),
	.w6(32'hbadecd9a),
	.w7(32'h3b6a58b6),
	.w8(32'h3987f498),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ca968),
	.w1(32'hba8991b9),
	.w2(32'hbb68c4b9),
	.w3(32'hba9adeb1),
	.w4(32'h3a386a7a),
	.w5(32'hba61531a),
	.w6(32'hbb67545b),
	.w7(32'h3ab19348),
	.w8(32'hbb005c79),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb13a),
	.w1(32'hbaf262ee),
	.w2(32'hbb130449),
	.w3(32'hbb55bcb2),
	.w4(32'h3985b659),
	.w5(32'hb91f9189),
	.w6(32'hbb56cf81),
	.w7(32'h3a84ebfb),
	.w8(32'hb9de5e88),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d68c2),
	.w1(32'hba924726),
	.w2(32'hbbb422c1),
	.w3(32'hbbb95977),
	.w4(32'hbb048785),
	.w5(32'hba8a1d23),
	.w6(32'hbbca292e),
	.w7(32'hbb9a996c),
	.w8(32'hba7b6f0b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fabef),
	.w1(32'hb9200040),
	.w2(32'h398a0bd5),
	.w3(32'h39f62d35),
	.w4(32'hb82f9445),
	.w5(32'h39a96149),
	.w6(32'hb9b7d721),
	.w7(32'hb974644e),
	.w8(32'h3839b64c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fec641),
	.w1(32'hba0d7dfa),
	.w2(32'hba0cd9f4),
	.w3(32'hba288d99),
	.w4(32'hb9fcfc89),
	.w5(32'hba137c22),
	.w6(32'hbaa4ee19),
	.w7(32'hbad14209),
	.w8(32'hba859a72),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883552f),
	.w1(32'h3a4420fc),
	.w2(32'h3a792564),
	.w3(32'h38daa5b5),
	.w4(32'h3a5f686a),
	.w5(32'h3a8de949),
	.w6(32'h3a528416),
	.w7(32'h3a4669ff),
	.w8(32'h3a510c4a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5373a),
	.w1(32'hb9a48bc4),
	.w2(32'hbb694481),
	.w3(32'hb96d2aaf),
	.w4(32'hba99bce5),
	.w5(32'hbafe8a31),
	.w6(32'hbaf23bfa),
	.w7(32'hba64ffc1),
	.w8(32'hbb15ec8d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8344a),
	.w1(32'h3a301c94),
	.w2(32'hba96a5ea),
	.w3(32'hba8eb297),
	.w4(32'h3a604676),
	.w5(32'hba65a701),
	.w6(32'h3a90194b),
	.w7(32'h3a4b36d1),
	.w8(32'h3a06bc11),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba45441),
	.w1(32'hbb5377a8),
	.w2(32'hbc12d3fe),
	.w3(32'hbb7c5e61),
	.w4(32'hb8eda366),
	.w5(32'hbb793676),
	.w6(32'hbb9a837d),
	.w7(32'hbaf28cc0),
	.w8(32'hbb51f743),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974fe86),
	.w1(32'hb92e67c8),
	.w2(32'hba55665d),
	.w3(32'h38513759),
	.w4(32'h38b4d068),
	.w5(32'hb9809ab0),
	.w6(32'h3a5245ca),
	.w7(32'h3a40df09),
	.w8(32'h39cba9e9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994412b),
	.w1(32'h3a4ca2e3),
	.w2(32'h3986b776),
	.w3(32'h3934d6b5),
	.w4(32'h3a2ab93b),
	.w5(32'h39992ec9),
	.w6(32'h3a507fc2),
	.w7(32'h39b3b425),
	.w8(32'h3a29a480),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e32b7),
	.w1(32'h3a245da0),
	.w2(32'h3a432d15),
	.w3(32'hb93cabfd),
	.w4(32'h3a28fcec),
	.w5(32'h3a349735),
	.w6(32'h3a38945a),
	.w7(32'h3a373f19),
	.w8(32'h39f456e8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e1d3a),
	.w1(32'h39ab53a9),
	.w2(32'hb9c41835),
	.w3(32'h3a7f6e9b),
	.w4(32'hb9b24e1c),
	.w5(32'hba22c288),
	.w6(32'hba4f0f6a),
	.w7(32'hba4f8f0b),
	.w8(32'hb9c04bf7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c2386e),
	.w1(32'h3a7057ed),
	.w2(32'h3a8dc629),
	.w3(32'hba43e91a),
	.w4(32'h3a0b72a7),
	.w5(32'h39c0e0b2),
	.w6(32'h39546178),
	.w7(32'h3a8244cb),
	.w8(32'h39a488ba),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9130dce),
	.w1(32'hba65c1a9),
	.w2(32'hba51283d),
	.w3(32'hb9243b4b),
	.w4(32'hba3e84f2),
	.w5(32'hba4f8dea),
	.w6(32'hba761ef6),
	.w7(32'hba8246d7),
	.w8(32'hba806182),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7907cf),
	.w1(32'hba833596),
	.w2(32'hbb15be44),
	.w3(32'hbb4a4212),
	.w4(32'hba022cb0),
	.w5(32'hba924d06),
	.w6(32'hbb002d50),
	.w7(32'h389af8de),
	.w8(32'hba5a6de0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb434d27),
	.w1(32'hbadf1ee9),
	.w2(32'hbb499a76),
	.w3(32'hbafdfdc4),
	.w4(32'h38739a54),
	.w5(32'hba87d514),
	.w6(32'hbb885a81),
	.w7(32'hb9be2f9a),
	.w8(32'hba8110a9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b51c4),
	.w1(32'hba860aa3),
	.w2(32'hbaa84cb7),
	.w3(32'hb9b6be48),
	.w4(32'hbac41593),
	.w5(32'hbabeef2d),
	.w6(32'hb9c19ffd),
	.w7(32'hba1c3c26),
	.w8(32'h3a4e2695),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d894d),
	.w1(32'h3a45e414),
	.w2(32'h3a49c5f1),
	.w3(32'h3861967b),
	.w4(32'h3a21f13e),
	.w5(32'h3a1cd3a6),
	.w6(32'h3a7271bd),
	.w7(32'h3a53192a),
	.w8(32'h3a96e23b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94e0c2),
	.w1(32'hb955b77d),
	.w2(32'h3821aca3),
	.w3(32'h3a71167f),
	.w4(32'hb9078962),
	.w5(32'hb79e5a30),
	.w6(32'hb95b16c8),
	.w7(32'hb8de215c),
	.w8(32'hb9b0235e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8093fdb),
	.w1(32'hb9546a8d),
	.w2(32'hb9665fe6),
	.w3(32'h36ace964),
	.w4(32'hb9d920c8),
	.w5(32'h38d9e00f),
	.w6(32'hba1f9ed9),
	.w7(32'hba029321),
	.w8(32'hba4854a3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccf537),
	.w1(32'hbbcb8998),
	.w2(32'hbc26f952),
	.w3(32'hbbc53042),
	.w4(32'hba40fdc6),
	.w5(32'hbaa49fa6),
	.w6(32'hbc0c0167),
	.w7(32'hbb525537),
	.w8(32'hba9cc2c7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad978a),
	.w1(32'hb9da0708),
	.w2(32'hbb554499),
	.w3(32'hbadeacb0),
	.w4(32'h3b1dd745),
	.w5(32'h38c12cf0),
	.w6(32'h3be10bc4),
	.w7(32'h3bdef111),
	.w8(32'h3a622cce),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7b241),
	.w1(32'hba9ffb17),
	.w2(32'hbb92b18c),
	.w3(32'hba597fd9),
	.w4(32'h3b06d40f),
	.w5(32'hb9d2d91c),
	.w6(32'h39821efa),
	.w7(32'h3b9a7b1e),
	.w8(32'h3abe5787),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba39206),
	.w1(32'h3bb5f489),
	.w2(32'h3aa6222f),
	.w3(32'hbbaae6cf),
	.w4(32'h3b7b89f7),
	.w5(32'hb9f9bec6),
	.w6(32'hbbd002f0),
	.w7(32'h3bc24ad9),
	.w8(32'hba9f7cff),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edc4eb),
	.w1(32'h39d0b0dc),
	.w2(32'h3a2acf96),
	.w3(32'h3aa6e71c),
	.w4(32'h3995a42b),
	.w5(32'h39b21484),
	.w6(32'h3a036f4f),
	.w7(32'h3a01a63d),
	.w8(32'h3996f459),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd72a3),
	.w1(32'hba230e0f),
	.w2(32'hba10a689),
	.w3(32'h39c29ce1),
	.w4(32'hba09efa2),
	.w5(32'hba24502a),
	.w6(32'hba24e1e5),
	.w7(32'hba5f13fb),
	.w8(32'hba2b44e4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4be7b),
	.w1(32'hba424d09),
	.w2(32'hba3241eb),
	.w3(32'hba0226b8),
	.w4(32'hba281782),
	.w5(32'hba4eb608),
	.w6(32'hba3d3c27),
	.w7(32'hba8a23a4),
	.w8(32'hba745bd8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2b343),
	.w1(32'hb9008c8d),
	.w2(32'hba6f067c),
	.w3(32'hbaaf4b04),
	.w4(32'h3a512ae3),
	.w5(32'h3a10dd9f),
	.w6(32'hba8b1f7f),
	.w7(32'h3a0d1c60),
	.w8(32'hb98cfc72),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99546ce),
	.w1(32'h39da551b),
	.w2(32'h3a1e598a),
	.w3(32'hb91a1564),
	.w4(32'h392b05e7),
	.w5(32'h3981cf95),
	.w6(32'h3981ff5b),
	.w7(32'h3987f938),
	.w8(32'h394bdaa5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b645f),
	.w1(32'hbb2a6132),
	.w2(32'hbb2efc1b),
	.w3(32'hbb24e448),
	.w4(32'hbab90e2d),
	.w5(32'h39c9558e),
	.w6(32'hbb3f148c),
	.w7(32'hbafc92ba),
	.w8(32'h39e441e6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ee90),
	.w1(32'hbb1b0513),
	.w2(32'hbb88c5b2),
	.w3(32'hbb93dc1e),
	.w4(32'hbb044ac0),
	.w5(32'hbb21d35e),
	.w6(32'hbb3c756b),
	.w7(32'h395084f2),
	.w8(32'hbacfe8b1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926ed8),
	.w1(32'hb9979cca),
	.w2(32'hbacfc0c2),
	.w3(32'hbbbb3f87),
	.w4(32'hbaea52db),
	.w5(32'hbacdc6b2),
	.w6(32'hbbec8e83),
	.w7(32'hbb3adecd),
	.w8(32'hbae9fc8b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab365b4),
	.w1(32'hba33ea44),
	.w2(32'hbb0261ca),
	.w3(32'hbab64393),
	.w4(32'h3a6e2038),
	.w5(32'h39e22939),
	.w6(32'hbae6edb8),
	.w7(32'hb9df99ad),
	.w8(32'hb9b00119),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba698e),
	.w1(32'hba8742dd),
	.w2(32'hbb3b160b),
	.w3(32'hbabf4ec6),
	.w4(32'h39ffaf8f),
	.w5(32'h389438d3),
	.w6(32'hbad82c43),
	.w7(32'hb941282a),
	.w8(32'hb9a2aa3c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81d9a1),
	.w1(32'h3a0da54d),
	.w2(32'hba97bd7d),
	.w3(32'h37cb1827),
	.w4(32'h3a8cc04d),
	.w5(32'hba0ce461),
	.w6(32'hb9ee2499),
	.w7(32'h3ac51ac4),
	.w8(32'h3961c216),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade4358),
	.w1(32'hb91d5464),
	.w2(32'hbb0eb4e9),
	.w3(32'hbaaa2d5f),
	.w4(32'hb99faa1e),
	.w5(32'hba6299e7),
	.w6(32'hba83daee),
	.w7(32'hba28cedd),
	.w8(32'hb765bc3b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fa985d),
	.w1(32'h398aaaf0),
	.w2(32'h378c39d3),
	.w3(32'hb97acf2a),
	.w4(32'h39c10bae),
	.w5(32'hb7152b9b),
	.w6(32'h3a0b427a),
	.w7(32'h394fc4e5),
	.w8(32'h3a22db62),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60c9c1f),
	.w1(32'h3921818c),
	.w2(32'h39b296d2),
	.w3(32'h3903388a),
	.w4(32'h38b8ed3f),
	.w5(32'h39690136),
	.w6(32'h38062427),
	.w7(32'h39140bc4),
	.w8(32'hb9285583),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b391f6),
	.w1(32'h3a977b9a),
	.w2(32'h3a9ef60c),
	.w3(32'hb963e647),
	.w4(32'hba00f914),
	.w5(32'hb7fb37b5),
	.w6(32'h3a3e05b3),
	.w7(32'h3a98ad71),
	.w8(32'h39bfeef5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d8787),
	.w1(32'h3ab99894),
	.w2(32'h3aacbad4),
	.w3(32'hb989f383),
	.w4(32'h3a8985ca),
	.w5(32'h3a91482f),
	.w6(32'h3a5166db),
	.w7(32'h3a54aee4),
	.w8(32'h3a698209),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb716d0c),
	.w1(32'hb9cd0ff4),
	.w2(32'h3a30f4f6),
	.w3(32'hbb320186),
	.w4(32'h3ac9fb16),
	.w5(32'h3ad36f3f),
	.w6(32'hbb17e498),
	.w7(32'h3b11de41),
	.w8(32'h3a1d07b9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920821c),
	.w1(32'h3a81ae03),
	.w2(32'h39e4ff2e),
	.w3(32'hb86a7c01),
	.w4(32'h3a5e1cab),
	.w5(32'h390924c0),
	.w6(32'h399ad051),
	.w7(32'h3a531977),
	.w8(32'h39f9f0ef),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa26106),
	.w1(32'h3979e437),
	.w2(32'hba8faa3b),
	.w3(32'hba03aed7),
	.w4(32'h3a6d75dd),
	.w5(32'hb9abe49a),
	.w6(32'hba255be8),
	.w7(32'h3aa06930),
	.w8(32'hba26c848),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87581c),
	.w1(32'hba0f9059),
	.w2(32'hbb8e013e),
	.w3(32'hbb79f403),
	.w4(32'h3932c0b5),
	.w5(32'h398e71ef),
	.w6(32'hbbabb2e2),
	.w7(32'hba192c42),
	.w8(32'h3a6d2d13),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15dc08),
	.w1(32'h3b467cb0),
	.w2(32'h3abb671e),
	.w3(32'hba1c93a9),
	.w4(32'h3b05d078),
	.w5(32'hba215347),
	.w6(32'hb9ddf525),
	.w7(32'h3b34c0c5),
	.w8(32'h391a3693),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04c9b5),
	.w1(32'hbb77d3e9),
	.w2(32'hbbb09511),
	.w3(32'hbb9e1306),
	.w4(32'hb9bc46e2),
	.w5(32'hbb18f5a7),
	.w6(32'h39d258f1),
	.w7(32'h3ad7a545),
	.w8(32'hba7275ce),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b187fcd),
	.w1(32'h3b950aa1),
	.w2(32'h3b0eacb7),
	.w3(32'h3b052ffb),
	.w4(32'h3b87ed98),
	.w5(32'h3ac519e8),
	.w6(32'h3b093fbc),
	.w7(32'h3b87df14),
	.w8(32'h3b1f0243),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8902a3),
	.w1(32'hbade9d7a),
	.w2(32'hbb951dca),
	.w3(32'hbb07ffe4),
	.w4(32'h3acce058),
	.w5(32'h3a23ae6a),
	.w6(32'hb91dc658),
	.w7(32'h3addc8d6),
	.w8(32'h399f3b77),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ea39c),
	.w1(32'hba79d511),
	.w2(32'hbac4db43),
	.w3(32'hbaa52cf6),
	.w4(32'h3afd1238),
	.w5(32'h39c5a306),
	.w6(32'hbaf25055),
	.w7(32'h3a3b4b09),
	.w8(32'hba99d1dd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1850ea),
	.w1(32'h39a99d6a),
	.w2(32'hba572767),
	.w3(32'hbb27eda3),
	.w4(32'h3ab52230),
	.w5(32'hba3cb7b9),
	.w6(32'hbbb60db4),
	.w7(32'hb9db6c31),
	.w8(32'hbaae3168),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e97160),
	.w1(32'h3aa766d6),
	.w2(32'h3aabf8a0),
	.w3(32'h3a3dd8c4),
	.w4(32'h3a8683e8),
	.w5(32'h3ac3d2c8),
	.w6(32'h3a7e4242),
	.w7(32'h3ae31fe7),
	.w8(32'h3a6cdc64),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb652f94),
	.w1(32'hbaa81d6d),
	.w2(32'hbbe50e08),
	.w3(32'hbb2fdd05),
	.w4(32'hb7a2bf58),
	.w5(32'hbb3c9417),
	.w6(32'hbb9df2a4),
	.w7(32'hbb04ad16),
	.w8(32'hbb5ba223),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3360d),
	.w1(32'hbb53cc36),
	.w2(32'hbb9fed0c),
	.w3(32'hbb703bd6),
	.w4(32'h3a2e0de6),
	.w5(32'h3916ad86),
	.w6(32'hba5bbab5),
	.w7(32'h3b0935ad),
	.w8(32'h39b179f3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1e3ae),
	.w1(32'h3b6fbb47),
	.w2(32'hbb46092a),
	.w3(32'hbbea43a5),
	.w4(32'h39888d61),
	.w5(32'hbb074d59),
	.w6(32'h3a1381be),
	.w7(32'h3ba0d5c0),
	.w8(32'h3b2624d6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ce2ec),
	.w1(32'h3bc4a13d),
	.w2(32'h3b88fc90),
	.w3(32'hbb32a7ce),
	.w4(32'h3be963f7),
	.w5(32'h3ba056f9),
	.w6(32'hba169995),
	.w7(32'h3bc9d822),
	.w8(32'h3b881943),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35869c),
	.w1(32'h3a5d2799),
	.w2(32'hbb151f86),
	.w3(32'hbb53536d),
	.w4(32'hba969ab7),
	.w5(32'hbb1cfd7a),
	.w6(32'hbbd67c7b),
	.w7(32'hbab223cc),
	.w8(32'hbb7bc1fa),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3477e),
	.w1(32'hbb340235),
	.w2(32'hbbc665e2),
	.w3(32'hbb623b41),
	.w4(32'h3aae6260),
	.w5(32'hba5a2a53),
	.w6(32'hba8d9abb),
	.w7(32'hb9b40010),
	.w8(32'hba8ba3ca),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a16a9),
	.w1(32'h38296a47),
	.w2(32'hb90226aa),
	.w3(32'h3a61b5ea),
	.w4(32'h3a38b2f4),
	.w5(32'hb846474f),
	.w6(32'h39a49792),
	.w7(32'h3a11d517),
	.w8(32'h3a04f29d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15eab5),
	.w1(32'hbbb40c78),
	.w2(32'hbb96b253),
	.w3(32'hbbd86914),
	.w4(32'h39d4f0a5),
	.w5(32'hba916976),
	.w6(32'hbbd27b48),
	.w7(32'h3a611ca7),
	.w8(32'hbb124520),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99cc91),
	.w1(32'hbb265ace),
	.w2(32'hbac0fff3),
	.w3(32'hbbb57cc1),
	.w4(32'hbb934f60),
	.w5(32'hbb694ac4),
	.w6(32'hbafccaab),
	.w7(32'hbadc7c0c),
	.w8(32'hbb4049df),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b463c),
	.w1(32'h39775510),
	.w2(32'h39cea9d5),
	.w3(32'hb92023ab),
	.w4(32'h390d7da6),
	.w5(32'hb93b8dae),
	.w6(32'h38b54f58),
	.w7(32'h390ad357),
	.w8(32'hba1fe03a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad524e9),
	.w1(32'hba824287),
	.w2(32'hbaa0127d),
	.w3(32'hba19d408),
	.w4(32'h39728ff7),
	.w5(32'hb9f24d26),
	.w6(32'h37b44d05),
	.w7(32'h3a34ed72),
	.w8(32'h3a4bdd92),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36c365),
	.w1(32'hbab73cd4),
	.w2(32'hbb7fdfe7),
	.w3(32'hbb6f29f0),
	.w4(32'hbb258b82),
	.w5(32'hbb32c5b0),
	.w6(32'hbbb22938),
	.w7(32'hbb995880),
	.w8(32'hbb870431),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00ac86),
	.w1(32'h3a11e632),
	.w2(32'hb9ebaa67),
	.w3(32'hbb162f2c),
	.w4(32'hba32287f),
	.w5(32'hbaf44fad),
	.w6(32'hbb9dafbb),
	.w7(32'hba9f2340),
	.w8(32'hbb18facd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8934b),
	.w1(32'hba6bde84),
	.w2(32'hbb278fab),
	.w3(32'hbb4b3ed7),
	.w4(32'hba99b05b),
	.w5(32'hbb4112a9),
	.w6(32'hbbb77caa),
	.w7(32'hbac9cb6c),
	.w8(32'hbb745dbe),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1169ff),
	.w1(32'hba126996),
	.w2(32'hbae7facd),
	.w3(32'hbb21fd29),
	.w4(32'hba2185fd),
	.w5(32'hbac8874e),
	.w6(32'hbb2a1a7b),
	.w7(32'hba64ada2),
	.w8(32'hba4f72b6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b58e0c),
	.w1(32'h3b1512be),
	.w2(32'h39d34634),
	.w3(32'hba4e74b5),
	.w4(32'h3a33f09a),
	.w5(32'hba61b710),
	.w6(32'h3b6f1336),
	.w7(32'h3ba6fd6f),
	.w8(32'h3b0896cf),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb456a1),
	.w1(32'hbb4f500d),
	.w2(32'hbbaf990a),
	.w3(32'hbb44a471),
	.w4(32'h397295ce),
	.w5(32'hbace49e8),
	.w6(32'hbb9da5bb),
	.w7(32'hbb35ff0b),
	.w8(32'hbb5bb479),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee95f4),
	.w1(32'h3873396d),
	.w2(32'hba778a60),
	.w3(32'hbb03d65d),
	.w4(32'h38f5f954),
	.w5(32'hba5568e3),
	.w6(32'hbaf24c9f),
	.w7(32'hb9817eb6),
	.w8(32'hb9ba6272),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a517bf0),
	.w1(32'hb935cc8e),
	.w2(32'hb9b18d3b),
	.w3(32'h3a24a04a),
	.w4(32'hb946c7a9),
	.w5(32'hba0d8f3c),
	.w6(32'hb93de44a),
	.w7(32'hb998d07e),
	.w8(32'hb87fbb2b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48d75a),
	.w1(32'hba229a2e),
	.w2(32'hba360c08),
	.w3(32'hba08f459),
	.w4(32'hba11d091),
	.w5(32'hba4044d5),
	.w6(32'hba0b2d25),
	.w7(32'hba3f3dc6),
	.w8(32'hba7c9237),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17fc66),
	.w1(32'hb88755dd),
	.w2(32'hb9a04824),
	.w3(32'hba323508),
	.w4(32'hb969834c),
	.w5(32'hba21d83d),
	.w6(32'hb9683fb0),
	.w7(32'hb9af40a5),
	.w8(32'hb9a9c5cb),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18fb06),
	.w1(32'hba84fcba),
	.w2(32'hba8fd174),
	.w3(32'hba2e7e14),
	.w4(32'hb9b038b3),
	.w5(32'hb9da393d),
	.w6(32'hb9d31e9a),
	.w7(32'hb9e8bc4b),
	.w8(32'hba823209),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e2c6f),
	.w1(32'h3a5ec157),
	.w2(32'hba319f8c),
	.w3(32'hba88a5d3),
	.w4(32'h3a8a1366),
	.w5(32'h3984fcb4),
	.w6(32'hbac721e0),
	.w7(32'h3ad138fd),
	.w8(32'hb994085c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0510a5),
	.w1(32'hb9c59365),
	.w2(32'hba5a234d),
	.w3(32'h399bfa4e),
	.w4(32'hb9be088c),
	.w5(32'hba8a8240),
	.w6(32'hba1060fd),
	.w7(32'hba28f0f4),
	.w8(32'hb9d8c08d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb255dbe),
	.w1(32'hb88e13a4),
	.w2(32'hbb1024b1),
	.w3(32'hbb386374),
	.w4(32'hba9d7100),
	.w5(32'hbaadee31),
	.w6(32'hb99cf7d5),
	.w7(32'hbabbf5f1),
	.w8(32'hba92c5c8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a4e90),
	.w1(32'h39b8dac0),
	.w2(32'hb99d3164),
	.w3(32'hbb701604),
	.w4(32'hb9a70032),
	.w5(32'hbaef55de),
	.w6(32'hbb9d0214),
	.w7(32'hba7a51c0),
	.w8(32'hbb5ff75c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d924c),
	.w1(32'hbaa54ce0),
	.w2(32'hbaa65fad),
	.w3(32'hba45e7b3),
	.w4(32'hb988dd0f),
	.w5(32'hb8afe89a),
	.w6(32'h36abce4c),
	.w7(32'h3a09b56c),
	.w8(32'hbae61d6c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bfa45),
	.w1(32'h3a2f6c1e),
	.w2(32'hb97f2a29),
	.w3(32'hb991dce3),
	.w4(32'h3a133a1f),
	.w5(32'hba1da292),
	.w6(32'h3ac20efe),
	.w7(32'h3a22d589),
	.w8(32'h3a932407),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8991c),
	.w1(32'hb81729f1),
	.w2(32'hb956c6bb),
	.w3(32'hb872bbe8),
	.w4(32'h39812668),
	.w5(32'h394b103a),
	.w6(32'h39bc5ad6),
	.w7(32'h396bc271),
	.w8(32'h399b477a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373405d2),
	.w1(32'hbc085b08),
	.w2(32'hbbea85ee),
	.w3(32'hba209a44),
	.w4(32'hbc67b0d5),
	.w5(32'hbc56e300),
	.w6(32'h3c5c0ca4),
	.w7(32'h3d22018e),
	.w8(32'h3c25caa7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01ead0),
	.w1(32'hbaf07ac9),
	.w2(32'hbcb8948f),
	.w3(32'hbb4b9b86),
	.w4(32'hbc222a6f),
	.w5(32'hbcf45ab0),
	.w6(32'h3c94bf0a),
	.w7(32'h3d3d9662),
	.w8(32'h3bf286b8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb08367),
	.w1(32'h3c4cc3ca),
	.w2(32'hba5f55d7),
	.w3(32'hbbefe591),
	.w4(32'h3c4704b5),
	.w5(32'h3c3e75c7),
	.w6(32'hbc3b379b),
	.w7(32'h3aeca433),
	.w8(32'h3a8a1178),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bf9d5),
	.w1(32'h39493083),
	.w2(32'h3c9bf408),
	.w3(32'hbbaab17c),
	.w4(32'hbbad2052),
	.w5(32'h3b43c6f6),
	.w6(32'h3b0b349c),
	.w7(32'hbc8f5121),
	.w8(32'hbbbae5bb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1daccc),
	.w1(32'hbc7d8488),
	.w2(32'hbbecc819),
	.w3(32'hbc83a69e),
	.w4(32'hbc630355),
	.w5(32'hbc7d938f),
	.w6(32'hbb0e338d),
	.w7(32'hbc2d5394),
	.w8(32'h3a632f71),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e74ed),
	.w1(32'hbc778bba),
	.w2(32'hbc7e51b7),
	.w3(32'hbc4cea24),
	.w4(32'h3c153723),
	.w5(32'h3a6a6e57),
	.w6(32'hbc8e93f4),
	.w7(32'hbb6f4b9d),
	.w8(32'hbb56c42d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc094a58),
	.w1(32'h3c208770),
	.w2(32'h3ab9ec3b),
	.w3(32'h3bc0c660),
	.w4(32'h3b4f535e),
	.w5(32'h39e6ccd6),
	.w6(32'h3c1d1bed),
	.w7(32'h3aa1d07a),
	.w8(32'hbbc8c076),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8683),
	.w1(32'h3b6ab6dc),
	.w2(32'hbcac08ba),
	.w3(32'h3b18d536),
	.w4(32'hbbafed0e),
	.w5(32'hbd07c0df),
	.w6(32'h3c623171),
	.w7(32'h3d27fd0b),
	.w8(32'h3beeb1a0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a59ad),
	.w1(32'hbbf5e13e),
	.w2(32'h3c35b047),
	.w3(32'hbc8e564f),
	.w4(32'hbbb6608e),
	.w5(32'h3a977f5c),
	.w6(32'hbb1f3a76),
	.w7(32'hbcd17de1),
	.w8(32'hbbfc35f3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf726f2),
	.w1(32'h3ab87971),
	.w2(32'hbcb991b8),
	.w3(32'hbc680f0c),
	.w4(32'hbc02a703),
	.w5(32'hbcdee643),
	.w6(32'h3c23fbb5),
	.w7(32'h3d4e28c2),
	.w8(32'h3c2411a6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bed16),
	.w1(32'hba0a22af),
	.w2(32'hbc0aa60d),
	.w3(32'hbae96b5a),
	.w4(32'hbb60a1ee),
	.w5(32'hbc5aa563),
	.w6(32'h3c67b131),
	.w7(32'h3cfc1ec3),
	.w8(32'hba05207e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f0a88),
	.w1(32'hbc1cffc1),
	.w2(32'h3ce409e9),
	.w3(32'h3b4a7ce9),
	.w4(32'h3bdd4b84),
	.w5(32'h3cfac92f),
	.w6(32'hbc911d88),
	.w7(32'hbd81b196),
	.w8(32'hbc86653d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc328e3c),
	.w1(32'hbc6f7152),
	.w2(32'hbcdeacbc),
	.w3(32'hba542de6),
	.w4(32'h3be98863),
	.w5(32'h3bb7e511),
	.w6(32'hbb64da8c),
	.w7(32'hbb73cb19),
	.w8(32'hbacb1e5a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89fd45),
	.w1(32'hbbca4dad),
	.w2(32'hbd0962fc),
	.w3(32'hbb828552),
	.w4(32'hbb7b418d),
	.w5(32'hbb0fdd4b),
	.w6(32'hba442f63),
	.w7(32'h3b739c02),
	.w8(32'hbbf865f4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc525262),
	.w1(32'h393b71a9),
	.w2(32'hbaff12e1),
	.w3(32'hba67ed2c),
	.w4(32'hbbfa09ca),
	.w5(32'hbc49b0ca),
	.w6(32'h3bcbd550),
	.w7(32'h3cc9032c),
	.w8(32'h3c0f2cdd),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ad864),
	.w1(32'h3b76eef5),
	.w2(32'hbca7a19d),
	.w3(32'hbbfac13e),
	.w4(32'hbae518b1),
	.w5(32'hbd0dae11),
	.w6(32'h3953d18e),
	.w7(32'h3d6b053c),
	.w8(32'h3c471138),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22fe98),
	.w1(32'h3a078255),
	.w2(32'hbcc6ead6),
	.w3(32'hb7c312ca),
	.w4(32'h3b37007c),
	.w5(32'h39052698),
	.w6(32'hb80b9cb0),
	.w7(32'hb992f7f9),
	.w8(32'hbace1f37),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc96dd5),
	.w1(32'h3ba85b3e),
	.w2(32'hbc1d0f84),
	.w3(32'hbc00aae9),
	.w4(32'hbb8b3bbb),
	.w5(32'hbc820978),
	.w6(32'h3c76ef59),
	.w7(32'h3cfcef4b),
	.w8(32'h3b3d05e7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dd1bc),
	.w1(32'hbb2fac66),
	.w2(32'hbbc4c77a),
	.w3(32'h39d59d55),
	.w4(32'hbc106129),
	.w5(32'hbc651d43),
	.w6(32'hbb62c82f),
	.w7(32'h3ba15268),
	.w8(32'h3b8d91da),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39352a),
	.w1(32'hbc1f0687),
	.w2(32'h3cd39dd9),
	.w3(32'hbbb9611e),
	.w4(32'hbafcf562),
	.w5(32'h3c8719e7),
	.w6(32'hbc75b3e1),
	.w7(32'hbd4a57ef),
	.w8(32'hbc5c3cda),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc473cf2),
	.w1(32'h3b3e4064),
	.w2(32'h3c0a18c6),
	.w3(32'hbc215d1f),
	.w4(32'h39d2fc31),
	.w5(32'h3ae2c711),
	.w6(32'hbaddaedb),
	.w7(32'hbc32cce1),
	.w8(32'hbb365c0f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f1c3d),
	.w1(32'h3b1ebc40),
	.w2(32'hbc248ca7),
	.w3(32'hbc2a9370),
	.w4(32'hbc1cffef),
	.w5(32'hbc76a29f),
	.w6(32'h3b99c9e5),
	.w7(32'h3c937e3c),
	.w8(32'hbb414c17),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1faf7),
	.w1(32'hbc13bc5d),
	.w2(32'hbce1fa34),
	.w3(32'hbb317136),
	.w4(32'h3b447f50),
	.w5(32'hbc7fe9d5),
	.w6(32'h3c1d29de),
	.w7(32'h3d2522c7),
	.w8(32'h3c0d395c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc829c78),
	.w1(32'hbcae512d),
	.w2(32'hbd318263),
	.w3(32'h3b653efb),
	.w4(32'h3b86a3d8),
	.w5(32'hbb0d6fcc),
	.w6(32'hbad9761b),
	.w7(32'hbba5ac16),
	.w8(32'hbbf1a8b2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5a17f),
	.w1(32'hba817159),
	.w2(32'h3b69d808),
	.w3(32'hbc243b46),
	.w4(32'h3bab1b07),
	.w5(32'h3b259091),
	.w6(32'hbc176c65),
	.w7(32'hbb4439ef),
	.w8(32'hbc007bf9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5af644),
	.w1(32'hbb1cde39),
	.w2(32'hbcf22f0d),
	.w3(32'h392d28e7),
	.w4(32'hbc089f80),
	.w5(32'hbce58f17),
	.w6(32'h3c2300a4),
	.w7(32'h3d43f99e),
	.w8(32'h3c21b3bd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a0b92a),
	.w1(32'h3b85896b),
	.w2(32'hbabd0e4d),
	.w3(32'hbb921015),
	.w4(32'hbb003be3),
	.w5(32'hbb3e373a),
	.w6(32'hbb57069a),
	.w7(32'h3b299e4f),
	.w8(32'hbade8552),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d8a5e),
	.w1(32'hbc474ee7),
	.w2(32'hbd171aad),
	.w3(32'h3ae364d9),
	.w4(32'hbbf78c0a),
	.w5(32'hbc5f6402),
	.w6(32'h39372ae7),
	.w7(32'hbb65844d),
	.w8(32'h3abb8783),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44b12b),
	.w1(32'hb9a9b40f),
	.w2(32'hbc8693ec),
	.w3(32'hb9e58467),
	.w4(32'hbbc6aebb),
	.w5(32'hbc86d2b1),
	.w6(32'h3c03bcf9),
	.w7(32'h3cb72a71),
	.w8(32'h3bd24d80),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd976d),
	.w1(32'h3c025c52),
	.w2(32'h3b5d3e41),
	.w3(32'hbbfd0953),
	.w4(32'h3b0703ba),
	.w5(32'h3a0482e5),
	.w6(32'hbad97d62),
	.w7(32'hbbd619ae),
	.w8(32'hbc448f6e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc179095),
	.w1(32'hba962b7f),
	.w2(32'h3bea48d8),
	.w3(32'hbb49b4f5),
	.w4(32'hba3b68ab),
	.w5(32'hbb82c763),
	.w6(32'hbc6d33be),
	.w7(32'h3bdd4823),
	.w8(32'hbbf82295),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b089622),
	.w1(32'h3b2e6fd2),
	.w2(32'h38dd9440),
	.w3(32'hba814b1b),
	.w4(32'h3c1bbd14),
	.w5(32'h3b825214),
	.w6(32'hbb9184aa),
	.w7(32'h3a7650f2),
	.w8(32'h3b0b3791),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45640),
	.w1(32'h39e5b85a),
	.w2(32'hbc6fd120),
	.w3(32'h3b1c3650),
	.w4(32'hb6ff4399),
	.w5(32'hbc46a5be),
	.w6(32'h3c2dc6f4),
	.w7(32'h3cd2f233),
	.w8(32'h3c1b1f7f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf07307),
	.w1(32'h3a944b2a),
	.w2(32'hbc523ffd),
	.w3(32'h3accbc11),
	.w4(32'h3938623b),
	.w5(32'hbc16de47),
	.w6(32'h3c0a58da),
	.w7(32'h3cce8232),
	.w8(32'h3c17c065),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb916988),
	.w1(32'h39b90cd9),
	.w2(32'hbb8d2632),
	.w3(32'h3856d8dc),
	.w4(32'hbbbe13ad),
	.w5(32'hbb8dea70),
	.w6(32'h3b8ae873),
	.w7(32'h3c89e34b),
	.w8(32'h3c403f6b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6f6ea),
	.w1(32'h3bb67f96),
	.w2(32'h39a64c3d),
	.w3(32'hbb8f2b81),
	.w4(32'hbad989c6),
	.w5(32'hbb0f8df6),
	.w6(32'h3bef1c49),
	.w7(32'h3af74880),
	.w8(32'hbaa7a016),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb222354),
	.w1(32'hb9e1a2d5),
	.w2(32'h3cb43d6c),
	.w3(32'hbc4f87ba),
	.w4(32'h3c365eab),
	.w5(32'h3cdc87a7),
	.w6(32'hbbd482f6),
	.w7(32'hbd1ab405),
	.w8(32'hbc7d6833),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08af7a),
	.w1(32'hbb4220fe),
	.w2(32'hbcb2601e),
	.w3(32'h3bc4775a),
	.w4(32'hbacaae64),
	.w5(32'hbba96713),
	.w6(32'h3b701196),
	.w7(32'h3c96b044),
	.w8(32'h3b8e3998),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcab1e4),
	.w1(32'h3b504334),
	.w2(32'h3c9c87ce),
	.w3(32'h3ab8d4cd),
	.w4(32'hbb10a3a0),
	.w5(32'h3bb48e5b),
	.w6(32'h3b381288),
	.w7(32'hbc8963d1),
	.w8(32'hbbb1b8f8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57d4bb),
	.w1(32'hbbce4fbc),
	.w2(32'h3c4df134),
	.w3(32'hbc22d4c0),
	.w4(32'hbbb37c7e),
	.w5(32'h3abdbfd7),
	.w6(32'hbba45e68),
	.w7(32'hbccc4b06),
	.w8(32'hbbd1ff9f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f9f8c),
	.w1(32'hbaf22569),
	.w2(32'hbcbfe03b),
	.w3(32'hbc448ef7),
	.w4(32'hbc14dd4c),
	.w5(32'hbcd99398),
	.w6(32'h3c228fd2),
	.w7(32'h3d2a0bb0),
	.w8(32'h3bed3688),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5cd0b),
	.w1(32'h3a313fbc),
	.w2(32'h3c79c52d),
	.w3(32'hbbaab331),
	.w4(32'hbb9e70b2),
	.w5(32'h3ae11658),
	.w6(32'h3aaab5b8),
	.w7(32'hbc2814b5),
	.w8(32'hba2d91e4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823811),
	.w1(32'hbb830b44),
	.w2(32'hbbea71e4),
	.w3(32'hbc0bcc43),
	.w4(32'h3ba3f051),
	.w5(32'hbb18968e),
	.w6(32'hbbc37454),
	.w7(32'h3b5d9af4),
	.w8(32'h3ad83bb2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0691a6),
	.w1(32'h3abd6baa),
	.w2(32'hbb0e4dc7),
	.w3(32'hb8fd42a0),
	.w4(32'hbbf5d18d),
	.w5(32'hbba29bcd),
	.w6(32'h3c58a024),
	.w7(32'h3bdba47c),
	.w8(32'h3b801310),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfac06),
	.w1(32'h3b75f146),
	.w2(32'hbc162d51),
	.w3(32'hbc4556d6),
	.w4(32'hbb8b0901),
	.w5(32'hbc9b69b4),
	.w6(32'h3bd3bef6),
	.w7(32'h3ce04c71),
	.w8(32'h3bf2f87e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a776b57),
	.w1(32'hbc5d1243),
	.w2(32'h3d3338ba),
	.w3(32'hbb93d29f),
	.w4(32'h3c9c3094),
	.w5(32'h3d44e9f7),
	.w6(32'hbcec2ec2),
	.w7(32'hbd9e8ab5),
	.w8(32'hbc505a3a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6946f0),
	.w1(32'hbc35ffe9),
	.w2(32'h3bc9522d),
	.w3(32'hbb91cade),
	.w4(32'h3c00bf6f),
	.w5(32'h3c8e7496),
	.w6(32'hbc961cc6),
	.w7(32'hbc507d97),
	.w8(32'h3c39b024),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892ec5),
	.w1(32'hbbde7714),
	.w2(32'h3a8f8fb5),
	.w3(32'hb95bc0f1),
	.w4(32'h3b8fa1e4),
	.w5(32'h3c5917dd),
	.w6(32'h3a7f2b21),
	.w7(32'hbc1fe6c7),
	.w8(32'hbb5b5f25),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c51c),
	.w1(32'hbb4e76e5),
	.w2(32'hbc647af9),
	.w3(32'h3b86b645),
	.w4(32'h3b13d3bb),
	.w5(32'h3bfdb569),
	.w6(32'h3b2fc630),
	.w7(32'hbb77feef),
	.w8(32'hbc618a7e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9c18c),
	.w1(32'hbb08d88a),
	.w2(32'hbb031503),
	.w3(32'h3bd6f101),
	.w4(32'h3ac5fc24),
	.w5(32'hbb8d906a),
	.w6(32'hbb74fdc9),
	.w7(32'hba83e571),
	.w8(32'h3b00f5fb),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc2c49),
	.w1(32'h3abea93c),
	.w2(32'hbc307eeb),
	.w3(32'hbb804243),
	.w4(32'hbba501fb),
	.w5(32'hbc7ee83e),
	.w6(32'h3bc323ec),
	.w7(32'h3cc117ff),
	.w8(32'h3bfe2f5b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a826088),
	.w1(32'h3b2f07e8),
	.w2(32'hbc96bf08),
	.w3(32'hbb741c92),
	.w4(32'hbb840dfd),
	.w5(32'hbcbdb674),
	.w6(32'h3c37aad6),
	.w7(32'h3d375b49),
	.w8(32'h3c301919),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b631371),
	.w1(32'hbabe92a1),
	.w2(32'h3cdd5d9f),
	.w3(32'hba8ac764),
	.w4(32'h3b6594ff),
	.w5(32'h3c6abda2),
	.w6(32'hbc39a8b7),
	.w7(32'hbcc76ea6),
	.w8(32'hbbe4d6d2),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec3580),
	.w1(32'hba522871),
	.w2(32'hbb9478ea),
	.w3(32'h3b4b216e),
	.w4(32'hbbcb8f61),
	.w5(32'h3b1cb0d0),
	.w6(32'h3a60e470),
	.w7(32'h3bc4af80),
	.w8(32'hbbec45e7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905ceb3),
	.w1(32'hba998f6b),
	.w2(32'hbca67be1),
	.w3(32'hbb7dec67),
	.w4(32'hbc7038ac),
	.w5(32'hbd15f050),
	.w6(32'h3bd5264a),
	.w7(32'h3d00a949),
	.w8(32'h3b87d808),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb980a45),
	.w1(32'hba4097d9),
	.w2(32'h3aeaf288),
	.w3(32'hbc84003b),
	.w4(32'h3b823fb6),
	.w5(32'h3a01941e),
	.w6(32'h3b8651a9),
	.w7(32'hbb34b9ac),
	.w8(32'h3bc89e0a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ca920),
	.w1(32'h3a9e0b25),
	.w2(32'h3bc463a6),
	.w3(32'hbc1b4d28),
	.w4(32'h3b286669),
	.w5(32'h3bcd04ec),
	.w6(32'hbaac1fb8),
	.w7(32'hbc20d9d4),
	.w8(32'h3b126575),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65e780),
	.w1(32'hbc0348fc),
	.w2(32'hbbd18f69),
	.w3(32'h3b082709),
	.w4(32'h3ae933f9),
	.w5(32'h3a9d1b55),
	.w6(32'hbc2f2e02),
	.w7(32'h385e7df6),
	.w8(32'h3b1973d9),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae715ab),
	.w1(32'h39d38123),
	.w2(32'h3b301fe7),
	.w3(32'hba94be83),
	.w4(32'hbb0076cf),
	.w5(32'hbbd84130),
	.w6(32'h3b0c9d7e),
	.w7(32'h3b718332),
	.w8(32'h3c2c0f9d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ca9b6),
	.w1(32'h3b80f0fd),
	.w2(32'hbbb501e2),
	.w3(32'hbbd8d1bc),
	.w4(32'h3ad1cb2c),
	.w5(32'h3a1fefab),
	.w6(32'hbb01561d),
	.w7(32'h3b7531dd),
	.w8(32'h3c226492),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9729a0),
	.w1(32'h38429c4c),
	.w2(32'h3ca76f12),
	.w3(32'hbc717715),
	.w4(32'hbb9dfac1),
	.w5(32'h3b2a6876),
	.w6(32'hbbdec702),
	.w7(32'hbca01240),
	.w8(32'h3b4879bc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc719680),
	.w1(32'hbb5ff90e),
	.w2(32'hbcee9ab2),
	.w3(32'hbc992c8c),
	.w4(32'hbc3719c4),
	.w5(32'hbd03c546),
	.w6(32'h3ba5c362),
	.w7(32'h3d38f29d),
	.w8(32'h3c0659b6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe02907),
	.w1(32'hbb22416a),
	.w2(32'h3c3f3bee),
	.w3(32'hbbc934a2),
	.w4(32'hbc371fb8),
	.w5(32'hbb969abb),
	.w6(32'hbb80b131),
	.w7(32'hbc33dd0c),
	.w8(32'hbbc1b01f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd9bb7),
	.w1(32'h3adc9bcd),
	.w2(32'hbc394a50),
	.w3(32'hbc78e325),
	.w4(32'hbbeda9f7),
	.w5(32'hbcb8c249),
	.w6(32'h3c22a21a),
	.w7(32'h3d0f6366),
	.w8(32'h3c14cbf0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fdb0e),
	.w1(32'h3b0ad37f),
	.w2(32'hbbaa7222),
	.w3(32'hba718ffa),
	.w4(32'hbc19c533),
	.w5(32'hbb0e680f),
	.w6(32'h3bc9b686),
	.w7(32'h3c17975d),
	.w8(32'h3b46187c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f9cf2),
	.w1(32'hbbffc732),
	.w2(32'h3d03694b),
	.w3(32'hbc5b8b86),
	.w4(32'h3c49c2ac),
	.w5(32'h3d0a787d),
	.w6(32'hbc92010a),
	.w7(32'hbd605e17),
	.w8(32'hbc1ff5a5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8bfe7),
	.w1(32'hbb1f599f),
	.w2(32'h3ba47186),
	.w3(32'hb92947dc),
	.w4(32'hbba43445),
	.w5(32'hbac11ae4),
	.w6(32'hbb866339),
	.w7(32'hbc4b367e),
	.w8(32'hba84032b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebbf75),
	.w1(32'hbb76772e),
	.w2(32'hbb8630f4),
	.w3(32'hbb65a247),
	.w4(32'hbb4c95e3),
	.w5(32'hbbf4697f),
	.w6(32'h3ab29db7),
	.w7(32'h3bf1bd77),
	.w8(32'h3bf6f31e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19bc9b),
	.w1(32'hbb407211),
	.w2(32'hbc08512a),
	.w3(32'hbbcc6466),
	.w4(32'h3bc020f7),
	.w5(32'h3b4de281),
	.w6(32'hbbc7cdef),
	.w7(32'hbc01e884),
	.w8(32'hbba2537e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3608b),
	.w1(32'hbbb57725),
	.w2(32'hba649788),
	.w3(32'hbbb4a2ae),
	.w4(32'h3c28b667),
	.w5(32'hbb0e5538),
	.w6(32'hbc279da3),
	.w7(32'h3a5d059c),
	.w8(32'h3a746aed),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b143833),
	.w1(32'h39c98f4b),
	.w2(32'hbceea396),
	.w3(32'hbb543fbf),
	.w4(32'hba8c5757),
	.w5(32'hbca1ef99),
	.w6(32'h3bf8812f),
	.w7(32'h3d04d9d5),
	.w8(32'h3bd05b97),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0329fa),
	.w1(32'h3b730349),
	.w2(32'h3c74dd75),
	.w3(32'hbbafb65d),
	.w4(32'h3c42db86),
	.w5(32'h3ce5e952),
	.w6(32'hbbfecdae),
	.w7(32'hbc79a582),
	.w8(32'hbc20955d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e1766),
	.w1(32'hbb971ac4),
	.w2(32'h3c8282c7),
	.w3(32'h3c7f63e4),
	.w4(32'hbb2a9b3c),
	.w5(32'h3c0099f2),
	.w6(32'hbbeb8fe1),
	.w7(32'hbcde600a),
	.w8(32'hbbbc75f1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf87914),
	.w1(32'hbb8fc90f),
	.w2(32'hbcc83f1c),
	.w3(32'hbc0f4f7d),
	.w4(32'hbbae76fe),
	.w5(32'hbcb84206),
	.w6(32'h3b835b74),
	.w7(32'h3d027ab0),
	.w8(32'h3bc05926),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5585c),
	.w1(32'hbb8562e3),
	.w2(32'hbcc5de43),
	.w3(32'hbb80d3f6),
	.w4(32'hbc118ec3),
	.w5(32'hbcc1f34f),
	.w6(32'h3bec6af7),
	.w7(32'h3d17a4ce),
	.w8(32'h3bc7a6d3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb546563),
	.w1(32'h3aa5d3b4),
	.w2(32'hbcc3e9a4),
	.w3(32'hbb44712a),
	.w4(32'h3b869ac6),
	.w5(32'hbc005292),
	.w6(32'h3be56307),
	.w7(32'h3ce4efdf),
	.w8(32'h3c1cfe6b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf7f65),
	.w1(32'h3b8f7a1a),
	.w2(32'h3c79f1a9),
	.w3(32'h3b881fb3),
	.w4(32'hbbef777f),
	.w5(32'hbba4b1ac),
	.w6(32'hba9d732a),
	.w7(32'hbc27a86b),
	.w8(32'hbabd6cfa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a7c12),
	.w1(32'hbc3d1164),
	.w2(32'hbce96516),
	.w3(32'hbc89ba8f),
	.w4(32'hbb2176fe),
	.w5(32'h3c00ba4e),
	.w6(32'h3c233cf0),
	.w7(32'h3a911950),
	.w8(32'hbc00ba0e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d589c),
	.w1(32'hbb3a6e3d),
	.w2(32'hbce16334),
	.w3(32'h3c2fe9e9),
	.w4(32'hba833706),
	.w5(32'hbcd22e51),
	.w6(32'h3bfb028b),
	.w7(32'h3d5b8999),
	.w8(32'h3c33582f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad9204),
	.w1(32'h3aab0742),
	.w2(32'h3c2cd59a),
	.w3(32'h3b8e66e7),
	.w4(32'hbbb93151),
	.w5(32'h3ad29e68),
	.w6(32'h3950a1f1),
	.w7(32'hbc9b5642),
	.w8(32'hb988ad5b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb80ba),
	.w1(32'hbaaf5b17),
	.w2(32'hbbc678ba),
	.w3(32'hbc6b52c2),
	.w4(32'hbb9c3c17),
	.w5(32'hbc1592fd),
	.w6(32'h3a76d9cd),
	.w7(32'h3c182313),
	.w8(32'h3c385899),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee818b),
	.w1(32'hbad6e2c5),
	.w2(32'hbc8baa66),
	.w3(32'h3b469487),
	.w4(32'hba371a68),
	.w5(32'hbc726cf8),
	.w6(32'h3c885680),
	.w7(32'h3d339409),
	.w8(32'h3c0c4874),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbf24d),
	.w1(32'hbb27d5b7),
	.w2(32'hbbab7435),
	.w3(32'h3ade1a98),
	.w4(32'h3bbd03f1),
	.w5(32'hbb95c7fa),
	.w6(32'hbbfa5b89),
	.w7(32'h3b46d0d6),
	.w8(32'hbb3bc7e9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e19d8),
	.w1(32'h3b81a4f7),
	.w2(32'h3ca1638a),
	.w3(32'hbc04e14c),
	.w4(32'hbc2e8cbb),
	.w5(32'h3ae0060f),
	.w6(32'h3bb7767d),
	.w7(32'hbabd2790),
	.w8(32'h3b7643f9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cefda),
	.w1(32'hba5e4ddf),
	.w2(32'hbc1650aa),
	.w3(32'hbbea5029),
	.w4(32'hb9ee0c0f),
	.w5(32'hbbb00cce),
	.w6(32'h3b3c770e),
	.w7(32'h3b6d2252),
	.w8(32'h3ba46e64),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26d723),
	.w1(32'hb863eed9),
	.w2(32'h3c5d3d53),
	.w3(32'hbb9aa83d),
	.w4(32'hbbaf9b2f),
	.w5(32'h3b1677d7),
	.w6(32'h3ba56783),
	.w7(32'hbbcc0e7e),
	.w8(32'h3aed2129),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21c43a),
	.w1(32'hba77133d),
	.w2(32'hbb39857b),
	.w3(32'hbc521806),
	.w4(32'h3a24e6b9),
	.w5(32'hbb61ee4f),
	.w6(32'hbc0f7ba8),
	.w7(32'hbafc0b3b),
	.w8(32'hbbbb72e7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812bb2),
	.w1(32'hbb3b4214),
	.w2(32'h3ac77d43),
	.w3(32'hbc1b7b86),
	.w4(32'hbc073e5d),
	.w5(32'hbc02d611),
	.w6(32'hbb88c132),
	.w7(32'hbb59ea22),
	.w8(32'h3b914baa),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb43d51),
	.w1(32'h3ac87c9d),
	.w2(32'h3bdb151a),
	.w3(32'hbc96ee99),
	.w4(32'h3c1aa615),
	.w5(32'h3c5e0135),
	.w6(32'hbb817873),
	.w7(32'hba07d4b4),
	.w8(32'h3c80a309),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c4ff4),
	.w1(32'h3990db47),
	.w2(32'hbc81225d),
	.w3(32'hbb3b6f9a),
	.w4(32'h3b8d9e53),
	.w5(32'hbbdb6c59),
	.w6(32'h3c1d2b26),
	.w7(32'h3cd50fee),
	.w8(32'h3c086f84),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dfd25),
	.w1(32'h3b7714f2),
	.w2(32'h3c134e70),
	.w3(32'h3ba55ca3),
	.w4(32'h3b7925a4),
	.w5(32'h3b9d543a),
	.w6(32'h3b5e5d05),
	.w7(32'hbb72e7ea),
	.w8(32'h3ba34944),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab42754),
	.w1(32'hbb1cf96d),
	.w2(32'hbcc33086),
	.w3(32'hbb1e7015),
	.w4(32'hbb90eb6d),
	.w5(32'hbcb1881f),
	.w6(32'h3c4e7bd3),
	.w7(32'h3d1a4185),
	.w8(32'h3bb20d46),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14ed5f),
	.w1(32'h3aff2818),
	.w2(32'hbc88971d),
	.w3(32'hbb043b63),
	.w4(32'h3b35151a),
	.w5(32'hbc17c347),
	.w6(32'h3b224759),
	.w7(32'h3caabe1a),
	.w8(32'h3b749880),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb680742),
	.w1(32'hbc20889e),
	.w2(32'h3c7d4a47),
	.w3(32'h3a5124b6),
	.w4(32'h3831487f),
	.w5(32'h3c8452e4),
	.w6(32'hbc70ea15),
	.w7(32'hbd28f6c0),
	.w8(32'hbc5357af),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7503a),
	.w1(32'h3be4ab38),
	.w2(32'h3c40913a),
	.w3(32'hbbd00d05),
	.w4(32'h3ba60291),
	.w5(32'h3bffff98),
	.w6(32'hba885ed2),
	.w7(32'hbc0265d1),
	.w8(32'hbb0b46af),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc267c3c),
	.w1(32'hbb2fba6b),
	.w2(32'hbb42d285),
	.w3(32'hbb86f811),
	.w4(32'h3b89dc35),
	.w5(32'hbba277d1),
	.w6(32'hbc468699),
	.w7(32'h3b4bd2af),
	.w8(32'hbb53a046),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc19ce8),
	.w1(32'hbc4be868),
	.w2(32'hbb8c37a8),
	.w3(32'hbb1475f5),
	.w4(32'hbc195b17),
	.w5(32'hbb4bd8a6),
	.w6(32'h3b2513d2),
	.w7(32'hbbc80c72),
	.w8(32'h3b093d5f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc487edb),
	.w1(32'h3b9fa04e),
	.w2(32'h3b48c789),
	.w3(32'hbc111d7f),
	.w4(32'h3af1cff7),
	.w5(32'hba684a93),
	.w6(32'h39a08b55),
	.w7(32'h3c04dd9a),
	.w8(32'hbabc29a5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcded85),
	.w1(32'h3b47fb9e),
	.w2(32'h3ba0382b),
	.w3(32'hbae4fffe),
	.w4(32'h3c204f6e),
	.w5(32'h3b5c8317),
	.w6(32'h39e3c5a0),
	.w7(32'hbbfb4edb),
	.w8(32'hbc238c42),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39061677),
	.w1(32'hbb16b062),
	.w2(32'h3bc03f00),
	.w3(32'h3a5270ca),
	.w4(32'hbb2be359),
	.w5(32'h3b0a6c40),
	.w6(32'hbb13f45f),
	.w7(32'h3ba9dad6),
	.w8(32'h3c437928),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b687959),
	.w1(32'h3b8a51f7),
	.w2(32'h3cc0e98f),
	.w3(32'h3b85088d),
	.w4(32'hbc075a88),
	.w5(32'hb8e32b86),
	.w6(32'h3c0f9934),
	.w7(32'hbbc3ccbb),
	.w8(32'h3b776827),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce62e),
	.w1(32'h3bb02d2e),
	.w2(32'hb9cf51ce),
	.w3(32'hbc0e657d),
	.w4(32'h3b4a0b09),
	.w5(32'hbb0cb38f),
	.w6(32'h3b563288),
	.w7(32'h3bc181dc),
	.w8(32'hbb7436f7),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb933f67),
	.w1(32'h3c086bbb),
	.w2(32'h3b49e4b6),
	.w3(32'hba299abb),
	.w4(32'h3b576755),
	.w5(32'hbbd98ad2),
	.w6(32'h3c00b437),
	.w7(32'hbbc9d219),
	.w8(32'h3c1834d8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab83992),
	.w1(32'hb9a3d318),
	.w2(32'hbb570aa9),
	.w3(32'hbaadcb1b),
	.w4(32'hbc137c1f),
	.w5(32'h3c3a4b3e),
	.w6(32'h3c219160),
	.w7(32'h3c10fdd6),
	.w8(32'hbb683e75),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66480f),
	.w1(32'hbba40160),
	.w2(32'hbd38ba82),
	.w3(32'hbba0f857),
	.w4(32'hbb6e8850),
	.w5(32'hbd216a9c),
	.w6(32'h3c4378d4),
	.w7(32'h3da23014),
	.w8(32'h3c866e54),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef2a04),
	.w1(32'hbba1a5f6),
	.w2(32'hbcf1e201),
	.w3(32'h3bcd38d1),
	.w4(32'hbbdcfbdb),
	.w5(32'hbce701f4),
	.w6(32'h3b6400ab),
	.w7(32'h3d077eaa),
	.w8(32'h3b7699ef),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc235d27),
	.w1(32'hbb17a6cd),
	.w2(32'hbca66c74),
	.w3(32'hbc19ad0d),
	.w4(32'hbab439a0),
	.w5(32'hbc987cdc),
	.w6(32'h3beeef36),
	.w7(32'h3d21a5b4),
	.w8(32'h3c0fef08),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dbead),
	.w1(32'hbae5d320),
	.w2(32'hbc523d50),
	.w3(32'h3b3926a8),
	.w4(32'hbc121071),
	.w5(32'hbc5fa03d),
	.w6(32'h3bd43718),
	.w7(32'h3cbf4fb5),
	.w8(32'h3be9e131),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b3e33),
	.w1(32'hbc9e6010),
	.w2(32'hbc0a60de),
	.w3(32'hbb64bf96),
	.w4(32'hbc70f897),
	.w5(32'hbc346c4f),
	.w6(32'hbbd82e23),
	.w7(32'hbc0ae949),
	.w8(32'h3c1172fe),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc940dd7),
	.w1(32'hbb99165e),
	.w2(32'hbcb65910),
	.w3(32'hbc8a9dce),
	.w4(32'h3bb0735b),
	.w5(32'hbc4b40ab),
	.w6(32'h3bbaa027),
	.w7(32'h3ce1e788),
	.w8(32'h3c036727),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104e8d),
	.w1(32'hbb1a6c35),
	.w2(32'hbca9532f),
	.w3(32'h3b3b5ba7),
	.w4(32'hbade518e),
	.w5(32'hbca79ce4),
	.w6(32'h3bed5dbc),
	.w7(32'h3d2d4813),
	.w8(32'h3c20ff80),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5275c),
	.w1(32'hbba33c2c),
	.w2(32'h3cd45a6d),
	.w3(32'h3b70d06c),
	.w4(32'hb99a6051),
	.w5(32'h3c2a8297),
	.w6(32'hbc022b35),
	.w7(32'hbc91408e),
	.w8(32'h3c0bfa56),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5ddfc),
	.w1(32'h39ea8f8d),
	.w2(32'hbcb5dc62),
	.w3(32'hbbb28b5a),
	.w4(32'hbb96b3b4),
	.w5(32'hbc9717b6),
	.w6(32'h3c082067),
	.w7(32'h3d057bf3),
	.w8(32'h3b2eda7e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d9af0),
	.w1(32'h3a9de970),
	.w2(32'hbc1d630b),
	.w3(32'hbbdd07ff),
	.w4(32'hbc024004),
	.w5(32'hbc08d04f),
	.w6(32'hbbe36fe3),
	.w7(32'h3b274d47),
	.w8(32'hbc0eeab1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7540b0),
	.w1(32'hbb08f09b),
	.w2(32'hbcdd677b),
	.w3(32'hbb7d26dc),
	.w4(32'hbb078c62),
	.w5(32'hbc99e4a1),
	.w6(32'h3c262a07),
	.w7(32'h3d044122),
	.w8(32'h3b40c88b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23eda7),
	.w1(32'hbb5df436),
	.w2(32'h3c01c94a),
	.w3(32'hbc064e13),
	.w4(32'hbc12195b),
	.w5(32'hbb5c8848),
	.w6(32'hbbb796ab),
	.w7(32'hbc2e9913),
	.w8(32'h3acfdfb2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb798f39),
	.w1(32'h3c3fe84d),
	.w2(32'hbb8a99f8),
	.w3(32'hbc51c930),
	.w4(32'h3a3701fb),
	.w5(32'hbcda552b),
	.w6(32'h3c72b140),
	.w7(32'h3d11ad51),
	.w8(32'h3c2ed175),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3aa96a),
	.w1(32'hbb610fdf),
	.w2(32'hbcf33c9e),
	.w3(32'hbb019942),
	.w4(32'hbb006535),
	.w5(32'hbce5dddd),
	.w6(32'h3c2df34c),
	.w7(32'h3d73977b),
	.w8(32'h3c5b3719),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdda975),
	.w1(32'hba2c7578),
	.w2(32'hbcafd420),
	.w3(32'h3bb48a5f),
	.w4(32'hbbe98739),
	.w5(32'hbcbbcb70),
	.w6(32'h3c2112a8),
	.w7(32'h3d24fee8),
	.w8(32'h3c232944),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75219c),
	.w1(32'hba70e725),
	.w2(32'hbcbebc15),
	.w3(32'hbb0a4733),
	.w4(32'hbbe40cd8),
	.w5(32'hbcc6dde2),
	.w6(32'h3c39a9a1),
	.w7(32'h3d2a9069),
	.w8(32'h3c1a83e9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb579192),
	.w1(32'hbb2a108d),
	.w2(32'hbca5cb25),
	.w3(32'hbb870c86),
	.w4(32'hbb837182),
	.w5(32'hbc85a20f),
	.w6(32'h3bda3b77),
	.w7(32'h3c6f4ec1),
	.w8(32'h39dfdee8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcee227),
	.w1(32'hbbad1308),
	.w2(32'h3b045dc5),
	.w3(32'hbb611767),
	.w4(32'hbbd57826),
	.w5(32'hbc015652),
	.w6(32'hbbe6726b),
	.w7(32'hbce857f9),
	.w8(32'hbb890462),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdf297),
	.w1(32'h3b3a8c18),
	.w2(32'hbc884f3c),
	.w3(32'hbae68fb9),
	.w4(32'hbb1309e7),
	.w5(32'hbc9ff697),
	.w6(32'h3bd3ff2e),
	.w7(32'h3caf9593),
	.w8(32'h3c36b71a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf59472),
	.w1(32'h3bc7d7d4),
	.w2(32'hba84837c),
	.w3(32'hbc694123),
	.w4(32'hbc17a63d),
	.w5(32'hbc8bb6c5),
	.w6(32'h3c3438c2),
	.w7(32'h3cbf1959),
	.w8(32'h38eaec60),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fb092),
	.w1(32'h3abc6431),
	.w2(32'hbcb49f2e),
	.w3(32'hbc33b4d9),
	.w4(32'hbc198233),
	.w5(32'hbce44355),
	.w6(32'h3c5173d5),
	.w7(32'h3d4ef82f),
	.w8(32'h3c243027),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79c456),
	.w1(32'h3b8ee7fe),
	.w2(32'hbc306ae6),
	.w3(32'hbb808a26),
	.w4(32'hba323570),
	.w5(32'hba8ffe2d),
	.w6(32'h3b69152b),
	.w7(32'h3a06025e),
	.w8(32'hbbd0eb9e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a2ea4),
	.w1(32'h3c13fb31),
	.w2(32'hbb867e84),
	.w3(32'hbb0429cd),
	.w4(32'hbb8bd68e),
	.w5(32'hbd10162e),
	.w6(32'h3c3e3af4),
	.w7(32'h3d06ae3a),
	.w8(32'h3b97df35),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1a7a3),
	.w1(32'hbb4fbc28),
	.w2(32'hbcf2bc2e),
	.w3(32'hbcc57b59),
	.w4(32'h3c03b8c6),
	.w5(32'hbc58c386),
	.w6(32'h3c313de6),
	.w7(32'h3d084f08),
	.w8(32'h3c3ac7c3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5911cc),
	.w1(32'h3766b3df),
	.w2(32'hb8b61f33),
	.w3(32'h3bef7995),
	.w4(32'h3969c837),
	.w5(32'h390b952a),
	.w6(32'h39b862cc),
	.w7(32'h39073de9),
	.w8(32'h39223db8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba731616),
	.w1(32'h3b0357bd),
	.w2(32'h3b2871b8),
	.w3(32'hba4d2fac),
	.w4(32'hb5c891a4),
	.w5(32'h3afc6c9a),
	.w6(32'h3a9caa6b),
	.w7(32'h3b8993d3),
	.w8(32'h3b760c73),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule