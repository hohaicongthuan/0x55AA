module layer_10_featuremap_466(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba70d6e),
	.w1(32'hbbf80cfa),
	.w2(32'hba909f4c),
	.w3(32'hbb96bd1d),
	.w4(32'hbb3fa219),
	.w5(32'h3b295221),
	.w6(32'hbbf873a2),
	.w7(32'hbb2dde01),
	.w8(32'h3b5354b5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd63c0),
	.w1(32'h3c4a70e1),
	.w2(32'h3c26d7d4),
	.w3(32'h39863ab9),
	.w4(32'h3c308ba5),
	.w5(32'h3cc4b749),
	.w6(32'h3b5f5f68),
	.w7(32'h3ba9cd2d),
	.w8(32'h3b76f0ce),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af13425),
	.w1(32'h3c1c880f),
	.w2(32'h3c1f67e7),
	.w3(32'hbb528ea3),
	.w4(32'h3bfb85f9),
	.w5(32'h3b867d01),
	.w6(32'h39ab6713),
	.w7(32'hba935cd2),
	.w8(32'h3c20cba2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085788),
	.w1(32'h3c1d9e12),
	.w2(32'h3c0a31bb),
	.w3(32'hbc06be78),
	.w4(32'h3bdf5f59),
	.w5(32'h3c0ac906),
	.w6(32'h3ad189c2),
	.w7(32'h3c853509),
	.w8(32'h3bc5b6b8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c980dd9),
	.w1(32'hbbeb6df5),
	.w2(32'hbaf920a3),
	.w3(32'h3c8af69b),
	.w4(32'hbbc86eb1),
	.w5(32'hbb102f91),
	.w6(32'h3c537e74),
	.w7(32'hbb754c97),
	.w8(32'hbb7577bf),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8928e),
	.w1(32'hbc01ae9e),
	.w2(32'hbbb98652),
	.w3(32'h3b1b90aa),
	.w4(32'hbb11674a),
	.w5(32'hbc814089),
	.w6(32'hbaa64902),
	.w7(32'hbc0b8408),
	.w8(32'hbc338e95),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadad356),
	.w1(32'hbc5f6671),
	.w2(32'hbafd7095),
	.w3(32'hbaa5f39a),
	.w4(32'hbc4eaa89),
	.w5(32'h3bc2b796),
	.w6(32'hb92085dd),
	.w7(32'hbb854b11),
	.w8(32'hbb91d666),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc211f26),
	.w1(32'hbbe0881f),
	.w2(32'hbb11d0f4),
	.w3(32'hbbe6c0fe),
	.w4(32'hbb93feec),
	.w5(32'hbc4d2dec),
	.w6(32'hbc2454a5),
	.w7(32'h3c126089),
	.w8(32'h39a50931),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c114d9c),
	.w1(32'hbc0b2fb6),
	.w2(32'h3af606ba),
	.w3(32'h3b8d8fec),
	.w4(32'hbc17c809),
	.w5(32'h3bb909bb),
	.w6(32'h3c3605e6),
	.w7(32'hbc08cdc7),
	.w8(32'h3b74bd89),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0df4a7),
	.w1(32'hba9c0fa7),
	.w2(32'hbb411fbb),
	.w3(32'hbabc585e),
	.w4(32'h3b116ee3),
	.w5(32'h3b737a31),
	.w6(32'h3b36a2c8),
	.w7(32'h3a83249a),
	.w8(32'h3b79e93c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ad79),
	.w1(32'hbba63260),
	.w2(32'hbba8832b),
	.w3(32'h3c487ca8),
	.w4(32'hbc1dcb24),
	.w5(32'hbb581796),
	.w6(32'h3b480c30),
	.w7(32'hbc840fb8),
	.w8(32'hbc47695f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04324b),
	.w1(32'hbb261aef),
	.w2(32'hbb8ea85f),
	.w3(32'hbb957004),
	.w4(32'hba0f2c74),
	.w5(32'hbb7b7faa),
	.w6(32'hbc043d11),
	.w7(32'h3b92b777),
	.w8(32'hb9bf3dd1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82996f),
	.w1(32'hbc511011),
	.w2(32'h3bccb725),
	.w3(32'h3b8eca18),
	.w4(32'hbc619edf),
	.w5(32'h3c651928),
	.w6(32'h3b7e4c54),
	.w7(32'hbc58ef27),
	.w8(32'h3aabe067),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31b94f),
	.w1(32'hbb54c1d1),
	.w2(32'hbb274426),
	.w3(32'hbc35cd62),
	.w4(32'hbc023794),
	.w5(32'hbad4c31e),
	.w6(32'hbc5fa378),
	.w7(32'hbbc4118c),
	.w8(32'h3aa91b49),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a3a5c),
	.w1(32'h3c2d58e1),
	.w2(32'hbc0a1516),
	.w3(32'hbb86ab7c),
	.w4(32'h3c6a02da),
	.w5(32'hbbeefc04),
	.w6(32'hbb182dff),
	.w7(32'h3c88c854),
	.w8(32'hbbb27c96),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e4877),
	.w1(32'h3ac19c3e),
	.w2(32'h389feb20),
	.w3(32'h3c19cd94),
	.w4(32'h39d0ccc7),
	.w5(32'hbb804cff),
	.w6(32'h3b3c978e),
	.w7(32'h398d2840),
	.w8(32'hba9fde37),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e5f47a),
	.w1(32'hbb8ea945),
	.w2(32'hbc12f3b2),
	.w3(32'h3c26af27),
	.w4(32'hbb82366b),
	.w5(32'hbc00dbf2),
	.w6(32'hb70698ae),
	.w7(32'h3aca3035),
	.w8(32'hbb8ffa64),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152309),
	.w1(32'hbbec09c8),
	.w2(32'h3b887425),
	.w3(32'hbb3c4451),
	.w4(32'hbc217d5d),
	.w5(32'h3bd862dc),
	.w6(32'hbb981528),
	.w7(32'hbb6b1906),
	.w8(32'h3c1dbda8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3f13c),
	.w1(32'h3b0f06bb),
	.w2(32'hbbfa2ff3),
	.w3(32'h3c07394a),
	.w4(32'h3bfc2e81),
	.w5(32'hbc237c60),
	.w6(32'h3c2642fc),
	.w7(32'h3b829db8),
	.w8(32'hbc0411d7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16dbf3),
	.w1(32'h3b363a66),
	.w2(32'hbb8be478),
	.w3(32'h3b7e01ca),
	.w4(32'h3b6b0f42),
	.w5(32'hbb0e4fef),
	.w6(32'h3bc67c4f),
	.w7(32'hbb4c0f5e),
	.w8(32'hb5b7b12f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4cef4),
	.w1(32'h3b64cf1b),
	.w2(32'hbab2de2b),
	.w3(32'hbc3dc218),
	.w4(32'h399293dc),
	.w5(32'hbc092c20),
	.w6(32'hbb4554aa),
	.w7(32'hbbafc7bb),
	.w8(32'hbc0489d6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b271b9),
	.w1(32'h3b22608f),
	.w2(32'hba8fcc6b),
	.w3(32'h39d39a39),
	.w4(32'h3bf03eca),
	.w5(32'h394d5db6),
	.w6(32'hbbdb1593),
	.w7(32'h3b81e5a7),
	.w8(32'hbb376ff0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81bdc9),
	.w1(32'hba22fc53),
	.w2(32'hbc1c3de2),
	.w3(32'hba38b35d),
	.w4(32'h3bbe9049),
	.w5(32'h3bb4658b),
	.w6(32'hbb682071),
	.w7(32'h3abd8ead),
	.w8(32'hbc330f04),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ddce0),
	.w1(32'hbabce886),
	.w2(32'hbac8d65b),
	.w3(32'hbaca4860),
	.w4(32'hbb8562f6),
	.w5(32'hbb83c4d4),
	.w6(32'hbbc1f8ec),
	.w7(32'h396790de),
	.w8(32'hbb93d955),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3863422c),
	.w1(32'hbb280459),
	.w2(32'h3c143c11),
	.w3(32'hb8ecc6b5),
	.w4(32'hbbcbc709),
	.w5(32'h3c9d2153),
	.w6(32'hbbb48bc3),
	.w7(32'hbc1b5f32),
	.w8(32'h3c2781e1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05c2ea),
	.w1(32'h3a41d1e6),
	.w2(32'h3b5f2263),
	.w3(32'h3a96915a),
	.w4(32'h3b20b76f),
	.w5(32'hb9eec234),
	.w6(32'h3b8d7df7),
	.w7(32'h3b978411),
	.w8(32'h3bdc2960),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ab01),
	.w1(32'hbbc43286),
	.w2(32'hbb4bba87),
	.w3(32'h3c4c4bd7),
	.w4(32'hbc2b36c8),
	.w5(32'h3b4a4159),
	.w6(32'h3bcd077f),
	.w7(32'hbbd7c8fd),
	.w8(32'hbb4d9a6a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0d937),
	.w1(32'hbb57c2cb),
	.w2(32'h3b1040e8),
	.w3(32'h3a0a9c1c),
	.w4(32'h3adb7c72),
	.w5(32'h3bdbe7f6),
	.w6(32'h3b3bbe70),
	.w7(32'h3b5eac30),
	.w8(32'h3bac45c9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c37d7),
	.w1(32'hbb3c6d89),
	.w2(32'h3a05a438),
	.w3(32'h39aaf927),
	.w4(32'h3c0e6c93),
	.w5(32'h3b5091c0),
	.w6(32'h3abc0931),
	.w7(32'hba2102b5),
	.w8(32'hbbefbbb8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba80d72),
	.w1(32'hbc113a8c),
	.w2(32'hbc0141ae),
	.w3(32'hbb7ed8b3),
	.w4(32'hbc4ebae5),
	.w5(32'hbc3df587),
	.w6(32'hbc05336a),
	.w7(32'hbbee5585),
	.w8(32'hbc0ef3af),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a171a4),
	.w1(32'hb9d83d7f),
	.w2(32'hbb441d0d),
	.w3(32'h3b0c2892),
	.w4(32'hbb2a3eda),
	.w5(32'h3b021830),
	.w6(32'hbb81c4d1),
	.w7(32'hbaca52ed),
	.w8(32'hba689857),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e2948),
	.w1(32'h3bd502fa),
	.w2(32'h3b292b82),
	.w3(32'hbb8ad07e),
	.w4(32'h3a79c9ff),
	.w5(32'h3c287f23),
	.w6(32'hbbcd40a6),
	.w7(32'h3aaa9fbd),
	.w8(32'h3ba0a995),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb254ad),
	.w1(32'h3bbff9e4),
	.w2(32'h3b96ca93),
	.w3(32'hbbab0a70),
	.w4(32'h3bcb63f6),
	.w5(32'h3c60ed97),
	.w6(32'hba9320dd),
	.w7(32'h3c019730),
	.w8(32'h3c32ca4f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f9650),
	.w1(32'hbb5661a6),
	.w2(32'hbb4b96b3),
	.w3(32'hbbd388b5),
	.w4(32'h3b03ce6a),
	.w5(32'h3b3a4f0c),
	.w6(32'hbb02d572),
	.w7(32'h3ba1dcd4),
	.w8(32'hbbcfef89),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1ea23),
	.w1(32'h3af341aa),
	.w2(32'hbabfaba5),
	.w3(32'hbc87ee5b),
	.w4(32'h3b20ecad),
	.w5(32'hbb27ebdb),
	.w6(32'hbc71ae31),
	.w7(32'h3a5dfddf),
	.w8(32'hbb930476),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5d885),
	.w1(32'h3b4af3ce),
	.w2(32'h3c03917d),
	.w3(32'hbb69b855),
	.w4(32'h3b1ea26b),
	.w5(32'h3bee6669),
	.w6(32'h39ea10fa),
	.w7(32'h3be230b1),
	.w8(32'h3b51819d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd268ce),
	.w1(32'hbc164dec),
	.w2(32'hbc2f875d),
	.w3(32'h3ba43a2c),
	.w4(32'hbc2a4579),
	.w5(32'h395cf495),
	.w6(32'h3be27211),
	.w7(32'hbc88e7ac),
	.w8(32'hbc29e8ab),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0f68),
	.w1(32'hbbebcca9),
	.w2(32'h3b79d1c3),
	.w3(32'hbb23aeca),
	.w4(32'hbba25558),
	.w5(32'h3c798a54),
	.w6(32'hbbc3bff7),
	.w7(32'h38cb5294),
	.w8(32'h3bbea4cb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb58b3e),
	.w1(32'hbb802fa2),
	.w2(32'h3c12cd3e),
	.w3(32'hbb1ca999),
	.w4(32'hbb92f1d7),
	.w5(32'h3cd8ee50),
	.w6(32'h3ae4a640),
	.w7(32'hbb8d301c),
	.w8(32'h3c3f5d3f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc168cfe),
	.w1(32'h3b366605),
	.w2(32'h3c11fb91),
	.w3(32'hbc877a1d),
	.w4(32'h3abbe9e2),
	.w5(32'h3c166965),
	.w6(32'hbad3edbc),
	.w7(32'h3c269ce6),
	.w8(32'h3c66faec),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3df21),
	.w1(32'hbb902866),
	.w2(32'hba868929),
	.w3(32'h3cb09a78),
	.w4(32'hbaf09b6a),
	.w5(32'h3b0df0aa),
	.w6(32'h3ca9c048),
	.w7(32'h3b91b99b),
	.w8(32'h3b5efd35),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecd507),
	.w1(32'h3bd1f2b5),
	.w2(32'hbb5e56b0),
	.w3(32'h3c106cda),
	.w4(32'h3bb13e26),
	.w5(32'hbc3e4f7d),
	.w6(32'h3b41c1af),
	.w7(32'h3ae937a7),
	.w8(32'hbb86fce6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae78417),
	.w1(32'h3c270706),
	.w2(32'h3c6a0d95),
	.w3(32'h3c8d81d6),
	.w4(32'h3c2200e6),
	.w5(32'h3cbb33f8),
	.w6(32'h3bc1ff18),
	.w7(32'h3c838a88),
	.w8(32'h3c2688a6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c617121),
	.w1(32'hbb341eaa),
	.w2(32'h3b12e585),
	.w3(32'hbbb9dfc7),
	.w4(32'hba9602e3),
	.w5(32'h3c031236),
	.w6(32'hb7d7b52a),
	.w7(32'h3b8ef54c),
	.w8(32'h3beb2035),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba314fed),
	.w1(32'h3be2d38f),
	.w2(32'hb9d7e7ff),
	.w3(32'hbb508f74),
	.w4(32'h3c1466ed),
	.w5(32'hbb498669),
	.w6(32'h3bc6187b),
	.w7(32'h3bdc728d),
	.w8(32'hbb2d5e35),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa4226),
	.w1(32'hb9bf0426),
	.w2(32'h3b06329d),
	.w3(32'hbae4f0fd),
	.w4(32'hbb286a83),
	.w5(32'hbaaf723c),
	.w6(32'h394d0db7),
	.w7(32'hb9b1c023),
	.w8(32'h3acca759),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cbfe8),
	.w1(32'hbb2a9266),
	.w2(32'hbb9cd444),
	.w3(32'h3c081d8a),
	.w4(32'hbc1295e9),
	.w5(32'hbc2dc614),
	.w6(32'hbb7bd678),
	.w7(32'hbc312730),
	.w8(32'hbc290fb1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5433a),
	.w1(32'h3b111a4d),
	.w2(32'h3c1f6274),
	.w3(32'hbc621d92),
	.w4(32'h3b5e83c9),
	.w5(32'h3c9482b7),
	.w6(32'hbc93076b),
	.w7(32'h3be56289),
	.w8(32'h3c3b7902),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a947557),
	.w1(32'hbba4b32e),
	.w2(32'hbb9f1913),
	.w3(32'h3bc65ce9),
	.w4(32'hbb9c374e),
	.w5(32'hbc15195a),
	.w6(32'h3b9b8473),
	.w7(32'hba0691f7),
	.w8(32'h39f2d677),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee047b),
	.w1(32'h3b6b7bb0),
	.w2(32'h3bf8e9da),
	.w3(32'hbab5a346),
	.w4(32'hbb134333),
	.w5(32'h3b806351),
	.w6(32'hbb412fe1),
	.w7(32'h3b852162),
	.w8(32'h3bddcd4f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b576520),
	.w1(32'h3c050a7a),
	.w2(32'hbba903ec),
	.w3(32'h3bc3cec6),
	.w4(32'h3c1a3c6c),
	.w5(32'hbc18a243),
	.w6(32'hb890e15d),
	.w7(32'h3a880941),
	.w8(32'hbb2604cd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49be05),
	.w1(32'hbb03428b),
	.w2(32'h3a827574),
	.w3(32'hbbaa8a43),
	.w4(32'hbba6c95c),
	.w5(32'h3c9b3b6e),
	.w6(32'hba359d72),
	.w7(32'hbb72b93a),
	.w8(32'h3baf0f01),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b5b33),
	.w1(32'h39f209c9),
	.w2(32'hba54365c),
	.w3(32'hbb7c6ac6),
	.w4(32'h3ac3d0f6),
	.w5(32'hbb8d1206),
	.w6(32'h39ba3d7f),
	.w7(32'h3a2450b4),
	.w8(32'hbc0db1f1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea6385),
	.w1(32'h3af79259),
	.w2(32'h3bf36ded),
	.w3(32'hbba91745),
	.w4(32'h3bce80ab),
	.w5(32'h3bf76988),
	.w6(32'hbba89544),
	.w7(32'h3ba9afa5),
	.w8(32'h3b17de8f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cab0a),
	.w1(32'hbb46172d),
	.w2(32'h3c3b7f49),
	.w3(32'hbba2b5e8),
	.w4(32'hbbe7a53e),
	.w5(32'h3c4b95fe),
	.w6(32'h3b3f559f),
	.w7(32'hbbab5b6f),
	.w8(32'h3c0c128c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba15adf),
	.w1(32'h3bfdaee4),
	.w2(32'h3c43cab9),
	.w3(32'h3bc43061),
	.w4(32'h3c6a6a2e),
	.w5(32'h3c4db278),
	.w6(32'h3a1ff984),
	.w7(32'h3c13e588),
	.w8(32'h3c3b1c7d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b349f),
	.w1(32'hbb5a586b),
	.w2(32'hbbcac606),
	.w3(32'hbb76efa6),
	.w4(32'hbb9ff651),
	.w5(32'hbbd2ff8e),
	.w6(32'h3c02e89f),
	.w7(32'hbb4ff800),
	.w8(32'hbbd48fca),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fea7d),
	.w1(32'hbb6093c5),
	.w2(32'hbb38ba63),
	.w3(32'hbb12193a),
	.w4(32'hbbf27fe8),
	.w5(32'hbba8a9c7),
	.w6(32'hbb5862bf),
	.w7(32'hbb76713e),
	.w8(32'hba8fbc0b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe8f6f),
	.w1(32'h3b3fc9ec),
	.w2(32'h3a3dbfc8),
	.w3(32'hbb84dfe4),
	.w4(32'hbb3ac90b),
	.w5(32'h3c34a1b1),
	.w6(32'hbbe923c2),
	.w7(32'h3b971e01),
	.w8(32'h3b3c89a3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6c28a),
	.w1(32'hbb8b2101),
	.w2(32'h3b3e5c76),
	.w3(32'h3b18a2cc),
	.w4(32'hbc1cd422),
	.w5(32'h3b02360c),
	.w6(32'h3b0ee4e2),
	.w7(32'hbc0d79e4),
	.w8(32'hbc12acaf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec82c9),
	.w1(32'h3c460e11),
	.w2(32'h3bcb6bc4),
	.w3(32'h3bd7cbcf),
	.w4(32'h3b14db6f),
	.w5(32'hbb664cdc),
	.w6(32'h3b2453d3),
	.w7(32'h3b1a9527),
	.w8(32'h3b081762),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2f55a),
	.w1(32'h3bae32ee),
	.w2(32'hbbf6a73f),
	.w3(32'h3c8b45a0),
	.w4(32'h3c1407a5),
	.w5(32'h3ada2c7b),
	.w6(32'h3beef3fe),
	.w7(32'h3c1e8667),
	.w8(32'hbb899d3c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1389fe),
	.w1(32'h3bd53796),
	.w2(32'h3bf986f4),
	.w3(32'hbbbf7e20),
	.w4(32'hb86b717b),
	.w5(32'h3bf6fcc8),
	.w6(32'hbb361c82),
	.w7(32'h3c06227d),
	.w8(32'h3c09109e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb01257),
	.w1(32'hbb34e8d0),
	.w2(32'hbbc993e2),
	.w3(32'h3be9d42f),
	.w4(32'hbb0683a3),
	.w5(32'hbc0eeaea),
	.w6(32'h3c66b84c),
	.w7(32'hbb90b3b7),
	.w8(32'h38d4be2d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e7393),
	.w1(32'h3b3a65de),
	.w2(32'h3b2abb80),
	.w3(32'hbb614d37),
	.w4(32'h385665d1),
	.w5(32'hbb92beff),
	.w6(32'h3ba2c29f),
	.w7(32'h3a1bbf74),
	.w8(32'h3ba3df62),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad54d3),
	.w1(32'hbc046060),
	.w2(32'hbb3dc360),
	.w3(32'h3c094e62),
	.w4(32'hbb0000a8),
	.w5(32'h39ae906b),
	.w6(32'h3c29526a),
	.w7(32'hbb138de0),
	.w8(32'hb94aa529),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1688c1),
	.w1(32'hbbe5106e),
	.w2(32'hbc391022),
	.w3(32'hbb503aeb),
	.w4(32'h3b7840dd),
	.w5(32'hbc2d9ee5),
	.w6(32'h3aca9932),
	.w7(32'hbc567ef7),
	.w8(32'hbba68375),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164c52),
	.w1(32'hbaae063d),
	.w2(32'hbae5ee9a),
	.w3(32'hba8069a3),
	.w4(32'h3b5e7cd1),
	.w5(32'hbc4cef62),
	.w6(32'hbb6357f5),
	.w7(32'hbab6497f),
	.w8(32'h3bf7ec9e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc60514),
	.w1(32'h3c6ce682),
	.w2(32'h3c2e93c9),
	.w3(32'h390b2c36),
	.w4(32'h3c751335),
	.w5(32'h3c79cea2),
	.w6(32'h3b3bb4ca),
	.w7(32'h3c2aca7c),
	.w8(32'h3c2b36ad),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b885242),
	.w1(32'hba935007),
	.w2(32'hbb7703bb),
	.w3(32'h3baeddaa),
	.w4(32'hbb7afd33),
	.w5(32'hbacf87b3),
	.w6(32'h3c060071),
	.w7(32'hbb58c48c),
	.w8(32'hbb3f74da),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1e0de),
	.w1(32'h3b50bb64),
	.w2(32'h3a74ccb9),
	.w3(32'h3bc2ee6d),
	.w4(32'h3b04dc79),
	.w5(32'hbbac840a),
	.w6(32'h3b38a978),
	.w7(32'h3bab4683),
	.w8(32'hbb870e20),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8b5b2),
	.w1(32'h3bd0a691),
	.w2(32'hbab32320),
	.w3(32'hba940563),
	.w4(32'h3a5efdbe),
	.w5(32'hbba4d7ee),
	.w6(32'h3b5caa0e),
	.w7(32'hbb96e82c),
	.w8(32'h3ab9f4ec),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e0c73),
	.w1(32'hbb311616),
	.w2(32'hbb0d2752),
	.w3(32'hbafdc5d8),
	.w4(32'hba71717d),
	.w5(32'h398faf27),
	.w6(32'hbb8726a5),
	.w7(32'h3b631fcc),
	.w8(32'h3a870f6e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf90f70),
	.w1(32'h3b55f6ca),
	.w2(32'h3be530f3),
	.w3(32'hbb5fdf6e),
	.w4(32'h3bb2df86),
	.w5(32'h3ba4a927),
	.w6(32'hbb2b4afa),
	.w7(32'hbb2d3ebe),
	.w8(32'hbbf629ec),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a477f),
	.w1(32'hbbac728d),
	.w2(32'h3ba670c9),
	.w3(32'hbbfc7908),
	.w4(32'hbc36e353),
	.w5(32'hbaeb1405),
	.w6(32'hbc5afdd0),
	.w7(32'h39c2fef4),
	.w8(32'h3c1e0ca5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8197d),
	.w1(32'hbbd3e8e2),
	.w2(32'hba18c9e7),
	.w3(32'hbbebeb79),
	.w4(32'hbb1ca9f1),
	.w5(32'h3bbbc673),
	.w6(32'h3aaae605),
	.w7(32'h3a22805e),
	.w8(32'h39e7b103),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb458e1),
	.w1(32'h3b86d3ac),
	.w2(32'h3a951e13),
	.w3(32'hbb7e6fe2),
	.w4(32'h3a071885),
	.w5(32'h39566bb6),
	.w6(32'hbb0c786d),
	.w7(32'hbaad3e0d),
	.w8(32'hbb440823),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3396d),
	.w1(32'h3b85a90c),
	.w2(32'h3bbfa292),
	.w3(32'h3bf2a424),
	.w4(32'h3a615774),
	.w5(32'h3b89d4ee),
	.w6(32'hbad1314e),
	.w7(32'hbc142904),
	.w8(32'hbba1b454),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f7185),
	.w1(32'hbb71bce9),
	.w2(32'hbb1379ba),
	.w3(32'h3b98ff92),
	.w4(32'hbbc60b3c),
	.w5(32'hbb16fe54),
	.w6(32'h3ba48f5b),
	.w7(32'hbb88f795),
	.w8(32'hba812d1a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68e742),
	.w1(32'h3b0b2f09),
	.w2(32'hbb1406a3),
	.w3(32'hbb983639),
	.w4(32'h3ba6a734),
	.w5(32'hbace6178),
	.w6(32'hbb44828c),
	.w7(32'h3bf62621),
	.w8(32'hb710e35b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c399718),
	.w1(32'h3bd85774),
	.w2(32'h3b3098f3),
	.w3(32'h3c05a5ff),
	.w4(32'h3b9db669),
	.w5(32'h3952957f),
	.w6(32'h3a69152c),
	.w7(32'h3afad6e3),
	.w8(32'hbb66d400),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba919f7c),
	.w1(32'h3a3c82a6),
	.w2(32'h3bc5b31c),
	.w3(32'hbba627f3),
	.w4(32'h3a0b3ef6),
	.w5(32'h3b8e0261),
	.w6(32'hb9e5c45b),
	.w7(32'hbb7b67c9),
	.w8(32'h3a4dec56),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55ccfa),
	.w1(32'hbb4c4dfd),
	.w2(32'hbb47bdf0),
	.w3(32'h3b85ed89),
	.w4(32'hbacaee95),
	.w5(32'h3b8a50a0),
	.w6(32'h3b41d80f),
	.w7(32'h3bdd4b91),
	.w8(32'h3c5cc908),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b996d10),
	.w1(32'h3b940368),
	.w2(32'h3adfd631),
	.w3(32'h3be2fcd8),
	.w4(32'h3aa21cd2),
	.w5(32'hbabbfdb6),
	.w6(32'h3bf2230c),
	.w7(32'hbb8c7a76),
	.w8(32'hb9ddce43),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e037e),
	.w1(32'h3a9ba411),
	.w2(32'hba73d7c5),
	.w3(32'h3c00099a),
	.w4(32'h3c1ca9cc),
	.w5(32'h3a0ce2a2),
	.w6(32'h3c3596e3),
	.w7(32'h3bb0f84a),
	.w8(32'h3b58677e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998ac5f),
	.w1(32'h3c24a270),
	.w2(32'h3a005098),
	.w3(32'hba8e2043),
	.w4(32'h3b1981ac),
	.w5(32'h3b39f2c3),
	.w6(32'hb9cfae4c),
	.w7(32'hbb277124),
	.w8(32'hba35d379),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae6e28),
	.w1(32'hbad8ac74),
	.w2(32'hbb80db7f),
	.w3(32'hbb6c3d2a),
	.w4(32'h3a623a75),
	.w5(32'hbb2117f7),
	.w6(32'hbb8226b0),
	.w7(32'h3bd8a1f9),
	.w8(32'hba5554d2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b067),
	.w1(32'hbc129063),
	.w2(32'hbc205644),
	.w3(32'h3b1f2d4f),
	.w4(32'hba86dc97),
	.w5(32'hba03b188),
	.w6(32'hbae6616b),
	.w7(32'h382f3cda),
	.w8(32'hbaa59848),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3937c1),
	.w1(32'hba5ae9fb),
	.w2(32'h39684cae),
	.w3(32'hbbecdae1),
	.w4(32'hbb97656b),
	.w5(32'h3ad052a0),
	.w6(32'hbbaeaee7),
	.w7(32'hbb4985ed),
	.w8(32'h3a2db5db),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718817),
	.w1(32'hbb43139d),
	.w2(32'h3b823777),
	.w3(32'h3b1ac43b),
	.w4(32'h3a8f7577),
	.w5(32'h3b493538),
	.w6(32'hbab735fe),
	.w7(32'hba558b54),
	.w8(32'h3b27ad9e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3b278),
	.w1(32'hbaf0a14b),
	.w2(32'h3b986bec),
	.w3(32'h3bb2558d),
	.w4(32'h3b8794cc),
	.w5(32'h3bb3759a),
	.w6(32'hba9c9e7c),
	.w7(32'h399ca55d),
	.w8(32'h3b0077d7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8ec4f),
	.w1(32'h3b04f33b),
	.w2(32'h3bd9ee8f),
	.w3(32'hba9788e7),
	.w4(32'h3af5d146),
	.w5(32'h3bb6b41f),
	.w6(32'hbaaa7a8f),
	.w7(32'hbb179ea5),
	.w8(32'hbb00b247),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba230098),
	.w1(32'hbb1bcf36),
	.w2(32'hbb6504fc),
	.w3(32'h39ab7ecc),
	.w4(32'h3a3c2f37),
	.w5(32'h3ba8f615),
	.w6(32'h3a395fdc),
	.w7(32'hbaaa7ea3),
	.w8(32'h3b02b28c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7b58f),
	.w1(32'h3b08a40f),
	.w2(32'h395e67df),
	.w3(32'h3b7f8137),
	.w4(32'hb8d35366),
	.w5(32'hb940c628),
	.w6(32'hbab85934),
	.w7(32'hbc12e6a6),
	.w8(32'hbc488cbe),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba013ee),
	.w1(32'h3ba03f32),
	.w2(32'h3c40d6ff),
	.w3(32'hbbd487b9),
	.w4(32'hbbc71f01),
	.w5(32'hbb781cb4),
	.w6(32'hbbe900e9),
	.w7(32'hbaf14211),
	.w8(32'hbb1892b0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86398b),
	.w1(32'h3bdf5e56),
	.w2(32'h3beb43a5),
	.w3(32'hbb9427ba),
	.w4(32'h3c4cd21a),
	.w5(32'h3c172572),
	.w6(32'h3b05a94d),
	.w7(32'h3b9ed579),
	.w8(32'h3a296f43),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4894f5),
	.w1(32'hb9732f26),
	.w2(32'h3ad8c0b4),
	.w3(32'hbbf6b976),
	.w4(32'h3bd1e40b),
	.w5(32'h3bacde0a),
	.w6(32'hbbec2bdc),
	.w7(32'h3a032a90),
	.w8(32'h3b3c5a29),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0972f),
	.w1(32'h39228ce4),
	.w2(32'hbb1c9d55),
	.w3(32'hbb4bdda5),
	.w4(32'hb92e5685),
	.w5(32'hba8b868d),
	.w6(32'hbb44b459),
	.w7(32'h3ba76a5c),
	.w8(32'h3b938434),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae50e70),
	.w1(32'hbbe29af5),
	.w2(32'hbab7e5ef),
	.w3(32'h3b806f53),
	.w4(32'hbb724c50),
	.w5(32'hbb8a9d68),
	.w6(32'h38a728e6),
	.w7(32'h3ab6a1b9),
	.w8(32'h3b5f4d4b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69afeb),
	.w1(32'hbb822760),
	.w2(32'hbb63433e),
	.w3(32'h3b1b5292),
	.w4(32'hbaf1e626),
	.w5(32'h3a705d8e),
	.w6(32'hbab5e57e),
	.w7(32'h3ba43780),
	.w8(32'h3c0c478c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c8f7),
	.w1(32'h3b89a7d1),
	.w2(32'h3c4ca779),
	.w3(32'hbabde416),
	.w4(32'h395b9532),
	.w5(32'h3bd5e885),
	.w6(32'hbaeeda48),
	.w7(32'hbb935ae8),
	.w8(32'hbbb6d312),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dca6f),
	.w1(32'hbbbec531),
	.w2(32'hbb7f022d),
	.w3(32'hbb055a91),
	.w4(32'hbb91d21a),
	.w5(32'h37a1674a),
	.w6(32'hbc166787),
	.w7(32'hbc06ee00),
	.w8(32'hbb9a9ee3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d4cc),
	.w1(32'hbc3e293a),
	.w2(32'hbc661036),
	.w3(32'h3a31c222),
	.w4(32'hbc10279d),
	.w5(32'hbc026832),
	.w6(32'hbaf51fb6),
	.w7(32'hbb61e86c),
	.w8(32'hbb0d9f3c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58eacb),
	.w1(32'hbb1a1f96),
	.w2(32'hbbf49cef),
	.w3(32'hbc0c9bc6),
	.w4(32'h3c01eadf),
	.w5(32'hbbe0ec09),
	.w6(32'hba7737c1),
	.w7(32'hbb114bd4),
	.w8(32'hbc1abb06),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc430840),
	.w1(32'hbb9c9f03),
	.w2(32'hbb0267eb),
	.w3(32'hbc5022a8),
	.w4(32'hbafc1e04),
	.w5(32'h3bca48ef),
	.w6(32'hbc54cc11),
	.w7(32'h3b52ae73),
	.w8(32'h3bf963a2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf6ca4),
	.w1(32'hbb73fc6d),
	.w2(32'h3b33b61f),
	.w3(32'h3b5a08fe),
	.w4(32'hbb887da6),
	.w5(32'h3b94ef90),
	.w6(32'h3a9fa10a),
	.w7(32'h3a83aaaf),
	.w8(32'h3baccdc8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b12f),
	.w1(32'h3afce8dd),
	.w2(32'h3ba76b83),
	.w3(32'h3baef8fc),
	.w4(32'h3af0a710),
	.w5(32'h3a34932e),
	.w6(32'h3b65bb9a),
	.w7(32'h3a8270a1),
	.w8(32'hbb5ff4dd),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7fd7f),
	.w1(32'hbb6fd9cb),
	.w2(32'h3afb9531),
	.w3(32'hbbb4cb7e),
	.w4(32'hbb63d904),
	.w5(32'hb99812b9),
	.w6(32'hbb572b20),
	.w7(32'hbbdcc72f),
	.w8(32'hba80f43b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50f2d0),
	.w1(32'hb9ff4806),
	.w2(32'hba11cc2a),
	.w3(32'h3b1ee4b7),
	.w4(32'hbb0c4b47),
	.w5(32'h394f25d3),
	.w6(32'h3b87d5fc),
	.w7(32'hbb9fc0c2),
	.w8(32'hbb0f1ab8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e753e),
	.w1(32'h39c23190),
	.w2(32'hbc1e2d99),
	.w3(32'hbb713e91),
	.w4(32'h3bca8294),
	.w5(32'h3bce40f6),
	.w6(32'hbbcfeed5),
	.w7(32'h3a29601b),
	.w8(32'h3c37e064),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7ba93),
	.w1(32'hbbf2b8f5),
	.w2(32'hbb85edee),
	.w3(32'hbb7e7854),
	.w4(32'hbba4adc3),
	.w5(32'h3b5ac07d),
	.w6(32'h3b87bd44),
	.w7(32'hb9f478a4),
	.w8(32'hb99eb672),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafd698),
	.w1(32'hba6f5777),
	.w2(32'h3b97153e),
	.w3(32'hbadb8dcd),
	.w4(32'hbb4ac617),
	.w5(32'h3b90a6b2),
	.w6(32'hbb476d7f),
	.w7(32'hba7e59d7),
	.w8(32'h3b722a6f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ddc681),
	.w1(32'hbc0d306b),
	.w2(32'hbb83fcf2),
	.w3(32'h3bae4e04),
	.w4(32'hbafd0eac),
	.w5(32'hbb04d828),
	.w6(32'h3b43a9eb),
	.w7(32'h3aa22f18),
	.w8(32'h3afd154f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892cc21),
	.w1(32'h3af7c8b5),
	.w2(32'h3c889934),
	.w3(32'h3aec785e),
	.w4(32'h3cb1631d),
	.w5(32'h3d1f9f7c),
	.w6(32'h3bceaaa4),
	.w7(32'h3b5a39b2),
	.w8(32'h3b233773),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbe3fe),
	.w1(32'hbb70f114),
	.w2(32'h39cf207b),
	.w3(32'hbb9f2240),
	.w4(32'hbc1cbecc),
	.w5(32'h3b2d27a1),
	.w6(32'hbb8d7042),
	.w7(32'hbc050cbc),
	.w8(32'hbaea76e4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7f3d7),
	.w1(32'h3b36f4e4),
	.w2(32'h3bf96d5c),
	.w3(32'h3bee4d48),
	.w4(32'h3ad318fc),
	.w5(32'h3c2f0e07),
	.w6(32'h3baebac9),
	.w7(32'h3b6622a1),
	.w8(32'h3c364e6f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64f8bd),
	.w1(32'h3b794c0b),
	.w2(32'hba12f34d),
	.w3(32'h3bb3faa5),
	.w4(32'h3bd17ebc),
	.w5(32'h3b19cb76),
	.w6(32'h3c1f4534),
	.w7(32'h3ab73b25),
	.w8(32'h3baa45e3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe02767),
	.w1(32'hbba91d52),
	.w2(32'hbc70cd8b),
	.w3(32'hbc274665),
	.w4(32'h3be2c9aa),
	.w5(32'hbb354af0),
	.w6(32'hbabd1ee1),
	.w7(32'h3ba72953),
	.w8(32'hba882212),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbda86a),
	.w1(32'hbbaf6246),
	.w2(32'h3ab945ce),
	.w3(32'hba5f5e69),
	.w4(32'h3b6bcdc0),
	.w5(32'h3c0be3e0),
	.w6(32'hbb67bf50),
	.w7(32'hbb6a3e81),
	.w8(32'hb9ac53a6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b9195),
	.w1(32'hbb79907b),
	.w2(32'hbb940bef),
	.w3(32'h38aebfba),
	.w4(32'hbb4936aa),
	.w5(32'h3bacc970),
	.w6(32'hbbcdd83e),
	.w7(32'hbb57a2af),
	.w8(32'h3944b5cd),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4559a4),
	.w1(32'hba4e33fb),
	.w2(32'hbade2fee),
	.w3(32'hbbc70928),
	.w4(32'hbbbb36b7),
	.w5(32'hba75ed0a),
	.w6(32'hbbc2b860),
	.w7(32'hbbf01bb1),
	.w8(32'hbb1326dc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c9707),
	.w1(32'hbbaffbac),
	.w2(32'h39fa406d),
	.w3(32'h3b6fbb0d),
	.w4(32'h3b85fe22),
	.w5(32'h3ab5b7ca),
	.w6(32'h3b023ee3),
	.w7(32'hbb8bafce),
	.w8(32'h3b22670e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944734f),
	.w1(32'hbae107d6),
	.w2(32'h3801fc8f),
	.w3(32'h3b48430f),
	.w4(32'h39e25393),
	.w5(32'hbbb4d633),
	.w6(32'h3be0ee5a),
	.w7(32'h39c8f247),
	.w8(32'hbb392343),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade4539),
	.w1(32'hbb7d0278),
	.w2(32'hb975d3ce),
	.w3(32'hbb82defc),
	.w4(32'hbbaa61af),
	.w5(32'hbb367f19),
	.w6(32'h3b32e44d),
	.w7(32'hbb3f67f4),
	.w8(32'hbb080898),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f8030),
	.w1(32'hba6eaae2),
	.w2(32'hba2096b7),
	.w3(32'hbb48fa2d),
	.w4(32'h3a16fe7d),
	.w5(32'hbb694a86),
	.w6(32'hbac94416),
	.w7(32'hbb85bb86),
	.w8(32'hba32fc25),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81fe43),
	.w1(32'hbb5d174d),
	.w2(32'h39ec8b57),
	.w3(32'hba9155d9),
	.w4(32'hbb101961),
	.w5(32'h3b57e069),
	.w6(32'hbb2821d7),
	.w7(32'hbbcdc933),
	.w8(32'hb9596d82),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f8c5f),
	.w1(32'h39cbd0b9),
	.w2(32'h3aefdc55),
	.w3(32'hba977b88),
	.w4(32'h3b20499b),
	.w5(32'h3916346d),
	.w6(32'hbb8ec4da),
	.w7(32'h3b00528a),
	.w8(32'h3a71ac56),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1ea00),
	.w1(32'h3c1d3a07),
	.w2(32'h3bdc0c83),
	.w3(32'hb8b00631),
	.w4(32'hbabcd844),
	.w5(32'h37b1a0a6),
	.w6(32'hbbbcde1b),
	.w7(32'hbc1701a2),
	.w8(32'hbadd1ac1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025959),
	.w1(32'hbaa51734),
	.w2(32'hbb28340a),
	.w3(32'hbb1fe126),
	.w4(32'hbb037c6c),
	.w5(32'hbb9f91ed),
	.w6(32'hbb820e74),
	.w7(32'h3b631822),
	.w8(32'h3aadd8b3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae72a98),
	.w1(32'h3bc1a229),
	.w2(32'h3bc607c8),
	.w3(32'h3a3dcd77),
	.w4(32'h3adcb850),
	.w5(32'h3c212a31),
	.w6(32'h3ae66172),
	.w7(32'h3961daab),
	.w8(32'h3c33e1fd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6e64e),
	.w1(32'hbbd7ba6b),
	.w2(32'h3c1f6347),
	.w3(32'h3c3890ab),
	.w4(32'hbb945344),
	.w5(32'h3c2ef4e3),
	.w6(32'h3b7dd0d1),
	.w7(32'hbc73530c),
	.w8(32'hbc25020a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84f571),
	.w1(32'h396b6cd3),
	.w2(32'hbb6cdc4e),
	.w3(32'hbae46fff),
	.w4(32'h3ac0cb7e),
	.w5(32'hbbd33aed),
	.w6(32'hbc650c65),
	.w7(32'hbbb8b426),
	.w8(32'hbbd2a764),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc6ea0),
	.w1(32'h3a1360d4),
	.w2(32'hba31b92c),
	.w3(32'hbbc3a4cb),
	.w4(32'h3b449c1c),
	.w5(32'h39da3774),
	.w6(32'hbc0b46ab),
	.w7(32'h3b879930),
	.w8(32'hb98b9a2c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa32ecc),
	.w1(32'h383d05a6),
	.w2(32'hbb0e0236),
	.w3(32'hba50ecba),
	.w4(32'hbb362b0d),
	.w5(32'hbb370055),
	.w6(32'hba50bdb3),
	.w7(32'hbb99b1fe),
	.w8(32'hbafcaa87),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857b33),
	.w1(32'h3a8acf3a),
	.w2(32'h3c18886b),
	.w3(32'hbad6c916),
	.w4(32'h3bc16874),
	.w5(32'h3c3dbc4f),
	.w6(32'hbb58288c),
	.w7(32'hb97cee5e),
	.w8(32'h3a1f47bc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeca8ce),
	.w1(32'h3c21495c),
	.w2(32'h3c4f3717),
	.w3(32'hbaf34f42),
	.w4(32'hbae5bf41),
	.w5(32'hb93a1027),
	.w6(32'hbb4312ba),
	.w7(32'hbc938c64),
	.w8(32'hbc8da425),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b287a6),
	.w1(32'hbc1242d2),
	.w2(32'hbc1cc413),
	.w3(32'hbb0745fe),
	.w4(32'h38d9513d),
	.w5(32'hbad48cf8),
	.w6(32'hbc11df89),
	.w7(32'hbbdd5d2a),
	.w8(32'hbc2cd335),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c0f1a),
	.w1(32'h3badfde8),
	.w2(32'h3b82b4cb),
	.w3(32'hbc4613a1),
	.w4(32'h3b896090),
	.w5(32'h3b5da6ca),
	.w6(32'hbc84e52e),
	.w7(32'h3b50f3ae),
	.w8(32'h3bb3a6b9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b493509),
	.w1(32'h3bffe697),
	.w2(32'h3c33e5d9),
	.w3(32'h3a982c01),
	.w4(32'hba8715ce),
	.w5(32'h3b8b9e13),
	.w6(32'h3a364e55),
	.w7(32'hbc169aaf),
	.w8(32'hbc1e85c8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f76ca),
	.w1(32'h38b50599),
	.w2(32'h3b4c444b),
	.w3(32'hbbd84eb9),
	.w4(32'hbbc6899f),
	.w5(32'h3b7d725f),
	.w6(32'hbc6129da),
	.w7(32'hbb96cf29),
	.w8(32'hb963f1d4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11eaba),
	.w1(32'hbc19fa4d),
	.w2(32'h3bbd678c),
	.w3(32'h3ac647c8),
	.w4(32'hbc3bfc79),
	.w5(32'h3c94b9a7),
	.w6(32'h3af1b75a),
	.w7(32'hbb319818),
	.w8(32'h3c86de5e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbeecc),
	.w1(32'h3b6f72f1),
	.w2(32'hbb7147ed),
	.w3(32'h3c77187a),
	.w4(32'h3c361967),
	.w5(32'h3a861318),
	.w6(32'h3c212664),
	.w7(32'h3c09c298),
	.w8(32'h3c0c0e86),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b6681),
	.w1(32'hbb904c0c),
	.w2(32'hbc112907),
	.w3(32'hba8ef1e6),
	.w4(32'h3a8d0356),
	.w5(32'hbc4aad7c),
	.w6(32'hbb32f9c6),
	.w7(32'h3ab0d7cd),
	.w8(32'hbb83a4e9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb419909),
	.w1(32'hbb77833c),
	.w2(32'hb990f17e),
	.w3(32'hbc008326),
	.w4(32'hba212897),
	.w5(32'h3a7dc0ab),
	.w6(32'hbb0096b6),
	.w7(32'hba4ca23b),
	.w8(32'hba451910),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f7bff),
	.w1(32'hbbbb9f33),
	.w2(32'hbb06c68c),
	.w3(32'hbae563bd),
	.w4(32'hbb009a2c),
	.w5(32'h3ba88593),
	.w6(32'h3ae73b9d),
	.w7(32'h3b29160d),
	.w8(32'h3c0919e3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7aa37),
	.w1(32'h386eb72e),
	.w2(32'hb992fc85),
	.w3(32'hbaf414ee),
	.w4(32'hbadda024),
	.w5(32'hbb644fcc),
	.w6(32'h3b892850),
	.w7(32'hbab347bb),
	.w8(32'hbb6ec1cc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f7544),
	.w1(32'h3a524447),
	.w2(32'h3b1cae2a),
	.w3(32'hbac9e165),
	.w4(32'h3a4cd175),
	.w5(32'h3b3aa2eb),
	.w6(32'hbb49a18e),
	.w7(32'h3a189abf),
	.w8(32'h39809a22),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5837e),
	.w1(32'h3ab5ecde),
	.w2(32'hbb9875dd),
	.w3(32'hbb93fcf3),
	.w4(32'h3b8e319d),
	.w5(32'hbaaed8dc),
	.w6(32'hbb3c2c36),
	.w7(32'h3c135890),
	.w8(32'hba89c259),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedc15f),
	.w1(32'h3bb445c1),
	.w2(32'h3af80851),
	.w3(32'h3bf95a30),
	.w4(32'h3bfce707),
	.w5(32'h3a6a10cc),
	.w6(32'hb91c99e2),
	.w7(32'h3bb40ab8),
	.w8(32'hb88e3e78),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5361c2),
	.w1(32'h3aa6776b),
	.w2(32'hbad4bbc6),
	.w3(32'hbb900bbe),
	.w4(32'h3b43a185),
	.w5(32'h3bb31d89),
	.w6(32'hbb18ca43),
	.w7(32'h3b0a555c),
	.w8(32'hba214f8f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66151d),
	.w1(32'h3adcdc16),
	.w2(32'hbb5ba0dc),
	.w3(32'h3b39bfe1),
	.w4(32'h3ac1f6c0),
	.w5(32'hbaa2b625),
	.w6(32'hbabbb812),
	.w7(32'hbb93a6f6),
	.w8(32'h3b784424),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb8bb),
	.w1(32'h3c04de54),
	.w2(32'h3bc1cd17),
	.w3(32'hb94c401b),
	.w4(32'h3b897c09),
	.w5(32'h3b12d612),
	.w6(32'h3bc97b4c),
	.w7(32'h3b379d5c),
	.w8(32'h3a006abe),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b078ad8),
	.w1(32'h38eee5d7),
	.w2(32'h3acdee3a),
	.w3(32'h3a7f80b3),
	.w4(32'h3a4c4564),
	.w5(32'h3abcd965),
	.w6(32'hbb3a65c2),
	.w7(32'hbb1bb4a2),
	.w8(32'hbaf5a2d8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dd526),
	.w1(32'h3b1d9c0e),
	.w2(32'h3a9a14c9),
	.w3(32'h3a779e26),
	.w4(32'hb98e4763),
	.w5(32'hbaa8e6c3),
	.w6(32'hbb2f8355),
	.w7(32'h39519f80),
	.w8(32'hbb99a1e0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb045849),
	.w1(32'h3b478d8c),
	.w2(32'h3bd1140c),
	.w3(32'hbb24d224),
	.w4(32'h3ba907fe),
	.w5(32'h3b5cf535),
	.w6(32'hba66f288),
	.w7(32'h3b34459d),
	.w8(32'h3b3ce340),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e7b9e),
	.w1(32'hbb6a5e14),
	.w2(32'h3b61118f),
	.w3(32'h37ce06ac),
	.w4(32'hba03da77),
	.w5(32'h39566154),
	.w6(32'h394436d0),
	.w7(32'hbbb08103),
	.w8(32'hba8936dd),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9990265),
	.w1(32'h3c15e67c),
	.w2(32'h3b57d57e),
	.w3(32'hba89bf31),
	.w4(32'h3a6dd33f),
	.w5(32'hbb2c304e),
	.w6(32'hbb7395c9),
	.w7(32'h3aee27cd),
	.w8(32'h3b576e42),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82bb66),
	.w1(32'hbae1d38b),
	.w2(32'h3acbcf03),
	.w3(32'h3b789c4d),
	.w4(32'hbb8ae275),
	.w5(32'h3abf278c),
	.w6(32'h3c1b8c9a),
	.w7(32'hbb806d4a),
	.w8(32'hba10a36a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929af41),
	.w1(32'h3aca506d),
	.w2(32'hbb2d2dd2),
	.w3(32'h3ab2257f),
	.w4(32'hbbb27c2e),
	.w5(32'hbbe4e22e),
	.w6(32'hba1214de),
	.w7(32'hbb0bf25f),
	.w8(32'h3b2fc1eb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba082dd6),
	.w1(32'hbb369d63),
	.w2(32'h3bcd7f08),
	.w3(32'hbba38dd9),
	.w4(32'hbb5cc557),
	.w5(32'h3c3a2833),
	.w6(32'h397c088e),
	.w7(32'hbb7dee01),
	.w8(32'h3a987904),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bce4c),
	.w1(32'h3aaba0ea),
	.w2(32'hba8df8ca),
	.w3(32'h3c003480),
	.w4(32'h3b22ac5e),
	.w5(32'h390bb038),
	.w6(32'h3b3604a8),
	.w7(32'h3b4c8db7),
	.w8(32'h383e81cc),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfec258),
	.w1(32'hb8b74608),
	.w2(32'h3b141737),
	.w3(32'hbb86953a),
	.w4(32'h3bb521e0),
	.w5(32'h3b253fad),
	.w6(32'hbbae9e8b),
	.w7(32'h3b7fa90c),
	.w8(32'hba35aabb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40543b),
	.w1(32'hbb1b90d4),
	.w2(32'hbc3f8c33),
	.w3(32'h3b490a31),
	.w4(32'h3c151fa2),
	.w5(32'h3ac356b7),
	.w6(32'hba910fdb),
	.w7(32'h3c8203bb),
	.w8(32'h3c311679),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa58e68),
	.w1(32'h3ab98588),
	.w2(32'h3aee5dc6),
	.w3(32'h38aac891),
	.w4(32'h3ade48a0),
	.w5(32'h3b3551cd),
	.w6(32'h3aa79873),
	.w7(32'hb9c4fd83),
	.w8(32'h39925491),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad125dd),
	.w1(32'hbb76cf4b),
	.w2(32'h3bdf4757),
	.w3(32'hba236039),
	.w4(32'hbc26d25d),
	.w5(32'h3bbbca08),
	.w6(32'hb8cb765c),
	.w7(32'hbb3f76f3),
	.w8(32'h3bdcdb65),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3eebcc),
	.w1(32'h3bc98d27),
	.w2(32'h3c39aa18),
	.w3(32'h3c285bf6),
	.w4(32'hbab6b071),
	.w5(32'h3c5e5196),
	.w6(32'h3c0a9c2b),
	.w7(32'hbb35825c),
	.w8(32'h3b6ef69b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c694),
	.w1(32'h3b823122),
	.w2(32'h3ad19a4a),
	.w3(32'h3bc54505),
	.w4(32'hb9e47e4a),
	.w5(32'h3a514fe5),
	.w6(32'h3b462177),
	.w7(32'hbb8ede37),
	.w8(32'h3b41e552),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86488a),
	.w1(32'h3b696f35),
	.w2(32'hba5d8af6),
	.w3(32'hba051ce1),
	.w4(32'h3b94053a),
	.w5(32'hbb131295),
	.w6(32'h3ba3ec7c),
	.w7(32'h3b5424eb),
	.w8(32'hb846da09),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fe684),
	.w1(32'h3bac885a),
	.w2(32'hbc1f9d99),
	.w3(32'hbb8d2d21),
	.w4(32'hba4013dd),
	.w5(32'hbc6a1e7d),
	.w6(32'hba9d1759),
	.w7(32'hbbbf9314),
	.w8(32'hbc0b014a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36c612),
	.w1(32'hbb480283),
	.w2(32'hbaecf816),
	.w3(32'hbc674e40),
	.w4(32'hba1d332d),
	.w5(32'h3ab2ca2c),
	.w6(32'hbc791c87),
	.w7(32'hbb50f865),
	.w8(32'h3a0f378d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea8c8b),
	.w1(32'hbbc9df56),
	.w2(32'hbb13765e),
	.w3(32'hbc1d1320),
	.w4(32'hbb90b11a),
	.w5(32'hbb8f8699),
	.w6(32'hbb9f4874),
	.w7(32'hbbffa149),
	.w8(32'hbb895afa),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cb802),
	.w1(32'h3ac553f1),
	.w2(32'hb954820b),
	.w3(32'h39485e51),
	.w4(32'h3a94c1a4),
	.w5(32'h3b5e5edb),
	.w6(32'hbad58781),
	.w7(32'h3b01494d),
	.w8(32'h3b9485c3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad53792),
	.w1(32'h3ba34409),
	.w2(32'hb8d418c3),
	.w3(32'hb9ff0621),
	.w4(32'h3bc76189),
	.w5(32'hbb377693),
	.w6(32'hbadb122b),
	.w7(32'h3a791967),
	.w8(32'hba9df2af),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7da535),
	.w1(32'hb9818539),
	.w2(32'hbaf93294),
	.w3(32'hbb368312),
	.w4(32'hba651c2b),
	.w5(32'hb9ff22cb),
	.w6(32'h3b4d942d),
	.w7(32'h3a878f79),
	.w8(32'hbb9c66be),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b1356),
	.w1(32'h3b4890d4),
	.w2(32'h3af9806d),
	.w3(32'hbb3e6367),
	.w4(32'h3b855b26),
	.w5(32'h3be469bf),
	.w6(32'h392ed0eb),
	.w7(32'hb8c59a15),
	.w8(32'h3b935394),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba53e46),
	.w1(32'h3bf34a65),
	.w2(32'hbb4e2cd1),
	.w3(32'h3b2a76e2),
	.w4(32'h3b9b436f),
	.w5(32'hbbb2ea8e),
	.w6(32'h3a23b917),
	.w7(32'h3b90898e),
	.w8(32'hbbd4cc4e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cdff2),
	.w1(32'h3b9b5171),
	.w2(32'hbac4feb4),
	.w3(32'hbb3dfcc0),
	.w4(32'h3c6ef3bf),
	.w5(32'h3b119387),
	.w6(32'hbb5bfa9e),
	.w7(32'h3ba7bb04),
	.w8(32'hba4301f2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5615ae),
	.w1(32'hbb405424),
	.w2(32'h3bc59960),
	.w3(32'hbc1ccc01),
	.w4(32'hbc36960e),
	.w5(32'h3c06ba3f),
	.w6(32'hbc0c194a),
	.w7(32'hbaddd495),
	.w8(32'h3baec7c9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a367d),
	.w1(32'hba409f91),
	.w2(32'hbbf0bf38),
	.w3(32'h3ba58dd9),
	.w4(32'hbb9249b0),
	.w5(32'hbb450079),
	.w6(32'h3c1b1e25),
	.w7(32'hbb121b4f),
	.w8(32'hbab3aec8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba343fe4),
	.w1(32'h3ba6f85e),
	.w2(32'hbbddf6e4),
	.w3(32'h3b08aea7),
	.w4(32'h3b777cd6),
	.w5(32'hba462dbc),
	.w6(32'h3b2a4292),
	.w7(32'h3bd0a536),
	.w8(32'h3aa266da),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd093a6),
	.w1(32'h3a81a2aa),
	.w2(32'h3aedb5d0),
	.w3(32'hbbafc0a8),
	.w4(32'hbab36dc6),
	.w5(32'hbaa5a3bf),
	.w6(32'h3a27d3e4),
	.w7(32'hbbd46367),
	.w8(32'hbc132f72),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affa825),
	.w1(32'h3afa835d),
	.w2(32'hbb7ce4bb),
	.w3(32'h398998f2),
	.w4(32'h3bedeadd),
	.w5(32'h39edf3ce),
	.w6(32'hbb58d0ce),
	.w7(32'h3aafa0ad),
	.w8(32'hbb94c30c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dc3e0),
	.w1(32'hbb583ad8),
	.w2(32'hbb7ecec3),
	.w3(32'hbb6bba5d),
	.w4(32'h3934d6f3),
	.w5(32'h3b3cca93),
	.w6(32'hbb10d050),
	.w7(32'h3b202c42),
	.w8(32'h3b60d0c9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86af0e),
	.w1(32'hbbb6816d),
	.w2(32'hbb5d0ae2),
	.w3(32'h3a562df3),
	.w4(32'hbb00f0ea),
	.w5(32'hbb9e93b1),
	.w6(32'hba4f3572),
	.w7(32'hbb458b7a),
	.w8(32'hbb50cf6f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc297ab2),
	.w1(32'hbb2090ff),
	.w2(32'h3b1ac656),
	.w3(32'hbbbc9ea6),
	.w4(32'hbbce323b),
	.w5(32'hbb772ef0),
	.w6(32'hbb888070),
	.w7(32'hbbb96e73),
	.w8(32'hb9560b09),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55f08b),
	.w1(32'hba27ac19),
	.w2(32'hbb170419),
	.w3(32'hbb8338e3),
	.w4(32'h3be38300),
	.w5(32'h3b43220d),
	.w6(32'hbada5285),
	.w7(32'h3b087e67),
	.w8(32'hbba081c7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9df6e),
	.w1(32'hbc303328),
	.w2(32'hbc18edcd),
	.w3(32'h3b3cf6e2),
	.w4(32'hbb9a13cb),
	.w5(32'h3ab1c173),
	.w6(32'hbbca91d1),
	.w7(32'hbbac03e4),
	.w8(32'hbb47a38c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac26335),
	.w1(32'hbb4600e4),
	.w2(32'h3b9765f6),
	.w3(32'h3c0e7b15),
	.w4(32'hbb4a65bb),
	.w5(32'hba6e6c12),
	.w6(32'hbac5a274),
	.w7(32'hbbd224cb),
	.w8(32'hbbb56093),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf117b3),
	.w1(32'hbb859c05),
	.w2(32'h3ad8f4f6),
	.w3(32'h3aa83f6d),
	.w4(32'hbb9e80a9),
	.w5(32'hbbc5ce07),
	.w6(32'hbabe3441),
	.w7(32'hbabbcae3),
	.w8(32'hbb96cb8b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be4a7d),
	.w1(32'hbb09e373),
	.w2(32'h3b5a7fc2),
	.w3(32'hba28320d),
	.w4(32'hbaa2b3ac),
	.w5(32'h3b910cca),
	.w6(32'h3936743d),
	.w7(32'hbb8cf3af),
	.w8(32'h3b260e71),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39684cbb),
	.w1(32'hbb8c48e1),
	.w2(32'hbb809ec6),
	.w3(32'h3a257430),
	.w4(32'hbb94243f),
	.w5(32'hbbe1b717),
	.w6(32'h3ae3d3d1),
	.w7(32'hbc1a4090),
	.w8(32'hbbb0eaae),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd56db2),
	.w1(32'hbb173b0d),
	.w2(32'h3b21cbc0),
	.w3(32'h3c3b515a),
	.w4(32'hbc0ff787),
	.w5(32'hba1ab886),
	.w6(32'h3ba5d196),
	.w7(32'hbb37d621),
	.w8(32'h3b40476d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514d5c),
	.w1(32'h3c30b8c9),
	.w2(32'h3b7794af),
	.w3(32'h3b5309d2),
	.w4(32'h3b9b1bf8),
	.w5(32'hbbce64ba),
	.w6(32'h3bc2f1cb),
	.w7(32'h3b85f8b4),
	.w8(32'hbb48f6f5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacf811),
	.w1(32'h39d4e082),
	.w2(32'hba8eaab9),
	.w3(32'hbbb5c7aa),
	.w4(32'h3b94a54b),
	.w5(32'h3bcb55e4),
	.w6(32'hbb184293),
	.w7(32'hb9dc3ab7),
	.w8(32'h3b6d2bb2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9560a),
	.w1(32'hbb0bdc2a),
	.w2(32'hbbf72364),
	.w3(32'hbc00b08a),
	.w4(32'hbc261432),
	.w5(32'hbc787d6a),
	.w6(32'hbba9a2e0),
	.w7(32'hbc68a746),
	.w8(32'hbc81ecb4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7a752),
	.w1(32'hbc1d7905),
	.w2(32'hbb6491a0),
	.w3(32'hbc4b33d5),
	.w4(32'hbb9d5e67),
	.w5(32'hbbd7b6a4),
	.w6(32'hbc96d2e7),
	.w7(32'hbb664fc7),
	.w8(32'h3b0941b1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc833ab),
	.w1(32'h3b6cf3c3),
	.w2(32'h3b0cc594),
	.w3(32'h3c52ddf4),
	.w4(32'h3add7c16),
	.w5(32'h3ab2eefd),
	.w6(32'h3c2f57fd),
	.w7(32'h3b284f25),
	.w8(32'h3b1e6cd3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53495b),
	.w1(32'hba171f55),
	.w2(32'h392fbc87),
	.w3(32'h3cabc13c),
	.w4(32'hb9e50eb8),
	.w5(32'hb8dc573b),
	.w6(32'h3c20d98c),
	.w7(32'h38bd1b5f),
	.w8(32'h395f329c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae61fff),
	.w1(32'h39891e66),
	.w2(32'hba1f3df4),
	.w3(32'h3b0018df),
	.w4(32'hb9de1cf6),
	.w5(32'hb9cee73b),
	.w6(32'h3b01f0fb),
	.w7(32'hb990c1b1),
	.w8(32'hb9bbb5f2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bf2a9),
	.w1(32'hb93f2237),
	.w2(32'h38ca1cff),
	.w3(32'hbab1b703),
	.w4(32'hb8ae1781),
	.w5(32'h3a6d7ab5),
	.w6(32'hba8968a6),
	.w7(32'hb980c796),
	.w8(32'hba2aa117),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb824e294),
	.w1(32'h3a0a2adc),
	.w2(32'h3a8d4b87),
	.w3(32'h39994259),
	.w4(32'h39b5922d),
	.w5(32'h3b1835f2),
	.w6(32'hbaaa2fb1),
	.w7(32'h392c4ea5),
	.w8(32'h3a577ea2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb6895),
	.w1(32'hba7f30c5),
	.w2(32'hba8069a6),
	.w3(32'h3b466405),
	.w4(32'hba52b1f7),
	.w5(32'hba03970d),
	.w6(32'h3b35455f),
	.w7(32'hb9beb9bf),
	.w8(32'hba1bb12a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb011810),
	.w1(32'hbb222ef9),
	.w2(32'hbb13d53c),
	.w3(32'hba7dbee1),
	.w4(32'hba945e14),
	.w5(32'hba832dd7),
	.w6(32'hba4a4d62),
	.w7(32'hbb27bcdd),
	.w8(32'hbab3479e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba642d2c),
	.w1(32'hbb1ee5d6),
	.w2(32'hbad05525),
	.w3(32'hbab12453),
	.w4(32'hbacef245),
	.w5(32'hba03a857),
	.w6(32'hbaae358c),
	.w7(32'hbb164fb8),
	.w8(32'hbac48c27),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba956752),
	.w1(32'hba7b2819),
	.w2(32'h3732c45b),
	.w3(32'hba3fbfd8),
	.w4(32'hb9a1df74),
	.w5(32'h3984eb4a),
	.w6(32'hbadc07f0),
	.w7(32'h39921b2c),
	.w8(32'h3acc4811),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa754e0),
	.w1(32'hb9d69b4b),
	.w2(32'hba41d8c6),
	.w3(32'h3aee144d),
	.w4(32'hbad02cba),
	.w5(32'hb9861687),
	.w6(32'h3b107d7a),
	.w7(32'h39e46cdb),
	.w8(32'hba1cc764),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d63125),
	.w1(32'h393a4fa1),
	.w2(32'h3a62fe4e),
	.w3(32'h384b9b1d),
	.w4(32'hb9536c75),
	.w5(32'h39dad7e5),
	.w6(32'hb93bdc89),
	.w7(32'h3a2e5b84),
	.w8(32'h3a9a0745),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af751b7),
	.w1(32'hbb03f18d),
	.w2(32'hba73c7e6),
	.w3(32'h3b2e9794),
	.w4(32'hba6f0bb7),
	.w5(32'h3995ea8e),
	.w6(32'h3a92da49),
	.w7(32'h39cc787e),
	.w8(32'h3ab1a31d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6302fa),
	.w1(32'h3bbd9436),
	.w2(32'h3ba57fe1),
	.w3(32'hba89e6d0),
	.w4(32'h3b7fb176),
	.w5(32'h3b3f5e1e),
	.w6(32'h3930d9f0),
	.w7(32'h3ba81bfc),
	.w8(32'h3b878cfc),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b892a01),
	.w1(32'hba5be702),
	.w2(32'h379f2f5f),
	.w3(32'h3b313b19),
	.w4(32'hba475bf9),
	.w5(32'h38967aa7),
	.w6(32'h3b21d55f),
	.w7(32'hba353e0d),
	.w8(32'hba2a377c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99a633),
	.w1(32'hba8fb1a6),
	.w2(32'hbaaa0dfd),
	.w3(32'h3a81a470),
	.w4(32'hb9df7c97),
	.w5(32'hbabce01a),
	.w6(32'h3a9a7473),
	.w7(32'hba0187b8),
	.w8(32'hba6439b1),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9df054),
	.w1(32'h39af072e),
	.w2(32'hba88e443),
	.w3(32'hbacaff63),
	.w4(32'hba005d95),
	.w5(32'h3942aac0),
	.w6(32'hba99b815),
	.w7(32'hba2fa91d),
	.w8(32'h3ad78f7d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992e4a7),
	.w1(32'hbab1bfe3),
	.w2(32'hbaf00a6b),
	.w3(32'h3a149517),
	.w4(32'hbae98122),
	.w5(32'hb8a55cae),
	.w6(32'h3b0ba0d3),
	.w7(32'hba6e053a),
	.w8(32'hb99a0e01),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80990),
	.w1(32'h3a931949),
	.w2(32'hb9e6b3cd),
	.w3(32'hba9c0c42),
	.w4(32'hba16d985),
	.w5(32'hb85b6633),
	.w6(32'h39545642),
	.w7(32'hbaafc3ce),
	.w8(32'hbb0cf0ff),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4621a),
	.w1(32'h3a94606e),
	.w2(32'hba97bcfa),
	.w3(32'hbaa0f1c4),
	.w4(32'hb8d06c6a),
	.w5(32'h39a6ba0d),
	.w6(32'hbb20491f),
	.w7(32'h38aabec1),
	.w8(32'hbad4aa57),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbe9b5),
	.w1(32'h3b0bbd89),
	.w2(32'h3a2313b1),
	.w3(32'h3914131f),
	.w4(32'h39fa2a7a),
	.w5(32'h3a947b22),
	.w6(32'hb95c8040),
	.w7(32'hba6e8041),
	.w8(32'hbb36b9ad),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ad5c9),
	.w1(32'hba66076d),
	.w2(32'hbac09127),
	.w3(32'h39fe871d),
	.w4(32'hbaa89c76),
	.w5(32'hbb0592a5),
	.w6(32'hba8ddc1b),
	.w7(32'hba2338aa),
	.w8(32'h399104cc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba637786),
	.w1(32'hba361346),
	.w2(32'h38b5298c),
	.w3(32'hb9ca33c4),
	.w4(32'h3a1c1d08),
	.w5(32'h3a659d68),
	.w6(32'hb94adb63),
	.w7(32'h3ad147ce),
	.w8(32'h3abb8906),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39535894),
	.w1(32'hbaefd3c7),
	.w2(32'hba8c552b),
	.w3(32'hb9a909b8),
	.w4(32'hbaf62c9a),
	.w5(32'hba454836),
	.w6(32'h3949d256),
	.w7(32'hbae45a3b),
	.w8(32'hbafff282),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b26df),
	.w1(32'h3b2c5b5e),
	.w2(32'h3afaf161),
	.w3(32'h3a2afacb),
	.w4(32'hb707127c),
	.w5(32'hb8bd0565),
	.w6(32'hb82fd1cf),
	.w7(32'hba45c1cc),
	.w8(32'hba601d7f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a4ff3),
	.w1(32'hba04c125),
	.w2(32'hbb2167b9),
	.w3(32'h39daf9b7),
	.w4(32'h3a84fecb),
	.w5(32'hba38b5c3),
	.w6(32'hba4186a1),
	.w7(32'h39393088),
	.w8(32'hba156697),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba885c5c),
	.w1(32'h3886f537),
	.w2(32'hba32328a),
	.w3(32'hb8f2d9a5),
	.w4(32'h3989130e),
	.w5(32'hba81b7c1),
	.w6(32'hba85e67e),
	.w7(32'hb9a99ce0),
	.w8(32'hb9d1b28d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d809cc),
	.w1(32'hb969a4a6),
	.w2(32'hba619548),
	.w3(32'h3a1f8f95),
	.w4(32'h3a8c6be2),
	.w5(32'h39e0dd9a),
	.w6(32'hb9f231b1),
	.w7(32'h39a4c670),
	.w8(32'h3ab78c92),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a5fa1),
	.w1(32'hb8206d07),
	.w2(32'hb9cad3af),
	.w3(32'hba9bfea3),
	.w4(32'hba9c8b64),
	.w5(32'hba6d6816),
	.w6(32'h3a8fb4e4),
	.w7(32'hbaafad12),
	.w8(32'hba6e6317),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b6626),
	.w1(32'hb87817b1),
	.w2(32'h3a27806f),
	.w3(32'hba28e153),
	.w4(32'hba8d5c43),
	.w5(32'h39581ea5),
	.w6(32'h39fded7c),
	.w7(32'hba2d52fe),
	.w8(32'hba2ed83b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89764d),
	.w1(32'hba831d5f),
	.w2(32'h3b0e49e5),
	.w3(32'h39a13cd4),
	.w4(32'hb944b58e),
	.w5(32'h3b5a3952),
	.w6(32'h3a2b5f35),
	.w7(32'h3960e165),
	.w8(32'h3b2862e0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b291ab0),
	.w1(32'h3b58a4a2),
	.w2(32'h3b461c54),
	.w3(32'h3b144be5),
	.w4(32'h3b87b982),
	.w5(32'h3b681a60),
	.w6(32'h3ae5616a),
	.w7(32'h3b867512),
	.w8(32'h3b85cf34),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b506cef),
	.w1(32'hbae9648f),
	.w2(32'hbb042c38),
	.w3(32'h3b479c2b),
	.w4(32'hb9b63fdf),
	.w5(32'h398c73af),
	.w6(32'h3b93b333),
	.w7(32'h3944f018),
	.w8(32'h3a6c70a2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b2722),
	.w1(32'h3ab6af30),
	.w2(32'h398904a0),
	.w3(32'hba24ac34),
	.w4(32'h3b170677),
	.w5(32'h3ae201bb),
	.w6(32'h3accb93e),
	.w7(32'h3af9a8d7),
	.w8(32'h3b190372),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cffbc),
	.w1(32'hb9b6239f),
	.w2(32'h393b5c88),
	.w3(32'h3af3dafd),
	.w4(32'hba0c971f),
	.w5(32'h39c2c56f),
	.w6(32'h3b079fd8),
	.w7(32'hba14478b),
	.w8(32'h38ef676f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f703b3),
	.w1(32'h38829801),
	.w2(32'hba2f9951),
	.w3(32'hba7200a5),
	.w4(32'hbad9fda7),
	.w5(32'hbaf76ac4),
	.w6(32'hba2db3fe),
	.w7(32'hbab8cd36),
	.w8(32'hbb1fcc17),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d01e0),
	.w1(32'h381c85a9),
	.w2(32'hb815dd35),
	.w3(32'hbb1f420f),
	.w4(32'hbaa7e02d),
	.w5(32'h39a8c9a1),
	.w6(32'hbaed3937),
	.w7(32'hba47bf05),
	.w8(32'hb9a23d2a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb6ef),
	.w1(32'hbb1f2b79),
	.w2(32'hbb4d4414),
	.w3(32'hbab14aec),
	.w4(32'h3926b16e),
	.w5(32'hba043f0e),
	.w6(32'hb9169b81),
	.w7(32'h3992fa99),
	.w8(32'h38b8c312),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170c43),
	.w1(32'hba3507ba),
	.w2(32'hba8457bc),
	.w3(32'hbafd794c),
	.w4(32'hb9aab9e3),
	.w5(32'hba854c8c),
	.w6(32'hbaa84bbb),
	.w7(32'h3a0a3e4e),
	.w8(32'h397ddcf2),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999106f),
	.w1(32'hba588f90),
	.w2(32'hbab39b30),
	.w3(32'h39fece0b),
	.w4(32'hbae6e622),
	.w5(32'hbb130ceb),
	.w6(32'h3a8eb688),
	.w7(32'hbafab7b4),
	.w8(32'hbb2336fb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cdff5),
	.w1(32'hb8e67746),
	.w2(32'hba0a4e7b),
	.w3(32'hbadeee64),
	.w4(32'hba5e0e91),
	.w5(32'hbaab80cb),
	.w6(32'hbaba72d0),
	.w7(32'h3a8a9d01),
	.w8(32'hb8c21572),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b751d),
	.w1(32'hbad00c81),
	.w2(32'hba4f42cc),
	.w3(32'hba63c72f),
	.w4(32'hbaa3acbf),
	.w5(32'hb9a850c1),
	.w6(32'hb9b3febe),
	.w7(32'hbb0aae3d),
	.w8(32'hbb013eeb),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12b7d9),
	.w1(32'hbb2921e6),
	.w2(32'hbb083219),
	.w3(32'hbb2e04fa),
	.w4(32'hb8ea64c4),
	.w5(32'hb9b872d7),
	.w6(32'hbb39fa4d),
	.w7(32'hba8634f5),
	.w8(32'hba196370),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab35c53),
	.w1(32'h3a1651e5),
	.w2(32'hb976213a),
	.w3(32'hbaad293c),
	.w4(32'hba283b2d),
	.w5(32'hb9d587f7),
	.w6(32'hba8d2152),
	.w7(32'hbafea964),
	.w8(32'hbab0cfbf),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9c54e),
	.w1(32'h3ab7f01b),
	.w2(32'h3adc3455),
	.w3(32'hbadbdc6f),
	.w4(32'h39f54a4e),
	.w5(32'h3a8992a2),
	.w6(32'hba28706f),
	.w7(32'h3a9f9b67),
	.w8(32'h3aa0ee6b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2182aa),
	.w1(32'h39b13d9f),
	.w2(32'h39bb6244),
	.w3(32'h3a924eb9),
	.w4(32'hb8ddb77d),
	.w5(32'hbab552c2),
	.w6(32'h3a4057aa),
	.w7(32'hb885e495),
	.w8(32'hbac615a9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9e133),
	.w1(32'hbb6eb60b),
	.w2(32'hbac9336b),
	.w3(32'hbaed8979),
	.w4(32'hbb6b2305),
	.w5(32'hbb0b7760),
	.w6(32'hbae67c59),
	.w7(32'hbb6533ea),
	.w8(32'hbb12c5a6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca0ac6),
	.w1(32'h39eea185),
	.w2(32'hb7f88849),
	.w3(32'hba03d6ed),
	.w4(32'h3adc16a6),
	.w5(32'h39a6b025),
	.w6(32'hbafa603a),
	.w7(32'h3ab325b4),
	.w8(32'h3a5789ec),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef57f3),
	.w1(32'h39aa69a6),
	.w2(32'h39837b7b),
	.w3(32'hba811c71),
	.w4(32'h39ef9523),
	.w5(32'h39a55dbe),
	.w6(32'hba8cfdba),
	.w7(32'h3a296c34),
	.w8(32'h3a57c809),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a085cad),
	.w1(32'hbad5e66d),
	.w2(32'hbb0c8679),
	.w3(32'h3a934f5a),
	.w4(32'hb96fc83d),
	.w5(32'hbb1e23ec),
	.w6(32'h3ab62246),
	.w7(32'hba97506e),
	.w8(32'hbad6f313),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba882a70),
	.w1(32'hba87a48a),
	.w2(32'hbac50d90),
	.w3(32'hba981252),
	.w4(32'h39ee637e),
	.w5(32'hb9512788),
	.w6(32'hba97c8a3),
	.w7(32'h38d83d7d),
	.w8(32'hb94c604a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba668ab6),
	.w1(32'hb9faa103),
	.w2(32'hba3ea182),
	.w3(32'h391ae6c2),
	.w4(32'hba93c908),
	.w5(32'h39d5b987),
	.w6(32'hba5e146a),
	.w7(32'hb9efe430),
	.w8(32'hbaa11d8c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a5ab3),
	.w1(32'h3a6efc7f),
	.w2(32'hbaad8b2d),
	.w3(32'h3a2e5e03),
	.w4(32'h3ac3767f),
	.w5(32'hba3679ce),
	.w6(32'hb9d8b0cb),
	.w7(32'h3aae4659),
	.w8(32'hb8d7d4f0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafe815),
	.w1(32'h3904c46b),
	.w2(32'h39d8144a),
	.w3(32'hbaa6bd30),
	.w4(32'h3a9aa2f5),
	.w5(32'h3a9e4bea),
	.w6(32'hbaad8500),
	.w7(32'h3a2947f6),
	.w8(32'h3a736c3e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5561a5),
	.w1(32'h3a798bde),
	.w2(32'hb95b7253),
	.w3(32'h3b26f990),
	.w4(32'h3a347c0a),
	.w5(32'hbab3925a),
	.w6(32'h3b150484),
	.w7(32'h3a398a0c),
	.w8(32'h3a13c76b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaccd7),
	.w1(32'h3817d86c),
	.w2(32'h3a0a4065),
	.w3(32'hbab09991),
	.w4(32'hba5bc10a),
	.w5(32'hba12f8d6),
	.w6(32'h3a284391),
	.w7(32'hba42ca3f),
	.w8(32'hba432e50),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a9526),
	.w1(32'h3b29af5e),
	.w2(32'h3ae689ed),
	.w3(32'hba8c69c4),
	.w4(32'h3ad438af),
	.w5(32'h3a3f98ff),
	.w6(32'hb819018f),
	.w7(32'h3ad27283),
	.w8(32'h3aa3bb42),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb5af7),
	.w1(32'hba2950fc),
	.w2(32'hbaa755a5),
	.w3(32'hbaa69f5c),
	.w4(32'hba093a47),
	.w5(32'h3a7ba5c6),
	.w6(32'hba163d66),
	.w7(32'hba8947a7),
	.w8(32'h38260572),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae81164),
	.w1(32'hbaa4ac95),
	.w2(32'hba0d91ae),
	.w3(32'hba34fcae),
	.w4(32'h391c0fbf),
	.w5(32'h3a85b83f),
	.w6(32'hb9f7e0f4),
	.w7(32'h3831a7d8),
	.w8(32'h38362eb3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e24fb1),
	.w1(32'hbb4cb354),
	.w2(32'hbb0ee23a),
	.w3(32'h3a167490),
	.w4(32'hbb4243d9),
	.w5(32'hbac6be92),
	.w6(32'hb9138f29),
	.w7(32'hbb858f27),
	.w8(32'hbaf68d8f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00b138),
	.w1(32'hba356a9d),
	.w2(32'hba66cf8b),
	.w3(32'hba57030c),
	.w4(32'hbae42afc),
	.w5(32'hbaec7d20),
	.w6(32'hbaa2802b),
	.w7(32'hbb183e24),
	.w8(32'hbb2625c0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule