module layer_10_featuremap_439(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947c75a),
	.w1(32'hba05e024),
	.w2(32'hba16df9f),
	.w3(32'h3a039a23),
	.w4(32'hba2bfb8a),
	.w5(32'hba506928),
	.w6(32'h39842ad7),
	.w7(32'hba26d4f6),
	.w8(32'hba2dbcaf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42a8c9),
	.w1(32'hb92e97bf),
	.w2(32'hbb53823e),
	.w3(32'h3a910e85),
	.w4(32'hbade6807),
	.w5(32'hbacd0b85),
	.w6(32'hba2930e1),
	.w7(32'hbb188d80),
	.w8(32'hbb038472),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff4855),
	.w1(32'hba17513b),
	.w2(32'hb91e2149),
	.w3(32'hb8dd089c),
	.w4(32'hba658fad),
	.w5(32'hba4a6a1c),
	.w6(32'hb9aad757),
	.w7(32'hba6ca203),
	.w8(32'hba210832),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79f106),
	.w1(32'hbaffc231),
	.w2(32'hba75526d),
	.w3(32'hba817f3c),
	.w4(32'hbabbce02),
	.w5(32'hb951c8df),
	.w6(32'hbac28d05),
	.w7(32'hbabaf1e2),
	.w8(32'hba3b2932),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e5f38),
	.w1(32'hb9f905f4),
	.w2(32'hb9cb6e93),
	.w3(32'hba00bf18),
	.w4(32'hb9da80a9),
	.w5(32'hb8d2f78c),
	.w6(32'hba2dedb9),
	.w7(32'hba03daae),
	.w8(32'hb98807e0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a6032),
	.w1(32'h3a0fbe5e),
	.w2(32'h3a6dc484),
	.w3(32'hb97f0593),
	.w4(32'h3a86b0bd),
	.w5(32'h3a94ffd5),
	.w6(32'hb8bd7968),
	.w7(32'h39e4e955),
	.w8(32'h3a3e31c7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63f3a1),
	.w1(32'hbb80c6dc),
	.w2(32'h3b935254),
	.w3(32'hbbaf19b1),
	.w4(32'hbb006783),
	.w5(32'h3be75c36),
	.w6(32'hbbfbd090),
	.w7(32'hb9d70c8b),
	.w8(32'h3c0cd556),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c334ece),
	.w1(32'h3b6f79e9),
	.w2(32'h3be2924e),
	.w3(32'h3c3cec5d),
	.w4(32'h3c124693),
	.w5(32'hbb030177),
	.w6(32'h3c2eacf4),
	.w7(32'h3bb88529),
	.w8(32'h3b45acfb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c8ab3),
	.w1(32'h3a9ac837),
	.w2(32'h3a270360),
	.w3(32'h3a15aae9),
	.w4(32'h3a8ea8e2),
	.w5(32'h39e5e084),
	.w6(32'hb94db2a4),
	.w7(32'h3a539bf0),
	.w8(32'h3a107d83),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a826981),
	.w1(32'h3ad05328),
	.w2(32'h3b38c2b1),
	.w3(32'hb9ce2061),
	.w4(32'hba0577d9),
	.w5(32'h3b33a7dc),
	.w6(32'h3980125a),
	.w7(32'hb9c48bf7),
	.w8(32'h3b44f340),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55754e),
	.w1(32'hb9812725),
	.w2(32'hba093cb2),
	.w3(32'hb9c567f6),
	.w4(32'h3979b2dc),
	.w5(32'h39917530),
	.w6(32'hb99f5294),
	.w7(32'h394de6c5),
	.w8(32'hb89ffbfc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac8a51),
	.w1(32'hbb903e57),
	.w2(32'h3bc422c0),
	.w3(32'hbbaccda6),
	.w4(32'hbb396fd0),
	.w5(32'h3b9955c4),
	.w6(32'hbbd73635),
	.w7(32'hbb89a475),
	.w8(32'h3ba7aea4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a986ae3),
	.w1(32'h3aa9f42d),
	.w2(32'h3bb0dda4),
	.w3(32'hbb1815c4),
	.w4(32'h3936f967),
	.w5(32'h3b719023),
	.w6(32'hba3f9bf1),
	.w7(32'h3a3ec13c),
	.w8(32'h3b77f667),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba3699),
	.w1(32'h3b4bef42),
	.w2(32'h3ae97c71),
	.w3(32'h3a745052),
	.w4(32'h3b3a0a2c),
	.w5(32'h3a25ce97),
	.w6(32'hba880b90),
	.w7(32'h3a123c73),
	.w8(32'hba00cca1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84f49b),
	.w1(32'hbaa2e992),
	.w2(32'hb9f48dc7),
	.w3(32'hb9b3a56f),
	.w4(32'hbb359103),
	.w5(32'hbaabd8c9),
	.w6(32'hba84583a),
	.w7(32'hbb3f8786),
	.w8(32'hbb1b0daf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b521fa6),
	.w1(32'h3ade68de),
	.w2(32'h392d1a0c),
	.w3(32'h3b53fcac),
	.w4(32'hba57ce50),
	.w5(32'hbb3c5a61),
	.w6(32'h3b3caf6a),
	.w7(32'h3b18daa5),
	.w8(32'h36b031e0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02eac6),
	.w1(32'h39cacda4),
	.w2(32'h3a0b8105),
	.w3(32'hba84728a),
	.w4(32'h39cd4c3a),
	.w5(32'h398b9e85),
	.w6(32'hba27db9e),
	.w7(32'h39ac36c1),
	.w8(32'h389b0fc6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9a1dc),
	.w1(32'h3bf3fbf6),
	.w2(32'h3c84b831),
	.w3(32'h3b64525d),
	.w4(32'h3c30f9b1),
	.w5(32'h3c049ee1),
	.w6(32'h3c0a3214),
	.w7(32'h3c662c3f),
	.w8(32'h3c36e343),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade8a57),
	.w1(32'h3b1d794a),
	.w2(32'h3be560b2),
	.w3(32'h3ace1f3a),
	.w4(32'h3b7eeac5),
	.w5(32'h3b6c51cc),
	.w6(32'h3b48d268),
	.w7(32'h3bb0eaf4),
	.w8(32'h3b9c66d9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d774c),
	.w1(32'hb997feb7),
	.w2(32'hba05ba8f),
	.w3(32'hba280a7b),
	.w4(32'hb9a1607f),
	.w5(32'hb9d3d7f0),
	.w6(32'hb9e8d686),
	.w7(32'hba1d0485),
	.w8(32'hb81d3bed),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56f817),
	.w1(32'h3a88878a),
	.w2(32'h3a0ea06f),
	.w3(32'hba1f5c7f),
	.w4(32'h3aa3059d),
	.w5(32'h3a901dfc),
	.w6(32'hb998262f),
	.w7(32'h3a9900d3),
	.w8(32'h3abed7bc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84fb8f),
	.w1(32'h3a719d49),
	.w2(32'hb8592a20),
	.w3(32'h3a665d67),
	.w4(32'h39ab2881),
	.w5(32'h38acdb49),
	.w6(32'h3a06b18c),
	.w7(32'hb98dfa4d),
	.w8(32'hb9366c3d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b488e41),
	.w1(32'h3ba0fb14),
	.w2(32'h3c93ab1b),
	.w3(32'h3b3e385d),
	.w4(32'hbbd973fc),
	.w5(32'h3c0f4379),
	.w6(32'h3c00b742),
	.w7(32'h3bf27a34),
	.w8(32'h3c657a83),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a138ae6),
	.w1(32'h39849f6b),
	.w2(32'hbb22a385),
	.w3(32'hbab6b86e),
	.w4(32'hbb3a208d),
	.w5(32'hbb0ab250),
	.w6(32'hb9348475),
	.w7(32'hbaf6be45),
	.w8(32'hbaa13664),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb066fc),
	.w1(32'h397b54f0),
	.w2(32'hbbb25ba4),
	.w3(32'h3b7d6519),
	.w4(32'hbb30d8d6),
	.w5(32'hbb269602),
	.w6(32'h3b603fce),
	.w7(32'hbb041d8a),
	.w8(32'hbba7f86b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aadd4),
	.w1(32'h3affc109),
	.w2(32'h3b156f67),
	.w3(32'hba51b4ac),
	.w4(32'h3b579874),
	.w5(32'h3b98293a),
	.w6(32'hb9fb6af5),
	.w7(32'h3b18e604),
	.w8(32'h3b5ceba8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a893689),
	.w1(32'hba4db509),
	.w2(32'hba995135),
	.w3(32'h3aeec10a),
	.w4(32'hbae2f085),
	.w5(32'hbaa23cb6),
	.w6(32'h3abc1faf),
	.w7(32'hbab03e8c),
	.w8(32'hba7f9c1a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a3ce7),
	.w1(32'hbb56b689),
	.w2(32'hba65dfd0),
	.w3(32'hbaa439c2),
	.w4(32'hbb950789),
	.w5(32'hbb63f224),
	.w6(32'hbc23be13),
	.w7(32'hbb64193d),
	.w8(32'hbb8fedf3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60d11a),
	.w1(32'hba13c746),
	.w2(32'h398d8751),
	.w3(32'hbab2fddb),
	.w4(32'hba2f3190),
	.w5(32'hb909047a),
	.w6(32'hbb0302f4),
	.w7(32'hba0855af),
	.w8(32'hb9d390aa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9c22e),
	.w1(32'hbb01a296),
	.w2(32'hbba9c220),
	.w3(32'h3aa5f90c),
	.w4(32'hbb32c23b),
	.w5(32'hbb4cf9e3),
	.w6(32'hbb80e4cd),
	.w7(32'hbb7268de),
	.w8(32'hbb46cea6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12422d),
	.w1(32'h39ff5801),
	.w2(32'h39098d02),
	.w3(32'h3a0b4f2a),
	.w4(32'h3a0a6c91),
	.w5(32'hb972360b),
	.w6(32'h39efc187),
	.w7(32'h39a361c7),
	.w8(32'hb974d577),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a079d29),
	.w1(32'hb988027f),
	.w2(32'hb9b508df),
	.w3(32'h3a493499),
	.w4(32'hb9e7946b),
	.w5(32'hb9e33fd5),
	.w6(32'h3a096c9d),
	.w7(32'hb9aea1ec),
	.w8(32'hb9de8a38),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f8795),
	.w1(32'hb97e3b1a),
	.w2(32'h3ac5d883),
	.w3(32'hba71b1e1),
	.w4(32'hb847124a),
	.w5(32'h3a8cdd54),
	.w6(32'hba2098d4),
	.w7(32'h391a8281),
	.w8(32'h3aa2454f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b746956),
	.w1(32'h3a45a526),
	.w2(32'hbaa37b11),
	.w3(32'h3ab06d92),
	.w4(32'hba17b13f),
	.w5(32'h38eb5c1c),
	.w6(32'h393abe51),
	.w7(32'hbaa08c65),
	.w8(32'hba6e8edc),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc1fa8),
	.w1(32'h3a905b04),
	.w2(32'h3a281433),
	.w3(32'hb9ab6393),
	.w4(32'h3aafd302),
	.w5(32'h3a4bb251),
	.w6(32'hbae7aeed),
	.w7(32'h3a1221bf),
	.w8(32'h3831d201),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e13575),
	.w1(32'hbb18c860),
	.w2(32'h39e85d0d),
	.w3(32'hbaafce9b),
	.w4(32'hbaf264af),
	.w5(32'h3a88be8d),
	.w6(32'hba2dcd5e),
	.w7(32'hbb6503a4),
	.w8(32'h3a222def),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0e97c),
	.w1(32'hbc90a03a),
	.w2(32'h3b023926),
	.w3(32'hb9694ea8),
	.w4(32'hbc8bd0cd),
	.w5(32'hbbbab74a),
	.w6(32'hbae089f0),
	.w7(32'hbc623858),
	.w8(32'h3a7b4ac1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bde28),
	.w1(32'h39342498),
	.w2(32'hbc0fe6aa),
	.w3(32'h3b18dbe1),
	.w4(32'hbbf8f5ff),
	.w5(32'hbc0c1334),
	.w6(32'h3af3ca77),
	.w7(32'hbbebe69a),
	.w8(32'hbbdfb005),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fb1a0),
	.w1(32'hbaee1012),
	.w2(32'hbb3d5bfd),
	.w3(32'h39dd3d48),
	.w4(32'hbb89de5d),
	.w5(32'hba609b70),
	.w6(32'hbbf2a44a),
	.w7(32'hbb75f21c),
	.w8(32'hbb5815ce),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399739e7),
	.w1(32'hbaec586d),
	.w2(32'hbb2bdfde),
	.w3(32'hb9e8e810),
	.w4(32'hbad77660),
	.w5(32'hbaead3d2),
	.w6(32'hb93514f0),
	.w7(32'hbb01f5f8),
	.w8(32'hbb1e240f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0aa012),
	.w1(32'h3a8f5fd5),
	.w2(32'h39ceb3a0),
	.w3(32'hb999fdf6),
	.w4(32'h3a02b0bb),
	.w5(32'h3713d400),
	.w6(32'hba11aed0),
	.w7(32'h3a80db08),
	.w8(32'h3a1724bf),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f735c),
	.w1(32'hba1141a1),
	.w2(32'hba790841),
	.w3(32'h39416fe1),
	.w4(32'hba76b839),
	.w5(32'hba75dbb5),
	.w6(32'h39a0cd14),
	.w7(32'hba44e8af),
	.w8(32'hba817fa8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36da5c),
	.w1(32'h39b8a204),
	.w2(32'hba4d6bbc),
	.w3(32'h3a65e992),
	.w4(32'h39459a72),
	.w5(32'hb8b732a0),
	.w6(32'h3a42c9ee),
	.w7(32'h399d0276),
	.w8(32'h386f0d32),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a453e88),
	.w1(32'h3acd13cd),
	.w2(32'h3bc8b0c4),
	.w3(32'h3b42db90),
	.w4(32'h3b895dd9),
	.w5(32'h3b8d34c6),
	.w6(32'h3b7cea12),
	.w7(32'h3bdfcc09),
	.w8(32'h3b331a00),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80bb43),
	.w1(32'h39cedcc2),
	.w2(32'hbb43ac31),
	.w3(32'h3ab6aad7),
	.w4(32'hbb59993c),
	.w5(32'hbb259087),
	.w6(32'h3a5255a8),
	.w7(32'hbb6cb7dd),
	.w8(32'hbb4b1c9c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d644f),
	.w1(32'h3a816ce3),
	.w2(32'hbae0a485),
	.w3(32'hbb164588),
	.w4(32'hbb4cf686),
	.w5(32'hba029198),
	.w6(32'hb99709e6),
	.w7(32'hbb879bdb),
	.w8(32'hbace16ab),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b993cfa),
	.w1(32'h3ab8dccf),
	.w2(32'hb8bbcd16),
	.w3(32'h3b600d82),
	.w4(32'hb9ca4c1e),
	.w5(32'hba677b26),
	.w6(32'h3b94615d),
	.w7(32'h3ab1daa5),
	.w8(32'h3a6a9018),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd2b8d),
	.w1(32'h3b897cf7),
	.w2(32'h3c9bada6),
	.w3(32'hba979432),
	.w4(32'h3bc64dcd),
	.w5(32'h3c343cc9),
	.w6(32'h3bd98875),
	.w7(32'h3c1a1835),
	.w8(32'h3c4f6692),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48efd9),
	.w1(32'h3aa4dc85),
	.w2(32'h3a8d5b28),
	.w3(32'h3a709d3e),
	.w4(32'h3a481fb8),
	.w5(32'h3a6ea9a1),
	.w6(32'h3a098349),
	.w7(32'h39aed352),
	.w8(32'h3a43afdb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a364be5),
	.w1(32'h3a6628cd),
	.w2(32'h3aa13fb7),
	.w3(32'h39d94762),
	.w4(32'h3a3c375c),
	.w5(32'h3acaf85f),
	.w6(32'h3a4e0aad),
	.w7(32'h3a88f1e0),
	.w8(32'h3aff68b7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929ef57),
	.w1(32'hb9c1ea4b),
	.w2(32'h38eec3a3),
	.w3(32'hba07f42b),
	.w4(32'hb9c34c84),
	.w5(32'hba0b7933),
	.w6(32'hba311470),
	.w7(32'hb7a6a5b8),
	.w8(32'hb94dbdf2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cdcef),
	.w1(32'h3af81d20),
	.w2(32'h3aebd4e8),
	.w3(32'h3b6462a2),
	.w4(32'hb9a02b5a),
	.w5(32'hba532482),
	.w6(32'h3b1a2353),
	.w7(32'h3a6906ac),
	.w8(32'h39b7a279),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeeeb0),
	.w1(32'h3a3d84af),
	.w2(32'h3a7b1441),
	.w3(32'h3a1c150c),
	.w4(32'h3a8df349),
	.w5(32'h3a712fb2),
	.w6(32'h3a96b576),
	.w7(32'h3a715b51),
	.w8(32'h3a7acfbc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995acf2),
	.w1(32'h3bd5aca3),
	.w2(32'h3c757099),
	.w3(32'h3ae2d91d),
	.w4(32'h3c03fbc9),
	.w5(32'h3c0a4fe5),
	.w6(32'h3b07e325),
	.w7(32'h3be80996),
	.w8(32'h3c1abce0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe4021),
	.w1(32'hb704fd4c),
	.w2(32'h3aaecd6a),
	.w3(32'h3a68bb27),
	.w4(32'h390c1041),
	.w5(32'hb98f6554),
	.w6(32'h3a1acbff),
	.w7(32'h386e27aa),
	.w8(32'h39b4ca0a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80ddc2),
	.w1(32'hb9ce0f89),
	.w2(32'hba247731),
	.w3(32'hba94f6b2),
	.w4(32'hba0b0b22),
	.w5(32'hba6dd101),
	.w6(32'hba95a763),
	.w7(32'hba01c405),
	.w8(32'hba8ccce2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cbc84),
	.w1(32'hba3f0408),
	.w2(32'hba15403b),
	.w3(32'hb8aef296),
	.w4(32'hba13e025),
	.w5(32'hba20f705),
	.w6(32'hba6caffe),
	.w7(32'hb9f8f368),
	.w8(32'hb9cca752),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a273d),
	.w1(32'h3a2e5a85),
	.w2(32'hb84ed15a),
	.w3(32'hba0f4bee),
	.w4(32'h3a2e3ee6),
	.w5(32'h39d69a45),
	.w6(32'hba56068e),
	.w7(32'h3a23fa8f),
	.w8(32'hb8d275bf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56aa28),
	.w1(32'hbaa53966),
	.w2(32'hba9d952f),
	.w3(32'hba1f322f),
	.w4(32'hbab7c77a),
	.w5(32'hbaa0a39c),
	.w6(32'hb9560541),
	.w7(32'hba969c5e),
	.w8(32'hba2081e0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59df06),
	.w1(32'hba2a7113),
	.w2(32'h39135626),
	.w3(32'hba4a5ecd),
	.w4(32'h38c4ba49),
	.w5(32'hb92d5715),
	.w6(32'hba101f83),
	.w7(32'hba38d0d4),
	.w8(32'hb9232a1b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399eb128),
	.w1(32'h3a2e4dd5),
	.w2(32'h3b97b134),
	.w3(32'hb9e50767),
	.w4(32'h3b0f8273),
	.w5(32'h3b8ee7d6),
	.w6(32'h39ac8ccf),
	.w7(32'h3b4a35b6),
	.w8(32'h3b890f0b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56e57f),
	.w1(32'h3b9f22c5),
	.w2(32'h3b13f589),
	.w3(32'h3b891e25),
	.w4(32'h3b8945f3),
	.w5(32'h3b122194),
	.w6(32'h3b44f842),
	.w7(32'h3b942997),
	.w8(32'h3ab72b50),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b5061),
	.w1(32'hb95916b4),
	.w2(32'hba1541c3),
	.w3(32'hb9b2d46b),
	.w4(32'h38e2b4e0),
	.w5(32'hba25ea82),
	.w6(32'hba045e60),
	.w7(32'h3956f94a),
	.w8(32'hb9a59f79),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9678bbe),
	.w1(32'h36a59d6e),
	.w2(32'hb93566cc),
	.w3(32'hb9dc53ff),
	.w4(32'hb847a173),
	.w5(32'hba40d597),
	.w6(32'hb8b2b47d),
	.w7(32'hb8c1f738),
	.w8(32'hb9dc2a95),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e1345),
	.w1(32'h396e77a2),
	.w2(32'h39441dbe),
	.w3(32'hba59d289),
	.w4(32'hb687e996),
	.w5(32'hb8f0b0b9),
	.w6(32'hba04b1ff),
	.w7(32'h3989472d),
	.w8(32'hb832e3f3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b5cb6),
	.w1(32'h39f25532),
	.w2(32'h3798226b),
	.w3(32'h3995241a),
	.w4(32'h3899a884),
	.w5(32'h37045641),
	.w6(32'h386ad678),
	.w7(32'h399005d3),
	.w8(32'h380bbc64),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc060af),
	.w1(32'h3aefc404),
	.w2(32'h3c078160),
	.w3(32'h3ab6be46),
	.w4(32'h3b18591b),
	.w5(32'hbaab6595),
	.w6(32'hbbd27189),
	.w7(32'h3a2eaa12),
	.w8(32'h3b272a56),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a534f),
	.w1(32'hb8b35047),
	.w2(32'hb9bab8aa),
	.w3(32'hbb2a7629),
	.w4(32'hbb190c94),
	.w5(32'h3bb00452),
	.w6(32'hb96ef0b2),
	.w7(32'hbba5d4ad),
	.w8(32'h37c8d2da),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d46d6),
	.w1(32'h3bbee7c1),
	.w2(32'h3bdae881),
	.w3(32'h3b697c57),
	.w4(32'h3b8ff814),
	.w5(32'h3bb84b36),
	.w6(32'h3bcd46fc),
	.w7(32'h3c04c4b7),
	.w8(32'h3c240edd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0250d6),
	.w1(32'hbc8d8bf8),
	.w2(32'hbc5915de),
	.w3(32'h3b55717f),
	.w4(32'hbbf3b2a9),
	.w5(32'hbc3f8566),
	.w6(32'h3b433379),
	.w7(32'hbb11b508),
	.w8(32'hbc2d1059),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aa1d6),
	.w1(32'hbb9005fc),
	.w2(32'hbb7a65e0),
	.w3(32'hbc59acf5),
	.w4(32'h3be24e0d),
	.w5(32'h3c440c05),
	.w6(32'hbbd612e1),
	.w7(32'h3c0451fb),
	.w8(32'h3b83530a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad43de5),
	.w1(32'hbb3995ca),
	.w2(32'h39e5352e),
	.w3(32'h3c0a7167),
	.w4(32'h3959dbf5),
	.w5(32'h3c2569d8),
	.w6(32'h3ad54fa1),
	.w7(32'hbbf5ea26),
	.w8(32'hbb8a0c28),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52531e),
	.w1(32'hbb956c2d),
	.w2(32'h3b2b8715),
	.w3(32'hbb333198),
	.w4(32'hbb31ff3c),
	.w5(32'hbbd0b0e9),
	.w6(32'hbc5d85bc),
	.w7(32'hbbb5d7a6),
	.w8(32'hbc8fcffa),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eda74),
	.w1(32'h38c3c7e3),
	.w2(32'h3c19eaf7),
	.w3(32'h3a1b2c78),
	.w4(32'h3b8beee4),
	.w5(32'h3b31438a),
	.w6(32'hbb017821),
	.w7(32'h3b849b74),
	.w8(32'h3b9b8b4b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a723336),
	.w1(32'hbbc6f2ca),
	.w2(32'hbbab0a07),
	.w3(32'h3b0ebcbe),
	.w4(32'h3c4f3e48),
	.w5(32'h3cc99b7a),
	.w6(32'h3b57bcba),
	.w7(32'h3b9164af),
	.w8(32'hbbc1b1e4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398af7ad),
	.w1(32'hbb347f69),
	.w2(32'h3bd48239),
	.w3(32'h3c4f4ef7),
	.w4(32'hb9897867),
	.w5(32'h3c180f39),
	.w6(32'h3b4cb67d),
	.w7(32'h3b27a07f),
	.w8(32'h3bf2d0bc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfaf92),
	.w1(32'h3bb72517),
	.w2(32'h3c48503c),
	.w3(32'h3b08ab8c),
	.w4(32'h3b879f34),
	.w5(32'h3c0975e8),
	.w6(32'h3bdd8f5d),
	.w7(32'hbb2c74df),
	.w8(32'h3bd7bf3c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92e351),
	.w1(32'h3c0af76b),
	.w2(32'h3ca7a89d),
	.w3(32'h3a1c22ec),
	.w4(32'hbbe82506),
	.w5(32'hbc5fcc8f),
	.w6(32'hba2c13b5),
	.w7(32'h3c2b09aa),
	.w8(32'h3cacf25e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b0488),
	.w1(32'hbb722fa2),
	.w2(32'h3b27cd44),
	.w3(32'hbbcbd11c),
	.w4(32'hbaf3baa1),
	.w5(32'h3c112be0),
	.w6(32'h3bb888a0),
	.w7(32'h3c1a4039),
	.w8(32'h3c4b91a3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14073c),
	.w1(32'hb98105bd),
	.w2(32'h3ba4c2da),
	.w3(32'h3c28655c),
	.w4(32'h3b1c6e64),
	.w5(32'h3ba93486),
	.w6(32'hbb2a85d4),
	.w7(32'hbb9dfc9b),
	.w8(32'hbb080d14),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f9c5b),
	.w1(32'h3b483e8b),
	.w2(32'h3a83393a),
	.w3(32'hbbde62ca),
	.w4(32'h3aa54009),
	.w5(32'hbac83d93),
	.w6(32'h3b1bf555),
	.w7(32'h3b999a7b),
	.w8(32'h3bd1d874),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6aadfe),
	.w1(32'hbb1f14ad),
	.w2(32'hb94de69e),
	.w3(32'h3c09c862),
	.w4(32'hbae89745),
	.w5(32'hbb01ea38),
	.w6(32'h3c441f71),
	.w7(32'h3b502c49),
	.w8(32'h3afedd0e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf11ab3),
	.w1(32'h3b65055c),
	.w2(32'hbba49afe),
	.w3(32'hbb8aa7fe),
	.w4(32'h3c1afc71),
	.w5(32'h3c63644b),
	.w6(32'hbbd48309),
	.w7(32'h3c0971cc),
	.w8(32'h3c2d9d90),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b107e36),
	.w1(32'h3ad723cb),
	.w2(32'h3a90a709),
	.w3(32'h3be4f716),
	.w4(32'h3bfb4e44),
	.w5(32'h3c31325c),
	.w6(32'h3ba71a64),
	.w7(32'h3ba2228d),
	.w8(32'h3aea3951),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8ff87),
	.w1(32'hbbb8df23),
	.w2(32'hbaaf6e08),
	.w3(32'h3ba0225f),
	.w4(32'hbc03aaca),
	.w5(32'hbb5dae5a),
	.w6(32'h3b9f1d83),
	.w7(32'hbbd30a89),
	.w8(32'hbc665a0c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8c3d0),
	.w1(32'hb98388f3),
	.w2(32'hbb8cc822),
	.w3(32'hbb851f7f),
	.w4(32'h3ae8268c),
	.w5(32'h3c2ee079),
	.w6(32'hbb03f4f7),
	.w7(32'hbbbc936e),
	.w8(32'h3a2748de),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b645980),
	.w1(32'hbc565966),
	.w2(32'hbc9904f9),
	.w3(32'hbbbee574),
	.w4(32'hbc45c951),
	.w5(32'hbc4dfe5a),
	.w6(32'h3b8518cd),
	.w7(32'hbc04cc3c),
	.w8(32'hbc5f4301),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76af24),
	.w1(32'hbc569d93),
	.w2(32'hbc25437c),
	.w3(32'hbbcd2f3a),
	.w4(32'hbb730985),
	.w5(32'hbbd8216d),
	.w6(32'hbc46f755),
	.w7(32'hbbc99267),
	.w8(32'hbc7c6ef8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc67573),
	.w1(32'h3b110beb),
	.w2(32'hbb650450),
	.w3(32'hbb113e09),
	.w4(32'hbb52350e),
	.w5(32'h3adcad13),
	.w6(32'hb4d8f9e8),
	.w7(32'h3aa22a93),
	.w8(32'h3be4887f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ca434),
	.w1(32'h3a7c2e90),
	.w2(32'h3c308a51),
	.w3(32'h3c1f9404),
	.w4(32'h3b1b696d),
	.w5(32'h3ba7099e),
	.w6(32'h3ca8b869),
	.w7(32'h3c2e2cf3),
	.w8(32'h3c343abf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b343c),
	.w1(32'hbb05d1f9),
	.w2(32'h3b618558),
	.w3(32'hbb38670f),
	.w4(32'hbb94efb1),
	.w5(32'h3b5d8898),
	.w6(32'hbb8f2435),
	.w7(32'hbba93493),
	.w8(32'h3a5881a6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab64e86),
	.w1(32'hbbd12de9),
	.w2(32'h3c367057),
	.w3(32'hbbbd409b),
	.w4(32'hbb5af481),
	.w5(32'h3c19517a),
	.w6(32'hbbca2fb9),
	.w7(32'hbb5635d6),
	.w8(32'h3c1a56dd),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f66ca),
	.w1(32'h3bafe1ac),
	.w2(32'hbc120d71),
	.w3(32'hbacee725),
	.w4(32'h3bbd725f),
	.w5(32'h3cbce2b5),
	.w6(32'h3bc753e7),
	.w7(32'hbb54fcf9),
	.w8(32'hbc4e851c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0315a),
	.w1(32'hb8136a3d),
	.w2(32'hbba443e4),
	.w3(32'h3c3c3a89),
	.w4(32'h3b0bd4bb),
	.w5(32'h3beee68b),
	.w6(32'h3bfdefe0),
	.w7(32'h3b0a1e71),
	.w8(32'h39dc3eda),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71e15c),
	.w1(32'h3b8414f6),
	.w2(32'hb8aadd24),
	.w3(32'h3a0b9e97),
	.w4(32'h3ba7ea33),
	.w5(32'h3c3d218a),
	.w6(32'hbadf27f2),
	.w7(32'h3a988ef9),
	.w8(32'h3bb832ec),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98f76a),
	.w1(32'h3ca33218),
	.w2(32'h3cbdf249),
	.w3(32'h3c1e101d),
	.w4(32'h39bf4926),
	.w5(32'hbc0da014),
	.w6(32'h3bba421a),
	.w7(32'h3b9c60af),
	.w8(32'h3c259d54),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc5bc2),
	.w1(32'hbbde7791),
	.w2(32'hbc671656),
	.w3(32'hb9c8dfcb),
	.w4(32'hb850635f),
	.w5(32'h3c1e35df),
	.w6(32'h3cf12e17),
	.w7(32'hb973a487),
	.w8(32'hbba5026a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc251480),
	.w1(32'h3b817499),
	.w2(32'h3be4f009),
	.w3(32'hbb5ca63e),
	.w4(32'hbb6e6d9f),
	.w5(32'h3ad1fa7a),
	.w6(32'hba0c2c9a),
	.w7(32'hbac0dd98),
	.w8(32'h3b27ac83),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfce28f),
	.w1(32'hbc083fd3),
	.w2(32'h3bbfc68c),
	.w3(32'hbb4556f3),
	.w4(32'hbbe33190),
	.w5(32'hbb587fa5),
	.w6(32'hbbfa004b),
	.w7(32'hbc019f96),
	.w8(32'h3c00b07a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d092),
	.w1(32'hbc16d633),
	.w2(32'h3c245735),
	.w3(32'h3c2b7349),
	.w4(32'hbc9605e3),
	.w5(32'hbb4a5362),
	.w6(32'h3a801b3e),
	.w7(32'hbc185d75),
	.w8(32'hbbcb1edc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4703f),
	.w1(32'hbb472f45),
	.w2(32'hbbe21c68),
	.w3(32'hbb0e3c18),
	.w4(32'hbbe532cb),
	.w5(32'h3afa851e),
	.w6(32'hbb692a48),
	.w7(32'hbb96f8e0),
	.w8(32'hbc0bf41d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a174975),
	.w1(32'h3b72f160),
	.w2(32'hbc995426),
	.w3(32'h3b06ebff),
	.w4(32'hb933ee71),
	.w5(32'h3b88fda9),
	.w6(32'h37c3240c),
	.w7(32'hbbbdc23e),
	.w8(32'hbc2b9d3f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7cce36),
	.w1(32'hbbc1ed24),
	.w2(32'h3a0a0521),
	.w3(32'hbc194c53),
	.w4(32'hbca2645c),
	.w5(32'hbc7e6314),
	.w6(32'h3bf41daa),
	.w7(32'hbbea81a6),
	.w8(32'h3b606bb0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f25c2),
	.w1(32'hbb4ba007),
	.w2(32'hbb6776ad),
	.w3(32'hbb5956d0),
	.w4(32'hbba7247c),
	.w5(32'hbc0cec87),
	.w6(32'h3b206952),
	.w7(32'hbb143384),
	.w8(32'hbbc4dda1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca986b8),
	.w1(32'h3cba5cfb),
	.w2(32'h3c656134),
	.w3(32'h3bd14524),
	.w4(32'h3be334f0),
	.w5(32'h3cb7b293),
	.w6(32'h3af5ba68),
	.w7(32'h3d0b6ad8),
	.w8(32'h3cf22f44),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4a6ce),
	.w1(32'hbb5dc827),
	.w2(32'h3b0e9536),
	.w3(32'h3c9bbc34),
	.w4(32'h3bc1b750),
	.w5(32'h3cae3665),
	.w6(32'h3c9e7744),
	.w7(32'h3b583388),
	.w8(32'h3b106537),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7357c),
	.w1(32'h3b26d552),
	.w2(32'hba9b9791),
	.w3(32'h3c08dd12),
	.w4(32'h3af8393f),
	.w5(32'h3bffe473),
	.w6(32'h3b9f6c98),
	.w7(32'h3b538f9d),
	.w8(32'h3bf2201b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d4718),
	.w1(32'h3b85a77f),
	.w2(32'h3bed8c28),
	.w3(32'hbaf876cc),
	.w4(32'hb9bd9ca6),
	.w5(32'hbabd50e4),
	.w6(32'hbab7152b),
	.w7(32'h3b954545),
	.w8(32'hbb2c0c69),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f0ec2),
	.w1(32'h3939c8bb),
	.w2(32'hbb471101),
	.w3(32'hb9d2a4ef),
	.w4(32'hbb4f7873),
	.w5(32'h3c819a86),
	.w6(32'hbaced4d0),
	.w7(32'h3b3d094b),
	.w8(32'h3ba1c2af),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab0b62),
	.w1(32'h3ca97356),
	.w2(32'h3b08dac1),
	.w3(32'h3b30b0c1),
	.w4(32'h3ca61741),
	.w5(32'h3d04ca2a),
	.w6(32'hbaa98538),
	.w7(32'h3c48a6ee),
	.w8(32'h3b162220),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b552847),
	.w1(32'h3ba20c02),
	.w2(32'h3c8fe77a),
	.w3(32'h3ca6407d),
	.w4(32'hba6ef365),
	.w5(32'hbb949bd3),
	.w6(32'h3cb90e10),
	.w7(32'hb9093df0),
	.w8(32'h3bd59f1a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf55413),
	.w1(32'hbb8be79f),
	.w2(32'hbbc18be2),
	.w3(32'h3bddc27c),
	.w4(32'hbbfbdbce),
	.w5(32'hbc440e6b),
	.w6(32'hb89a9dfa),
	.w7(32'hbb9ccfdb),
	.w8(32'h3ae2ba11),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75755e),
	.w1(32'hbc59be62),
	.w2(32'hbb69fcff),
	.w3(32'hbbd1e45d),
	.w4(32'hbb6618b2),
	.w5(32'h3b858dea),
	.w6(32'hb98fc9ea),
	.w7(32'hbc2a1b2e),
	.w8(32'hbc3de6de),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c0383),
	.w1(32'h3cb3be4b),
	.w2(32'h3c28cd25),
	.w3(32'h3a67c2cd),
	.w4(32'h3923cc9f),
	.w5(32'h3c26e2d3),
	.w6(32'hbc26bbcd),
	.w7(32'h3ab24cc6),
	.w8(32'h3af1952f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae9499),
	.w1(32'h3b781386),
	.w2(32'hbc1a7ccc),
	.w3(32'h3aef1022),
	.w4(32'h37efa7fe),
	.w5(32'h3ac1b3a3),
	.w6(32'hbb100243),
	.w7(32'hbac94e5d),
	.w8(32'h39bb7217),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4edde8),
	.w1(32'hbbb427d7),
	.w2(32'h3a45f204),
	.w3(32'hba5d7ae7),
	.w4(32'h3b040a1a),
	.w5(32'h3be85eda),
	.w6(32'hb9e16cdd),
	.w7(32'h3b67d86c),
	.w8(32'hbb0f8813),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2fd05),
	.w1(32'hbb46792e),
	.w2(32'hbafb7369),
	.w3(32'hbb10eb28),
	.w4(32'hbbd9d846),
	.w5(32'h3c73a2db),
	.w6(32'h3a22992d),
	.w7(32'hbbd197ec),
	.w8(32'hba983009),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9426980),
	.w1(32'hbbbca541),
	.w2(32'hbc85bc29),
	.w3(32'hb995d76f),
	.w4(32'h3b79c38c),
	.w5(32'h3ba46cd2),
	.w6(32'h3c26f8b8),
	.w7(32'hbb166591),
	.w8(32'h3ab42bed),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7df64a),
	.w1(32'h3c2390ca),
	.w2(32'h3cae95a6),
	.w3(32'hbb032bb0),
	.w4(32'h3b41289e),
	.w5(32'hbcb64806),
	.w6(32'h3b102b36),
	.w7(32'h3c19eb05),
	.w8(32'h3cde1b53),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64d4a8),
	.w1(32'hba1da9b7),
	.w2(32'hbbb7b79e),
	.w3(32'h3aa7d9f5),
	.w4(32'h399972f7),
	.w5(32'hbbd463f0),
	.w6(32'h3c930541),
	.w7(32'hbbf43d93),
	.w8(32'hbbc69d2b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5cbb5),
	.w1(32'h3aefd151),
	.w2(32'hbac2cb86),
	.w3(32'hbbd397f5),
	.w4(32'h3a5a29e6),
	.w5(32'h3b9e41de),
	.w6(32'hbb97156d),
	.w7(32'hbb7de796),
	.w8(32'hbb062c7e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c501b59),
	.w1(32'hbbf188b5),
	.w2(32'hbb8444ce),
	.w3(32'hb9d6cadf),
	.w4(32'hbbbd6e39),
	.w5(32'hbacde7c5),
	.w6(32'hbb356e6e),
	.w7(32'hbc0e6c2d),
	.w8(32'hbbd8bde2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3275b),
	.w1(32'hbbfbe0e4),
	.w2(32'hbc6eea42),
	.w3(32'hbc0f783a),
	.w4(32'hbafdb4ee),
	.w5(32'h3c106e4b),
	.w6(32'hbae2385e),
	.w7(32'hbbd5c04e),
	.w8(32'hbc96f15d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12ba55),
	.w1(32'h3b97f4dc),
	.w2(32'hbbd7c99a),
	.w3(32'hbbe46026),
	.w4(32'h39c22e52),
	.w5(32'hbb19d463),
	.w6(32'hbc333524),
	.w7(32'h3bd9efb3),
	.w8(32'hbbf1bcf8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba246f0f),
	.w1(32'hbbc55f9d),
	.w2(32'hbc119467),
	.w3(32'hbbd84117),
	.w4(32'hbc63a8ab),
	.w5(32'hb8ebc2d1),
	.w6(32'h3b01e880),
	.w7(32'hbc47070a),
	.w8(32'hbc444375),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc584a9f),
	.w1(32'h3ba0d17f),
	.w2(32'hba5fe286),
	.w3(32'hbafe5224),
	.w4(32'h3c28cbc0),
	.w5(32'h3c65ffb2),
	.w6(32'hbbc32cbf),
	.w7(32'h3b88c862),
	.w8(32'hbbff9295),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cafe9),
	.w1(32'h3c213078),
	.w2(32'h3bb96636),
	.w3(32'h3bcf374f),
	.w4(32'h3b84c093),
	.w5(32'h3bff32f4),
	.w6(32'hbc91a778),
	.w7(32'h3b8e74be),
	.w8(32'h3b2f27ac),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56a866),
	.w1(32'hbb00e457),
	.w2(32'h3c54b3e3),
	.w3(32'hbbb10429),
	.w4(32'h3b896027),
	.w5(32'h3cab0405),
	.w6(32'hbbfc49ea),
	.w7(32'h3a393030),
	.w8(32'h3a2b44f9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b66097),
	.w1(32'h3b0b5199),
	.w2(32'h3b3fd958),
	.w3(32'hbbfa6fb6),
	.w4(32'h3c28b2d8),
	.w5(32'h3bc00c93),
	.w6(32'hbac15690),
	.w7(32'h3b58936f),
	.w8(32'h3bbf1e49),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93fc8b),
	.w1(32'h39cd43b4),
	.w2(32'h3c039edb),
	.w3(32'h3c239451),
	.w4(32'hbb395f15),
	.w5(32'h3b162c29),
	.w6(32'h3bede6b1),
	.w7(32'hbb496330),
	.w8(32'h3b8240bc),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed974f),
	.w1(32'h3b66204d),
	.w2(32'h3b2c5d1e),
	.w3(32'hbb3e1f27),
	.w4(32'h3ad5b903),
	.w5(32'h3c2143d8),
	.w6(32'hbb2e771c),
	.w7(32'h3b041f0a),
	.w8(32'hbaf93e01),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb150360),
	.w1(32'hbc3de907),
	.w2(32'hbc5882af),
	.w3(32'h3a8e4c18),
	.w4(32'hbc198314),
	.w5(32'hbc46a018),
	.w6(32'h3ad28880),
	.w7(32'hbbab267d),
	.w8(32'hbbff2893),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47bc3f),
	.w1(32'h3bbe18c6),
	.w2(32'hbbd414e5),
	.w3(32'hbc11cc6f),
	.w4(32'h3c1d8937),
	.w5(32'h3c1abb7c),
	.w6(32'hbc8b2942),
	.w7(32'h3b514fad),
	.w8(32'h3c0df009),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7e7f),
	.w1(32'hba7785fd),
	.w2(32'hbc44395b),
	.w3(32'h3b59caa1),
	.w4(32'hbb5e689c),
	.w5(32'hbbdcdcc6),
	.w6(32'h3bebcf5f),
	.w7(32'h3bc1949e),
	.w8(32'h3bdd5db2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd68d79),
	.w1(32'h3c3c75e4),
	.w2(32'h3cf775a0),
	.w3(32'hbb7e0016),
	.w4(32'h38cabb14),
	.w5(32'hbc43bab6),
	.w6(32'hb8e44bf0),
	.w7(32'h3c955f61),
	.w8(32'h3cdb1f2e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4448e8),
	.w1(32'h3b289bc0),
	.w2(32'h39c31ae5),
	.w3(32'hbb2edf82),
	.w4(32'h3ab9fa02),
	.w5(32'hbb235cfa),
	.w6(32'h3c760a08),
	.w7(32'hbb221903),
	.w8(32'hb9426046),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e9640),
	.w1(32'hbc3542b7),
	.w2(32'hba34af80),
	.w3(32'h3b916ff7),
	.w4(32'hbbeba582),
	.w5(32'h3b9277ac),
	.w6(32'h3b665e8e),
	.w7(32'hbb6d58d4),
	.w8(32'h3b9fe378),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20a732),
	.w1(32'h3b437a74),
	.w2(32'h3c0b291e),
	.w3(32'hbbd58022),
	.w4(32'h3bad08b6),
	.w5(32'h3ccc7962),
	.w6(32'hbaff95c4),
	.w7(32'h3c197777),
	.w8(32'h3c8f2f9e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becd9df),
	.w1(32'h3b92b42d),
	.w2(32'hbb08e781),
	.w3(32'h3c2be95d),
	.w4(32'hba14bd2b),
	.w5(32'h3c1d7422),
	.w6(32'hba6a2c33),
	.w7(32'hbbbf9470),
	.w8(32'hbb8e13f5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826fcc),
	.w1(32'h3b98a171),
	.w2(32'h3beeb1d0),
	.w3(32'h3b9581b5),
	.w4(32'h3a4ff78e),
	.w5(32'hbb09f024),
	.w6(32'h3a8b38b6),
	.w7(32'hba8e98d2),
	.w8(32'hbb6c3c6a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed7677),
	.w1(32'h3a3907f1),
	.w2(32'h3c6d3510),
	.w3(32'h3bb2d424),
	.w4(32'h3bb74781),
	.w5(32'h3cd87e29),
	.w6(32'h3bc83edd),
	.w7(32'h3caf58e2),
	.w8(32'h3cc7b8c6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3da10),
	.w1(32'h3bd2e6be),
	.w2(32'hbbce3026),
	.w3(32'h3c3db2a8),
	.w4(32'hbb4889f7),
	.w5(32'h3c44d048),
	.w6(32'h3b810a66),
	.w7(32'h3b81706a),
	.w8(32'h3a904813),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0b4a9),
	.w1(32'hbc73f6c6),
	.w2(32'hbca13990),
	.w3(32'h3c27d6d1),
	.w4(32'hbc4c7f92),
	.w5(32'hbca9e12e),
	.w6(32'h3c392740),
	.w7(32'hbbb5c224),
	.w8(32'hbc153e5e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80c304),
	.w1(32'hbc121bb4),
	.w2(32'hb9d3f0f1),
	.w3(32'hbc8c6130),
	.w4(32'hbb955737),
	.w5(32'hbb0a4ff4),
	.w6(32'hbc4c78b3),
	.w7(32'hbb1a786a),
	.w8(32'hbbc14691),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae22496),
	.w1(32'hbc1af7d3),
	.w2(32'hbc08a06e),
	.w3(32'hbb817115),
	.w4(32'hbc3b6261),
	.w5(32'hbc6b461a),
	.w6(32'hbba0516a),
	.w7(32'hbc337f2a),
	.w8(32'hbc1c3d22),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc237d3e),
	.w1(32'hb7aca84a),
	.w2(32'hbbc478c1),
	.w3(32'hbc59e935),
	.w4(32'hbb9a7013),
	.w5(32'hbb75ef72),
	.w6(32'hbc067e9b),
	.w7(32'hbbc1f25b),
	.w8(32'hba4bd178),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb905270),
	.w1(32'hbbb643bd),
	.w2(32'hbbba5736),
	.w3(32'hb7f3c186),
	.w4(32'hbb948c58),
	.w5(32'hbbc301a9),
	.w6(32'h3c31d915),
	.w7(32'hba99e6c6),
	.w8(32'hbabd7517),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56548c),
	.w1(32'h3b63c04e),
	.w2(32'hbb8d8347),
	.w3(32'hbc01bb75),
	.w4(32'h3b8ec22b),
	.w5(32'hbbb76b84),
	.w6(32'hba6dc2ed),
	.w7(32'hbae1d64d),
	.w8(32'h3b05a803),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee8394),
	.w1(32'h3bb1f106),
	.w2(32'hbb8d78e5),
	.w3(32'hbbf90c0d),
	.w4(32'h3af80a87),
	.w5(32'h3b6a8a2a),
	.w6(32'hbb9c07b5),
	.w7(32'h3b7ceb3a),
	.w8(32'h3a239232),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabbc59),
	.w1(32'h3bbb765d),
	.w2(32'hbb66021d),
	.w3(32'h3baa49f9),
	.w4(32'h3924e669),
	.w5(32'h3b7af88a),
	.w6(32'h3b2d8a04),
	.w7(32'hbb94e968),
	.w8(32'h3baa1b8e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac344f),
	.w1(32'hbc1866b8),
	.w2(32'hbbe15f5c),
	.w3(32'hbc4c8e1d),
	.w4(32'h37ca026a),
	.w5(32'hbab2c875),
	.w6(32'hbbe8fb90),
	.w7(32'hbab2ab9c),
	.w8(32'h3b85db13),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a094cb1),
	.w1(32'h3a9135e2),
	.w2(32'h3b7f9093),
	.w3(32'hbc01b892),
	.w4(32'h3c13c1ec),
	.w5(32'h3b87e88f),
	.w6(32'hbad842bd),
	.w7(32'hb90691b2),
	.w8(32'h3a7457e5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1081ca),
	.w1(32'hbbacd20e),
	.w2(32'hbb833eb0),
	.w3(32'hbb46ba25),
	.w4(32'hbc28715e),
	.w5(32'hbbfc6afc),
	.w6(32'hbc65f378),
	.w7(32'hbb855ebe),
	.w8(32'hbb2c8f1e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c12a77),
	.w1(32'hbb423419),
	.w2(32'hbbf21073),
	.w3(32'hbb5f7d5c),
	.w4(32'h3b00f969),
	.w5(32'h3b9156f2),
	.w6(32'hbb16b0e3),
	.w7(32'h3aa925db),
	.w8(32'h3b6e2123),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85d418),
	.w1(32'h3ba4458d),
	.w2(32'h3bb73fff),
	.w3(32'hbb8092d7),
	.w4(32'hbae4019f),
	.w5(32'h3bd0c07b),
	.w6(32'h39674014),
	.w7(32'h3b72d59f),
	.w8(32'h3a8bf98a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7388ea),
	.w1(32'hbad484b2),
	.w2(32'hba01232a),
	.w3(32'h3bba53fc),
	.w4(32'hbb4ebaa6),
	.w5(32'hbbda6967),
	.w6(32'h3c0839ec),
	.w7(32'hbad8dc04),
	.w8(32'hba9ed81e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dfd70f),
	.w1(32'hbc1ff35e),
	.w2(32'hbc1059f8),
	.w3(32'hbb030f30),
	.w4(32'hbc291572),
	.w5(32'hbbea2bb3),
	.w6(32'h3ba69d67),
	.w7(32'hbbbf67a0),
	.w8(32'hbb4787db),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fe9eb),
	.w1(32'hb947b769),
	.w2(32'h3b1805fc),
	.w3(32'h398cef99),
	.w4(32'hbb0be0c5),
	.w5(32'hbbc2f79c),
	.w6(32'hbbabe8b5),
	.w7(32'hb8cfd388),
	.w8(32'hbb86e043),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b500e59),
	.w1(32'hb9366d6b),
	.w2(32'h3bc4e98f),
	.w3(32'hbb292f9e),
	.w4(32'hbbf2708a),
	.w5(32'hbc63a0f5),
	.w6(32'hb93b6266),
	.w7(32'h3b17c9f7),
	.w8(32'h3b33cea5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01e68a),
	.w1(32'hbbdd0adf),
	.w2(32'h398a81f1),
	.w3(32'hbb019cfb),
	.w4(32'hbbcb24f5),
	.w5(32'hbb944102),
	.w6(32'h3a43536b),
	.w7(32'hb99314f9),
	.w8(32'hba459820),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb469083),
	.w1(32'h3afd0d58),
	.w2(32'h3b5c9c60),
	.w3(32'hbc28fba9),
	.w4(32'hbbcc81ca),
	.w5(32'h3a17318a),
	.w6(32'hb943e63c),
	.w7(32'hbc2b762c),
	.w8(32'hbc07a0e6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbad86f),
	.w1(32'h3a0dcf93),
	.w2(32'h3beeb269),
	.w3(32'hba4b6054),
	.w4(32'hbbc37b6b),
	.w5(32'hbc0bf4ea),
	.w6(32'hbbc36484),
	.w7(32'hbb8e7f12),
	.w8(32'hbad25923),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf1be1),
	.w1(32'hba4bcd2b),
	.w2(32'hbbaff9ac),
	.w3(32'hbbb61b14),
	.w4(32'h3c0882d7),
	.w5(32'h3c16d00d),
	.w6(32'h3bfd3f29),
	.w7(32'h3af22c92),
	.w8(32'h3b98383b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4fb5f),
	.w1(32'hbbc86309),
	.w2(32'hbb9a0faf),
	.w3(32'h3c5151f7),
	.w4(32'h3a75e96e),
	.w5(32'hbbc1861d),
	.w6(32'h3bac5064),
	.w7(32'hbbbc897a),
	.w8(32'hbb8d8210),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27b81c),
	.w1(32'hbb2a3106),
	.w2(32'hbaa7909b),
	.w3(32'h3b106da2),
	.w4(32'hbc12101f),
	.w5(32'h3c678483),
	.w6(32'hbbad9ff5),
	.w7(32'hbc64da54),
	.w8(32'hbb141b07),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0da9f),
	.w1(32'h3a470d3c),
	.w2(32'h3b5ab61c),
	.w3(32'h3ab9e218),
	.w4(32'hbb0eb367),
	.w5(32'h3c573c1b),
	.w6(32'h3a4d52cb),
	.w7(32'h3be16224),
	.w8(32'h3ccdb5fa),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbd414),
	.w1(32'h3c3df5ae),
	.w2(32'h3c9226c4),
	.w3(32'h3b812991),
	.w4(32'h3c1226bc),
	.w5(32'h3cbc8900),
	.w6(32'h3c229f2b),
	.w7(32'h3bbb2a13),
	.w8(32'h3bc154a0),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3027a),
	.w1(32'hbbf47c05),
	.w2(32'hbc34ff95),
	.w3(32'h3c17f2c8),
	.w4(32'hbc22c312),
	.w5(32'hbbec89cc),
	.w6(32'h3c9d7aa9),
	.w7(32'hbbe8ff00),
	.w8(32'h3b8a0da9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf78fb9),
	.w1(32'h38d55000),
	.w2(32'h3b130ab4),
	.w3(32'hbba40365),
	.w4(32'h3bc3a9ff),
	.w5(32'h3b3f3f0e),
	.w6(32'h3afb2b13),
	.w7(32'h3b94fefd),
	.w8(32'h3c2dd2e5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02ccb7),
	.w1(32'hb9ef47d1),
	.w2(32'hbc3e1501),
	.w3(32'h3aaf0166),
	.w4(32'hbc1243f9),
	.w5(32'hbb90a1a1),
	.w6(32'h398edb34),
	.w7(32'hbb9aceb1),
	.w8(32'h3aa6611c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099dc2),
	.w1(32'hbb8e4a53),
	.w2(32'h3bb34d11),
	.w3(32'hbc2b55a0),
	.w4(32'h3b106290),
	.w5(32'h3c6cf7f2),
	.w6(32'h3901a083),
	.w7(32'hb8cf1f56),
	.w8(32'h38831257),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1458f6),
	.w1(32'hbb5e4fcf),
	.w2(32'hbbfc835c),
	.w3(32'hbb848535),
	.w4(32'hbc227401),
	.w5(32'hbc20856a),
	.w6(32'hbc2d98d6),
	.w7(32'hbc65f8bd),
	.w8(32'hbc0760ea),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ef7e),
	.w1(32'hbb1dd72d),
	.w2(32'h3b846bd9),
	.w3(32'hba5be81b),
	.w4(32'h3c168a6d),
	.w5(32'h3bc488c6),
	.w6(32'hbb65d4df),
	.w7(32'h3b529afe),
	.w8(32'hbc234504),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71818c),
	.w1(32'hbb1debf0),
	.w2(32'h3c8541ee),
	.w3(32'hba56d50e),
	.w4(32'h3b02baaf),
	.w5(32'h3bbc42fb),
	.w6(32'hbc0c3b33),
	.w7(32'h3b43f48d),
	.w8(32'hbb201500),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b884d1b),
	.w1(32'h3c6641c8),
	.w2(32'h3b8920a9),
	.w3(32'h3bddcf33),
	.w4(32'h3c538e67),
	.w5(32'h3ca0756d),
	.w6(32'h3c0cc4ae),
	.w7(32'h3c8edefc),
	.w8(32'h3c037147),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c240c93),
	.w1(32'hbbe21520),
	.w2(32'hbbce1749),
	.w3(32'h3c11290b),
	.w4(32'hbb27c041),
	.w5(32'hbbca4590),
	.w6(32'h3bef2d94),
	.w7(32'hbb8cc0d1),
	.w8(32'hbbaacfb0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc191ff6),
	.w1(32'h3b9ea414),
	.w2(32'h3b58a821),
	.w3(32'hbbd05c99),
	.w4(32'h3bbc09ba),
	.w5(32'hb9f7c5a6),
	.w6(32'hbb8dae9e),
	.w7(32'h38c3f0c0),
	.w8(32'h3ba873bf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac29be0),
	.w1(32'h3b0db371),
	.w2(32'h38909f39),
	.w3(32'h3be22838),
	.w4(32'h3b9581b0),
	.w5(32'h3aa2297b),
	.w6(32'h3c5d76cc),
	.w7(32'hba29abed),
	.w8(32'h3bbe75f7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5830fb),
	.w1(32'hbb266124),
	.w2(32'hbbdbcc0e),
	.w3(32'h3bb6d1ea),
	.w4(32'hbb9d77c0),
	.w5(32'h3bb88c06),
	.w6(32'h39ce97e5),
	.w7(32'h3aa624e2),
	.w8(32'h3c27fd2c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf2525),
	.w1(32'h3bdc9d48),
	.w2(32'hba9ce186),
	.w3(32'hbb6a5565),
	.w4(32'h3b8ebbbe),
	.w5(32'hbb608676),
	.w6(32'hbb82e7bc),
	.w7(32'h3b2ac306),
	.w8(32'hbbb711c5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1b242),
	.w1(32'h3b649d16),
	.w2(32'h3b542a5c),
	.w3(32'h3b4ccf87),
	.w4(32'h39ef8da9),
	.w5(32'hbc54efe2),
	.w6(32'h3bbee6d7),
	.w7(32'h3bfe1432),
	.w8(32'h3c2158bb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f13c),
	.w1(32'h3ac2b4dc),
	.w2(32'h3b898432),
	.w3(32'h3b4c597f),
	.w4(32'h3b83b875),
	.w5(32'h3ba95107),
	.w6(32'h3be88199),
	.w7(32'h3bb5d29e),
	.w8(32'h3a49614a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0db3d),
	.w1(32'hbb33ae0e),
	.w2(32'h3ba53b44),
	.w3(32'h3b571e30),
	.w4(32'hbab01d93),
	.w5(32'h3a94f8ca),
	.w6(32'h3bd09946),
	.w7(32'h3c165342),
	.w8(32'h3c60004f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c307a9b),
	.w1(32'hba97e9e5),
	.w2(32'h3af3c921),
	.w3(32'h3b3dcd08),
	.w4(32'hba03900a),
	.w5(32'hbb5d56eb),
	.w6(32'h3bf0a2ee),
	.w7(32'h3bec1ab7),
	.w8(32'h3b0431cd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b4e0d),
	.w1(32'h3b02f158),
	.w2(32'hb936b36d),
	.w3(32'hbc85bf4b),
	.w4(32'hbb05a7ff),
	.w5(32'h3be6303f),
	.w6(32'hbc30f58c),
	.w7(32'h3b8555a9),
	.w8(32'h3bb92a8e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8756f),
	.w1(32'hbb66a65b),
	.w2(32'hbc087a22),
	.w3(32'h397a28f6),
	.w4(32'hbc48e8b0),
	.w5(32'hbc5f2ebd),
	.w6(32'hbb5450b6),
	.w7(32'hbc277ac8),
	.w8(32'hbc0d917f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc96d9),
	.w1(32'h3af5d6dd),
	.w2(32'h3c0c51a4),
	.w3(32'h3a265c9f),
	.w4(32'hb89386c5),
	.w5(32'h3b9c8c89),
	.w6(32'hbb443603),
	.w7(32'h3ad77f0e),
	.w8(32'hbb444b29),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c586017),
	.w1(32'h3b168387),
	.w2(32'h3c82c5ff),
	.w3(32'hba96fcb9),
	.w4(32'h3b7999fd),
	.w5(32'h3c1c8b65),
	.w6(32'hb997bdde),
	.w7(32'h3bfa3a91),
	.w8(32'h3bf870dc),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2122d7),
	.w1(32'h3c212dc9),
	.w2(32'h3c70c638),
	.w3(32'h3c247f8b),
	.w4(32'hbbb8c709),
	.w5(32'hbc96fe38),
	.w6(32'hbc44d2f7),
	.w7(32'h3a980978),
	.w8(32'h3b8975d9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08eb05),
	.w1(32'hbb3820d9),
	.w2(32'h3b54afc0),
	.w3(32'h3b4bab5e),
	.w4(32'hbbe77339),
	.w5(32'hbaee7841),
	.w6(32'hbb8a974c),
	.w7(32'hbb87567c),
	.w8(32'h3a24d4bb),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b530d2b),
	.w1(32'hbc117caf),
	.w2(32'hbb6b5585),
	.w3(32'hb9659b51),
	.w4(32'hbb049b77),
	.w5(32'h3bc7d699),
	.w6(32'h3b57df42),
	.w7(32'h3a9f558b),
	.w8(32'h3a16eaec),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95958f),
	.w1(32'hbaacc626),
	.w2(32'hb97e03f7),
	.w3(32'h3b83a209),
	.w4(32'h3c086a14),
	.w5(32'h3be094f4),
	.w6(32'hbc16f6a8),
	.w7(32'h3b1f3570),
	.w8(32'h3a517058),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bf9d5),
	.w1(32'hbc0c7892),
	.w2(32'hbc1afe9c),
	.w3(32'h3b8c847e),
	.w4(32'h3b106d97),
	.w5(32'h3b855848),
	.w6(32'h3ab6b74f),
	.w7(32'h3bda8cff),
	.w8(32'h3c40bf77),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e454c),
	.w1(32'h3b7f331c),
	.w2(32'h3bf8b868),
	.w3(32'h3b9e30ae),
	.w4(32'h3a0aed23),
	.w5(32'h3c3e1a0e),
	.w6(32'h3bb5eaf7),
	.w7(32'h3989d5e7),
	.w8(32'h3bd9a96e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1c2e2),
	.w1(32'h3c5164ff),
	.w2(32'h3c2a0a1a),
	.w3(32'h3b3f79a1),
	.w4(32'h3ac20a5b),
	.w5(32'h3c562a93),
	.w6(32'h3c95bb77),
	.w7(32'hba3bc8b6),
	.w8(32'h3ac63c1f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19e81a),
	.w1(32'hbb80bab6),
	.w2(32'h3bcf14ab),
	.w3(32'h3c07a60c),
	.w4(32'h3b023c56),
	.w5(32'h3b767e76),
	.w6(32'h3b6ea316),
	.w7(32'hbb10fffd),
	.w8(32'hbb9de489),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7a26a),
	.w1(32'hbb6edc6e),
	.w2(32'hbbd477e8),
	.w3(32'h3a85e301),
	.w4(32'hbc0bba41),
	.w5(32'hbc15d6af),
	.w6(32'h3ba1b9a9),
	.w7(32'hbc46ff1a),
	.w8(32'hbba70154),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904f75),
	.w1(32'hbac6feaa),
	.w2(32'h3b9c4fb7),
	.w3(32'hbc4db052),
	.w4(32'hbaca2521),
	.w5(32'h3b894b43),
	.w6(32'hbc24f49b),
	.w7(32'hb96318ca),
	.w8(32'h3b7e1279),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c9fe8),
	.w1(32'h3a100d07),
	.w2(32'hb7e42555),
	.w3(32'h39a3533a),
	.w4(32'hbae4c1f4),
	.w5(32'h3add4dd0),
	.w6(32'h3b00cec4),
	.w7(32'hba9a178a),
	.w8(32'h3a67c9a3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63904c),
	.w1(32'hba450333),
	.w2(32'hba391414),
	.w3(32'h3a93b9aa),
	.w4(32'hba0fb4da),
	.w5(32'hb971812b),
	.w6(32'h3a71a984),
	.w7(32'hbab62007),
	.w8(32'hbad04141),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb29e21),
	.w1(32'h3b2aa957),
	.w2(32'h3aa7b3c2),
	.w3(32'h3b497292),
	.w4(32'h3a72ba81),
	.w5(32'h3a97adf0),
	.w6(32'h3aef2132),
	.w7(32'h3ac563fb),
	.w8(32'hba8230d8),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41c964),
	.w1(32'h38977d41),
	.w2(32'h389f5d89),
	.w3(32'h3b28fd4a),
	.w4(32'hb9c24b76),
	.w5(32'h396d7b08),
	.w6(32'h3b20ba7b),
	.w7(32'h38bbd13f),
	.w8(32'hb88811c7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba686da3),
	.w1(32'hbb0a6347),
	.w2(32'h37a591c1),
	.w3(32'h39ee995f),
	.w4(32'hba954d80),
	.w5(32'h3a2a243a),
	.w6(32'h3a4e5098),
	.w7(32'hbb3bcdda),
	.w8(32'hba81a294),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9b77),
	.w1(32'h3a5abf11),
	.w2(32'hbb342dec),
	.w3(32'h3a243b5d),
	.w4(32'hbb66bc13),
	.w5(32'hbb63a712),
	.w6(32'hba84de15),
	.w7(32'hbaff463c),
	.w8(32'hbb1c2aca),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c1978),
	.w1(32'h38772aae),
	.w2(32'h3997eb6d),
	.w3(32'hb9f9f645),
	.w4(32'hbb09f347),
	.w5(32'h39eb3554),
	.w6(32'hbaa38aea),
	.w7(32'hbb588e98),
	.w8(32'hb80afd81),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980dae7),
	.w1(32'h3a20aef7),
	.w2(32'h3a6ec14a),
	.w3(32'h39cd0965),
	.w4(32'hbaad8650),
	.w5(32'hba4d05aa),
	.w6(32'h3a80a649),
	.w7(32'h3921d21f),
	.w8(32'hba834741),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8189f8),
	.w1(32'h3992fbaf),
	.w2(32'hbb45e3a6),
	.w3(32'h3af3203c),
	.w4(32'hbb1babd9),
	.w5(32'hbb4514d7),
	.w6(32'hbb1a9b22),
	.w7(32'hbb76c028),
	.w8(32'hbb84ac8b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0f048),
	.w1(32'h3a9c3c0b),
	.w2(32'h3b414c4b),
	.w3(32'h3a8908af),
	.w4(32'h3a209a58),
	.w5(32'h3b609d3d),
	.w6(32'h3a183681),
	.w7(32'h3b10ec33),
	.w8(32'h3b6c8807),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78d0fb),
	.w1(32'h3afb2e80),
	.w2(32'h3b71c0b0),
	.w3(32'h3a2e1729),
	.w4(32'h3ab3b69f),
	.w5(32'h3ade6a49),
	.w6(32'h3a1503f7),
	.w7(32'h3a73d568),
	.w8(32'h3aea315e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f6a85),
	.w1(32'hbab8fa2a),
	.w2(32'hba7d2d56),
	.w3(32'h3a73edab),
	.w4(32'hbaf1f0c3),
	.w5(32'hbaa68aef),
	.w6(32'h3a730c69),
	.w7(32'hbaace6ee),
	.w8(32'hbaa7fc16),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ee9c2),
	.w1(32'h3a09e106),
	.w2(32'h392213c0),
	.w3(32'hba8d1be4),
	.w4(32'h3a514b7c),
	.w5(32'h38fcb615),
	.w6(32'hba7d5ab5),
	.w7(32'h3aabbf94),
	.w8(32'h3a255a51),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa1666),
	.w1(32'hbb7de565),
	.w2(32'hba8773b0),
	.w3(32'hbba1785f),
	.w4(32'hbb9fa2e4),
	.w5(32'h3be4529c),
	.w6(32'hbb739c88),
	.w7(32'hbbcd5e8e),
	.w8(32'h3b43650e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2bbf9),
	.w1(32'h3adea9a9),
	.w2(32'h3b35bcc1),
	.w3(32'h39df340b),
	.w4(32'hb8818586),
	.w5(32'h3b268967),
	.w6(32'h3bbe479b),
	.w7(32'h3b8115d8),
	.w8(32'h3bb59d1a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5657d2),
	.w1(32'hbb0c8ecb),
	.w2(32'hbb87edd4),
	.w3(32'h39937395),
	.w4(32'hbb52d8cc),
	.w5(32'hbb0bc8dc),
	.w6(32'h3a4fec75),
	.w7(32'hbb567c58),
	.w8(32'hbb63f1a8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd5d2f),
	.w1(32'hbb8e0f79),
	.w2(32'h3b5aa2fa),
	.w3(32'hbb05d021),
	.w4(32'hbb68c040),
	.w5(32'hbb7e627b),
	.w6(32'hbc35eadc),
	.w7(32'hbb34c6db),
	.w8(32'h3a82f26a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07ed36),
	.w1(32'h3af56093),
	.w2(32'hb964208b),
	.w3(32'hba193dc1),
	.w4(32'hba293707),
	.w5(32'hb9816545),
	.w6(32'hb9979e2f),
	.w7(32'h3993d36f),
	.w8(32'h38caa5fd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7740f5),
	.w1(32'h3ac44d82),
	.w2(32'h3ac01a13),
	.w3(32'h38d50450),
	.w4(32'h3a319449),
	.w5(32'h39d7887f),
	.w6(32'hb884ae97),
	.w7(32'h39392c1b),
	.w8(32'h3ae69ed7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d317bd),
	.w1(32'hbc3a528f),
	.w2(32'h3b8ed2aa),
	.w3(32'hbab7f4b6),
	.w4(32'hbc21432b),
	.w5(32'h3ba4b0ce),
	.w6(32'h3b190646),
	.w7(32'hbc1e9e24),
	.w8(32'h38a78ed6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6526a),
	.w1(32'h3b42c2c4),
	.w2(32'h3c12f611),
	.w3(32'hbac6d9d8),
	.w4(32'h3b89f8e7),
	.w5(32'h3bbe8775),
	.w6(32'h3b0de506),
	.w7(32'h3baab1c0),
	.w8(32'h3be8c92e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3be4e),
	.w1(32'hbbf056c4),
	.w2(32'h39caa5a8),
	.w3(32'hbb7c1a2f),
	.w4(32'hbbc68222),
	.w5(32'h3a82046c),
	.w6(32'h3ae58869),
	.w7(32'hbb61f128),
	.w8(32'h3b5584c4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2592f),
	.w1(32'h3aad000e),
	.w2(32'hbacb8a0f),
	.w3(32'h3aa4f6e0),
	.w4(32'h387751e0),
	.w5(32'hbb473bca),
	.w6(32'h3a85fb75),
	.w7(32'hb9cea6f4),
	.w8(32'hbb2b0ed9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf2cb6),
	.w1(32'h3ac1d2e2),
	.w2(32'hbb3ff08f),
	.w3(32'h3b85f747),
	.w4(32'hbb22e6a9),
	.w5(32'hbb9376b9),
	.w6(32'h3b0f0649),
	.w7(32'hbabebf47),
	.w8(32'hbb30c3e9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922fa7b),
	.w1(32'hba6385c2),
	.w2(32'hba571f4c),
	.w3(32'hb998ada1),
	.w4(32'hba7f9299),
	.w5(32'hb921f6bb),
	.w6(32'h39a7b8d3),
	.w7(32'h380b61a1),
	.w8(32'hba993952),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba470fee),
	.w1(32'h399fcdcc),
	.w2(32'h3a502257),
	.w3(32'hb9ac44fb),
	.w4(32'hb93fbeb2),
	.w5(32'h3aebaa03),
	.w6(32'hba3cb33c),
	.w7(32'hba8daa46),
	.w8(32'h384566ad),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb039b8a),
	.w1(32'hbadef653),
	.w2(32'hbae9ac8b),
	.w3(32'hbb4b3dbf),
	.w4(32'hbb1418ae),
	.w5(32'h3a44734f),
	.w6(32'hbaf44c5f),
	.w7(32'hbaacdc17),
	.w8(32'hb94d8b16),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a54bb),
	.w1(32'h3ad09f43),
	.w2(32'h3ac7b941),
	.w3(32'hba911053),
	.w4(32'h3aeafc21),
	.w5(32'h3aa0e4de),
	.w6(32'hb9b2dd15),
	.w7(32'h3acd9433),
	.w8(32'h3acddd0d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba052159),
	.w1(32'h393601ec),
	.w2(32'h3b2dba06),
	.w3(32'hbab05c20),
	.w4(32'h3a6ed4aa),
	.w5(32'h3b92fd3d),
	.w6(32'hbb2f19ba),
	.w7(32'hbac947e6),
	.w8(32'h3b08c010),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93fd16d),
	.w1(32'h3a07031f),
	.w2(32'h3b599849),
	.w3(32'hba994e5d),
	.w4(32'hbb1b4432),
	.w5(32'h3ab7567a),
	.w6(32'h3a46fca1),
	.w7(32'hbb897d59),
	.w8(32'h394ee2e6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac653be),
	.w1(32'h38203f83),
	.w2(32'hba3c5e7e),
	.w3(32'hba691c58),
	.w4(32'hbac74549),
	.w5(32'h39fdf089),
	.w6(32'hbb052b1b),
	.w7(32'hba9070bd),
	.w8(32'h3ac35103),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952388f),
	.w1(32'h39d38e9d),
	.w2(32'h39c891c2),
	.w3(32'hb3f7138c),
	.w4(32'h3a1c9433),
	.w5(32'hb89f5c14),
	.w6(32'h39a24dbe),
	.w7(32'hb9773dbd),
	.w8(32'h393248be),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51f0ab),
	.w1(32'hbba45a20),
	.w2(32'h3c01d769),
	.w3(32'hba2168ea),
	.w4(32'hbbc6da27),
	.w5(32'h3b57bb8d),
	.w6(32'h3b0e3c1b),
	.w7(32'hbbca9c55),
	.w8(32'h3b7da481),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba258e3d),
	.w1(32'h3a6efec2),
	.w2(32'h3b82cc90),
	.w3(32'hba443e78),
	.w4(32'h3abf2c16),
	.w5(32'h3b1cc0a6),
	.w6(32'hb9abcb7d),
	.w7(32'h3b3ed528),
	.w8(32'h3b0d5c8e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc9fbd),
	.w1(32'hba8e4e83),
	.w2(32'hbaad12fb),
	.w3(32'h3a14e068),
	.w4(32'hba064cbf),
	.w5(32'h39ee4e11),
	.w6(32'h3861c07c),
	.w7(32'hb99f4e34),
	.w8(32'hb919a3ed),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9503788),
	.w1(32'h3a466bf6),
	.w2(32'h3b65ee11),
	.w3(32'hba1b73e6),
	.w4(32'h3a81dc25),
	.w5(32'h3b0c40c2),
	.w6(32'hb971e941),
	.w7(32'h3b0b6dd3),
	.w8(32'h3b57fcfa),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba533b15),
	.w1(32'h3a3ff73c),
	.w2(32'h3aa65490),
	.w3(32'hba272607),
	.w4(32'h3aa3e54c),
	.w5(32'h3a73e984),
	.w6(32'hb90cc940),
	.w7(32'h3aa1e517),
	.w8(32'h391fe513),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a645b1f),
	.w1(32'hbac1848b),
	.w2(32'hba905950),
	.w3(32'h3a0cacf8),
	.w4(32'hba694716),
	.w5(32'hba74ad51),
	.w6(32'h3990dbb6),
	.w7(32'hb95c1fd9),
	.w8(32'hba1fe652),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb945d0c4),
	.w1(32'hba19b0e7),
	.w2(32'hba3c6a4e),
	.w3(32'hba81fa31),
	.w4(32'hb9a90ab9),
	.w5(32'hba9d7fe6),
	.w6(32'h39c9f494),
	.w7(32'hbacb9ff6),
	.w8(32'hbad70d02),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32a25b),
	.w1(32'h3a059bc7),
	.w2(32'h3a8e2e52),
	.w3(32'hbb01f302),
	.w4(32'h39c0298a),
	.w5(32'h3a8f09b9),
	.w6(32'hbb0600de),
	.w7(32'h3915660c),
	.w8(32'h3a4b8855),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3bc39),
	.w1(32'hbb059af7),
	.w2(32'hbb6f8cac),
	.w3(32'h3af73f82),
	.w4(32'hbb0a8917),
	.w5(32'hbb388edd),
	.w6(32'h3a8e6be3),
	.w7(32'hbb0330a8),
	.w8(32'hbb55ba16),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbf0f5),
	.w1(32'h3a09de0f),
	.w2(32'h3b72c41b),
	.w3(32'hba85e417),
	.w4(32'hbb1d246a),
	.w5(32'hba4f0f5d),
	.w6(32'hba1d3414),
	.w7(32'h3af28fca),
	.w8(32'h3b7d8e2b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a418fee),
	.w1(32'h3b21170a),
	.w2(32'h3b8bb023),
	.w3(32'hbab34778),
	.w4(32'h3ad82f45),
	.w5(32'h3b74937e),
	.w6(32'hbb12c8ff),
	.w7(32'h3a59bf08),
	.w8(32'h3b4f7ba9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cee254),
	.w1(32'h3a37e49e),
	.w2(32'h3bcadec9),
	.w3(32'hb987e557),
	.w4(32'h3afe8f6e),
	.w5(32'h3b39495d),
	.w6(32'hbacac4e9),
	.w7(32'h3ae9c111),
	.w8(32'h3b3fbca2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db706f),
	.w1(32'hba02a756),
	.w2(32'hba73af50),
	.w3(32'h395cb9ee),
	.w4(32'hba5ceb8d),
	.w5(32'hbafa1048),
	.w6(32'hba259989),
	.w7(32'hb9aca1a7),
	.w8(32'hbade9092),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38b8d9),
	.w1(32'hb9a115bc),
	.w2(32'hba39836e),
	.w3(32'hba5cae12),
	.w4(32'h39f6b1c8),
	.w5(32'h3790967e),
	.w6(32'hbabc7edf),
	.w7(32'h3a5a6eba),
	.w8(32'h37d20139),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979d09c),
	.w1(32'hba653140),
	.w2(32'hba07af12),
	.w3(32'h39e04dbe),
	.w4(32'hba49cfb8),
	.w5(32'hbb05f8e9),
	.w6(32'h3a09c974),
	.w7(32'hba855bcd),
	.w8(32'hbab9d70b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba275ddf),
	.w1(32'h3ac31c08),
	.w2(32'hb957c994),
	.w3(32'hba9c1e9e),
	.w4(32'h3a3b69a4),
	.w5(32'hba928dcb),
	.w6(32'hbab9933f),
	.w7(32'hb9c61e1a),
	.w8(32'hb9f07cd6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddcfc4),
	.w1(32'h3b0c3fbf),
	.w2(32'h3b937a57),
	.w3(32'hbaa0fd9d),
	.w4(32'h3a82f2b6),
	.w5(32'h3b159a27),
	.w6(32'hb8ba8b2b),
	.w7(32'h3a1faba9),
	.w8(32'h3aadc3af),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901659b),
	.w1(32'hb9d12a9d),
	.w2(32'h398d6c5e),
	.w3(32'h38a8aedc),
	.w4(32'h3a17f29b),
	.w5(32'h3af230c4),
	.w6(32'h395321d3),
	.w7(32'h3a9cf607),
	.w8(32'h3aee7799),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39432849),
	.w1(32'h39403fe3),
	.w2(32'h39ec1405),
	.w3(32'hba3b369b),
	.w4(32'hb797dad4),
	.w5(32'h3a101f84),
	.w6(32'hba7c3b39),
	.w7(32'h38161514),
	.w8(32'h3aa16760),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09ee7b),
	.w1(32'h3840f3ee),
	.w2(32'hba83f2b0),
	.w3(32'h3b364ac6),
	.w4(32'hba0485c2),
	.w5(32'hbad2631c),
	.w6(32'h3ab998f3),
	.w7(32'hbac4cb8f),
	.w8(32'hbabc202a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4115ab),
	.w1(32'h3a072ea7),
	.w2(32'hb9c6fae5),
	.w3(32'hb92e47fc),
	.w4(32'hba0d3211),
	.w5(32'h3ab3b46b),
	.w6(32'hba580d11),
	.w7(32'hb70999d5),
	.w8(32'h3a2295be),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bf82d),
	.w1(32'hbaa9f40e),
	.w2(32'h3a33389d),
	.w3(32'hbb0dd83d),
	.w4(32'hba756f8e),
	.w5(32'hb9f86986),
	.w6(32'hba3d1089),
	.w7(32'hbab48f11),
	.w8(32'h39d9f2e9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a528f86),
	.w1(32'h3888b208),
	.w2(32'hb9aa9b75),
	.w3(32'hb96a0a5e),
	.w4(32'h39c058fe),
	.w5(32'hb9d36bc7),
	.w6(32'hba3c47bd),
	.w7(32'hba46d8f9),
	.w8(32'hb9ac83f7),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a843f7a),
	.w1(32'h3b973464),
	.w2(32'h3bcf907f),
	.w3(32'h3a19db6e),
	.w4(32'h3aeff7ed),
	.w5(32'h3b249a4d),
	.w6(32'h3acbd209),
	.w7(32'h3bd34f9c),
	.w8(32'h3a13cc9a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b7b4e),
	.w1(32'hba90fb4c),
	.w2(32'hbafa1d1d),
	.w3(32'hba5bf3f7),
	.w4(32'hba578241),
	.w5(32'hbaa8f7e7),
	.w6(32'hbaba2d3f),
	.w7(32'hb92e6fd4),
	.w8(32'hbab5d75c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40ce5a),
	.w1(32'hbaf6ed47),
	.w2(32'hbba9e43f),
	.w3(32'hbb0acbe3),
	.w4(32'hbaefe1ea),
	.w5(32'hba306b9a),
	.w6(32'h3b2b3a0a),
	.w7(32'hb94ce63a),
	.w8(32'hba00427e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule