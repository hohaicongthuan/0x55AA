module layer_10_featuremap_269(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb036ddd),
	.w1(32'hbb98f44e),
	.w2(32'hbb19e3c2),
	.w3(32'hba9d8376),
	.w4(32'hba8197c3),
	.w5(32'h3acd1339),
	.w6(32'hbb91d206),
	.w7(32'hbb2247bd),
	.w8(32'hb993e967),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba541ca5),
	.w1(32'hb95122dd),
	.w2(32'hbb20c4b4),
	.w3(32'hbaac8075),
	.w4(32'h3989348a),
	.w5(32'hbb44c204),
	.w6(32'hbb0c8029),
	.w7(32'hbb2f1fa4),
	.w8(32'h3bec9f66),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21e7bc),
	.w1(32'h37d7198b),
	.w2(32'h3b85da1e),
	.w3(32'h3a7e4291),
	.w4(32'h3bc195e7),
	.w5(32'h3b028e1e),
	.w6(32'h3c639bf6),
	.w7(32'h3bf5a9a4),
	.w8(32'h3ac96dac),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8da807),
	.w1(32'h3b3c4f91),
	.w2(32'h3ba9223b),
	.w3(32'h3b8d5c3d),
	.w4(32'h3b130d6d),
	.w5(32'h395ae091),
	.w6(32'h3b137ee8),
	.w7(32'h3bac8e88),
	.w8(32'h3ba52b12),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bb633),
	.w1(32'h3ade8b74),
	.w2(32'h3b3800c9),
	.w3(32'h3a7af77c),
	.w4(32'h3a0264da),
	.w5(32'h3a25f032),
	.w6(32'h3bb7552a),
	.w7(32'h3ba5311e),
	.w8(32'h3a114073),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab65b60),
	.w1(32'h3a90c91b),
	.w2(32'h3a90d415),
	.w3(32'h3a6a5d3d),
	.w4(32'h3a8848b8),
	.w5(32'h3a6eb428),
	.w6(32'hb94c7cae),
	.w7(32'hba646382),
	.w8(32'hb9a42974),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba928601),
	.w1(32'hbba47804),
	.w2(32'hbbdf5a38),
	.w3(32'h3b007b99),
	.w4(32'hbb0e17c6),
	.w5(32'hbb8a2701),
	.w6(32'h3b15d183),
	.w7(32'hbb22d93c),
	.w8(32'hbb97900f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cd541),
	.w1(32'hbc10eb79),
	.w2(32'hbbbec23b),
	.w3(32'hbb6fcd9d),
	.w4(32'hbbe83454),
	.w5(32'hbbdd784b),
	.w6(32'hbc2c4189),
	.w7(32'hbc0b1710),
	.w8(32'hbb9c95b1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08a01d),
	.w1(32'hbaac9d5f),
	.w2(32'hbaa013b3),
	.w3(32'hbac38dbe),
	.w4(32'hbaeb26c7),
	.w5(32'h3ac4a603),
	.w6(32'hbb2a60f3),
	.w7(32'hbafbeb58),
	.w8(32'h3a412442),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac66371),
	.w1(32'h39ad74fe),
	.w2(32'hbbb8146b),
	.w3(32'h3b37d5e3),
	.w4(32'h3b604502),
	.w5(32'hbb41806f),
	.w6(32'hbb68bfa0),
	.w7(32'hbad83ea7),
	.w8(32'hbb84bc54),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a2076),
	.w1(32'h3b498c2d),
	.w2(32'h3b89fbf4),
	.w3(32'h3b3665ff),
	.w4(32'h3aa5df00),
	.w5(32'hbb37721d),
	.w6(32'h3aaab9da),
	.w7(32'h3a456c94),
	.w8(32'h3b4a10c6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea5c42),
	.w1(32'hbaaa98ae),
	.w2(32'hbba265be),
	.w3(32'h3a55748b),
	.w4(32'h3a8db36b),
	.w5(32'hba90e20a),
	.w6(32'h3c72a335),
	.w7(32'h3b13ee64),
	.w8(32'hbb8e2bba),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb454f5e),
	.w1(32'hba306251),
	.w2(32'hbbb9918e),
	.w3(32'h3b822408),
	.w4(32'h3b36438c),
	.w5(32'hbab4283e),
	.w6(32'h3a057ec4),
	.w7(32'h3bc97f7e),
	.w8(32'hbbd6773d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cae7a6),
	.w1(32'hbb93c8ca),
	.w2(32'hbbac2682),
	.w3(32'h3b60f3db),
	.w4(32'h3b2ffb4c),
	.w5(32'hbb03afcb),
	.w6(32'hbaa46306),
	.w7(32'hba56ecec),
	.w8(32'hbb47b256),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25ccef),
	.w1(32'hbb0803d3),
	.w2(32'hba9c66be),
	.w3(32'hbaa85894),
	.w4(32'h3a489315),
	.w5(32'hbb9f67a6),
	.w6(32'hbb26b4cd),
	.w7(32'hbb060d15),
	.w8(32'hbbb53233),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c02b9),
	.w1(32'hbbd49a84),
	.w2(32'hbc33774b),
	.w3(32'hbbd89a20),
	.w4(32'hb9c08066),
	.w5(32'hbb74a620),
	.w6(32'hbc199944),
	.w7(32'hbbdc93a4),
	.w8(32'hbc180642),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae76605),
	.w1(32'hbb027b2d),
	.w2(32'hbb25eb54),
	.w3(32'hbb5b6719),
	.w4(32'hbaa16994),
	.w5(32'h3a41cee5),
	.w6(32'h39a5df8a),
	.w7(32'hbab83ce9),
	.w8(32'h3b2f2ba3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0059c0),
	.w1(32'hbaf93993),
	.w2(32'hbbf7af08),
	.w3(32'hb935b1a6),
	.w4(32'h3b7c7c7f),
	.w5(32'h3ae641b5),
	.w6(32'hbad00c00),
	.w7(32'h3a6d27aa),
	.w8(32'hbb498a17),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e61ea),
	.w1(32'h3b7d8a11),
	.w2(32'hbafb0c16),
	.w3(32'h3c19c002),
	.w4(32'h3b95a792),
	.w5(32'hbb85b6b4),
	.w6(32'hbbc33630),
	.w7(32'hbaa4fb8f),
	.w8(32'hbb4b424c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5a7f8),
	.w1(32'h3a6b9dbc),
	.w2(32'hba4d5073),
	.w3(32'hbad78db2),
	.w4(32'h36dc7140),
	.w5(32'hbab97881),
	.w6(32'hbac56cf3),
	.w7(32'h3af40db5),
	.w8(32'hbaa20752),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a44c5),
	.w1(32'hba5cb71d),
	.w2(32'hbb3da2e5),
	.w3(32'hbade9cc8),
	.w4(32'hb5510300),
	.w5(32'h3b366b54),
	.w6(32'hbb552bf2),
	.w7(32'h37d892c7),
	.w8(32'h3ab6129e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977491),
	.w1(32'h3b62ab5a),
	.w2(32'h3b335033),
	.w3(32'h3b86df13),
	.w4(32'h3b5e03a4),
	.w5(32'hba798e77),
	.w6(32'hbaebe9be),
	.w7(32'h3b022d9d),
	.w8(32'h3aadca1a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef4188),
	.w1(32'hbc0aa055),
	.w2(32'hbc3a07dd),
	.w3(32'hbb8e6c65),
	.w4(32'h3b4d48da),
	.w5(32'h39fd4cc5),
	.w6(32'hbc030ffb),
	.w7(32'hbb3bd96d),
	.w8(32'hbc1d6d05),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cb629),
	.w1(32'hbaa25498),
	.w2(32'hbb3d284a),
	.w3(32'h3b1f3243),
	.w4(32'h3b37c665),
	.w5(32'hbbc5bc61),
	.w6(32'hbbd82b3e),
	.w7(32'hbafa1d8a),
	.w8(32'hbb9c2889),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72fdd3),
	.w1(32'h3b899329),
	.w2(32'h3ae5386f),
	.w3(32'hbb994648),
	.w4(32'hbb227b64),
	.w5(32'hbada5635),
	.w6(32'hbb50d110),
	.w7(32'hbb86b0e6),
	.w8(32'hbbca37b1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e3555),
	.w1(32'h39baa69a),
	.w2(32'h3a2675f7),
	.w3(32'hbae467c2),
	.w4(32'hba3d126f),
	.w5(32'h3b85bd54),
	.w6(32'hb9de0a54),
	.w7(32'h3a0ca761),
	.w8(32'h3a979a78),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac599ab),
	.w1(32'h3b5ecd9b),
	.w2(32'hb82a123b),
	.w3(32'h3a820a1d),
	.w4(32'h3b3c4884),
	.w5(32'h385ede8a),
	.w6(32'h3b329fe0),
	.w7(32'h3a205178),
	.w8(32'hbb10cf66),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be07447),
	.w1(32'hbb678183),
	.w2(32'hbb61dd36),
	.w3(32'h3b4f46a6),
	.w4(32'hbb53e864),
	.w5(32'hbb91671c),
	.w6(32'h3b83e729),
	.w7(32'hbb4e1958),
	.w8(32'hba99d3fd),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05c0ef),
	.w1(32'hba525574),
	.w2(32'h398323e3),
	.w3(32'hb89978e7),
	.w4(32'hba0e8394),
	.w5(32'hbaa9e354),
	.w6(32'h3a48e658),
	.w7(32'hba27047b),
	.w8(32'h3a979e7b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3761d3),
	.w1(32'h3bd50c02),
	.w2(32'h3bd3f959),
	.w3(32'h3af81581),
	.w4(32'h3b3540c2),
	.w5(32'hbbd109b2),
	.w6(32'h3b2a37df),
	.w7(32'h3b1639b2),
	.w8(32'hbb804c6c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc51d49),
	.w1(32'h3b50aa15),
	.w2(32'hbba87ac9),
	.w3(32'h39a1e822),
	.w4(32'h3a28e555),
	.w5(32'h3a0e921e),
	.w6(32'hbb6a1d27),
	.w7(32'h3a343721),
	.w8(32'h3bcc83fe),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec85c),
	.w1(32'hbbdd577f),
	.w2(32'hbb386cd9),
	.w3(32'hb9f2d9b9),
	.w4(32'h3a7eef3a),
	.w5(32'h3c1e07f9),
	.w6(32'h3c7afca0),
	.w7(32'h3b628bc1),
	.w8(32'h3b002686),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b7bf67),
	.w1(32'h3c27dd93),
	.w2(32'hbab7fd99),
	.w3(32'h3be09be9),
	.w4(32'h3b4b180a),
	.w5(32'hbb9f747c),
	.w6(32'hba57fb2a),
	.w7(32'h3ba3a191),
	.w8(32'hbb355ad3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99dc47),
	.w1(32'hbaeaca96),
	.w2(32'hbb87e103),
	.w3(32'hbba30391),
	.w4(32'h37379176),
	.w5(32'hbabc23f3),
	.w6(32'hbb6545da),
	.w7(32'hba7793f5),
	.w8(32'hbb688086),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a046f5a),
	.w1(32'hba219093),
	.w2(32'hb98ca6db),
	.w3(32'h390c0585),
	.w4(32'hbb18267c),
	.w5(32'h39e83978),
	.w6(32'h3a2ca567),
	.w7(32'hbae3f728),
	.w8(32'hbb7dba16),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35323c),
	.w1(32'hbad7f3d6),
	.w2(32'hbb08096e),
	.w3(32'hbabbc8cd),
	.w4(32'hba039476),
	.w5(32'hbaf0f25b),
	.w6(32'hbb989683),
	.w7(32'hba679716),
	.w8(32'h3b766636),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e444f),
	.w1(32'hba7f980b),
	.w2(32'hbbc7091c),
	.w3(32'hbb9e4c32),
	.w4(32'h3974a257),
	.w5(32'h3b12098e),
	.w6(32'hbbdf74e6),
	.w7(32'h3a59b542),
	.w8(32'hba9326fe),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb1472),
	.w1(32'h3c224da3),
	.w2(32'h3b9a20fb),
	.w3(32'hba8e3aec),
	.w4(32'h3ba00285),
	.w5(32'hbb0fd88d),
	.w6(32'hbbb49965),
	.w7(32'hbb30e95f),
	.w8(32'hbbe1d274),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33f223),
	.w1(32'h3b872e2d),
	.w2(32'h3a1066f5),
	.w3(32'h3979ad82),
	.w4(32'hbbd2fa74),
	.w5(32'hbb5732a3),
	.w6(32'h3ba1ec20),
	.w7(32'hbb6d595b),
	.w8(32'hbbfa1ea3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f530a),
	.w1(32'hbb256dac),
	.w2(32'h3a33554c),
	.w3(32'h3c013b05),
	.w4(32'h3c1256c3),
	.w5(32'h386893fd),
	.w6(32'hbbecab0a),
	.w7(32'h3b3d98c2),
	.w8(32'hbb2a0d65),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f19f7),
	.w1(32'hb8e38d44),
	.w2(32'hbb309f90),
	.w3(32'hbb21880a),
	.w4(32'hbb16fd1e),
	.w5(32'h3a971484),
	.w6(32'hbaf180a7),
	.w7(32'hbaf41342),
	.w8(32'h3aab7618),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80c1dc),
	.w1(32'hba98933e),
	.w2(32'h39054ab1),
	.w3(32'h3a179f32),
	.w4(32'h3af2ce9f),
	.w5(32'hba9c8c3f),
	.w6(32'h3b296f53),
	.w7(32'h3b8bc86c),
	.w8(32'hba9f58c0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedefa0),
	.w1(32'hba92ef35),
	.w2(32'hba688e7d),
	.w3(32'h3b0005f6),
	.w4(32'h3b909466),
	.w5(32'hbb5001a9),
	.w6(32'hbb0439c8),
	.w7(32'hbb288b5b),
	.w8(32'hbab8eb28),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38d281),
	.w1(32'h3a8d1636),
	.w2(32'hbc4192aa),
	.w3(32'hbc1e8d35),
	.w4(32'hbb78917d),
	.w5(32'h3c0758cb),
	.w6(32'h3b8750bd),
	.w7(32'hbbfe0cdc),
	.w8(32'hbbd3f16d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c9d57),
	.w1(32'hb973f522),
	.w2(32'hbb71ffa9),
	.w3(32'h3c7851f4),
	.w4(32'h3c799e4a),
	.w5(32'hbada891a),
	.w6(32'hbb1ef359),
	.w7(32'h397685c3),
	.w8(32'hbbe7a77b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc26bcb),
	.w1(32'hbb5e5fd9),
	.w2(32'hbbd77964),
	.w3(32'h3a0c2bd4),
	.w4(32'h3aeea8fd),
	.w5(32'h3b021569),
	.w6(32'hbbd94e3e),
	.w7(32'hbbbf4549),
	.w8(32'hbb97ad36),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad19988),
	.w1(32'hbb3d80f0),
	.w2(32'hbb4f8936),
	.w3(32'h3b4ab21a),
	.w4(32'h3b420118),
	.w5(32'hbb35101e),
	.w6(32'hbb0036cf),
	.w7(32'hbbe96734),
	.w8(32'hbbe65862),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f766c3),
	.w1(32'h3a8459eb),
	.w2(32'hbb41ce94),
	.w3(32'h3b28b88e),
	.w4(32'h399ec485),
	.w5(32'hbae33447),
	.w6(32'hbb508eb7),
	.w7(32'h39decc51),
	.w8(32'hbbe02530),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae07d52),
	.w1(32'h3a9a179a),
	.w2(32'hba4726c8),
	.w3(32'h3b6e0a59),
	.w4(32'h3b3f744f),
	.w5(32'h3ab979d5),
	.w6(32'h3b0bbd37),
	.w7(32'h3b488a46),
	.w8(32'hb99ef863),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d6ff8),
	.w1(32'h39c6daf3),
	.w2(32'h39b0220d),
	.w3(32'h3a28c14c),
	.w4(32'hb7a82c2d),
	.w5(32'hbb92789f),
	.w6(32'hbb3451f6),
	.w7(32'hbaab252d),
	.w8(32'hba9d0dd8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf865),
	.w1(32'hbbb57d16),
	.w2(32'hba6aa956),
	.w3(32'h3b93908a),
	.w4(32'hbb26d52d),
	.w5(32'h3b1ed1d6),
	.w6(32'hbbda89c4),
	.w7(32'hb99d663f),
	.w8(32'h3aefd9fb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9b278),
	.w1(32'h3b8d4c2c),
	.w2(32'hbb78f392),
	.w3(32'h3a608263),
	.w4(32'h3a220f3b),
	.w5(32'h3ab73944),
	.w6(32'hbae15dee),
	.w7(32'hb9388ba3),
	.w8(32'hba8885cc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e86f8),
	.w1(32'hbb39f800),
	.w2(32'hba68797a),
	.w3(32'h3aae7b2b),
	.w4(32'h3b1a88e0),
	.w5(32'hbb147f93),
	.w6(32'hba0438c6),
	.w7(32'hbb497a71),
	.w8(32'hbbd88707),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d675b),
	.w1(32'hbba5f5e8),
	.w2(32'hbc12e75d),
	.w3(32'h3b31f701),
	.w4(32'h3b7b91a3),
	.w5(32'hbc1f5a9f),
	.w6(32'hbb110181),
	.w7(32'hbb3c858f),
	.w8(32'hbc45deee),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d17ca3),
	.w1(32'h3a81b6ce),
	.w2(32'h392cc11e),
	.w3(32'hbb617b60),
	.w4(32'hbb208fe8),
	.w5(32'hbada8a3d),
	.w6(32'hbad162d9),
	.w7(32'hba154714),
	.w8(32'hba5c65d1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3b13b),
	.w1(32'hba681984),
	.w2(32'hba9e5bdc),
	.w3(32'h38c108e0),
	.w4(32'h3a32d9fa),
	.w5(32'hbb1a1748),
	.w6(32'h3b32e9aa),
	.w7(32'h39156cf6),
	.w8(32'hbb3a2291),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34efca),
	.w1(32'h3abdcad1),
	.w2(32'hba795a3e),
	.w3(32'hba9fdefb),
	.w4(32'hbadb28fa),
	.w5(32'hba83a095),
	.w6(32'hbb241b7d),
	.w7(32'h3a0c60fd),
	.w8(32'hb9fa8aa7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399da04e),
	.w1(32'hbb420134),
	.w2(32'hbb4ce993),
	.w3(32'h3b12f7cc),
	.w4(32'h3b38d94d),
	.w5(32'h399c2946),
	.w6(32'h3a9b5b24),
	.w7(32'hba4a3170),
	.w8(32'hbaa0e96c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a497180),
	.w1(32'h3a5ea890),
	.w2(32'h3a9ba851),
	.w3(32'hba9fe792),
	.w4(32'h38342675),
	.w5(32'h3ae05001),
	.w6(32'hba6adb85),
	.w7(32'h38ffa397),
	.w8(32'h3ba85a97),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6fed2),
	.w1(32'h3b751335),
	.w2(32'h3a970d24),
	.w3(32'h39de1ab1),
	.w4(32'hbb236fce),
	.w5(32'hb9bfd21d),
	.w6(32'hb9a61c08),
	.w7(32'hbb700955),
	.w8(32'hbb41a20e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4bcfa),
	.w1(32'hbb470929),
	.w2(32'hbb18b0a5),
	.w3(32'hbb1310c3),
	.w4(32'h39293d6d),
	.w5(32'hba3f624d),
	.w6(32'hbb0ab056),
	.w7(32'h3a6cbd1e),
	.w8(32'hbb92e56c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba890ed),
	.w1(32'hbbbf8124),
	.w2(32'hbb8fa7ce),
	.w3(32'hbba5354a),
	.w4(32'hb8cfda6d),
	.w5(32'hb9a92867),
	.w6(32'h39177b99),
	.w7(32'h3917209c),
	.w8(32'hbb65eebc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a55ed),
	.w1(32'h3a9b487f),
	.w2(32'h3a5de5a0),
	.w3(32'hbac4f2ea),
	.w4(32'hba3229c7),
	.w5(32'hbaeecda7),
	.w6(32'h3ac5648a),
	.w7(32'h392c8ca4),
	.w8(32'hbb56a9c2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ae5f3),
	.w1(32'hba25dea2),
	.w2(32'hbae34f5a),
	.w3(32'h39f59c28),
	.w4(32'h3a89daaf),
	.w5(32'h3aa76f1a),
	.w6(32'hbb20f367),
	.w7(32'hba9e02c6),
	.w8(32'hbb6b75b2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a514fa8),
	.w1(32'hbadcffdc),
	.w2(32'h3b4db86c),
	.w3(32'h3b1e8435),
	.w4(32'h3afd7ca5),
	.w5(32'hbaa85748),
	.w6(32'hbb507e06),
	.w7(32'h3a8cf947),
	.w8(32'hbb3e7c2c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816d51),
	.w1(32'h3b90da38),
	.w2(32'h3ac52484),
	.w3(32'hba9d11d3),
	.w4(32'hba0e9231),
	.w5(32'h3aba30fe),
	.w6(32'h3bc48d93),
	.w7(32'hbb1f2304),
	.w8(32'h39e65cee),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe42896),
	.w1(32'hbbb011bc),
	.w2(32'hbbe13628),
	.w3(32'h3b951356),
	.w4(32'h3ad1b7c9),
	.w5(32'hbb0586b2),
	.w6(32'hbaf8e324),
	.w7(32'hbb959336),
	.w8(32'hbbfc0fbb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3bc76),
	.w1(32'h3baf2a06),
	.w2(32'h3a6588e8),
	.w3(32'h3b1a2f6b),
	.w4(32'hba950607),
	.w5(32'hbc07b0ac),
	.w6(32'h3985ab42),
	.w7(32'hb80306e6),
	.w8(32'hbc6716c9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc7c28),
	.w1(32'hba5bfd93),
	.w2(32'hb9d7bca7),
	.w3(32'hbb82349f),
	.w4(32'h3b6c2368),
	.w5(32'hbacafaf2),
	.w6(32'hbc09bc46),
	.w7(32'h3b7070ff),
	.w8(32'hbaf49efc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8be7da),
	.w1(32'h3c2c2e97),
	.w2(32'h3a672f4f),
	.w3(32'h3b17ef17),
	.w4(32'h3c0e0bab),
	.w5(32'h3b91c637),
	.w6(32'hbb3c909a),
	.w7(32'h3aa10375),
	.w8(32'hbba1ca6d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ce856),
	.w1(32'h3baa583f),
	.w2(32'hb9c8dd12),
	.w3(32'h3b921229),
	.w4(32'h3b2f9655),
	.w5(32'hbb2ab1be),
	.w6(32'hbb273ca6),
	.w7(32'hba2ef8bd),
	.w8(32'hbb17d2ab),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3c74e),
	.w1(32'h3a9f2173),
	.w2(32'h39a2151e),
	.w3(32'hbb242989),
	.w4(32'hbb031780),
	.w5(32'hbb9f6498),
	.w6(32'h3afbeac6),
	.w7(32'h3b2bba36),
	.w8(32'h3a5ea5a1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad34b3f),
	.w1(32'hb93d8b0a),
	.w2(32'hbb25a308),
	.w3(32'hbbd0cbd3),
	.w4(32'hbb39f0b0),
	.w5(32'hbb9d24cf),
	.w6(32'h3b2b5311),
	.w7(32'hba849006),
	.w8(32'hbba0997f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd7bec),
	.w1(32'hbb35f8e7),
	.w2(32'h3a8af74a),
	.w3(32'hba578b5d),
	.w4(32'h3b44a2b2),
	.w5(32'hbaf64cfb),
	.w6(32'hbb946c99),
	.w7(32'h3a87f77e),
	.w8(32'hba81cab8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68590b),
	.w1(32'hbae7fcb2),
	.w2(32'h3a63de3a),
	.w3(32'hbb603502),
	.w4(32'hbb92cabd),
	.w5(32'hbb604d39),
	.w6(32'hb9022795),
	.w7(32'hbadb5783),
	.w8(32'hb89f15bc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41bc8b),
	.w1(32'hba7fa5ff),
	.w2(32'hba854d3b),
	.w3(32'h3a1bf2eb),
	.w4(32'hb92b1780),
	.w5(32'hbb34ac9a),
	.w6(32'hba9d843b),
	.w7(32'h3b0d684b),
	.w8(32'hbb755c3b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c78e),
	.w1(32'hbaccd853),
	.w2(32'hbb0b9be0),
	.w3(32'h385c96db),
	.w4(32'hba84cb41),
	.w5(32'hbac878c1),
	.w6(32'hbb919193),
	.w7(32'hbb519778),
	.w8(32'hbb80c251),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72c30d),
	.w1(32'hbac53e42),
	.w2(32'hbbe34ea2),
	.w3(32'h3b8c7541),
	.w4(32'h3bbacf14),
	.w5(32'hbbc799f1),
	.w6(32'hba94114b),
	.w7(32'h3a92310a),
	.w8(32'hbbdacd09),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c9a06),
	.w1(32'hbba2cf71),
	.w2(32'hbbd7ffa3),
	.w3(32'hba989215),
	.w4(32'hbb3df6c7),
	.w5(32'hbb16efc2),
	.w6(32'hbc101e3d),
	.w7(32'hbb99b3b9),
	.w8(32'hbb917936),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a44bd),
	.w1(32'hbb39ac16),
	.w2(32'hbb840483),
	.w3(32'h3b15e4a4),
	.w4(32'hb9a9f4f7),
	.w5(32'hbb4490f8),
	.w6(32'h39ab6d99),
	.w7(32'hb99153ac),
	.w8(32'hbbd1a488),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba987e0d),
	.w1(32'h392701f3),
	.w2(32'h3b081e45),
	.w3(32'hb9f49023),
	.w4(32'h3b6c8513),
	.w5(32'hbb4cfb40),
	.w6(32'hbc162d95),
	.w7(32'h3b432afd),
	.w8(32'hbb9cc35c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8356de),
	.w1(32'hbb1b7256),
	.w2(32'hbba46529),
	.w3(32'h3a879a7c),
	.w4(32'h3ac02c77),
	.w5(32'hbb56fea2),
	.w6(32'hbb71ac41),
	.w7(32'hbaf7310d),
	.w8(32'hbbaaa821),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1911da),
	.w1(32'hbb24ceb6),
	.w2(32'h3b2309c4),
	.w3(32'hbab1f86a),
	.w4(32'h39bc32f0),
	.w5(32'hbb4be865),
	.w6(32'hbbb82282),
	.w7(32'h3a50a46d),
	.w8(32'h3a23c39b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d37a3),
	.w1(32'h3b94fd6a),
	.w2(32'h3bbd01c1),
	.w3(32'hbafbbb1f),
	.w4(32'hba9cfe3f),
	.w5(32'hbaa3ec7f),
	.w6(32'hbab51028),
	.w7(32'h3bc38c53),
	.w8(32'hbb29b496),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4b903),
	.w1(32'hb9bce249),
	.w2(32'h3a291341),
	.w3(32'h39d0791b),
	.w4(32'h39f72e7e),
	.w5(32'h3ae3d912),
	.w6(32'hbb7bd2d4),
	.w7(32'hbb0fd1b8),
	.w8(32'h3a9fe114),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4f07b),
	.w1(32'hbaae0eb5),
	.w2(32'hbadcda6c),
	.w3(32'h3b9966a1),
	.w4(32'h3ba9e4a2),
	.w5(32'hba15bf12),
	.w6(32'h3a4d677b),
	.w7(32'hbb09f70b),
	.w8(32'hbacc22cb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72eec8),
	.w1(32'h3a45c8f7),
	.w2(32'hbb8a0632),
	.w3(32'hbb2f16cd),
	.w4(32'h3c1158ad),
	.w5(32'h39e00986),
	.w6(32'h3b8e4fda),
	.w7(32'hbb4111cc),
	.w8(32'hba55c568),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68c111),
	.w1(32'h3b081d29),
	.w2(32'h3ad4832f),
	.w3(32'h3ab4ebd4),
	.w4(32'h392a6fbe),
	.w5(32'hba7ef205),
	.w6(32'h3b5adff1),
	.w7(32'h3a4f1217),
	.w8(32'hbb23ee0a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2be8),
	.w1(32'hbaf83092),
	.w2(32'hbab43fd2),
	.w3(32'hba18ef6a),
	.w4(32'hba3c8042),
	.w5(32'hbb560c38),
	.w6(32'hbb9d788f),
	.w7(32'hbb44b714),
	.w8(32'hbb64cf40),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ac0aa),
	.w1(32'h3951c8cb),
	.w2(32'h39fa4bbe),
	.w3(32'hbb3e11d7),
	.w4(32'hbad39537),
	.w5(32'hbaad38bd),
	.w6(32'hbc03c1a7),
	.w7(32'hbb8be45f),
	.w8(32'hbb9d0048),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e3dea),
	.w1(32'h3b4f596b),
	.w2(32'h3b707d99),
	.w3(32'h3b5af216),
	.w4(32'h3a354155),
	.w5(32'h3b867240),
	.w6(32'h3aaf2f35),
	.w7(32'h391c6810),
	.w8(32'hbb0136b6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee699e),
	.w1(32'hbb85a978),
	.w2(32'h3adf5069),
	.w3(32'h3abb96aa),
	.w4(32'hba886a67),
	.w5(32'h3c433ab6),
	.w6(32'hbba7d8ff),
	.w7(32'h3a4b1a25),
	.w8(32'hbbbfa577),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab11e40),
	.w1(32'hb9231153),
	.w2(32'hbb0c365a),
	.w3(32'h3b343ef1),
	.w4(32'h3b31faae),
	.w5(32'h3aea6800),
	.w6(32'h3c9a39bb),
	.w7(32'hb9404675),
	.w8(32'hbb22a83e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb705f08),
	.w1(32'hbb02ec9b),
	.w2(32'hbc1b336d),
	.w3(32'h3b941de1),
	.w4(32'h3b7c7d2c),
	.w5(32'hba626aef),
	.w6(32'hbbcd311c),
	.w7(32'hbbdc2ce3),
	.w8(32'hbbf8cc84),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11fd7a),
	.w1(32'hbb294a34),
	.w2(32'hbb9e68c7),
	.w3(32'hba84b9bd),
	.w4(32'hba2ac395),
	.w5(32'h3b7be23b),
	.w6(32'hbb582c87),
	.w7(32'hbb52185d),
	.w8(32'h3c0f4e81),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d030f),
	.w1(32'hbb6fbce2),
	.w2(32'hbb8f65a0),
	.w3(32'hb908d1ba),
	.w4(32'h3ae7b1aa),
	.w5(32'hbc0efc06),
	.w6(32'h3cb8dd73),
	.w7(32'h3b4164d9),
	.w8(32'hbbfae1e0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f7dc2),
	.w1(32'hbba1062c),
	.w2(32'h3a8c96b5),
	.w3(32'h393709f3),
	.w4(32'hba8dd2e7),
	.w5(32'h3b544079),
	.w6(32'hbc3456c4),
	.w7(32'hbb406808),
	.w8(32'hbb578882),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48a20b),
	.w1(32'h3a9208a8),
	.w2(32'hbc0075a3),
	.w3(32'h3b27a243),
	.w4(32'h3b96c066),
	.w5(32'hbb59e867),
	.w6(32'hbbf431fb),
	.w7(32'hbaa66a34),
	.w8(32'hbbf47183),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e7654),
	.w1(32'hb9d6d43a),
	.w2(32'hbb876cdd),
	.w3(32'h3a7560d5),
	.w4(32'h39d869c2),
	.w5(32'hbb297f6b),
	.w6(32'hbb3d0a5d),
	.w7(32'hbb392f2a),
	.w8(32'hbb9fc5af),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03d81f),
	.w1(32'hbbd2260b),
	.w2(32'hbbe0625d),
	.w3(32'hbc0dd220),
	.w4(32'hbb9d7bbc),
	.w5(32'h3be7957a),
	.w6(32'hbc49b4be),
	.w7(32'h3a29cdec),
	.w8(32'h3b7eaa4d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49e697),
	.w1(32'h3bf381ff),
	.w2(32'h3bee7188),
	.w3(32'hba8e5337),
	.w4(32'h3bc64a93),
	.w5(32'h3b32d47a),
	.w6(32'hbb4d728a),
	.w7(32'h3b1e669c),
	.w8(32'hbb5a7718),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d1b1e),
	.w1(32'hbb93b591),
	.w2(32'hbbd01843),
	.w3(32'hbaec5059),
	.w4(32'h3a14d6bd),
	.w5(32'hbba31306),
	.w6(32'hbb8a28ae),
	.w7(32'hbb737452),
	.w8(32'hbbe6ac15),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb6ba3),
	.w1(32'hbb78c957),
	.w2(32'hbbc10abf),
	.w3(32'hbaca08d9),
	.w4(32'h3a8095f6),
	.w5(32'h3bb358b8),
	.w6(32'hbba608fd),
	.w7(32'h3aa9ef59),
	.w8(32'h3b18dbd6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a472b41),
	.w1(32'hbab6d001),
	.w2(32'h3a729924),
	.w3(32'hba925fde),
	.w4(32'h3adbc5de),
	.w5(32'hbb067cfc),
	.w6(32'hba347680),
	.w7(32'h3a4c6609),
	.w8(32'hb8b1944d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82e886),
	.w1(32'hbc34a0ec),
	.w2(32'hbbbd3e67),
	.w3(32'hbc00c15e),
	.w4(32'hbb183e63),
	.w5(32'hbb7b027a),
	.w6(32'hbbb9d536),
	.w7(32'h3ad23ec8),
	.w8(32'hbb8e2bb6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1a0e8),
	.w1(32'hba301fca),
	.w2(32'hbb21945c),
	.w3(32'hbb49f660),
	.w4(32'hbb867733),
	.w5(32'hbb8ac8dd),
	.w6(32'hba8f3f3b),
	.w7(32'hba7451e6),
	.w8(32'hbb87bbe8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e3c4c),
	.w1(32'hbaf1bb21),
	.w2(32'hbbb3577e),
	.w3(32'hbb1a6a17),
	.w4(32'hba952ee0),
	.w5(32'hb9c93616),
	.w6(32'hba927c0a),
	.w7(32'hbb703276),
	.w8(32'h39ec131a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb184a4c),
	.w1(32'h3a9f170e),
	.w2(32'hbb2bacc4),
	.w3(32'hb7a7e867),
	.w4(32'h3a63282f),
	.w5(32'h39a52ff5),
	.w6(32'h3ae6e1fa),
	.w7(32'hba3326ca),
	.w8(32'hbb0cfde7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891666),
	.w1(32'hbac889b7),
	.w2(32'hbbf9566a),
	.w3(32'h3af678e2),
	.w4(32'h3b0d2259),
	.w5(32'h3a258af3),
	.w6(32'hbaa6428f),
	.w7(32'hbad9a090),
	.w8(32'hbb4e7653),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b655674),
	.w1(32'h3b86ce4d),
	.w2(32'h3b311b1c),
	.w3(32'h3b7a7aee),
	.w4(32'h3be8dec4),
	.w5(32'hbb4627db),
	.w6(32'h3b86fa9d),
	.w7(32'h3bd17e36),
	.w8(32'hbb46618f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2b6b2),
	.w1(32'h3b2a4f42),
	.w2(32'hbb312424),
	.w3(32'hba1b6c31),
	.w4(32'h384d6fe1),
	.w5(32'hbabea05d),
	.w6(32'h388007d4),
	.w7(32'hbb26b899),
	.w8(32'hbb63ce93),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a21e3),
	.w1(32'h3b24f2c6),
	.w2(32'h3a41a076),
	.w3(32'h3b12027e),
	.w4(32'h3b36b66a),
	.w5(32'hba8bfec4),
	.w6(32'h39ac48d2),
	.w7(32'h3aedad48),
	.w8(32'hbb72c7b7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ae15e),
	.w1(32'h3b40291e),
	.w2(32'h3bc6d220),
	.w3(32'hba8d9b33),
	.w4(32'h3a80f9bf),
	.w5(32'h39bfa15b),
	.w6(32'hbbd6e2a3),
	.w7(32'h3a65f512),
	.w8(32'hba576d3a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab27e5),
	.w1(32'hbb97e152),
	.w2(32'hbbd89734),
	.w3(32'hbb531e44),
	.w4(32'hbb4a76f3),
	.w5(32'hbbe665ca),
	.w6(32'hbbc868ca),
	.w7(32'hbbc1d381),
	.w8(32'hbc101276),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb5a73),
	.w1(32'hba034b61),
	.w2(32'hbb3e1ece),
	.w3(32'hbb49979c),
	.w4(32'hbb6bc1af),
	.w5(32'hb9cafc36),
	.w6(32'hbb84410a),
	.w7(32'hbb997a21),
	.w8(32'hbb2c29fc),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa07f),
	.w1(32'hba611cc5),
	.w2(32'hba79b155),
	.w3(32'h3a09abb8),
	.w4(32'hb9f4c7d0),
	.w5(32'h3b2efd7a),
	.w6(32'hb9fa7e73),
	.w7(32'h3a144af8),
	.w8(32'h3aa55463),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cf647),
	.w1(32'h3814c523),
	.w2(32'hba8dc11c),
	.w3(32'h3b5f713d),
	.w4(32'h3b364e6f),
	.w5(32'hba1dfc9b),
	.w6(32'h39c6dd15),
	.w7(32'hba4f4d0e),
	.w8(32'hbb1500b5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4497d9),
	.w1(32'hbb598922),
	.w2(32'h38c77df1),
	.w3(32'hbabe1a20),
	.w4(32'hbb111e6c),
	.w5(32'h3a44272b),
	.w6(32'h3ae591e6),
	.w7(32'h3a520199),
	.w8(32'h3a8d67ab),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b068880),
	.w1(32'h3aa14e60),
	.w2(32'h39f4b790),
	.w3(32'hba045b04),
	.w4(32'hbae4d814),
	.w5(32'hb9832e70),
	.w6(32'hb94390b1),
	.w7(32'hbad4f088),
	.w8(32'hbb4fafae),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e9e5),
	.w1(32'hbb6ede1e),
	.w2(32'hbb9e3597),
	.w3(32'hbb01bf65),
	.w4(32'h394fa547),
	.w5(32'hbb38bc75),
	.w6(32'hbbcbd948),
	.w7(32'hbb99f073),
	.w8(32'hbb4a19c2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e052a),
	.w1(32'hb94c96e7),
	.w2(32'h39c488db),
	.w3(32'hba9b4638),
	.w4(32'hbac050fc),
	.w5(32'hbb380446),
	.w6(32'hbae1128e),
	.w7(32'hb90e02ca),
	.w8(32'hb9ba8d22),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb010408),
	.w1(32'h3915fb30),
	.w2(32'h3a7c401f),
	.w3(32'h399da2cd),
	.w4(32'hbacf779d),
	.w5(32'hb992bb4d),
	.w6(32'hb90fe7c4),
	.w7(32'h3ab85acc),
	.w8(32'hbb882a88),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d8225),
	.w1(32'hba5b194a),
	.w2(32'hba9b8986),
	.w3(32'hbae7f619),
	.w4(32'h38bdb614),
	.w5(32'hbba0d339),
	.w6(32'hbb9a5ac6),
	.w7(32'hbb0a81ce),
	.w8(32'hbbdc6705),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dae3b3),
	.w1(32'h3b72972d),
	.w2(32'h3aae1179),
	.w3(32'hba19b5af),
	.w4(32'hba627f89),
	.w5(32'h3a9b2711),
	.w6(32'h3b55432c),
	.w7(32'h3a356b1b),
	.w8(32'hba4ade96),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe3418),
	.w1(32'hb8d0e31d),
	.w2(32'h39e5654f),
	.w3(32'h3b452b6f),
	.w4(32'h39ca0c3f),
	.w5(32'hbb310a6f),
	.w6(32'h3a78b432),
	.w7(32'h3b0f034d),
	.w8(32'hbb64951b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8327c),
	.w1(32'hbbad513b),
	.w2(32'hbb2e8e01),
	.w3(32'hba84a11f),
	.w4(32'hb910687d),
	.w5(32'hb80941ed),
	.w6(32'hba7f73eb),
	.w7(32'hba459fd7),
	.w8(32'hb99bf316),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb796698),
	.w1(32'hbb0294b1),
	.w2(32'hbae2985d),
	.w3(32'h3b32871a),
	.w4(32'h3b124178),
	.w5(32'hb9d5aef7),
	.w6(32'h3a8360e2),
	.w7(32'hb9ba0f8c),
	.w8(32'hba0f9412),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948451),
	.w1(32'h3b4dff59),
	.w2(32'h3b10e3a6),
	.w3(32'h3b7784c6),
	.w4(32'h3af3c6ae),
	.w5(32'hbb139f0f),
	.w6(32'hb92d03e9),
	.w7(32'h39bd9807),
	.w8(32'hbb83bcbc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af4735),
	.w1(32'hbb324075),
	.w2(32'hbb632557),
	.w3(32'hbae68323),
	.w4(32'h3ac44384),
	.w5(32'hbbf172d8),
	.w6(32'hbb66ae55),
	.w7(32'h3addc96a),
	.w8(32'hbc2b7636),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d220b),
	.w1(32'hbb90a561),
	.w2(32'hbaeb7b3b),
	.w3(32'hba827e94),
	.w4(32'hbb4913b1),
	.w5(32'h397bc267),
	.w6(32'hbb558d15),
	.w7(32'hbb623f83),
	.w8(32'hbb868cbf),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dce48c),
	.w1(32'h39c2c32d),
	.w2(32'h3a3d13b9),
	.w3(32'hbaab6397),
	.w4(32'hbaea13f1),
	.w5(32'hbafad66a),
	.w6(32'hbbcdfb5c),
	.w7(32'hbb7f66a2),
	.w8(32'hbb955b84),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812f5d),
	.w1(32'hbb61bcd5),
	.w2(32'hbb1a9f7b),
	.w3(32'h39e60a82),
	.w4(32'hb90cb8e7),
	.w5(32'hbb8675f5),
	.w6(32'hbb15123c),
	.w7(32'hbb1e2a6d),
	.w8(32'hbb970700),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7d114),
	.w1(32'hbba20867),
	.w2(32'h3b2a155c),
	.w3(32'hbb480454),
	.w4(32'h3bff20bf),
	.w5(32'h3a3e48b0),
	.w6(32'hbbb5dbd6),
	.w7(32'h3bf149b9),
	.w8(32'hbb27fa6b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a299c),
	.w1(32'hbb588001),
	.w2(32'hbb20866e),
	.w3(32'h3b04bcae),
	.w4(32'h3b9b31f4),
	.w5(32'hb9fa4aa4),
	.w6(32'hba79ddbb),
	.w7(32'h3b07784e),
	.w8(32'hbbbb9108),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2323a),
	.w1(32'hbb8a1da3),
	.w2(32'hbbeb7fd7),
	.w3(32'h3b7cff90),
	.w4(32'h3b323ddb),
	.w5(32'hbb709e18),
	.w6(32'hbb2f2d0f),
	.w7(32'hbb42dd2f),
	.w8(32'hbbe60b94),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77356f),
	.w1(32'hbb9e594f),
	.w2(32'hbbafd547),
	.w3(32'hbb90c069),
	.w4(32'h39de9564),
	.w5(32'hba2995c7),
	.w6(32'hbbef3d3e),
	.w7(32'hbb91c739),
	.w8(32'hbae401cd),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb644),
	.w1(32'hba2bca8d),
	.w2(32'hba8ff6fa),
	.w3(32'h3a17b7c5),
	.w4(32'h3b9269a0),
	.w5(32'h3b241101),
	.w6(32'hbab3c7ed),
	.w7(32'h3b4d7f83),
	.w8(32'hbb25ca73),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb923172),
	.w1(32'hbb276e9d),
	.w2(32'hbb2de8cc),
	.w3(32'h3b4b3a48),
	.w4(32'h3ba01b14),
	.w5(32'h3907bc6f),
	.w6(32'hbb1ce9ba),
	.w7(32'h3b0c5c3c),
	.w8(32'hbb9637e7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdd4ad),
	.w1(32'hba8d400f),
	.w2(32'h3b04f2ab),
	.w3(32'hba9cd937),
	.w4(32'h3b004210),
	.w5(32'h3af62c94),
	.w6(32'hbbafb390),
	.w7(32'h3a7299d1),
	.w8(32'hbb6167a1),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af35531),
	.w1(32'h3b0a5c00),
	.w2(32'hba78c5de),
	.w3(32'h3a1550ac),
	.w4(32'hbaab05c1),
	.w5(32'hbbbeee08),
	.w6(32'hbb952fba),
	.w7(32'hbba40bfb),
	.w8(32'hbba443d2),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ea999),
	.w1(32'h39efa670),
	.w2(32'h3a4e4b64),
	.w3(32'hbb105410),
	.w4(32'h3abe9b50),
	.w5(32'hbb2e44b2),
	.w6(32'hba37d093),
	.w7(32'h3a916457),
	.w8(32'hbb503758),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd456c4),
	.w1(32'h3aecf5ca),
	.w2(32'h3bfc2616),
	.w3(32'h39cd8f7e),
	.w4(32'h3a8a9905),
	.w5(32'hbb1f8671),
	.w6(32'h3a81ab46),
	.w7(32'h39f95de8),
	.w8(32'hbb8f203a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0695e8),
	.w1(32'h3b0d1194),
	.w2(32'h3a7eb957),
	.w3(32'h3b1318eb),
	.w4(32'h3b455cf8),
	.w5(32'hbb111323),
	.w6(32'hb9a6998f),
	.w7(32'hba061b21),
	.w8(32'hbb3c88d6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb090511),
	.w1(32'hbb6e329b),
	.w2(32'hba376fa5),
	.w3(32'hbba887ce),
	.w4(32'hbb07f77d),
	.w5(32'hb9e01b81),
	.w6(32'hbb4b1723),
	.w7(32'h3a1cd586),
	.w8(32'hbae3f175),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bddb7),
	.w1(32'h3a4c4814),
	.w2(32'h3b41de78),
	.w3(32'h3a1397e1),
	.w4(32'h3b086e73),
	.w5(32'hbb1f2963),
	.w6(32'h3a5b58fb),
	.w7(32'h3a7fdfb8),
	.w8(32'hbaa4bbad),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb275bf1),
	.w1(32'hbac441a3),
	.w2(32'hbb04b785),
	.w3(32'hbb426b41),
	.w4(32'hbb14acc9),
	.w5(32'hbabd5bf5),
	.w6(32'hbb09c2a4),
	.w7(32'hbab48f95),
	.w8(32'h3b583aa9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c54f6),
	.w1(32'h3b69195d),
	.w2(32'h3ad20cd4),
	.w3(32'hbb98651a),
	.w4(32'hbac67743),
	.w5(32'hbb97f678),
	.w6(32'hb903968d),
	.w7(32'h3a3eb15e),
	.w8(32'hbc0a3d08),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc31f44),
	.w1(32'hba07d787),
	.w2(32'hbb3ddbe7),
	.w3(32'hba8b5736),
	.w4(32'h3ab7afff),
	.w5(32'hbaf20882),
	.w6(32'hbba2ed9e),
	.w7(32'hbab47269),
	.w8(32'hbb79c5a9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b7a0f),
	.w1(32'hba2fdbc8),
	.w2(32'hba8b2ec0),
	.w3(32'hbb852659),
	.w4(32'hbb816991),
	.w5(32'h3b98096b),
	.w6(32'hbb1280c0),
	.w7(32'hbafe3002),
	.w8(32'h3b425eb6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95d847),
	.w1(32'hba996572),
	.w2(32'hbba70fac),
	.w3(32'h3bddfb3a),
	.w4(32'h3ba86abe),
	.w5(32'hbb4ba5ae),
	.w6(32'hba080b55),
	.w7(32'hbaed8d49),
	.w8(32'hbbdbb3f2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76c20f),
	.w1(32'hba5f7930),
	.w2(32'hbb6977ee),
	.w3(32'hbaed75f4),
	.w4(32'hbb0f73df),
	.w5(32'hbb9798c1),
	.w6(32'hbb0836dc),
	.w7(32'hbb518d08),
	.w8(32'hbb0cc322),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf35841),
	.w1(32'hbbe12e44),
	.w2(32'hbbf9adba),
	.w3(32'hbbd0c0d8),
	.w4(32'hbb8d37c9),
	.w5(32'h39b08142),
	.w6(32'hbb906f76),
	.w7(32'hbade74b8),
	.w8(32'hbb9816c6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5af38c),
	.w1(32'hb892a086),
	.w2(32'hb96a1de5),
	.w3(32'h3a00a26e),
	.w4(32'h3894c5f6),
	.w5(32'hb90e1aae),
	.w6(32'h39f0a7b3),
	.w7(32'hbbc55f4d),
	.w8(32'hbb0b5c2d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b05a5),
	.w1(32'h3b750d1c),
	.w2(32'hb8e6aa15),
	.w3(32'h39b3088e),
	.w4(32'h3b5b5296),
	.w5(32'hb9e3b219),
	.w6(32'h3b4980ef),
	.w7(32'h3aeb7dfe),
	.w8(32'hbb2785ce),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6b4c2),
	.w1(32'hbb3e201d),
	.w2(32'hba4db2d1),
	.w3(32'hb8c1744a),
	.w4(32'h3af25712),
	.w5(32'h3a739f61),
	.w6(32'h3956b7f4),
	.w7(32'h3b22b96a),
	.w8(32'h3b0d56e2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073ca2),
	.w1(32'h3b71bc65),
	.w2(32'h3bb2e93b),
	.w3(32'h39db1731),
	.w4(32'h3b859903),
	.w5(32'hbb118985),
	.w6(32'h39b8e16c),
	.w7(32'h3b88f751),
	.w8(32'hbbb22d86),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f6445),
	.w1(32'hb8a558c0),
	.w2(32'hbb12dd33),
	.w3(32'hb9f45f2d),
	.w4(32'h3a72155c),
	.w5(32'hb9585261),
	.w6(32'hbb49fb5d),
	.w7(32'hba1e60e0),
	.w8(32'hba7fb1dd),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3169f),
	.w1(32'h3b76162f),
	.w2(32'h3b4d60e6),
	.w3(32'hbb11c0e1),
	.w4(32'hbb04909f),
	.w5(32'h3aa36295),
	.w6(32'hba9cb29a),
	.w7(32'hb62db3fa),
	.w8(32'h3ba4e6f9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b41a85),
	.w1(32'h3a803b4d),
	.w2(32'h3a9b46d1),
	.w3(32'h3b38db49),
	.w4(32'h3ae83c3a),
	.w5(32'hbae8e89c),
	.w6(32'h3c2089a0),
	.w7(32'h3bddad95),
	.w8(32'hbb08f566),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e657),
	.w1(32'h3be78dd4),
	.w2(32'h3bd31c67),
	.w3(32'hbac6abd8),
	.w4(32'hbb893109),
	.w5(32'h39cd233b),
	.w6(32'hbb2669c1),
	.w7(32'hbba46be6),
	.w8(32'h3bd48c76),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af30005),
	.w1(32'h3a04b720),
	.w2(32'hbb69b769),
	.w3(32'h3b44ad3a),
	.w4(32'h3b547af1),
	.w5(32'hbb99995a),
	.w6(32'h3b5ef89b),
	.w7(32'h3ba79ae7),
	.w8(32'hbbd73ed0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad29166),
	.w1(32'hbb25634f),
	.w2(32'hbb1533a5),
	.w3(32'hbb2b054d),
	.w4(32'hbacd0398),
	.w5(32'hbafd33d8),
	.w6(32'hbafcf6ad),
	.w7(32'hbaa78fa1),
	.w8(32'hba424c9f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fdd24),
	.w1(32'h3b618f40),
	.w2(32'h3b241f5d),
	.w3(32'hbb35665c),
	.w4(32'hbb1addde),
	.w5(32'hbb689106),
	.w6(32'hba547f8d),
	.w7(32'hbb2df638),
	.w8(32'hbb9004b6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5c419),
	.w1(32'hbb14fae3),
	.w2(32'hbb10f4fd),
	.w3(32'hbbaf2192),
	.w4(32'hbb9a154c),
	.w5(32'hbb2578b4),
	.w6(32'hbb1703f7),
	.w7(32'h3a1dbbbc),
	.w8(32'h3a870e84),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66cace),
	.w1(32'hb8c51304),
	.w2(32'hb9d549d1),
	.w3(32'h3a486214),
	.w4(32'hb9eba806),
	.w5(32'h3b98695c),
	.w6(32'h3be16e08),
	.w7(32'h3b70cb09),
	.w8(32'h398eeceb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac90ead),
	.w1(32'h399165c2),
	.w2(32'h3b95c461),
	.w3(32'h3b02d884),
	.w4(32'h3bcf2626),
	.w5(32'h397ab3ea),
	.w6(32'hb9cc6a5d),
	.w7(32'h3bf36546),
	.w8(32'hb95b7714),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9d83f),
	.w1(32'hbab7985a),
	.w2(32'h3a3f5d83),
	.w3(32'h3af354de),
	.w4(32'hba2a5391),
	.w5(32'h3b765b73),
	.w6(32'h3a4124f7),
	.w7(32'hb8f9c16d),
	.w8(32'h3b7b1c53),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f036),
	.w1(32'hba4ed6f6),
	.w2(32'h3ab248bf),
	.w3(32'h3b7cbdf6),
	.w4(32'h3bad555a),
	.w5(32'hbb223fcc),
	.w6(32'h3a454378),
	.w7(32'h3b7b8867),
	.w8(32'hbb615e02),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882a0cd),
	.w1(32'h3acd3432),
	.w2(32'hbaa4c0ae),
	.w3(32'hbae46759),
	.w4(32'hbb4abe37),
	.w5(32'hba7d77b9),
	.w6(32'hbbee0b5b),
	.w7(32'hbb496551),
	.w8(32'hbb7907a3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d78eec),
	.w1(32'h3ab95a07),
	.w2(32'h3ab41b8a),
	.w3(32'h3b178223),
	.w4(32'h3b687d35),
	.w5(32'h3b43aaf1),
	.w6(32'h39896a04),
	.w7(32'h39b54dc6),
	.w8(32'h3b9d99c1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19dbeb),
	.w1(32'h3b5981a5),
	.w2(32'hb97a0e7a),
	.w3(32'h392c26b5),
	.w4(32'h37b4253a),
	.w5(32'hbbf87627),
	.w6(32'h3b9e5ac6),
	.w7(32'h3b772b45),
	.w8(32'hbc46b9b4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bd19d),
	.w1(32'hbb734426),
	.w2(32'h3aab4b49),
	.w3(32'hbb9169d0),
	.w4(32'hbb63de5a),
	.w5(32'hba5b2395),
	.w6(32'hbbbf60a1),
	.w7(32'hbae46b02),
	.w8(32'hb931c6a0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb5fa0),
	.w1(32'hbb7efe00),
	.w2(32'hbc27c1f9),
	.w3(32'hbba8aa80),
	.w4(32'hb9fad96f),
	.w5(32'hbb8c0917),
	.w6(32'hbbd12f6b),
	.w7(32'hbb8495b3),
	.w8(32'hbba48b52),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2119),
	.w1(32'h3aa5421d),
	.w2(32'hbae90d5e),
	.w3(32'h3bddb285),
	.w4(32'h3bbce9c7),
	.w5(32'hbb3d448f),
	.w6(32'h3b7a1967),
	.w7(32'h3b78dae1),
	.w8(32'hbba8c8c8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb406f6),
	.w1(32'hbb3de535),
	.w2(32'hbbd90c1a),
	.w3(32'hbaf9f6a6),
	.w4(32'h3ab2ee4e),
	.w5(32'hb98032ab),
	.w6(32'hbb7adfa8),
	.w7(32'hba9b0b37),
	.w8(32'hbb6da582),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae14fa3),
	.w1(32'h3aa8d94f),
	.w2(32'h39134e8d),
	.w3(32'h3ba883bb),
	.w4(32'h3b4f682f),
	.w5(32'hbb26c01e),
	.w6(32'h3b3854e0),
	.w7(32'h3af281f4),
	.w8(32'hb783cd2b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8381d9),
	.w1(32'hbb2c9c5b),
	.w2(32'hbb848d5d),
	.w3(32'hbb1dcd39),
	.w4(32'hbb254937),
	.w5(32'h3b99963b),
	.w6(32'hba982b9a),
	.w7(32'hba8b6f04),
	.w8(32'h3ab59edd),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b6068),
	.w1(32'hba2d1503),
	.w2(32'h3aabf542),
	.w3(32'h3b8fe5e6),
	.w4(32'h3bb99d96),
	.w5(32'hbba81255),
	.w6(32'hb88c1cdd),
	.w7(32'h3a9906b9),
	.w8(32'hbb58e7d2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb400be7),
	.w1(32'hbae15c0a),
	.w2(32'hbb7f26f0),
	.w3(32'hbb56ceb7),
	.w4(32'hbb8555af),
	.w5(32'hbb181ebf),
	.w6(32'hbb443dde),
	.w7(32'hbb752055),
	.w8(32'hbbbebf16),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ffbb),
	.w1(32'hbb2bb39a),
	.w2(32'h3ad2a663),
	.w3(32'hbb357dc6),
	.w4(32'hbb4eb122),
	.w5(32'h39ff957a),
	.w6(32'hbb1177d1),
	.w7(32'hbaa6cdf1),
	.w8(32'h3a0a34f9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0aa40),
	.w1(32'hbb291d31),
	.w2(32'hbbc059bc),
	.w3(32'hbae22b00),
	.w4(32'hbaa6b55e),
	.w5(32'hbb9a7040),
	.w6(32'hbb8b35f2),
	.w7(32'hbb350707),
	.w8(32'hbbff0133),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85224f),
	.w1(32'hbb2f14ef),
	.w2(32'hbb4671e4),
	.w3(32'hbb5a319c),
	.w4(32'hbb219868),
	.w5(32'hbb494308),
	.w6(32'hbb865705),
	.w7(32'hbb110ccc),
	.w8(32'hbb22ba7e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b246a),
	.w1(32'hb9052239),
	.w2(32'h394dd45b),
	.w3(32'hbad11c7b),
	.w4(32'hba048899),
	.w5(32'hbb944eb5),
	.w6(32'hbaab177f),
	.w7(32'hba575151),
	.w8(32'hbb69b984),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ecaea),
	.w1(32'h390ceb97),
	.w2(32'h3ab52bd5),
	.w3(32'hbbbe2059),
	.w4(32'hbb8aa895),
	.w5(32'hba80bdc2),
	.w6(32'hbb842792),
	.w7(32'hbb80c954),
	.w8(32'hbaf61884),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e5055),
	.w1(32'h3a64c974),
	.w2(32'hbb771cdd),
	.w3(32'hbbd68f71),
	.w4(32'hbb481270),
	.w5(32'hbb8095ee),
	.w6(32'hbb7be7f7),
	.w7(32'hbb2a05de),
	.w8(32'hbb9e31c1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04b88e),
	.w1(32'hbbd0cba6),
	.w2(32'hbb75bcda),
	.w3(32'hbba319b2),
	.w4(32'hbb3cd1f2),
	.w5(32'h3b977614),
	.w6(32'hbbc09c75),
	.w7(32'hbb3b16d6),
	.w8(32'h3b0c4e25),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a403fca),
	.w1(32'hb984cb0f),
	.w2(32'h3a041164),
	.w3(32'h3b4e7fa8),
	.w4(32'h3b8c0367),
	.w5(32'h3bbe4d0c),
	.w6(32'h3980e42a),
	.w7(32'h3a7c324a),
	.w8(32'h3ab63a82),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbae496),
	.w1(32'hbb8a39f4),
	.w2(32'hbc06a4f0),
	.w3(32'h3bf38681),
	.w4(32'h3c43c011),
	.w5(32'hbbb05b36),
	.w6(32'hbb12b8c2),
	.w7(32'h3b94d053),
	.w8(32'hbbe00066),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b009b85),
	.w1(32'h3a188f83),
	.w2(32'hba12f3dd),
	.w3(32'h3b5207cc),
	.w4(32'h3b53e4ac),
	.w5(32'hba86a7c6),
	.w6(32'hb8d6e925),
	.w7(32'hbb29b7f3),
	.w8(32'hbb84e0f3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6c98d),
	.w1(32'hba910767),
	.w2(32'hbb0a43c3),
	.w3(32'h3ac07734),
	.w4(32'h3a935200),
	.w5(32'hbb5f6e5b),
	.w6(32'h3b1aad15),
	.w7(32'h3a387171),
	.w8(32'hbac5a8ee),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0079),
	.w1(32'hb93a59bb),
	.w2(32'h3ad5f3a2),
	.w3(32'hbb10e5db),
	.w4(32'hba8224b1),
	.w5(32'hbb32ffd1),
	.w6(32'h3a3038e0),
	.w7(32'h3978eea9),
	.w8(32'hbb33591e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1d24),
	.w1(32'hbadde74c),
	.w2(32'hba93b670),
	.w3(32'hbba42b44),
	.w4(32'hbb26b24b),
	.w5(32'hbbbaa5a0),
	.w6(32'hbb7680a5),
	.w7(32'hbb1dfa40),
	.w8(32'hbbbd3820),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb913770),
	.w1(32'hbb0b5653),
	.w2(32'hba76e730),
	.w3(32'hbbafd679),
	.w4(32'hbb5c48b6),
	.w5(32'hba52af56),
	.w6(32'hbbb4b415),
	.w7(32'hbb5109b4),
	.w8(32'hba6c45fc),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4598ca),
	.w1(32'hbaa86d64),
	.w2(32'hbae28aa7),
	.w3(32'h39d7c00b),
	.w4(32'hbb20f156),
	.w5(32'hbb267a33),
	.w6(32'h3a8a643a),
	.w7(32'hb9af1360),
	.w8(32'hbb281b3d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53961a),
	.w1(32'hbb43d2d6),
	.w2(32'hbb5a7ffd),
	.w3(32'hba81a12e),
	.w4(32'h3a20c1d1),
	.w5(32'hbb0fbc50),
	.w6(32'hbb8badd3),
	.w7(32'hbb2a7b14),
	.w8(32'hbb90f935),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807d0b),
	.w1(32'hbb05724a),
	.w2(32'hbbc3b3c4),
	.w3(32'hbac0d20c),
	.w4(32'h39dc4f79),
	.w5(32'hbbb06eed),
	.w6(32'hba97bd6f),
	.w7(32'h3a734562),
	.w8(32'hbbb1fdad),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb342c46),
	.w1(32'hb9258b6a),
	.w2(32'h3abd281e),
	.w3(32'hbb4bb590),
	.w4(32'h3a188c7f),
	.w5(32'hb99dba39),
	.w6(32'hbb6c4774),
	.w7(32'h3a35b898),
	.w8(32'hba279bc1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e6810),
	.w1(32'h3b1f551f),
	.w2(32'hbaa5d3f0),
	.w3(32'h38db33da),
	.w4(32'h3a9eaaca),
	.w5(32'h39de3cf2),
	.w6(32'hba5eb0d8),
	.w7(32'h3b32cc8c),
	.w8(32'hbab60857),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e55db),
	.w1(32'hb9d3c1fd),
	.w2(32'hbac67380),
	.w3(32'hba2a65e8),
	.w4(32'hba382469),
	.w5(32'h3a17cad2),
	.w6(32'h3b7a8b51),
	.w7(32'h3b58b394),
	.w8(32'h3b1fb4a7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905d67a),
	.w1(32'hba6e5faa),
	.w2(32'hbaf93b52),
	.w3(32'h3ab3bfa4),
	.w4(32'hba4fe7a9),
	.w5(32'h3b048cd8),
	.w6(32'h3ab4f8c8),
	.w7(32'hba5501cc),
	.w8(32'h3a3566ce),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e4ea7),
	.w1(32'hbba80cd1),
	.w2(32'hbb6ab030),
	.w3(32'hb989246c),
	.w4(32'hbb208f73),
	.w5(32'hbb77c9be),
	.w6(32'h3b331e52),
	.w7(32'h3b389ef9),
	.w8(32'hbb48f977),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb283569),
	.w1(32'hba642487),
	.w2(32'h3aea8674),
	.w3(32'hbad97bce),
	.w4(32'hbae94539),
	.w5(32'hb9b27a70),
	.w6(32'hba5c6d90),
	.w7(32'h3a917297),
	.w8(32'hbaf3b617),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c7b22),
	.w1(32'hba2cdb99),
	.w2(32'h3af110a1),
	.w3(32'hbaa814f2),
	.w4(32'h3ae26d0a),
	.w5(32'hbb968672),
	.w6(32'hbbaaa1a7),
	.w7(32'h3b504642),
	.w8(32'hbb908881),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54e65f),
	.w1(32'h3b14c54c),
	.w2(32'h3b229dc2),
	.w3(32'hbbbbbc89),
	.w4(32'hbb02a849),
	.w5(32'hb9ea2fd6),
	.w6(32'hbb98ba1f),
	.w7(32'hba954e0b),
	.w8(32'hbb141eb3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d169c),
	.w1(32'h38b85ce5),
	.w2(32'hbae46c41),
	.w3(32'hbb065b0a),
	.w4(32'hba1d49c9),
	.w5(32'hbb613a8a),
	.w6(32'hbb294209),
	.w7(32'hbb0097f7),
	.w8(32'hbbba5c97),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8074ad),
	.w1(32'hbb01d96c),
	.w2(32'h3a332f11),
	.w3(32'hbb9157ad),
	.w4(32'hbac5871e),
	.w5(32'h3a1b9fbb),
	.w6(32'hbb6e18b2),
	.w7(32'hbafdbb5b),
	.w8(32'h3a82c7aa),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5109ed),
	.w1(32'h3a4118e7),
	.w2(32'hb97b4a5a),
	.w3(32'h3ad574b1),
	.w4(32'h3b3efa54),
	.w5(32'hbb40cdad),
	.w6(32'hbabc6d2d),
	.w7(32'h3623e638),
	.w8(32'hbbaf256a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85e0f6),
	.w1(32'hbaaa3079),
	.w2(32'hbb013db9),
	.w3(32'h3ab2b891),
	.w4(32'h3b07b47d),
	.w5(32'hba9ff927),
	.w6(32'hba662905),
	.w7(32'h3aa00a7d),
	.w8(32'hbb80ddae),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a5468),
	.w1(32'hbb33dd5b),
	.w2(32'hbbf5cd9a),
	.w3(32'hbb462f85),
	.w4(32'hba360311),
	.w5(32'hbb67a58f),
	.w6(32'hbc1ba700),
	.w7(32'hbba89c1b),
	.w8(32'hbb8aad6f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c92da7),
	.w1(32'h3a593153),
	.w2(32'h3a2427b4),
	.w3(32'hba8d3f34),
	.w4(32'hba956d94),
	.w5(32'hbb0a4c51),
	.w6(32'h3ac54a9e),
	.w7(32'h3b39aed0),
	.w8(32'hbb005cd2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa1db),
	.w1(32'hbb68ff42),
	.w2(32'hba8852e0),
	.w3(32'hbae181da),
	.w4(32'hb940c018),
	.w5(32'h3b534aab),
	.w6(32'hbb4a96b9),
	.w7(32'hb92e9813),
	.w8(32'h3b36e3b3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3009bc),
	.w1(32'h3a56098a),
	.w2(32'h3703a344),
	.w3(32'h3b650b37),
	.w4(32'h3b40634b),
	.w5(32'hbb33f6d0),
	.w6(32'hb87d095a),
	.w7(32'h3b369c69),
	.w8(32'hbbb03269),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dc7f4),
	.w1(32'hbaa4729d),
	.w2(32'hbb8ffd4c),
	.w3(32'hba05e9ab),
	.w4(32'h39e8bac5),
	.w5(32'hbb984bf0),
	.w6(32'hbb8b69e9),
	.w7(32'hba9cbedd),
	.w8(32'hbc0857b6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3107d),
	.w1(32'hbaef5ae6),
	.w2(32'hbb1bc3d9),
	.w3(32'h39964127),
	.w4(32'h3b018745),
	.w5(32'h3a88fcee),
	.w6(32'hbafdca51),
	.w7(32'hb9b8979b),
	.w8(32'hbbb19983),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad72871),
	.w1(32'hbb0d7060),
	.w2(32'h39d2c30d),
	.w3(32'h3b380fbd),
	.w4(32'h39e2672e),
	.w5(32'hbb22fa70),
	.w6(32'hbba02383),
	.w7(32'hbb026c24),
	.w8(32'hbb658a67),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53ee17),
	.w1(32'hbb6cd683),
	.w2(32'hbb099119),
	.w3(32'hbb07a0e1),
	.w4(32'hbaf35215),
	.w5(32'h3a178e47),
	.w6(32'hbad83289),
	.w7(32'hba88939a),
	.w8(32'hb9e22cd2),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dd3bc),
	.w1(32'hbab38c53),
	.w2(32'h3a091fe0),
	.w3(32'h3b16352a),
	.w4(32'h3b9e91a9),
	.w5(32'hbb61b528),
	.w6(32'h3a4540b4),
	.w7(32'h3af46ecc),
	.w8(32'hbac4c101),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89d78b),
	.w1(32'h3ba61f7f),
	.w2(32'hba08d16f),
	.w3(32'hbbb121e8),
	.w4(32'hbb93d213),
	.w5(32'hbc09b56a),
	.w6(32'hb9d19a6f),
	.w7(32'h3b327ecf),
	.w8(32'hbb5a97c3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3fbd8),
	.w1(32'hbb066725),
	.w2(32'hbaf7b0fc),
	.w3(32'hbb2a24d0),
	.w4(32'hba50cb04),
	.w5(32'hbbd59ebe),
	.w6(32'hbb80d7d9),
	.w7(32'h3b3c415a),
	.w8(32'hbbdff864),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17cc9),
	.w1(32'hbb70d0d3),
	.w2(32'hbba4b5ac),
	.w3(32'h3985dd11),
	.w4(32'hba23cd22),
	.w5(32'hbb9cf249),
	.w6(32'hbba45faf),
	.w7(32'hbb19a5cf),
	.w8(32'hbbabd81e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e12b84),
	.w1(32'h3b22785a),
	.w2(32'h3bc519e9),
	.w3(32'hbbd9a8d4),
	.w4(32'hbb6360d5),
	.w5(32'hbae4199e),
	.w6(32'hbbb2d206),
	.w7(32'hbb80b8b0),
	.w8(32'hbb5a3a80),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea91ad),
	.w1(32'h3a934ba9),
	.w2(32'hba98c3e0),
	.w3(32'hbb4dd2fc),
	.w4(32'hbad05f46),
	.w5(32'h3a93b165),
	.w6(32'hbb94e87f),
	.w7(32'hbbaf0ee7),
	.w8(32'hb99cc65d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fe1ee),
	.w1(32'hbac96fb6),
	.w2(32'h3a44b9dc),
	.w3(32'hbad76642),
	.w4(32'h3ab150c0),
	.w5(32'h3b42b9ec),
	.w6(32'hba615e81),
	.w7(32'h3b16f6b7),
	.w8(32'hbb20b751),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f0cd1),
	.w1(32'h3b93bb96),
	.w2(32'h3ba38ccf),
	.w3(32'h3aefdb6a),
	.w4(32'h3b24b3f1),
	.w5(32'h3b1581c4),
	.w6(32'hbb83ce16),
	.w7(32'h3a24e178),
	.w8(32'h3b07da15),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39c282),
	.w1(32'h3b48a0ba),
	.w2(32'h3bb185d0),
	.w3(32'h3bba2d42),
	.w4(32'h3b2f346f),
	.w5(32'hbb2ca339),
	.w6(32'h3b9f09c7),
	.w7(32'h3b95338b),
	.w8(32'h3b34c1d4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24c340),
	.w1(32'h3ac28dcf),
	.w2(32'hba413585),
	.w3(32'hbb0b4ff7),
	.w4(32'h3a833bc3),
	.w5(32'hbb87029b),
	.w6(32'h3b148b2f),
	.w7(32'h3ac91792),
	.w8(32'hbc0e9a5a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf6dcb),
	.w1(32'hbbedff29),
	.w2(32'hb99ec405),
	.w3(32'hbc270de9),
	.w4(32'hbbf15cff),
	.w5(32'h3bca86d3),
	.w6(32'hbcad4992),
	.w7(32'hbbf5ff57),
	.w8(32'h3b6c20d1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c454a),
	.w1(32'h3c489719),
	.w2(32'h3b41bd1a),
	.w3(32'h3c12ae5f),
	.w4(32'h3b15da1e),
	.w5(32'hbb3dc704),
	.w6(32'hbbfa4045),
	.w7(32'h3c8d2d10),
	.w8(32'hbc5f6f9e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0252dd),
	.w1(32'hbbee82a1),
	.w2(32'h3a9ebc0b),
	.w3(32'hbc47ca1f),
	.w4(32'h3a81ab47),
	.w5(32'h3b1ef9f8),
	.w6(32'hbcdf70bf),
	.w7(32'hbc8401d6),
	.w8(32'h3b5a3dd2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29aefe),
	.w1(32'hbc027c11),
	.w2(32'hbb2a6438),
	.w3(32'h3c150253),
	.w4(32'h3b14b4ce),
	.w5(32'h3a927f8a),
	.w6(32'h3ba2ffd4),
	.w7(32'h3b68450d),
	.w8(32'h3aa2c043),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85d8ff),
	.w1(32'hbaa7fb51),
	.w2(32'hbb60910e),
	.w3(32'hbb800b94),
	.w4(32'hbb3dcece),
	.w5(32'h3b25d349),
	.w6(32'hbc1a2d30),
	.w7(32'h3b9c241a),
	.w8(32'h3b447692),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dd51b),
	.w1(32'h3ce1ed2b),
	.w2(32'h3ca3fee9),
	.w3(32'h3c9f0a61),
	.w4(32'h3c3d3e07),
	.w5(32'hbc45406d),
	.w6(32'h3bb856c8),
	.w7(32'h3cff34bf),
	.w8(32'hbc37c9e9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4c7b0),
	.w1(32'hb8adf9ff),
	.w2(32'h3b1874b8),
	.w3(32'hbbad16df),
	.w4(32'h3bf975a8),
	.w5(32'h3c4fa520),
	.w6(32'hbc53752e),
	.w7(32'hbc032c9c),
	.w8(32'h3c1389c3),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60dac5),
	.w1(32'h3be4e8d5),
	.w2(32'h3c3a67a7),
	.w3(32'h3c2c5777),
	.w4(32'h3c308957),
	.w5(32'h3c27a98a),
	.w6(32'hbc899ec1),
	.w7(32'h3b483c0f),
	.w8(32'h3c219a8d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850937),
	.w1(32'hbbc9b6ba),
	.w2(32'hbb2a5a82),
	.w3(32'h3c57ce8b),
	.w4(32'h38bee7fc),
	.w5(32'h3b9a48e7),
	.w6(32'hbbfee682),
	.w7(32'hbb7ba5ec),
	.w8(32'h3b1e1030),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d09c6a),
	.w1(32'hbb2451ec),
	.w2(32'hbb3b80f7),
	.w3(32'hb9718955),
	.w4(32'hba1285a8),
	.w5(32'hbb1c9637),
	.w6(32'hbafd6934),
	.w7(32'hbb14b4b2),
	.w8(32'hbc2f50f7),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadacf12),
	.w1(32'hbbce9e9c),
	.w2(32'h3c09de4c),
	.w3(32'hbc172c06),
	.w4(32'h3a69ee0f),
	.w5(32'hbb28f752),
	.w6(32'hbcb2f9b2),
	.w7(32'hbb1b553b),
	.w8(32'hbb01397c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac824e8),
	.w1(32'hbb9001c0),
	.w2(32'h3a90606e),
	.w3(32'hbb969dfc),
	.w4(32'h3a173153),
	.w5(32'h3b39effc),
	.w6(32'hb9fe9391),
	.w7(32'h39a4f690),
	.w8(32'h3a01cfb2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8a0d6),
	.w1(32'hba5a1bc2),
	.w2(32'h3bc78d8b),
	.w3(32'hbb139479),
	.w4(32'hbbb6ce44),
	.w5(32'hbbdf5fa5),
	.w6(32'hbb9e26c5),
	.w7(32'hbb805ae0),
	.w8(32'hbb200846),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d419a),
	.w1(32'hbbc2d815),
	.w2(32'hbbf98569),
	.w3(32'hbace8f1f),
	.w4(32'hbb97d995),
	.w5(32'hbc60f22a),
	.w6(32'hbc2fd145),
	.w7(32'hbbce4fca),
	.w8(32'hbc8c85e0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95cb63),
	.w1(32'hbcc0110f),
	.w2(32'hbcad5b42),
	.w3(32'hbc851fa2),
	.w4(32'hbc6c4546),
	.w5(32'hbb1c3bf8),
	.w6(32'hbc28ea21),
	.w7(32'hbcb3836b),
	.w8(32'hbbba4ef5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5e27),
	.w1(32'h38eb87aa),
	.w2(32'hbbcf4745),
	.w3(32'hbb336e21),
	.w4(32'hbb868adb),
	.w5(32'hbb0f00c4),
	.w6(32'hb9dfc1be),
	.w7(32'hbba82810),
	.w8(32'hbaa4d304),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34f8ef),
	.w1(32'h3aaaa8c3),
	.w2(32'h3bc01fe2),
	.w3(32'h3c099cf8),
	.w4(32'h3c8fa737),
	.w5(32'h39d2d312),
	.w6(32'hbc77640d),
	.w7(32'h3c642d1d),
	.w8(32'h3bc6945d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993b80f),
	.w1(32'hbbdeef61),
	.w2(32'h3b100d01),
	.w3(32'h3b8a73c5),
	.w4(32'hba87a090),
	.w5(32'hbae75e34),
	.w6(32'hbae8beef),
	.w7(32'hbab6a46c),
	.w8(32'hbba62bf7),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91feac),
	.w1(32'hbb74be1d),
	.w2(32'hbbad2787),
	.w3(32'hbaa1f430),
	.w4(32'hbb8ad25c),
	.w5(32'hbb4b334f),
	.w6(32'hbb2e8e58),
	.w7(32'hbbb3f052),
	.w8(32'h3c053565),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f1352),
	.w1(32'h3b80fb20),
	.w2(32'hbbed40bd),
	.w3(32'h3aa6bf12),
	.w4(32'h3c09bdde),
	.w5(32'h3bb25389),
	.w6(32'hbc731759),
	.w7(32'hb7868f48),
	.w8(32'h3ba7f1c6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a469b),
	.w1(32'h3c1cacda),
	.w2(32'h3c2f7d11),
	.w3(32'h38ac32e3),
	.w4(32'h3c1f2c20),
	.w5(32'h3bb7dbec),
	.w6(32'hbbcac428),
	.w7(32'h3c48a365),
	.w8(32'hbc45d8d5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf8d71),
	.w1(32'hb9ebd029),
	.w2(32'h3be7eb11),
	.w3(32'hbc0a784e),
	.w4(32'h3b79e399),
	.w5(32'hbb14eff4),
	.w6(32'hbd41d619),
	.w7(32'hbbd276f4),
	.w8(32'hbb20ba62),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398db3ab),
	.w1(32'hb8629c2a),
	.w2(32'h3c305370),
	.w3(32'h3bef1dae),
	.w4(32'hbb3f4c4a),
	.w5(32'hbb364ec1),
	.w6(32'h3a3d6918),
	.w7(32'hbbfd9950),
	.w8(32'hbb9fbb01),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5c6f),
	.w1(32'hbb74a19a),
	.w2(32'hbb8c3151),
	.w3(32'hbb43b582),
	.w4(32'hbb6e1fa1),
	.w5(32'h3a1f56ec),
	.w6(32'h3b305818),
	.w7(32'h3b742c45),
	.w8(32'h3b999178),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98b786),
	.w1(32'hbb4c8f66),
	.w2(32'hbc10334d),
	.w3(32'h3b2caaf0),
	.w4(32'hbb6d7bf2),
	.w5(32'hb91f6c66),
	.w6(32'h3c305785),
	.w7(32'hbc1cbe0e),
	.w8(32'h3ba045bb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d4faa),
	.w1(32'hbbb82498),
	.w2(32'hbc41eef8),
	.w3(32'h3b009700),
	.w4(32'hbbccaee3),
	.w5(32'hbb8ec46e),
	.w6(32'h3c68f70e),
	.w7(32'hbc19fbe5),
	.w8(32'hbb6a636d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8e0da),
	.w1(32'hbbea623f),
	.w2(32'hbc384f3f),
	.w3(32'hbac2c747),
	.w4(32'hbacfb5de),
	.w5(32'hbaed126e),
	.w6(32'h3b06af19),
	.w7(32'hbbb2bb5c),
	.w8(32'h3a73581e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1dbfb),
	.w1(32'h3aa07595),
	.w2(32'hbc29e1da),
	.w3(32'hbc1ecac2),
	.w4(32'hbbd6c535),
	.w5(32'h3b38d7c5),
	.w6(32'hbb892bdd),
	.w7(32'hbc20787f),
	.w8(32'hbbfcdaf8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad476ba),
	.w1(32'hbab88b51),
	.w2(32'h3a847538),
	.w3(32'h399ff550),
	.w4(32'h3b191014),
	.w5(32'hbaa1818c),
	.w6(32'hba499aea),
	.w7(32'hbb160c53),
	.w8(32'hbb200bc3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bc559),
	.w1(32'hbb03cf70),
	.w2(32'h3c1bb9ae),
	.w3(32'hbb0b842f),
	.w4(32'h3c1ae857),
	.w5(32'hbbec20de),
	.w6(32'hbc84ab49),
	.w7(32'h3b88f1d6),
	.w8(32'hbb8ebb4e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule