module layer_8_featuremap_133(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa5b2),
	.w1(32'h397d9a0a),
	.w2(32'h3b1b74e1),
	.w3(32'hbc62a16b),
	.w4(32'hbb553237),
	.w5(32'hba93bb0e),
	.w6(32'hbb5443aa),
	.w7(32'hbb4c3a6c),
	.w8(32'hbc0a19ed),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8954539),
	.w1(32'h3be40ec0),
	.w2(32'h3a9a97cb),
	.w3(32'h3ad53c5c),
	.w4(32'hbba11793),
	.w5(32'h3b709132),
	.w6(32'h3b0fd3ab),
	.w7(32'hbbb11dc1),
	.w8(32'h3bcb30ed),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ee8d5),
	.w1(32'h3bc5e6ba),
	.w2(32'hba673788),
	.w3(32'h3b29e320),
	.w4(32'hbbcaa40a),
	.w5(32'hbc01eb95),
	.w6(32'h3b5e67c8),
	.w7(32'hbb8716f9),
	.w8(32'hbc2c42fb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f0a5f),
	.w1(32'hbaa3d3e7),
	.w2(32'h3ab15b04),
	.w3(32'hbb245578),
	.w4(32'hbc14db68),
	.w5(32'h3b5e0469),
	.w6(32'hbc03ea08),
	.w7(32'hbc07d6e1),
	.w8(32'hbb8cdc2f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9e699),
	.w1(32'h3bdfc37c),
	.w2(32'h3b09f0d8),
	.w3(32'h3a7465b9),
	.w4(32'hbb894a81),
	.w5(32'h3bb16f5b),
	.w6(32'h3ad8c731),
	.w7(32'h3b29c489),
	.w8(32'hba6066a1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f37e3),
	.w1(32'h3c2bbd32),
	.w2(32'h3b898fc6),
	.w3(32'h3c246664),
	.w4(32'h3b8608d0),
	.w5(32'h3a5892fb),
	.w6(32'h3b66ed29),
	.w7(32'hbaafb734),
	.w8(32'hbb79d584),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb041),
	.w1(32'hbb994819),
	.w2(32'hbbceadb7),
	.w3(32'h3b88c290),
	.w4(32'hbbbbe352),
	.w5(32'hbbe829ef),
	.w6(32'hb94afc16),
	.w7(32'hbc046f2b),
	.w8(32'hbc2cf063),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd1d57),
	.w1(32'hbb9b97fc),
	.w2(32'h3b96cc37),
	.w3(32'h3a0467b8),
	.w4(32'h3aa39c5a),
	.w5(32'h3c501d8b),
	.w6(32'hbbc6406d),
	.w7(32'hbb564d00),
	.w8(32'h3c18d1c8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07ee4),
	.w1(32'hbb30c62d),
	.w2(32'h3b3eb76d),
	.w3(32'hbc9021ca),
	.w4(32'hbbd8f3a6),
	.w5(32'hbb658eb2),
	.w6(32'hbbf977dd),
	.w7(32'hbb6aa8c6),
	.w8(32'hbb7f0867),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42859e),
	.w1(32'h3bfdca3e),
	.w2(32'h3c8a4669),
	.w3(32'hbb2aa432),
	.w4(32'hbb7fb573),
	.w5(32'h3aa829b2),
	.w6(32'h3b2deff4),
	.w7(32'hba885512),
	.w8(32'h3bb3a774),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cda84),
	.w1(32'hbc29884e),
	.w2(32'hbbc6af37),
	.w3(32'hbbe7d104),
	.w4(32'hbc2e207e),
	.w5(32'hbc34b078),
	.w6(32'hbc4ec0a1),
	.w7(32'hbc3e52ed),
	.w8(32'hbc724963),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb570b0f),
	.w1(32'h3b8c5cb1),
	.w2(32'h3b27787e),
	.w3(32'h3b8d097b),
	.w4(32'hbb87da19),
	.w5(32'h3bca24c4),
	.w6(32'h3b803ba5),
	.w7(32'hbad376fc),
	.w8(32'hbb0ff803),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd101b),
	.w1(32'h3a9cbfcc),
	.w2(32'h3b7094a6),
	.w3(32'h3aa257ea),
	.w4(32'hbb030292),
	.w5(32'hbb2cecb3),
	.w6(32'h3a6b5aea),
	.w7(32'h382ab318),
	.w8(32'hbb15accc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30a06f),
	.w1(32'hbb0b9a38),
	.w2(32'h39e024c4),
	.w3(32'hbb4a689b),
	.w4(32'h3b0868a6),
	.w5(32'hbb467b1a),
	.w6(32'hbb92af3c),
	.w7(32'h3ae8c565),
	.w8(32'hbb13fa2a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fda730),
	.w1(32'hbb4cefc9),
	.w2(32'hba0adeec),
	.w3(32'hba8bc0a3),
	.w4(32'h3a958f4b),
	.w5(32'hba6b3aa0),
	.w6(32'hba96cec3),
	.w7(32'h3aba396f),
	.w8(32'h3a20dad7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e61db),
	.w1(32'hbb165ae4),
	.w2(32'h3bead456),
	.w3(32'hbabb82a6),
	.w4(32'h39de3337),
	.w5(32'h3c083ac6),
	.w6(32'hb86aa166),
	.w7(32'h3b31ac49),
	.w8(32'h3b09f3ca),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b564f),
	.w1(32'h38918a6e),
	.w2(32'hbc580201),
	.w3(32'h3aa0d668),
	.w4(32'hbbe967c8),
	.w5(32'hbb895e70),
	.w6(32'h3abe0bd6),
	.w7(32'hbc385a0f),
	.w8(32'hbc07db63),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba5ce0),
	.w1(32'hbb4c5712),
	.w2(32'h3bc244f0),
	.w3(32'h3a16db3e),
	.w4(32'hb9b1def4),
	.w5(32'h3c1ce249),
	.w6(32'hbc162d35),
	.w7(32'hbbcfe516),
	.w8(32'h3b4b8be5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabcf07),
	.w1(32'hbb955f6d),
	.w2(32'h3cb1447f),
	.w3(32'hbc293300),
	.w4(32'hbc2d304a),
	.w5(32'h3cc81863),
	.w6(32'hbc3fc72c),
	.w7(32'hbbf838b3),
	.w8(32'h3c21f3fd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb4ee9),
	.w1(32'h3ca4deef),
	.w2(32'h3bed9377),
	.w3(32'h3c1bda54),
	.w4(32'h3b2beba2),
	.w5(32'hbba83328),
	.w6(32'h3b125ea5),
	.w7(32'h3ba280ec),
	.w8(32'h3bbb12f1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbabb34),
	.w1(32'hb99dde67),
	.w2(32'h3c1663af),
	.w3(32'hba9a0320),
	.w4(32'hbb566349),
	.w5(32'hbc01c143),
	.w6(32'h3c4f9b4f),
	.w7(32'h3c06b246),
	.w8(32'hbc18860d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1921f),
	.w1(32'h3c4df743),
	.w2(32'h3c5b5f4f),
	.w3(32'h3c1cb439),
	.w4(32'h3c9d915a),
	.w5(32'h3c3d5184),
	.w6(32'h3c4a0e3d),
	.w7(32'h3c9e3734),
	.w8(32'h3cfadab6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c628bc6),
	.w1(32'h3c495e47),
	.w2(32'h3c625f23),
	.w3(32'hbc337a75),
	.w4(32'hbcd5111d),
	.w5(32'h3b5437ef),
	.w6(32'hbc6d84f2),
	.w7(32'hbc384d94),
	.w8(32'hbb52edb2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2efbba),
	.w1(32'h3a38d5c5),
	.w2(32'hbb3a9e3b),
	.w3(32'hbbcb2c19),
	.w4(32'hbae78da7),
	.w5(32'hbb4f9663),
	.w6(32'hbb3be1d3),
	.w7(32'hbb8ce480),
	.w8(32'hbb91ff34),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba29cea),
	.w1(32'hbb88540d),
	.w2(32'h3b9fc207),
	.w3(32'hbb3dbc03),
	.w4(32'h3bd95b40),
	.w5(32'h3b53fe51),
	.w6(32'hbb58c07b),
	.w7(32'h3befb920),
	.w8(32'h3c030880),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdc52b),
	.w1(32'h3b90cb9a),
	.w2(32'h3b941062),
	.w3(32'hbbb48c31),
	.w4(32'h3bbdba41),
	.w5(32'hbbb09e4d),
	.w6(32'hbc1ebbcf),
	.w7(32'hbbfd869c),
	.w8(32'hbbe00199),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc63673),
	.w1(32'hbac5728d),
	.w2(32'hbba4354e),
	.w3(32'hb9fc4efc),
	.w4(32'h3a7f5bdd),
	.w5(32'hbbb082b4),
	.w6(32'hbb9d55ad),
	.w7(32'h3be0fae8),
	.w8(32'hbbd560ac),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7981d6),
	.w1(32'hbd804c51),
	.w2(32'h3cc0ff9b),
	.w3(32'hbcbcc647),
	.w4(32'hbd117136),
	.w5(32'h3cb327ba),
	.w6(32'hbd8147f7),
	.w7(32'hbc589d90),
	.w8(32'h3d1f5d76),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08e1e3),
	.w1(32'h3c0cd57e),
	.w2(32'h3bb2e833),
	.w3(32'h3b6081ca),
	.w4(32'hbc319ebb),
	.w5(32'hbbe8a5b0),
	.w6(32'h3c612cbe),
	.w7(32'hbc11f1ab),
	.w8(32'hbbab48e8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc057455),
	.w1(32'h3b9c4da4),
	.w2(32'h3c94c232),
	.w3(32'h39fdbb92),
	.w4(32'hbaae6852),
	.w5(32'hbb596f83),
	.w6(32'hbbf48a1b),
	.w7(32'h3c7392d4),
	.w8(32'hbb29df7f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a481190),
	.w1(32'hbc1949f8),
	.w2(32'h3b006d7b),
	.w3(32'h38380ff4),
	.w4(32'h3ba4c9d6),
	.w5(32'h3c0c6c46),
	.w6(32'hbc25fb51),
	.w7(32'h3bec6437),
	.w8(32'h3c1b1859),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c133eca),
	.w1(32'h3b59e36e),
	.w2(32'hbb9d8952),
	.w3(32'h3ba46a28),
	.w4(32'hbc1dbe0a),
	.w5(32'hbbd7d9b0),
	.w6(32'h3c0c2d0e),
	.w7(32'hbb2ebd2a),
	.w8(32'hbc576fd8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe322a4),
	.w1(32'h3a66da32),
	.w2(32'hbbc09c6a),
	.w3(32'h393e7c34),
	.w4(32'hbbfce749),
	.w5(32'hbbae6e03),
	.w6(32'hb821180c),
	.w7(32'hbbf87773),
	.w8(32'hbab8a1cd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc072749),
	.w1(32'hb947842c),
	.w2(32'h3bb307fb),
	.w3(32'h39f8922f),
	.w4(32'hbbd56ec0),
	.w5(32'hb95c99c7),
	.w6(32'hbb08718e),
	.w7(32'hbbb764ee),
	.w8(32'hbb79749f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b48a),
	.w1(32'hbb15f48e),
	.w2(32'h3b9081cb),
	.w3(32'h3b9e83d8),
	.w4(32'h3becaa84),
	.w5(32'h3b9c90ec),
	.w6(32'h3ba80c63),
	.w7(32'h3bd9eba8),
	.w8(32'h3b87717d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bd3a5),
	.w1(32'hbb5edd5a),
	.w2(32'h3c099b84),
	.w3(32'hba8d4705),
	.w4(32'h3bd756ec),
	.w5(32'h3c3fd8c5),
	.w6(32'hbb258685),
	.w7(32'h3bf16978),
	.w8(32'h3c77c1a8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3810b7),
	.w1(32'h3c8884a8),
	.w2(32'hbb4792b6),
	.w3(32'h3b8005b1),
	.w4(32'h3ae4d5ec),
	.w5(32'h3b0b5980),
	.w6(32'h3badf7f5),
	.w7(32'hbb645d0b),
	.w8(32'hbb8e2e6b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25815d),
	.w1(32'h3bb22892),
	.w2(32'h3bdd6a67),
	.w3(32'h3beca7f7),
	.w4(32'h3c084583),
	.w5(32'h3c58c7e2),
	.w6(32'hbb0f7a2f),
	.w7(32'h3bd6d5ea),
	.w8(32'h3c8a5c32),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f7a00),
	.w1(32'h3b2cb6cf),
	.w2(32'h38853f86),
	.w3(32'hba952623),
	.w4(32'h38e7931f),
	.w5(32'hbb561a08),
	.w6(32'hb9902a1b),
	.w7(32'hbbb9a296),
	.w8(32'h39fad9ac),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dac64),
	.w1(32'h3b57fffc),
	.w2(32'h3c0a6b80),
	.w3(32'h39d19c66),
	.w4(32'hbb5ed388),
	.w5(32'hbbfad4cb),
	.w6(32'h3ae0d750),
	.w7(32'h3c57b673),
	.w8(32'h3c5ce4f1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda7338),
	.w1(32'h3cc0cb39),
	.w2(32'h3cf07e0f),
	.w3(32'hbc6bfc9c),
	.w4(32'hbab69d30),
	.w5(32'h3cb0a324),
	.w6(32'h39cbb1ef),
	.w7(32'hbbe823ed),
	.w8(32'h3b9f9e0c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c163b),
	.w1(32'hbb4e6515),
	.w2(32'h3ab08e2f),
	.w3(32'h3b9ee287),
	.w4(32'hbc457d9b),
	.w5(32'h3b915064),
	.w6(32'hb797d4ea),
	.w7(32'h3b2720ca),
	.w8(32'h3b930cca),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af0f91),
	.w1(32'h3bd36a7b),
	.w2(32'h3c65dd46),
	.w3(32'h38e6906d),
	.w4(32'h3c508423),
	.w5(32'hbbb41c65),
	.w6(32'h3c1c32d5),
	.w7(32'h3be5ed42),
	.w8(32'hbc09ea8f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bdb85),
	.w1(32'hbab6666b),
	.w2(32'hb9830b44),
	.w3(32'hbaa9be68),
	.w4(32'hbb494836),
	.w5(32'hbbba9ea4),
	.w6(32'hbc195676),
	.w7(32'hbb4a4ac6),
	.w8(32'hbbc1f9a2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf8fe9),
	.w1(32'hbbfac3cc),
	.w2(32'h3b7fe496),
	.w3(32'hbc741d38),
	.w4(32'hbc3cf1d0),
	.w5(32'hbbe14685),
	.w6(32'hbca23f72),
	.w7(32'hbc4bc969),
	.w8(32'hbb7c7db3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc701f69),
	.w1(32'hbb4cdbfb),
	.w2(32'hbaa84f90),
	.w3(32'hbbd3fe4b),
	.w4(32'h3ac9307f),
	.w5(32'h3c2b3271),
	.w6(32'hbba289bc),
	.w7(32'h3c100593),
	.w8(32'h3c67e29c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69fe26),
	.w1(32'h3ba3ae80),
	.w2(32'h3aed973c),
	.w3(32'h3b2e0652),
	.w4(32'h3b77d4a3),
	.w5(32'hbb48f453),
	.w6(32'h3bba90f4),
	.w7(32'h3c18942e),
	.w8(32'h3c271e9d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc30e8c),
	.w1(32'h3c154910),
	.w2(32'h3a212995),
	.w3(32'h3b2c0dba),
	.w4(32'h3c9d6b51),
	.w5(32'h3c2c91c1),
	.w6(32'h3b9c51cc),
	.w7(32'h3b82a5df),
	.w8(32'h3cb97580),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8483d5),
	.w1(32'h3c2f9bc2),
	.w2(32'hbad9b5ef),
	.w3(32'h3b10af65),
	.w4(32'hbbf85465),
	.w5(32'h3b8e25a6),
	.w6(32'hbaafc27e),
	.w7(32'hbb279418),
	.w8(32'hbb5a21bd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae0fc0),
	.w1(32'h3b18fedf),
	.w2(32'h3c1686cb),
	.w3(32'h3b12de26),
	.w4(32'hbc21b600),
	.w5(32'hbba01ef1),
	.w6(32'h3a01eefc),
	.w7(32'hbc05f1d2),
	.w8(32'hbb2b0f20),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ae8df),
	.w1(32'h3c4937db),
	.w2(32'h3b90977e),
	.w3(32'h3bfa575d),
	.w4(32'h3c705931),
	.w5(32'h3cafd2c2),
	.w6(32'h3c0e2154),
	.w7(32'hb8d9b19a),
	.w8(32'h3c355d77),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b2034),
	.w1(32'hb9f842dd),
	.w2(32'h3a4341b6),
	.w3(32'h3b37c467),
	.w4(32'hbb6fe843),
	.w5(32'h3bac990e),
	.w6(32'hbcccdfb8),
	.w7(32'hbd084ffe),
	.w8(32'hbc1344e4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefaaf2),
	.w1(32'hbb32ab93),
	.w2(32'h3c179811),
	.w3(32'h3b9f6ee1),
	.w4(32'hbc31cee5),
	.w5(32'hbba8af07),
	.w6(32'hbc1e9dea),
	.w7(32'hbc2c5796),
	.w8(32'hbc08fb04),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8402cf),
	.w1(32'h3a8340d1),
	.w2(32'h3be20435),
	.w3(32'hbbc884d2),
	.w4(32'hbbdb251d),
	.w5(32'hbb49de8c),
	.w6(32'h3b40b536),
	.w7(32'hba45a4ab),
	.w8(32'h3a86ca92),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49dd46),
	.w1(32'hbac476b4),
	.w2(32'hbb8eefe7),
	.w3(32'hbb23a1ca),
	.w4(32'h3bdc6536),
	.w5(32'hbc18a3bc),
	.w6(32'hbb23d0c8),
	.w7(32'h3bb23921),
	.w8(32'h3c26d236),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3cd9),
	.w1(32'h3b4866b0),
	.w2(32'h3c1adf27),
	.w3(32'hbc866002),
	.w4(32'hbab8cd81),
	.w5(32'h3c8a2517),
	.w6(32'h3bd7d654),
	.w7(32'h3b1adec4),
	.w8(32'h3c400f83),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6be7e6),
	.w1(32'h3b2f878e),
	.w2(32'h3ba1d49c),
	.w3(32'h3b8d1b49),
	.w4(32'hbbdf3388),
	.w5(32'hbbd15e74),
	.w6(32'h3b136f06),
	.w7(32'h3c1eff26),
	.w8(32'h3bbc3da0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80938b),
	.w1(32'hbb17c927),
	.w2(32'h3c98de83),
	.w3(32'hbc1ebbb1),
	.w4(32'h3cc70b70),
	.w5(32'h3cd70230),
	.w6(32'hbbb8cb08),
	.w7(32'h3c31bd1b),
	.w8(32'h3cd311f8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c889b16),
	.w1(32'h3c059a77),
	.w2(32'h3ab6d579),
	.w3(32'h3c330339),
	.w4(32'hb9c4d547),
	.w5(32'hbb59c15b),
	.w6(32'h3c41da30),
	.w7(32'h3ae22ac3),
	.w8(32'hba9fe7a1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52c99b),
	.w1(32'hba805998),
	.w2(32'h3bcc452c),
	.w3(32'hbbd50cfd),
	.w4(32'hbbd07882),
	.w5(32'h3ad1cbfb),
	.w6(32'hbbd7f369),
	.w7(32'hba8df730),
	.w8(32'hbb88c768),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda374b),
	.w1(32'hbb9f1c3d),
	.w2(32'h3bd7099b),
	.w3(32'h3be60121),
	.w4(32'h3bc18563),
	.w5(32'h3abde2f5),
	.w6(32'h3af10e20),
	.w7(32'hbb723a41),
	.w8(32'hbb98a0b5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7cbc8),
	.w1(32'hbb8f6406),
	.w2(32'hbb6454fe),
	.w3(32'hbaf8d077),
	.w4(32'hbaf71af0),
	.w5(32'hba8fbb22),
	.w6(32'hbb6d95d3),
	.w7(32'hbba69cb6),
	.w8(32'hbb19cfa1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c5e06),
	.w1(32'h3be7a747),
	.w2(32'h3c501905),
	.w3(32'hbab63902),
	.w4(32'hba95d2b2),
	.w5(32'h3c1769e8),
	.w6(32'hbc06f65e),
	.w7(32'hbc3a51ef),
	.w8(32'hbbaa7c2d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8668d8d),
	.w1(32'hbc135882),
	.w2(32'h3b31c228),
	.w3(32'h3c018322),
	.w4(32'hbb98e63e),
	.w5(32'hbbbaa0d8),
	.w6(32'hbbd303b7),
	.w7(32'hbb73f596),
	.w8(32'hbbbce408),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0557ec),
	.w1(32'hbbc7ac82),
	.w2(32'h3b8f9f74),
	.w3(32'hbbc04a57),
	.w4(32'hbbf620d9),
	.w5(32'hbbdeaf7a),
	.w6(32'hbbcef578),
	.w7(32'h3bdee360),
	.w8(32'hbb0944e0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e8106),
	.w1(32'h3a774260),
	.w2(32'h3c14ec83),
	.w3(32'hbacb30b6),
	.w4(32'h3b771bbc),
	.w5(32'h3bc8beb4),
	.w6(32'hba7dad4d),
	.w7(32'hba3c2e52),
	.w8(32'h3bc7beec),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8834a),
	.w1(32'hbb0de50b),
	.w2(32'h3b129a6b),
	.w3(32'hbb537897),
	.w4(32'hbbd1b0cb),
	.w5(32'h3b5bf042),
	.w6(32'hbbea8c92),
	.w7(32'hbc0f930b),
	.w8(32'hbb3d6c2e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0c695),
	.w1(32'hbc1893e0),
	.w2(32'h3bf977d1),
	.w3(32'hbb841a2d),
	.w4(32'hbbf020fc),
	.w5(32'h3b270a07),
	.w6(32'hbb5a5235),
	.w7(32'hbb79c2c3),
	.w8(32'hbad8f1a1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba921163),
	.w1(32'hbb911698),
	.w2(32'h3b028b58),
	.w3(32'hb9257c57),
	.w4(32'h3a4a444f),
	.w5(32'h3b8641c2),
	.w6(32'h3b7d38bf),
	.w7(32'h3aa7056f),
	.w8(32'hbaca38b1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89ebb8),
	.w1(32'hbc31e51e),
	.w2(32'h3a8ddedd),
	.w3(32'hbbce316d),
	.w4(32'hbc7aeac9),
	.w5(32'hbc4b05c3),
	.w6(32'hbc85868b),
	.w7(32'hbccf77cf),
	.w8(32'hbcf9e403),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2d380),
	.w1(32'hbc27d511),
	.w2(32'h3bd82489),
	.w3(32'h392d69fe),
	.w4(32'hbb916afb),
	.w5(32'h38d3bbbf),
	.w6(32'hbacdb8e6),
	.w7(32'h3b294bef),
	.w8(32'hbc0eda5e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92827e),
	.w1(32'hbb8ff287),
	.w2(32'h3beb3475),
	.w3(32'hba41cb04),
	.w4(32'h3be842c6),
	.w5(32'h3b4fea81),
	.w6(32'hbbb3ecf7),
	.w7(32'h3a78c546),
	.w8(32'hb96462b0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb8a1),
	.w1(32'hbbc7547a),
	.w2(32'hba550d2b),
	.w3(32'hbadf996e),
	.w4(32'hbb876a80),
	.w5(32'hbb7fb965),
	.w6(32'hbb07e90b),
	.w7(32'hbad3c414),
	.w8(32'hbb9c6bc5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993324a),
	.w1(32'h3beafaf6),
	.w2(32'h3c75a77d),
	.w3(32'hbc138bdd),
	.w4(32'h3a828047),
	.w5(32'h3c999420),
	.w6(32'h3a7e6c15),
	.w7(32'h3c41b2d7),
	.w8(32'h3b118f97),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb900820),
	.w1(32'h3b824b2a),
	.w2(32'h3b9d4041),
	.w3(32'h3c8c8ac5),
	.w4(32'h3c1ccb79),
	.w5(32'h3be2eab9),
	.w6(32'h3c8035f9),
	.w7(32'h3c787929),
	.w8(32'h3c86db92),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2f68a),
	.w1(32'h3c51ce36),
	.w2(32'h3bfaa974),
	.w3(32'h3b75a76e),
	.w4(32'h3b73e157),
	.w5(32'h3b90ef66),
	.w6(32'h38e229b0),
	.w7(32'h3b2c1572),
	.w8(32'h3b3f4c12),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c38f5c),
	.w1(32'hbb0249e5),
	.w2(32'hbb100468),
	.w3(32'h3b0ae036),
	.w4(32'hba438b23),
	.w5(32'hba8b3f3a),
	.w6(32'h3b88df07),
	.w7(32'hb8114b32),
	.w8(32'h3b7595d2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8c73e),
	.w1(32'h3ae50635),
	.w2(32'h3a97b09e),
	.w3(32'hbc2ca2ef),
	.w4(32'hbc1b6d5d),
	.w5(32'hbbce31f9),
	.w6(32'hbbf41f04),
	.w7(32'hbc2ffe7d),
	.w8(32'hbc2f8064),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe340ac),
	.w1(32'h3aa14aca),
	.w2(32'h3bc0197f),
	.w3(32'h3b94e5c0),
	.w4(32'h3bc12d6f),
	.w5(32'h3c205569),
	.w6(32'hbb4347a2),
	.w7(32'h3b8498b7),
	.w8(32'h3be81b5a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870d32),
	.w1(32'h3bcb9245),
	.w2(32'hbb5b4e5b),
	.w3(32'h3bcdc903),
	.w4(32'h3b94c5f8),
	.w5(32'hbb8c939f),
	.w6(32'h3b1147fa),
	.w7(32'h3bb8539d),
	.w8(32'hbaebf942),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bd025),
	.w1(32'hbc5b90ba),
	.w2(32'hbbcbe061),
	.w3(32'h3bb6edbc),
	.w4(32'hbca4ddf9),
	.w5(32'h3cd61a2c),
	.w6(32'hbb1f6db4),
	.w7(32'hbc865d40),
	.w8(32'hb8bc0dad),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb23f62),
	.w1(32'hbb8d0cef),
	.w2(32'hbc0f9aea),
	.w3(32'hbb645be8),
	.w4(32'hbc2a74df),
	.w5(32'hbc393ec1),
	.w6(32'hba8a963a),
	.w7(32'hbc98cac8),
	.w8(32'h3b8caf6f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd3edf6),
	.w1(32'h3c404754),
	.w2(32'h3c643869),
	.w3(32'hbc0d1846),
	.w4(32'hbb41e4af),
	.w5(32'hbc33d983),
	.w6(32'hbd0336fc),
	.w7(32'hbb5f7d76),
	.w8(32'hbcf0167e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeaec4),
	.w1(32'h3ca62c52),
	.w2(32'h3cf83d79),
	.w3(32'h3c893dc1),
	.w4(32'h3c5706b2),
	.w5(32'h3d03c390),
	.w6(32'hbcd20b92),
	.w7(32'hbac75ad2),
	.w8(32'hbb57f088),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd58424),
	.w1(32'h3c1f0c56),
	.w2(32'h3cf7bcbd),
	.w3(32'hbc5891bf),
	.w4(32'hbc529d11),
	.w5(32'hbc5de576),
	.w6(32'hbcdac019),
	.w7(32'hb8e7694b),
	.w8(32'hbd210958),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f9bac),
	.w1(32'hbb36f76b),
	.w2(32'h3c28766d),
	.w3(32'h3b881e94),
	.w4(32'hbcbcc633),
	.w5(32'h3bd2a268),
	.w6(32'h3c9a4ec0),
	.w7(32'hbcb39806),
	.w8(32'hbbb45f7b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcde02f7),
	.w1(32'h3c206970),
	.w2(32'h3986cd45),
	.w3(32'h3b91b45f),
	.w4(32'h3bd8d7b2),
	.w5(32'hbbe05917),
	.w6(32'h3c05230a),
	.w7(32'h3c43ed92),
	.w8(32'hbc261f18),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ff85f),
	.w1(32'h3b057f42),
	.w2(32'hbbc0e26a),
	.w3(32'hbc3381f5),
	.w4(32'h398acf23),
	.w5(32'hbbf32b37),
	.w6(32'hbc07988e),
	.w7(32'hba853734),
	.w8(32'h3be57c2b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1b968),
	.w1(32'h3b723a99),
	.w2(32'h3b0f6688),
	.w3(32'h3bc090e6),
	.w4(32'h3c125f5c),
	.w5(32'h3ab8064d),
	.w6(32'h3c308067),
	.w7(32'h3ba82423),
	.w8(32'h3a8b8531),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2c228),
	.w1(32'hbc302d80),
	.w2(32'h3c4bdf6e),
	.w3(32'hbb909cc9),
	.w4(32'h3bf93a07),
	.w5(32'hbaaaf071),
	.w6(32'hbbc0a82f),
	.w7(32'hbab97d6b),
	.w8(32'h3c6d32cd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2fbf6),
	.w1(32'hbb822930),
	.w2(32'hbb887c49),
	.w3(32'hbc73dde2),
	.w4(32'hbb67a50f),
	.w5(32'hbc07b3a4),
	.w6(32'h3c0c7dbe),
	.w7(32'hb9442d39),
	.w8(32'h39c91394),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7a4c5),
	.w1(32'hba94658b),
	.w2(32'h3b19a737),
	.w3(32'h3ba5963d),
	.w4(32'h394a5555),
	.w5(32'h3cdb3d71),
	.w6(32'hbb15846f),
	.w7(32'hbaa9f5d5),
	.w8(32'hbafe43af),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd3dc6),
	.w1(32'hbc658da7),
	.w2(32'h3bde21ad),
	.w3(32'hbc251058),
	.w4(32'hbc477ac6),
	.w5(32'hba727d3f),
	.w6(32'hba65cd7f),
	.w7(32'h3a1ce75e),
	.w8(32'hbc7b7d12),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84b6c0),
	.w1(32'hbc0d7324),
	.w2(32'h3c1b9d9c),
	.w3(32'hbc7050ec),
	.w4(32'hba9d3425),
	.w5(32'hbd0d817a),
	.w6(32'hbc32cb79),
	.w7(32'hb92333bb),
	.w8(32'hbb65a35c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1def5a),
	.w1(32'hbd06e7e1),
	.w2(32'h3b41f4fe),
	.w3(32'h3cef2dae),
	.w4(32'h3c05f390),
	.w5(32'h3bd695dc),
	.w6(32'h3c8fc041),
	.w7(32'h3b816a30),
	.w8(32'h3b9a91a1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79fc6e),
	.w1(32'hbb264ce6),
	.w2(32'hbc2117e1),
	.w3(32'hbbc3eb0c),
	.w4(32'hba0de137),
	.w5(32'h3b3c61ee),
	.w6(32'hbb9e3778),
	.w7(32'h3b960c71),
	.w8(32'hbc789a9d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89227d),
	.w1(32'hbb32ed63),
	.w2(32'hbb9fb7d7),
	.w3(32'h3b052ba0),
	.w4(32'hbc44473b),
	.w5(32'hbc0e5f5b),
	.w6(32'h3c1553ff),
	.w7(32'hbc6ca2bc),
	.w8(32'h3b07d3f3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c0592),
	.w1(32'h3cf4463f),
	.w2(32'h3c596e22),
	.w3(32'h3ca814d1),
	.w4(32'hbc4ed51b),
	.w5(32'hbc800823),
	.w6(32'h3ca1427c),
	.w7(32'hbb51b03a),
	.w8(32'hbc6e3ef3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ef467),
	.w1(32'h3cb0a93a),
	.w2(32'h3b138a5b),
	.w3(32'h3c62a206),
	.w4(32'h3c1e7448),
	.w5(32'hbbf819d9),
	.w6(32'h3d26c7bb),
	.w7(32'h3b95cefa),
	.w8(32'hbc59cbbb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5236a),
	.w1(32'h3b4079ca),
	.w2(32'h39812795),
	.w3(32'h3a97ec8f),
	.w4(32'h3c5652c5),
	.w5(32'hbcde996e),
	.w6(32'h3b810bb6),
	.w7(32'h3caa02a3),
	.w8(32'h3cdfe67f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b619d),
	.w1(32'h3b4a9a6f),
	.w2(32'h3b8d6773),
	.w3(32'hbce54c6f),
	.w4(32'h3a991598),
	.w5(32'hbb91fb2f),
	.w6(32'hbc919265),
	.w7(32'h3a18eb04),
	.w8(32'hbacb35d5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1286db),
	.w1(32'h3c1d6a04),
	.w2(32'h3affdc4f),
	.w3(32'h3b942784),
	.w4(32'h3af0773b),
	.w5(32'h3c99b7e5),
	.w6(32'hbc23dc27),
	.w7(32'h3ba75320),
	.w8(32'h3c9d1378),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb117d6f),
	.w1(32'h3c9884dc),
	.w2(32'hba809e2f),
	.w3(32'h3c07f859),
	.w4(32'hbc840656),
	.w5(32'hbbe10e99),
	.w6(32'h3ca9e52c),
	.w7(32'hbb89dc28),
	.w8(32'hbbdf5a78),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4751f9),
	.w1(32'h3cf357d8),
	.w2(32'hbbc17627),
	.w3(32'hbcacf8ad),
	.w4(32'hbb6dce71),
	.w5(32'hbab69c72),
	.w6(32'h3d028228),
	.w7(32'hba70204e),
	.w8(32'h3b35017d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b8c71),
	.w1(32'hbb2c66a3),
	.w2(32'hba1076f1),
	.w3(32'h3b99cbf2),
	.w4(32'h3c337712),
	.w5(32'hbbffa000),
	.w6(32'h3b1da9e8),
	.w7(32'h3c77231f),
	.w8(32'hbc8ed49e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdce6ea),
	.w1(32'hbba868c0),
	.w2(32'h3bb5c23a),
	.w3(32'h3c3fca54),
	.w4(32'h3c7aced2),
	.w5(32'hbcfa1aef),
	.w6(32'hbcb375af),
	.w7(32'h3b3bf7ce),
	.w8(32'h3bb92582),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2baba),
	.w1(32'hbbf35fc5),
	.w2(32'h39bdf3e6),
	.w3(32'h3b82f4ad),
	.w4(32'hbc28bf62),
	.w5(32'hbc99a6d8),
	.w6(32'hbd117e6a),
	.w7(32'hbc1ed6db),
	.w8(32'hbb99c833),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21ae4a),
	.w1(32'h3c6c6440),
	.w2(32'hbb1f7e96),
	.w3(32'hba00d5dc),
	.w4(32'hba0931fc),
	.w5(32'hbaceacd0),
	.w6(32'h3d03f244),
	.w7(32'hba486f58),
	.w8(32'h3c0e3ea5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23fbc8),
	.w1(32'h3b88f689),
	.w2(32'h3ae5fa43),
	.w3(32'h38b41739),
	.w4(32'hbc21ee07),
	.w5(32'h3a00bb6a),
	.w6(32'h3b412e58),
	.w7(32'hbb4f461b),
	.w8(32'hbad494d2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38a0da),
	.w1(32'h3ad2223c),
	.w2(32'hbbc99480),
	.w3(32'hbbb9ac12),
	.w4(32'h3bcec71e),
	.w5(32'hbb917748),
	.w6(32'hba925b5d),
	.w7(32'h3c8593e4),
	.w8(32'h3d407bc0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b268a),
	.w1(32'hbb0f3715),
	.w2(32'h3c2a9638),
	.w3(32'hbc900ec0),
	.w4(32'h3c04f1d9),
	.w5(32'hbafc1488),
	.w6(32'hbd1de8c6),
	.w7(32'hbab1c2f9),
	.w8(32'hbb3ef84f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a1777),
	.w1(32'h3b9464ed),
	.w2(32'h3c119d90),
	.w3(32'h3c22509f),
	.w4(32'hbc2eab72),
	.w5(32'h3ca2ece9),
	.w6(32'hbc1e5898),
	.w7(32'hba3e8054),
	.w8(32'h3d04eecf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc843e2),
	.w1(32'h3c101e4d),
	.w2(32'hbc4043ec),
	.w3(32'h3b4dfa68),
	.w4(32'hbb0a7782),
	.w5(32'hbc24c054),
	.w6(32'h3cc1c0fd),
	.w7(32'hbb46d093),
	.w8(32'hbb2f2db3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf29d0),
	.w1(32'hbae10d89),
	.w2(32'hbcc66e2c),
	.w3(32'h3bbd3ed9),
	.w4(32'hbc9a34f4),
	.w5(32'hbc8b9229),
	.w6(32'hbb5b1dc9),
	.w7(32'hbc70d9cb),
	.w8(32'hbc6bb48d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9bfb0),
	.w1(32'hbc049baa),
	.w2(32'h39bc4889),
	.w3(32'hbbad2277),
	.w4(32'h3b7b1254),
	.w5(32'h3c69d3ad),
	.w6(32'hbc024365),
	.w7(32'h3c738f13),
	.w8(32'h3c724f46),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0cd73),
	.w1(32'hbc804c80),
	.w2(32'h3af054b2),
	.w3(32'hbcc3e6e0),
	.w4(32'hbc3d39c1),
	.w5(32'h3c8aedd8),
	.w6(32'hbcf4b757),
	.w7(32'hbbf6d959),
	.w8(32'h3c3f9483),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7a553),
	.w1(32'hbc0b337b),
	.w2(32'hba92ab6f),
	.w3(32'h3d08ab56),
	.w4(32'h3b24e240),
	.w5(32'h3be59cc9),
	.w6(32'h3c877af8),
	.w7(32'h3b538b82),
	.w8(32'hbc7394f8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cff66),
	.w1(32'hbc4f157b),
	.w2(32'hbb9f2bf1),
	.w3(32'h3bf73348),
	.w4(32'hbb48612b),
	.w5(32'hba9b5f0d),
	.w6(32'hbab77928),
	.w7(32'hbbdaadb5),
	.w8(32'hbae8305d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf4962),
	.w1(32'h3adaafeb),
	.w2(32'hbb0acc13),
	.w3(32'hbaf4fc35),
	.w4(32'hbc1c976b),
	.w5(32'hbb195f84),
	.w6(32'hbb8c92ad),
	.w7(32'hbb1bd96d),
	.w8(32'hbc9e80cd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5ecb0),
	.w1(32'hbc494309),
	.w2(32'hbbb06107),
	.w3(32'h3c1615cc),
	.w4(32'hbbf06ec4),
	.w5(32'h3c4810e9),
	.w6(32'hbb13c4b9),
	.w7(32'h3b0d935d),
	.w8(32'hbc66a8c2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96b149),
	.w1(32'h3b8cdb5d),
	.w2(32'h3c483fdb),
	.w3(32'hbbe610f5),
	.w4(32'h3bd03c4a),
	.w5(32'hba1a22d8),
	.w6(32'h3b45340b),
	.w7(32'h3bcf3863),
	.w8(32'h3bbde7cf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5e626),
	.w1(32'h3c73d90b),
	.w2(32'h3ca56809),
	.w3(32'hba75cbad),
	.w4(32'h3a6a69b4),
	.w5(32'h3c371f91),
	.w6(32'h3b8e957b),
	.w7(32'hbb148d85),
	.w8(32'h3cd239c9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c932358),
	.w1(32'hbc0e0cfb),
	.w2(32'hbb96619c),
	.w3(32'hbcc56bc8),
	.w4(32'hb9ed4d89),
	.w5(32'hba911b08),
	.w6(32'hbb2581ae),
	.w7(32'hbb083b41),
	.w8(32'h3bd27dab),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77c0f),
	.w1(32'h3b0853ca),
	.w2(32'hbb9527a9),
	.w3(32'hbb00b503),
	.w4(32'h3b768657),
	.w5(32'hb8970ea7),
	.w6(32'hb9c24c49),
	.w7(32'h3ade503c),
	.w8(32'hbb9ec0a4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c2818),
	.w1(32'h3c025a40),
	.w2(32'h3ba2cb51),
	.w3(32'hbc16c140),
	.w4(32'h3c295165),
	.w5(32'hbcd89670),
	.w6(32'hbb21cb0f),
	.w7(32'h3c1f0787),
	.w8(32'h3cf5d0c9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf5209f),
	.w1(32'hbd1e872c),
	.w2(32'h39f5d314),
	.w3(32'hbbb286ca),
	.w4(32'hbc094cbd),
	.w5(32'hbb454b85),
	.w6(32'hbd202ab7),
	.w7(32'hbb3ef132),
	.w8(32'h3b82090e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f4982),
	.w1(32'h3c00e9d8),
	.w2(32'h3c09f133),
	.w3(32'h3c5ed576),
	.w4(32'hbc9b8395),
	.w5(32'h3b58b3eb),
	.w6(32'h3c9a2a7d),
	.w7(32'h3c1254f6),
	.w8(32'hbc2cc14b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3a0ca),
	.w1(32'hbc3d5870),
	.w2(32'hba6ed167),
	.w3(32'h3c71d030),
	.w4(32'h3b17ba4a),
	.w5(32'hbba7adbf),
	.w6(32'h3cc4cb86),
	.w7(32'h3b6d6e2f),
	.w8(32'hbbcf16f6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule