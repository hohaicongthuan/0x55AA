module layer_10_featuremap_224(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2acca),
	.w1(32'hbbc75554),
	.w2(32'h3b023fe3),
	.w3(32'hbc009566),
	.w4(32'hba90608a),
	.w5(32'hbc182aab),
	.w6(32'h3a29150b),
	.w7(32'h3b400227),
	.w8(32'hbbf9e6c6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af748f7),
	.w1(32'h3b23da43),
	.w2(32'hbbdd95d4),
	.w3(32'hbc0301a6),
	.w4(32'h3a7d7f43),
	.w5(32'hbbc46e1a),
	.w6(32'h3c1e49b8),
	.w7(32'hbbbfcde2),
	.w8(32'hb9443939),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0acab3),
	.w1(32'h38ba5997),
	.w2(32'hbad2cab9),
	.w3(32'hbb05d0c0),
	.w4(32'hbbdccbff),
	.w5(32'hbbd24ae1),
	.w6(32'h392c16bf),
	.w7(32'h3cc0669a),
	.w8(32'h3c015b82),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01b7b),
	.w1(32'hbc36b355),
	.w2(32'hbab7f027),
	.w3(32'h3c24c998),
	.w4(32'h3ca591b7),
	.w5(32'hbc4901a5),
	.w6(32'hbc0a1c10),
	.w7(32'hbc06703a),
	.w8(32'h3a8a6e03),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ca32b),
	.w1(32'hbb8fed5e),
	.w2(32'h3b91b809),
	.w3(32'hbb5748e5),
	.w4(32'h3c027e05),
	.w5(32'hba6ae5db),
	.w6(32'hbc369824),
	.w7(32'hbbc9355d),
	.w8(32'hbba8d480),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc7a36),
	.w1(32'hbad86534),
	.w2(32'h3b836eab),
	.w3(32'hbc3830fc),
	.w4(32'h3ad5e5d6),
	.w5(32'h3c0941f8),
	.w6(32'hbb9882d2),
	.w7(32'hbbebb144),
	.w8(32'hbc7beb0d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b460397),
	.w1(32'hbc83f211),
	.w2(32'hbc177c4f),
	.w3(32'h3c850748),
	.w4(32'hbb159a30),
	.w5(32'hbb92f6ce),
	.w6(32'hbb4f9d79),
	.w7(32'hbbe87148),
	.w8(32'hbb9624f9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38e2a4),
	.w1(32'hbb980544),
	.w2(32'h3b440780),
	.w3(32'hba9744e3),
	.w4(32'h3b63055f),
	.w5(32'hbb539f74),
	.w6(32'h3bc67ac4),
	.w7(32'hbb933439),
	.w8(32'hbb005368),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0eca6),
	.w1(32'h3bc189db),
	.w2(32'h3b4d75ca),
	.w3(32'hbbc7e691),
	.w4(32'hbc91cc42),
	.w5(32'hbc124a96),
	.w6(32'h3cb1531e),
	.w7(32'hbbc2be9e),
	.w8(32'hba6ab195),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75e9fe),
	.w1(32'h394006dd),
	.w2(32'hbc73201d),
	.w3(32'hbb88b39f),
	.w4(32'h3b83b6e5),
	.w5(32'hbb4b9a8e),
	.w6(32'h3b3cbb1a),
	.w7(32'h3b065622),
	.w8(32'h3aaa7750),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c115070),
	.w1(32'h3b884b1b),
	.w2(32'hbafa9fbf),
	.w3(32'hbc105c5b),
	.w4(32'hbb2219e3),
	.w5(32'h3b7f7a18),
	.w6(32'h3c159df3),
	.w7(32'hbb8f6fe0),
	.w8(32'h3b5be0c4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caaa63),
	.w1(32'hbb2d569d),
	.w2(32'hbbbb7cd9),
	.w3(32'hbadc8e38),
	.w4(32'hba887497),
	.w5(32'h39066d05),
	.w6(32'hbb08738d),
	.w7(32'h3805eb3e),
	.w8(32'h3c2e17eb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89e2e3),
	.w1(32'h3b1e441e),
	.w2(32'h3c24cf5e),
	.w3(32'hbb50f19e),
	.w4(32'hbbccac51),
	.w5(32'h3b46bc84),
	.w6(32'hbc0a29e3),
	.w7(32'hbb990e22),
	.w8(32'hbb0af6d6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58e244),
	.w1(32'h3bb84e2a),
	.w2(32'hbc9982e6),
	.w3(32'hbbd15e03),
	.w4(32'h3c0ed9c6),
	.w5(32'hbb7fd8b5),
	.w6(32'h3bc4e3d3),
	.w7(32'h3b4b611f),
	.w8(32'h3a58da39),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95d9f0),
	.w1(32'h3a940b3f),
	.w2(32'hbbe8a12c),
	.w3(32'hbb2325fd),
	.w4(32'hbbc03503),
	.w5(32'h3aee637b),
	.w6(32'h39d1f234),
	.w7(32'hbbc3a80b),
	.w8(32'h36cfb36a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5477a5),
	.w1(32'hbb5afc02),
	.w2(32'hba966d77),
	.w3(32'hbb35189d),
	.w4(32'h3a12c376),
	.w5(32'hbaebb63b),
	.w6(32'hbc769807),
	.w7(32'h3c248754),
	.w8(32'hbc063bc7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b4011),
	.w1(32'h3ad864f6),
	.w2(32'hbc6d5759),
	.w3(32'hb912faeb),
	.w4(32'h384f0a12),
	.w5(32'h3b5ed3b7),
	.w6(32'hbb33e387),
	.w7(32'hbc22c41a),
	.w8(32'hbb840af3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a033c),
	.w1(32'hba54960c),
	.w2(32'hbb9bed42),
	.w3(32'h3c6b4155),
	.w4(32'hba3d2498),
	.w5(32'hb923e57f),
	.w6(32'hbbcd38fa),
	.w7(32'hba6b102a),
	.w8(32'hba046a98),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2126e),
	.w1(32'h3b9b53ae),
	.w2(32'h3b951219),
	.w3(32'hbc4557b3),
	.w4(32'hbbabe4fa),
	.w5(32'hbc1e667f),
	.w6(32'h3c19c469),
	.w7(32'h3c885330),
	.w8(32'hba4d7e5a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb00200),
	.w1(32'h3c9456af),
	.w2(32'h3b94a865),
	.w3(32'h3ae04296),
	.w4(32'hb9ca3bb9),
	.w5(32'hbb480cb6),
	.w6(32'h3c2fdef8),
	.w7(32'hbaa8c191),
	.w8(32'hbb1b7336),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f813),
	.w1(32'h3b6858e2),
	.w2(32'hba97367c),
	.w3(32'h3cf0f638),
	.w4(32'h3bf7a444),
	.w5(32'h3a5535f3),
	.w6(32'hbb2b5e2d),
	.w7(32'h3af54723),
	.w8(32'h3abe5f49),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c176364),
	.w1(32'h3c381642),
	.w2(32'h3b836cd3),
	.w3(32'hba4d27fe),
	.w4(32'hbb60cf4e),
	.w5(32'h3bb24636),
	.w6(32'hbb0063c8),
	.w7(32'hb981f1f8),
	.w8(32'hbb11980d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ff9ab),
	.w1(32'hb9fce953),
	.w2(32'h3c11ccf9),
	.w3(32'hbae88a0f),
	.w4(32'h3a6749c7),
	.w5(32'h3bbe137d),
	.w6(32'hba71c696),
	.w7(32'h38e3dab4),
	.w8(32'hbab21d8f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f81db),
	.w1(32'hbb2cfa13),
	.w2(32'h3c072479),
	.w3(32'h3b9c41f3),
	.w4(32'hbab333c9),
	.w5(32'h3c50dbb3),
	.w6(32'h3ab7b86b),
	.w7(32'h3813c4b3),
	.w8(32'hb95659b7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c70f5),
	.w1(32'hbbd9eded),
	.w2(32'hbb51cd50),
	.w3(32'h3bc304c4),
	.w4(32'h3b093fdf),
	.w5(32'h3a4a112d),
	.w6(32'hbc328421),
	.w7(32'h3b274b8a),
	.w8(32'hbb96d114),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f8dbb),
	.w1(32'h3b0da6e4),
	.w2(32'hbc1c283d),
	.w3(32'h3c525f20),
	.w4(32'hb9edc3cd),
	.w5(32'hbbf7eb70),
	.w6(32'hbaa24ce3),
	.w7(32'hbace41a0),
	.w8(32'h390dc9fd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61b113),
	.w1(32'hbb9be6f9),
	.w2(32'h3c843f63),
	.w3(32'hbc8d8957),
	.w4(32'hbb24e9c4),
	.w5(32'hbb119161),
	.w6(32'hbc3ee89f),
	.w7(32'hbb563ffa),
	.w8(32'hbb5f5c1f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85281d),
	.w1(32'h3b416e7a),
	.w2(32'hbbcc4a09),
	.w3(32'hba6b4a3b),
	.w4(32'h3a8d371a),
	.w5(32'hbbde8c26),
	.w6(32'h39db2210),
	.w7(32'hbb34ef27),
	.w8(32'h3a8c11f2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c103322),
	.w1(32'h3b913886),
	.w2(32'hbc02b3f5),
	.w3(32'hba40e111),
	.w4(32'hb9536754),
	.w5(32'h39bd41d7),
	.w6(32'h3ab5fa01),
	.w7(32'hbac36790),
	.w8(32'hba6afd1b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfeea61),
	.w1(32'hbb05d7d8),
	.w2(32'hbc3db847),
	.w3(32'hb9b7f48e),
	.w4(32'hbabd5a19),
	.w5(32'hbc0ab819),
	.w6(32'hba97b7f3),
	.w7(32'hbbba96d0),
	.w8(32'h3b365521),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053021),
	.w1(32'hbbcf90a5),
	.w2(32'h3adc1bde),
	.w3(32'hbba95d62),
	.w4(32'h3cf2c396),
	.w5(32'h3bc94c07),
	.w6(32'h3a8304f2),
	.w7(32'hbb9c0490),
	.w8(32'hbbbc73a6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b21a1),
	.w1(32'h3bd8355c),
	.w2(32'hbb5f2bf9),
	.w3(32'h3baa8993),
	.w4(32'hbaf8ee21),
	.w5(32'h3b53b833),
	.w6(32'hbb28f838),
	.w7(32'hbc86c18e),
	.w8(32'hbc305766),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1fcd4),
	.w1(32'hbb1c96a2),
	.w2(32'hbb0dc7f9),
	.w3(32'h3aee3805),
	.w4(32'hbc179e63),
	.w5(32'hbb35ca40),
	.w6(32'h3abee3cf),
	.w7(32'hbb8d8aab),
	.w8(32'h3c2a3910),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be473),
	.w1(32'h3c05eecc),
	.w2(32'h3bf1456c),
	.w3(32'h3bdca68f),
	.w4(32'h3ce2e282),
	.w5(32'h3ad3347f),
	.w6(32'hbab57b68),
	.w7(32'h3c370efe),
	.w8(32'h3adbd473),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fef98),
	.w1(32'h3b64bf84),
	.w2(32'h3ad91b91),
	.w3(32'h3b8946e1),
	.w4(32'h3b115e3a),
	.w5(32'hbc843fb3),
	.w6(32'h3c9cb10a),
	.w7(32'hbc2e1ee1),
	.w8(32'h3c29a938),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b861e5d),
	.w1(32'hbbb2098e),
	.w2(32'h3bce79bf),
	.w3(32'h3c2f0916),
	.w4(32'h3a476e16),
	.w5(32'h3a98c467),
	.w6(32'h3b9e5cfd),
	.w7(32'hbb529f13),
	.w8(32'h3ada0cb7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ed33),
	.w1(32'h39629a89),
	.w2(32'hbc13f403),
	.w3(32'h3b8c0dad),
	.w4(32'hbba84a73),
	.w5(32'h3b44a801),
	.w6(32'h3b8887de),
	.w7(32'hbb96fc99),
	.w8(32'hbc64e1f5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28a8e4),
	.w1(32'h3a812d20),
	.w2(32'hbb6e3a4f),
	.w3(32'h3c137fd5),
	.w4(32'hbbbd3a98),
	.w5(32'hb66dc61d),
	.w6(32'hba6b26b9),
	.w7(32'h3c5173b9),
	.w8(32'hbbff7fe2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacdd87),
	.w1(32'hbb37ac4c),
	.w2(32'h39fcb550),
	.w3(32'hbbb2f028),
	.w4(32'hbb3858de),
	.w5(32'hbbcacefc),
	.w6(32'h3bb700b7),
	.w7(32'hbc334106),
	.w8(32'hbbe781d7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ac203),
	.w1(32'hb95276ea),
	.w2(32'hbb2c2f27),
	.w3(32'hbb8522ab),
	.w4(32'h3b93b8a9),
	.w5(32'hbbbb7746),
	.w6(32'h39d324c5),
	.w7(32'h3aa1c782),
	.w8(32'h3be59c50),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89ff1d6),
	.w1(32'h3c73d8b1),
	.w2(32'hba868f1f),
	.w3(32'hbc12f8f9),
	.w4(32'hbc3e3c7d),
	.w5(32'h3b8069cb),
	.w6(32'hb8e64bbe),
	.w7(32'hbba3c099),
	.w8(32'hba17807d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c87c8d),
	.w1(32'hbbb9aa29),
	.w2(32'hbc72551b),
	.w3(32'hba8542f6),
	.w4(32'h3b071a7f),
	.w5(32'h3c06dfc3),
	.w6(32'h3bc5d694),
	.w7(32'h3bcc1132),
	.w8(32'h3b65be62),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae68022),
	.w1(32'hba62fbdb),
	.w2(32'hba4cc4e1),
	.w3(32'hbc0852c7),
	.w4(32'hbbc19d81),
	.w5(32'hbbac0d42),
	.w6(32'hbb08a0ef),
	.w7(32'hbbbaea38),
	.w8(32'hbb91bc97),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5c082),
	.w1(32'h3b465de0),
	.w2(32'hbb0fbf60),
	.w3(32'h3aaff28c),
	.w4(32'hbabdca2c),
	.w5(32'hb9e06ca9),
	.w6(32'hbb086653),
	.w7(32'hba884819),
	.w8(32'hbb099ee4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04b9dc),
	.w1(32'hbaca9bd6),
	.w2(32'hbb9f6eb2),
	.w3(32'h3b421779),
	.w4(32'hbb03ad89),
	.w5(32'hbc1d63ab),
	.w6(32'h3a8929fa),
	.w7(32'hbb436d35),
	.w8(32'hb84ba5f5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4803a7),
	.w1(32'h3ab1093a),
	.w2(32'hbc307b6a),
	.w3(32'h3cd809bc),
	.w4(32'h3c040354),
	.w5(32'hbb36fd4d),
	.w6(32'h3b2715fe),
	.w7(32'hbb62b701),
	.w8(32'h39d8a85d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb596ea),
	.w1(32'h3b50a299),
	.w2(32'hbca2a004),
	.w3(32'hbbc07c6b),
	.w4(32'hbb47707e),
	.w5(32'h3aa1fcd1),
	.w6(32'hb86adc46),
	.w7(32'h3bcd3669),
	.w8(32'hbbc10837),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a498c51),
	.w1(32'h3c0be3d4),
	.w2(32'hbc326565),
	.w3(32'hbb3f1e39),
	.w4(32'hba238881),
	.w5(32'hbb3e81ad),
	.w6(32'h3c84c156),
	.w7(32'hbb8ea9ed),
	.w8(32'hbb8ad867),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb496bba),
	.w1(32'h3bbcb186),
	.w2(32'h3b0c228e),
	.w3(32'h3bafd97f),
	.w4(32'hbbdc3542),
	.w5(32'h3b6f8818),
	.w6(32'hbc834b4e),
	.w7(32'hbc5e1553),
	.w8(32'hbb617f07),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10d89f),
	.w1(32'h3b6068bd),
	.w2(32'h3bbc0b22),
	.w3(32'hbbe21345),
	.w4(32'hbc2e90dd),
	.w5(32'hbc36e5e5),
	.w6(32'hba7fb8f7),
	.w7(32'hba4ef5de),
	.w8(32'hbad07a42),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ae9081),
	.w1(32'hbbeb1e5a),
	.w2(32'hbb38ad07),
	.w3(32'hbbe94903),
	.w4(32'hbc29c0bb),
	.w5(32'hb9906880),
	.w6(32'h3bce3986),
	.w7(32'hba792dff),
	.w8(32'hbb86be9b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce41afc),
	.w1(32'h3967dce6),
	.w2(32'hb97a6b63),
	.w3(32'hbb8eea6e),
	.w4(32'h3a53ddd3),
	.w5(32'h3b5231ee),
	.w6(32'h3c811d73),
	.w7(32'h3bfef54e),
	.w8(32'hbc30426d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b426f),
	.w1(32'h3a8bada9),
	.w2(32'hbbeb953e),
	.w3(32'h3c1aceda),
	.w4(32'hb9e3cfd0),
	.w5(32'h3a230644),
	.w6(32'hbb209bc5),
	.w7(32'hbc01ac37),
	.w8(32'h3c7ffa96),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc97b5),
	.w1(32'h3b88d158),
	.w2(32'hbadaaa2a),
	.w3(32'hba9b3302),
	.w4(32'h3bfd1fca),
	.w5(32'h3c2b0741),
	.w6(32'h3bdb0ed4),
	.w7(32'hbc22526a),
	.w8(32'h3bbf782a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab94b81),
	.w1(32'h3bbf1bd2),
	.w2(32'hbaaa0eee),
	.w3(32'hbb102466),
	.w4(32'h3b55e1c1),
	.w5(32'hbb303ec4),
	.w6(32'hbb437569),
	.w7(32'h3b4cb18c),
	.w8(32'hbb54df00),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5002d),
	.w1(32'hbbb3da60),
	.w2(32'hbb4bab71),
	.w3(32'hbbc27750),
	.w4(32'h3a768265),
	.w5(32'hbb8c2188),
	.w6(32'hbac9e6f5),
	.w7(32'hbb7c898a),
	.w8(32'hb97ec1c0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc830850),
	.w1(32'h3ba02522),
	.w2(32'hbb31d9d4),
	.w3(32'hbba10d39),
	.w4(32'h3a93e060),
	.w5(32'hba9d2f1c),
	.w6(32'h3d0bad3e),
	.w7(32'h3afb8bf1),
	.w8(32'hba044bcb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbae0d2),
	.w1(32'hba9d7ca4),
	.w2(32'h3bf6c459),
	.w3(32'hbcc89dec),
	.w4(32'hbb1ceea8),
	.w5(32'hbb51ae8c),
	.w6(32'hbc231621),
	.w7(32'hbb1719a1),
	.w8(32'hbd98758b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2b2ce),
	.w1(32'hbb0d92c0),
	.w2(32'h3b1e0223),
	.w3(32'h3c0005c0),
	.w4(32'hbbd3b83a),
	.w5(32'h39c94b96),
	.w6(32'h3c11c7b9),
	.w7(32'h3c30586d),
	.w8(32'h3bad50a6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10b5f5),
	.w1(32'hbca71065),
	.w2(32'hbb55991f),
	.w3(32'h3aae36ad),
	.w4(32'h3b4e11d5),
	.w5(32'hbbd386d5),
	.w6(32'hbada7f02),
	.w7(32'hbb33b8ec),
	.w8(32'hba827d6c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adba9ee),
	.w1(32'h3c84788d),
	.w2(32'h3b50b715),
	.w3(32'h3ab32d30),
	.w4(32'h3b3d4aee),
	.w5(32'h3ad4417d),
	.w6(32'h3b5c1d11),
	.w7(32'hbaada4cc),
	.w8(32'hb9b3a35f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf6e43),
	.w1(32'h3b8f45ca),
	.w2(32'h38e9108f),
	.w3(32'h3b2465d8),
	.w4(32'h3c030567),
	.w5(32'h3c5b15b4),
	.w6(32'h3bfebb99),
	.w7(32'hbafc78e4),
	.w8(32'h3b048967),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc9fc2),
	.w1(32'hbb818986),
	.w2(32'h3b922731),
	.w3(32'hbb477570),
	.w4(32'hbb255ff6),
	.w5(32'hbadf194f),
	.w6(32'hbc9d6e93),
	.w7(32'hbbecb64b),
	.w8(32'hbb5f3677),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86ef46),
	.w1(32'hbb63c5af),
	.w2(32'hbbfc63ff),
	.w3(32'hbbca7554),
	.w4(32'hbba7f805),
	.w5(32'h3a85d90c),
	.w6(32'h3b3d2fef),
	.w7(32'h3c08d5ef),
	.w8(32'h38011442),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b851b37),
	.w1(32'h3a948ec5),
	.w2(32'hba57d203),
	.w3(32'hbc8c4254),
	.w4(32'h38883240),
	.w5(32'hbc0851cd),
	.w6(32'h3b1df252),
	.w7(32'h3b58ab07),
	.w8(32'hbc5dbaac),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc406ce0),
	.w1(32'hbb6b8090),
	.w2(32'h3c1176db),
	.w3(32'hbbfcc1e3),
	.w4(32'hbb86e7c0),
	.w5(32'hbaef7a92),
	.w6(32'h3a0413a0),
	.w7(32'hbc75d999),
	.w8(32'hbc552f5e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dfeb0),
	.w1(32'h3b10c2dd),
	.w2(32'hbc0e992a),
	.w3(32'h3a99817c),
	.w4(32'hbc3fca50),
	.w5(32'hbc3cb734),
	.w6(32'h38a1e5c7),
	.w7(32'hbae92c08),
	.w8(32'hbbd95bb5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8a68f),
	.w1(32'hbadbfa03),
	.w2(32'h3c8773f4),
	.w3(32'h3baff4e3),
	.w4(32'hbc0e632a),
	.w5(32'h3bab3f96),
	.w6(32'h3b85541b),
	.w7(32'hbbbffce2),
	.w8(32'hbb0c6b3c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b996c1b),
	.w1(32'hbadcd1e9),
	.w2(32'h3ac20b07),
	.w3(32'h3c044abd),
	.w4(32'hb71787bb),
	.w5(32'hba635f8a),
	.w6(32'h3afc44e5),
	.w7(32'h3bf12715),
	.w8(32'hbc2f3684),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8ad2f),
	.w1(32'hba865c06),
	.w2(32'hbbd51133),
	.w3(32'h39f5087a),
	.w4(32'hbbe0842a),
	.w5(32'hba80429e),
	.w6(32'hbba6a473),
	.w7(32'hbb954055),
	.w8(32'h3d27a375),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf32b2),
	.w1(32'hbbc2744c),
	.w2(32'hbc8ea262),
	.w3(32'hbd00715d),
	.w4(32'hbc0e010c),
	.w5(32'hbba08277),
	.w6(32'h3c05dc28),
	.w7(32'h3bf59d11),
	.w8(32'h3bfc0ff0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace6e9f),
	.w1(32'hbbed3bbf),
	.w2(32'hbb900b29),
	.w3(32'hbb3898fa),
	.w4(32'hbb5fd8aa),
	.w5(32'hb9b6d986),
	.w6(32'hba6e76df),
	.w7(32'hbb5b1f2c),
	.w8(32'hbbbe3fdd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82526c),
	.w1(32'hbaefd34b),
	.w2(32'hbb95d335),
	.w3(32'h3a3ffec5),
	.w4(32'h3baa75ff),
	.w5(32'hbd1f6fc6),
	.w6(32'hba311012),
	.w7(32'hbaba5b28),
	.w8(32'h3b8611a7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa07b9a),
	.w1(32'h37f1f984),
	.w2(32'hbbb441d4),
	.w3(32'hbae4d504),
	.w4(32'hbbb5bf35),
	.w5(32'h3b6bf1ac),
	.w6(32'h3baebae0),
	.w7(32'hb9bde065),
	.w8(32'h3affaaf1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4071f9),
	.w1(32'hbb90a50e),
	.w2(32'h39833244),
	.w3(32'hbbbcc77f),
	.w4(32'hb9cb34fc),
	.w5(32'hbadc4f93),
	.w6(32'h3d78d325),
	.w7(32'hbcf29176),
	.w8(32'h3b2b8aaa),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64e4aa),
	.w1(32'hbb8fa927),
	.w2(32'h3ce6fb13),
	.w3(32'hbb918825),
	.w4(32'hbbdb80d0),
	.w5(32'hbbda17dc),
	.w6(32'hbc8a60da),
	.w7(32'hbb0c7cf5),
	.w8(32'h3c473da0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c4ab7),
	.w1(32'h3c267513),
	.w2(32'h3bbb5573),
	.w3(32'h3b5c3455),
	.w4(32'hbba400d6),
	.w5(32'hbbce0549),
	.w6(32'hb950a633),
	.w7(32'h3c9d5c9a),
	.w8(32'h3bda272b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace633d),
	.w1(32'h3a1f4f54),
	.w2(32'h3a57563b),
	.w3(32'hbc34ebbf),
	.w4(32'hbb788333),
	.w5(32'h3afde394),
	.w6(32'hba9cda3d),
	.w7(32'hbca34305),
	.w8(32'hbcb85122),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade54d6),
	.w1(32'hbaaadba5),
	.w2(32'hba1b778f),
	.w3(32'hbc11e2f3),
	.w4(32'hb6d99be9),
	.w5(32'h3c0177fa),
	.w6(32'h3cb55e14),
	.w7(32'hbc018a7c),
	.w8(32'h3b7c9226),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d2c0c),
	.w1(32'hb9c75660),
	.w2(32'h3ba20e88),
	.w3(32'h3a6eff8b),
	.w4(32'hba84e3bf),
	.w5(32'hbc8f33e7),
	.w6(32'h39117d93),
	.w7(32'hbd3e621d),
	.w8(32'h3b803a9b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8383e0),
	.w1(32'hbbdc3e34),
	.w2(32'hb9f74c6b),
	.w3(32'h3b8969f9),
	.w4(32'h3cdd7807),
	.w5(32'h3b5a7aed),
	.w6(32'hbb13d7e5),
	.w7(32'hbad85018),
	.w8(32'hbacc09ff),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa28e76),
	.w1(32'hbd03aa06),
	.w2(32'hbb42e7f3),
	.w3(32'h3b820250),
	.w4(32'hbb409ec1),
	.w5(32'hbcebce84),
	.w6(32'hbbc9704c),
	.w7(32'h3c0ed1a8),
	.w8(32'h3bfebbb4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35b67c),
	.w1(32'hbc339eb4),
	.w2(32'hb9d1c723),
	.w3(32'hbb79218e),
	.w4(32'h3a2cde71),
	.w5(32'hb9c4deb1),
	.w6(32'hbc814df3),
	.w7(32'h3c868afc),
	.w8(32'hbc43cf42),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed4675),
	.w1(32'hbb3c6fd4),
	.w2(32'hbb63025a),
	.w3(32'hbbbf15a1),
	.w4(32'hbb5bbcab),
	.w5(32'hbbcaeb00),
	.w6(32'hbbf62be7),
	.w7(32'h3bce5669),
	.w8(32'hbbe9fb03),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba832b4f),
	.w1(32'h3b82d0a4),
	.w2(32'h39d473d3),
	.w3(32'hbacb898f),
	.w4(32'h3a81cb93),
	.w5(32'h3c4feae6),
	.w6(32'hbb24b54a),
	.w7(32'h3a951523),
	.w8(32'hba0fda9c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd792f9),
	.w1(32'h3a5d28e1),
	.w2(32'hbc0093bc),
	.w3(32'hbc0ff590),
	.w4(32'hb94359d6),
	.w5(32'h3bbba980),
	.w6(32'hbbf57961),
	.w7(32'hb85a58f4),
	.w8(32'h3c4692f6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba505fe),
	.w1(32'h3b9d3005),
	.w2(32'h3cd3b82b),
	.w3(32'h3c4c9e75),
	.w4(32'hbb00e01f),
	.w5(32'h3bfd895f),
	.w6(32'h3a2deed0),
	.w7(32'hbbcf3a40),
	.w8(32'h3c5982c3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba8b4f),
	.w1(32'h3c130858),
	.w2(32'hbb2e6210),
	.w3(32'h39b36a65),
	.w4(32'h3b8bf396),
	.w5(32'hbc27c72d),
	.w6(32'hb9ae5a58),
	.w7(32'h3b8aa40c),
	.w8(32'hbbf8b709),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54fb73),
	.w1(32'hbbc3aca9),
	.w2(32'hbc01355f),
	.w3(32'h3c263384),
	.w4(32'h3c36b3d9),
	.w5(32'h3b4ab648),
	.w6(32'h37e39c03),
	.w7(32'hbba424ea),
	.w8(32'hbac01ba8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f9815),
	.w1(32'h3ca7151f),
	.w2(32'hbbfb8256),
	.w3(32'h3b66f304),
	.w4(32'hbb6860e0),
	.w5(32'hbafeaebb),
	.w6(32'h3bd6e59e),
	.w7(32'h3bddd643),
	.w8(32'h3a907171),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5518d7),
	.w1(32'h3ab031d4),
	.w2(32'h3b7e597b),
	.w3(32'h3b4d719e),
	.w4(32'hbba8de6c),
	.w5(32'h3af0c12c),
	.w6(32'hbbc51f0e),
	.w7(32'hbabb280d),
	.w8(32'h3a8d5b59),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b845acb),
	.w1(32'hb9f23e3d),
	.w2(32'hbc3771e5),
	.w3(32'h3abf97f9),
	.w4(32'h3c0bc190),
	.w5(32'hbc0d6be9),
	.w6(32'hbbaebf4a),
	.w7(32'h3aed156e),
	.w8(32'h3c050cb8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cd063),
	.w1(32'h3c9cedfe),
	.w2(32'h3bd9d4b6),
	.w3(32'hbb889927),
	.w4(32'hbbcdb627),
	.w5(32'h3b14e8e6),
	.w6(32'hbb10c249),
	.w7(32'h3bc8d7ed),
	.w8(32'h3b0bd71f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11c026),
	.w1(32'hbb1203d7),
	.w2(32'hbc096d49),
	.w3(32'hba375050),
	.w4(32'h3c24de48),
	.w5(32'hb95d1d16),
	.w6(32'hbc326e96),
	.w7(32'h3af2d1f9),
	.w8(32'hbb296e2b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967ebbf),
	.w1(32'h39a9d1bf),
	.w2(32'hb8c5ffcc),
	.w3(32'h3b0781dc),
	.w4(32'hbaf86c3c),
	.w5(32'h3a6fb1cb),
	.w6(32'h3a8208ce),
	.w7(32'h3ba0025e),
	.w8(32'hbb95f132),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5db2b),
	.w1(32'h3cec31ea),
	.w2(32'h3ad6cb65),
	.w3(32'h381cca3e),
	.w4(32'hbbed7d95),
	.w5(32'h3af0b784),
	.w6(32'h3ca284fe),
	.w7(32'hbc2c80b5),
	.w8(32'h3af8b086),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc393be3),
	.w1(32'hb9b898b5),
	.w2(32'hbb831dc4),
	.w3(32'h3b2c1b8c),
	.w4(32'h3c249d92),
	.w5(32'hbbda7da2),
	.w6(32'hbbc5e0b7),
	.w7(32'h3a9a5a63),
	.w8(32'h382f2eb3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c49f9),
	.w1(32'hbc189411),
	.w2(32'h3aa64b3b),
	.w3(32'h39edb3ec),
	.w4(32'hbb1e3076),
	.w5(32'h39f2c5c9),
	.w6(32'hbbe24a5a),
	.w7(32'h3ba53a86),
	.w8(32'h3bef8919),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5325c9),
	.w1(32'hba68a2b8),
	.w2(32'h3bb2847c),
	.w3(32'hbb369dfd),
	.w4(32'h3b276d37),
	.w5(32'hb8bad0b9),
	.w6(32'h3b1526b0),
	.w7(32'h3bb6133a),
	.w8(32'h3bc36ca2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc139807),
	.w1(32'h3c6cda94),
	.w2(32'hbb885912),
	.w3(32'h3b363d89),
	.w4(32'hba0862d4),
	.w5(32'hbba37e7e),
	.w6(32'h39dec900),
	.w7(32'hbb1b93f1),
	.w8(32'h3a3d37a9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7b8e),
	.w1(32'hbba84813),
	.w2(32'h3b53234c),
	.w3(32'h3c89350e),
	.w4(32'hb9fcc3f5),
	.w5(32'h3b1c93ea),
	.w6(32'h3b974a2e),
	.w7(32'hbba88891),
	.w8(32'h3c3695b5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06f18c),
	.w1(32'hbc3a935b),
	.w2(32'hbb7c453a),
	.w3(32'hb91045d4),
	.w4(32'hbaaa524e),
	.w5(32'h38d7281b),
	.w6(32'hbb1e6ef2),
	.w7(32'hbb4a7f6d),
	.w8(32'h3b8f405c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7dd01),
	.w1(32'hbbb156b0),
	.w2(32'hba4ba7f6),
	.w3(32'hbb21fa94),
	.w4(32'hbab4613d),
	.w5(32'hbb1911d0),
	.w6(32'h3b4f39c1),
	.w7(32'hbb74dfd1),
	.w8(32'hbc2f4641),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcee08d),
	.w1(32'h39d03537),
	.w2(32'h3bc1ba08),
	.w3(32'hb9d0d42b),
	.w4(32'hbba5ff0c),
	.w5(32'h3ae63f48),
	.w6(32'h3be8debe),
	.w7(32'h38b526ba),
	.w8(32'hbb136150),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34d5bb),
	.w1(32'h3bb1ac4d),
	.w2(32'h3c5a1331),
	.w3(32'h3c7c5e95),
	.w4(32'hbb81f6ba),
	.w5(32'hbc07d596),
	.w6(32'h3b8ff43f),
	.w7(32'hbb870518),
	.w8(32'h3bf396b0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e45cd),
	.w1(32'h3b26d685),
	.w2(32'hbb5a3902),
	.w3(32'hbb1979ac),
	.w4(32'h3c08226f),
	.w5(32'h3a8df47e),
	.w6(32'hb963ba22),
	.w7(32'hba88d435),
	.w8(32'h3c43fb13),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6c526),
	.w1(32'hbc4d879e),
	.w2(32'h3bdf4e48),
	.w3(32'hbb2f2460),
	.w4(32'hbaaf9b17),
	.w5(32'h3a8b0733),
	.w6(32'h3bc80af1),
	.w7(32'h3b703348),
	.w8(32'hb781d616),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf92e86),
	.w1(32'h3a94ba93),
	.w2(32'hb9d40fc5),
	.w3(32'h3aa1bfc5),
	.w4(32'h3abd846e),
	.w5(32'hbbcbf3f2),
	.w6(32'h3ac07797),
	.w7(32'hbaac4cbf),
	.w8(32'hbb619fe8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e2517),
	.w1(32'h3a3dfb35),
	.w2(32'h3c7f0166),
	.w3(32'h3c387133),
	.w4(32'h3b405dd0),
	.w5(32'hbbb7c3f6),
	.w6(32'h3bd06726),
	.w7(32'hbbafae59),
	.w8(32'h3c21ebb6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c556f41),
	.w1(32'h3ba803fb),
	.w2(32'hb79a7375),
	.w3(32'hbc3b3ba0),
	.w4(32'h3c739d50),
	.w5(32'h3b60d1b8),
	.w6(32'h39d0a408),
	.w7(32'hbb9d3fb9),
	.w8(32'hbb9c09ec),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e097b),
	.w1(32'hbc9bfe8a),
	.w2(32'hbc30709c),
	.w3(32'h3a0993c3),
	.w4(32'h3b5e005a),
	.w5(32'hbb96daee),
	.w6(32'h3abb9024),
	.w7(32'h3be86c21),
	.w8(32'h3c1b03bd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb8e10),
	.w1(32'hbb8e8abb),
	.w2(32'hbb44d09a),
	.w3(32'h3b4cee68),
	.w4(32'hb9e83894),
	.w5(32'h3bdceeb4),
	.w6(32'h3b08f116),
	.w7(32'h3cd28993),
	.w8(32'h3b187889),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2fd83),
	.w1(32'hbc62bc42),
	.w2(32'hbb9ce842),
	.w3(32'h3a4a2daf),
	.w4(32'h3af9a8de),
	.w5(32'hbc1a7c2f),
	.w6(32'h3afa3ee0),
	.w7(32'h3ae874d3),
	.w8(32'h3c23c251),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1e8ef),
	.w1(32'h3bb78ab2),
	.w2(32'hbb1d8483),
	.w3(32'h3bfb5143),
	.w4(32'h3b56b52c),
	.w5(32'hbbab9e6c),
	.w6(32'hbb2c8d65),
	.w7(32'h3c5824fb),
	.w8(32'hbb827f81),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7025c0),
	.w1(32'hbc05c07b),
	.w2(32'hbbdd6d1b),
	.w3(32'hba55a274),
	.w4(32'h3b6a05dd),
	.w5(32'hbc82a4ac),
	.w6(32'h3ac17f57),
	.w7(32'h3bd6efdf),
	.w8(32'hba958825),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c082a31),
	.w1(32'h3c2d7986),
	.w2(32'hbc1d7876),
	.w3(32'hbc8aa4ed),
	.w4(32'h3b634b9c),
	.w5(32'hbb1c969b),
	.w6(32'hba220c3e),
	.w7(32'hbb8e8941),
	.w8(32'h3bcae24d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6e15e),
	.w1(32'h3c6e546c),
	.w2(32'h3c2c2e3f),
	.w3(32'h3b48c754),
	.w4(32'hbbae7b57),
	.w5(32'hb9b0d5be),
	.w6(32'h3c312882),
	.w7(32'h3a94dd58),
	.w8(32'hbc43c142),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0efb79),
	.w1(32'h3c944cc5),
	.w2(32'hbc74b8c9),
	.w3(32'hbc357749),
	.w4(32'hbc0c57ab),
	.w5(32'hbc47d7c0),
	.w6(32'hbbab94b1),
	.w7(32'hbaefe10c),
	.w8(32'hbc094bfe),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb838ba8),
	.w1(32'h3bf005a9),
	.w2(32'h3b407091),
	.w3(32'h3bd18d86),
	.w4(32'hbb547b8c),
	.w5(32'hbbc35b23),
	.w6(32'hbb150651),
	.w7(32'hb77edb9f),
	.w8(32'hbbe25d70),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb053dc9),
	.w1(32'hbabb0bb3),
	.w2(32'hbbea6a21),
	.w3(32'hbb12183f),
	.w4(32'hbaad674b),
	.w5(32'h3961fd06),
	.w6(32'h3b050896),
	.w7(32'h3afb082d),
	.w8(32'hbc91e133),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c9849),
	.w1(32'hbbdd41cf),
	.w2(32'h3c94e0ec),
	.w3(32'hb8efc7d1),
	.w4(32'h3b014261),
	.w5(32'hbc094d64),
	.w6(32'hbc1205e8),
	.w7(32'h3c16ef52),
	.w8(32'h3ba356b7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac81259),
	.w1(32'h3bc1a914),
	.w2(32'hb9cd1a6d),
	.w3(32'hba41a7a1),
	.w4(32'h3c87fbad),
	.w5(32'h3c19192d),
	.w6(32'h3af788ec),
	.w7(32'hba2abeb1),
	.w8(32'h3b0bf2e4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae61a5),
	.w1(32'hbc16e641),
	.w2(32'h3a7d30e2),
	.w3(32'hbb575bac),
	.w4(32'hbb98d3dd),
	.w5(32'hbc2fb7d5),
	.w6(32'h3b609a67),
	.w7(32'hb990181c),
	.w8(32'hbb100a48),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab2616),
	.w1(32'hbbb153e6),
	.w2(32'h3c232221),
	.w3(32'hb71eab4f),
	.w4(32'h3c1cac57),
	.w5(32'hba40ff07),
	.w6(32'hb98e8841),
	.w7(32'hbbe4a4e0),
	.w8(32'hbc1df8cf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2b76b),
	.w1(32'h3af40d12),
	.w2(32'h3ad62704),
	.w3(32'h3bf484b3),
	.w4(32'hbb337ef2),
	.w5(32'h3a0279ee),
	.w6(32'hb8796c2a),
	.w7(32'h3b0bc66d),
	.w8(32'h3b5cd2db),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94c3c1),
	.w1(32'h36c1f8d9),
	.w2(32'h3c64e645),
	.w3(32'hbb8a6ed1),
	.w4(32'h3b73ab6e),
	.w5(32'h3b5babeb),
	.w6(32'h3bedbe69),
	.w7(32'h3ad420aa),
	.w8(32'hbb171f96),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc016210),
	.w1(32'hbc0c51e0),
	.w2(32'h3a3fc910),
	.w3(32'h38bae39c),
	.w4(32'hb9bda4cd),
	.w5(32'hbb60b8d8),
	.w6(32'h3ad91a41),
	.w7(32'h3c3a6b3d),
	.w8(32'hbc2efe36),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba68794),
	.w1(32'h3b718c63),
	.w2(32'hbac5e336),
	.w3(32'hba6b546f),
	.w4(32'hbcb399fd),
	.w5(32'hbc68031f),
	.w6(32'hbc18b266),
	.w7(32'hbc0420b1),
	.w8(32'h3b98d1b1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb254db2),
	.w1(32'hbc6375bd),
	.w2(32'h3a66e8cc),
	.w3(32'hbc03a9c4),
	.w4(32'h3b6e9ce9),
	.w5(32'h3c3bb002),
	.w6(32'hbaeac4da),
	.w7(32'hbc3798e1),
	.w8(32'h3c927cff),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67238a),
	.w1(32'hbaba5579),
	.w2(32'h3c93aeb3),
	.w3(32'h3ae53bd7),
	.w4(32'h3a0f8d76),
	.w5(32'h3bbb1913),
	.w6(32'hbb5a3340),
	.w7(32'hbb5f3b94),
	.w8(32'h391e3d1c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a746f79),
	.w1(32'h3b4d5b09),
	.w2(32'hba957c38),
	.w3(32'h3b8cfa24),
	.w4(32'hbbb5663f),
	.w5(32'hb8c1c162),
	.w6(32'h3846f45f),
	.w7(32'hbca5a7b7),
	.w8(32'hbbfd471f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ec8a7),
	.w1(32'h3c5a62eb),
	.w2(32'hbb97509e),
	.w3(32'h3c2f4649),
	.w4(32'hba63e462),
	.w5(32'h3bd053cc),
	.w6(32'hbbdd04a8),
	.w7(32'h3a08d6a6),
	.w8(32'hba316600),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40f841),
	.w1(32'hbb9a1ac0),
	.w2(32'hba05429a),
	.w3(32'h3c6f8e6d),
	.w4(32'h3aee3200),
	.w5(32'h38d6c1da),
	.w6(32'h3ba21c97),
	.w7(32'hbbc1a724),
	.w8(32'hbb2f09ad),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d7dc7),
	.w1(32'hbb33e1d2),
	.w2(32'hbbb1a133),
	.w3(32'hbc0967e9),
	.w4(32'hbc3a67e9),
	.w5(32'h3c085545),
	.w6(32'h3c4e25c9),
	.w7(32'hb8c0fe5d),
	.w8(32'hbb6b74f1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36ac90),
	.w1(32'hbbe5406e),
	.w2(32'h3b894df7),
	.w3(32'h3b99cf92),
	.w4(32'h3bd8ad77),
	.w5(32'hbb8218b5),
	.w6(32'hbc2b4069),
	.w7(32'hba9fec9b),
	.w8(32'h3b79c690),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad7e24),
	.w1(32'hb9655c2a),
	.w2(32'h3b298a77),
	.w3(32'hbc9a241a),
	.w4(32'hbb343a72),
	.w5(32'hba4cf5bb),
	.w6(32'h38bbdcd8),
	.w7(32'h3a9c3a80),
	.w8(32'hbb355248),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a7e58),
	.w1(32'hbb219cea),
	.w2(32'hbc49f62e),
	.w3(32'hb94a1a6b),
	.w4(32'hbcc8deeb),
	.w5(32'h3a4fc33d),
	.w6(32'hb9709024),
	.w7(32'h3adb652f),
	.w8(32'hbbdc3dc9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2194e9),
	.w1(32'hbc1d2e15),
	.w2(32'h3b056107),
	.w3(32'hbbe8b654),
	.w4(32'hbae87a4b),
	.w5(32'h3b5171aa),
	.w6(32'hbb8ff191),
	.w7(32'h3a58cd4c),
	.w8(32'hbc9a8017),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46422d),
	.w1(32'h3bed6f56),
	.w2(32'hbba65ddd),
	.w3(32'h3b829b95),
	.w4(32'h3b89de40),
	.w5(32'h3984fc02),
	.w6(32'hbc13a20c),
	.w7(32'h3c4b3f02),
	.w8(32'h3bc3c1d2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7bf6d),
	.w1(32'h3b0edec0),
	.w2(32'hbc13d286),
	.w3(32'h3b0546ec),
	.w4(32'h3cc6fe6d),
	.w5(32'hbb0da15b),
	.w6(32'hbb1a5474),
	.w7(32'hbb501094),
	.w8(32'h3b654396),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa7e46),
	.w1(32'hbb088dd6),
	.w2(32'hba733167),
	.w3(32'h3c088138),
	.w4(32'h3bf4120f),
	.w5(32'hbbad80a4),
	.w6(32'h3a6622ce),
	.w7(32'hbaa89962),
	.w8(32'hbc466280),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80c5f9),
	.w1(32'hbbc2b927),
	.w2(32'h3c1a2424),
	.w3(32'h3cb31d62),
	.w4(32'hbbe1b1a9),
	.w5(32'hbba405be),
	.w6(32'h3c1f93f8),
	.w7(32'h3c356a6a),
	.w8(32'h3caa1653),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44e3e1),
	.w1(32'h3c4e8a52),
	.w2(32'hbc1d69b6),
	.w3(32'hbb881c06),
	.w4(32'h3ba5b739),
	.w5(32'hbb58d47c),
	.w6(32'hbb8c8dbb),
	.w7(32'h3cc657aa),
	.w8(32'h3d0433fc),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfde124),
	.w1(32'h3c19735a),
	.w2(32'h3c5e9438),
	.w3(32'hbbcdc556),
	.w4(32'hb9b8068a),
	.w5(32'hbbabced9),
	.w6(32'hbaa36ced),
	.w7(32'h3b81ca71),
	.w8(32'h3c59bab2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fff42),
	.w1(32'h3c706caa),
	.w2(32'hbc970c56),
	.w3(32'hbc4e1a67),
	.w4(32'hbbbc51ca),
	.w5(32'h3b414452),
	.w6(32'h3b3bba27),
	.w7(32'hbc601d9c),
	.w8(32'hbb92ad44),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a2c8e),
	.w1(32'hbb94bec8),
	.w2(32'hbc250572),
	.w3(32'hbc102a51),
	.w4(32'hbc0158de),
	.w5(32'hbc9386da),
	.w6(32'hbc72bb7a),
	.w7(32'hbbf8a2f3),
	.w8(32'hbb1ae01a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d1618),
	.w1(32'h3995b993),
	.w2(32'hbb7048e2),
	.w3(32'hbcbf569c),
	.w4(32'h3bf10ce5),
	.w5(32'h3ba2f097),
	.w6(32'h3c038940),
	.w7(32'h3c8df6b0),
	.w8(32'h3a37f4c7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b178f94),
	.w1(32'hbc51378b),
	.w2(32'hb94f17ea),
	.w3(32'hbbae24a7),
	.w4(32'h3c47fe12),
	.w5(32'h3a93fff4),
	.w6(32'h3c88bc0a),
	.w7(32'h3c7f5e6e),
	.w8(32'hbc7ab636),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e5fc6),
	.w1(32'h3a6f0268),
	.w2(32'hbbcdae2e),
	.w3(32'h3b5256c2),
	.w4(32'hbb7d21bc),
	.w5(32'h3cbdc521),
	.w6(32'h3a3252b0),
	.w7(32'hbc984484),
	.w8(32'h3d0d7163),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1560d7),
	.w1(32'hbbb9c235),
	.w2(32'h3ad8723d),
	.w3(32'hbc060e3e),
	.w4(32'hbb4730e4),
	.w5(32'hba74add2),
	.w6(32'h3d57c8c4),
	.w7(32'h3bbe91f4),
	.w8(32'h3a880ec0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba698ad0),
	.w1(32'hbb01829c),
	.w2(32'hbc9da932),
	.w3(32'h3c0b20ef),
	.w4(32'h3af8692d),
	.w5(32'hbb62dadc),
	.w6(32'hbb4591ce),
	.w7(32'hbc85c1f2),
	.w8(32'h3ab9ad11),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a254ab8),
	.w1(32'h3c2ced78),
	.w2(32'h3c336295),
	.w3(32'h3b4c2422),
	.w4(32'h3c4a3abe),
	.w5(32'h3a713007),
	.w6(32'h3b8922f3),
	.w7(32'h392652a8),
	.w8(32'h3ca7fa4f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c91c1),
	.w1(32'hbc0fbb33),
	.w2(32'hbb6332f0),
	.w3(32'hbb1ff334),
	.w4(32'h3bc1a2c5),
	.w5(32'h3c1a3730),
	.w6(32'hbccecc6a),
	.w7(32'hbb2bc23a),
	.w8(32'hbb84dec6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90b347),
	.w1(32'hbb9f9f40),
	.w2(32'hbb90cb17),
	.w3(32'hbb26cfb2),
	.w4(32'hbc0b07c1),
	.w5(32'hb8900963),
	.w6(32'hbbf7ab88),
	.w7(32'h3af743b3),
	.w8(32'hbc4a79eb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e6009),
	.w1(32'hbc2b1f0f),
	.w2(32'h3c061df1),
	.w3(32'h3c0d4953),
	.w4(32'h3c062147),
	.w5(32'hbc1cb452),
	.w6(32'h3abff172),
	.w7(32'hbb582e50),
	.w8(32'hbbb4d499),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaed0f2),
	.w1(32'hbbc05362),
	.w2(32'hbca1f0fe),
	.w3(32'hbbf2b747),
	.w4(32'hbbb75da9),
	.w5(32'h3bc943fd),
	.w6(32'h3bc80162),
	.w7(32'h3b1644d3),
	.w8(32'h3c3f1dec),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5de8fa),
	.w1(32'h3c0d779b),
	.w2(32'hbc65641b),
	.w3(32'h3c2fa486),
	.w4(32'h3b8d4e35),
	.w5(32'hbc47284c),
	.w6(32'h3cc041f3),
	.w7(32'h3c35f743),
	.w8(32'hbc9419b6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11ef6e),
	.w1(32'hbba3df4f),
	.w2(32'hbbac6f5e),
	.w3(32'hbbb2d843),
	.w4(32'h3c051407),
	.w5(32'h3ae0f69e),
	.w6(32'hbc6be241),
	.w7(32'hbb09b0f5),
	.w8(32'hbb623250),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0d8d),
	.w1(32'hbaec4132),
	.w2(32'hb74b4e85),
	.w3(32'h3c34bc8e),
	.w4(32'hbc730544),
	.w5(32'hbb820ec5),
	.w6(32'hbbfabd7b),
	.w7(32'h3b1fc3f2),
	.w8(32'h3bcdf4bb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb456fa8),
	.w1(32'hbb9ad269),
	.w2(32'h3bf14d46),
	.w3(32'hbb2d8cd9),
	.w4(32'hbbc51051),
	.w5(32'hbc4ff0c3),
	.w6(32'h3c8240e8),
	.w7(32'h3b9f8c7d),
	.w8(32'hbcaaa28a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf83e3d),
	.w1(32'hbb392c06),
	.w2(32'hba41b2f3),
	.w3(32'hbb8956cb),
	.w4(32'h3c14ef0d),
	.w5(32'h3c81d7ef),
	.w6(32'h3c94324f),
	.w7(32'h3b5c04c9),
	.w8(32'hbc0a8691),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a181b),
	.w1(32'hbc289039),
	.w2(32'hbc590dba),
	.w3(32'hbbb1c8eb),
	.w4(32'hbc36bea3),
	.w5(32'h3c036b74),
	.w6(32'h3b9f36c1),
	.w7(32'h3b609e32),
	.w8(32'h3be84fdb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf684b1),
	.w1(32'h3adc9b34),
	.w2(32'hbbaed7ec),
	.w3(32'h3c1c7d85),
	.w4(32'hbbbd6b13),
	.w5(32'hbb0e4be7),
	.w6(32'hbc3281cb),
	.w7(32'hbc2e31bd),
	.w8(32'hbc1eec44),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09b6e7),
	.w1(32'hbbcb678f),
	.w2(32'hbbce4826),
	.w3(32'h3c2482f7),
	.w4(32'h3b726404),
	.w5(32'hb94f388f),
	.w6(32'hbb1bf774),
	.w7(32'hbbab9b88),
	.w8(32'hbbdf41f7),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39987343),
	.w1(32'hbc0e1fda),
	.w2(32'hbaee7e2b),
	.w3(32'hbc4b63b2),
	.w4(32'hba5c161c),
	.w5(32'hba991d7b),
	.w6(32'hbc628aab),
	.w7(32'hba1f5bcb),
	.w8(32'h3c320ccd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58f95a),
	.w1(32'h3a862ea0),
	.w2(32'h3bb31174),
	.w3(32'h3c78d3d7),
	.w4(32'h3c175b54),
	.w5(32'h3c412530),
	.w6(32'h397e63af),
	.w7(32'h3c8ae0d7),
	.w8(32'h3ca3c167),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306516),
	.w1(32'hbc3aa9f7),
	.w2(32'h3c65d33f),
	.w3(32'hbc0806f9),
	.w4(32'h3c78987e),
	.w5(32'hbc06ed0b),
	.w6(32'h3b135303),
	.w7(32'h3c1a951f),
	.w8(32'h3b710967),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d5103),
	.w1(32'h3c386b9c),
	.w2(32'h3da964b4),
	.w3(32'h3ce394c0),
	.w4(32'h38495e42),
	.w5(32'h3cded33f),
	.w6(32'hbce59258),
	.w7(32'h3d1156ef),
	.w8(32'h3cc5806a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0309),
	.w1(32'hbc2f31cb),
	.w2(32'h3acafc6b),
	.w3(32'h3b6bc396),
	.w4(32'h3cb17b17),
	.w5(32'hbc05afeb),
	.w6(32'h3cb93d83),
	.w7(32'h3c862aa1),
	.w8(32'h3bbf4e8f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4da76),
	.w1(32'h3b8ff44c),
	.w2(32'h38d7a2c1),
	.w3(32'hbc103bed),
	.w4(32'h3c03edf3),
	.w5(32'hbaa013ef),
	.w6(32'hbbce570a),
	.w7(32'h3afa8936),
	.w8(32'h39eb9f85),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d73a5),
	.w1(32'hbb39b218),
	.w2(32'h39a6f9eb),
	.w3(32'h3c120f8e),
	.w4(32'h398eb528),
	.w5(32'hb84ab349),
	.w6(32'h3cd098b0),
	.w7(32'hbb221126),
	.w8(32'h3b68e1a3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae9938),
	.w1(32'hb8df393e),
	.w2(32'h3b2cb361),
	.w3(32'hb9adbb31),
	.w4(32'h37e005bf),
	.w5(32'hbcda6c97),
	.w6(32'h3badaf84),
	.w7(32'h3c104378),
	.w8(32'h3ba42871),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0facf),
	.w1(32'h3b32ed14),
	.w2(32'h3af5d32f),
	.w3(32'h3bc9db3f),
	.w4(32'h3bb460f3),
	.w5(32'hbb101e51),
	.w6(32'hbbf01ec4),
	.w7(32'hbb1c0389),
	.w8(32'hbb9e1019),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7df1cf),
	.w1(32'hbc479ae3),
	.w2(32'hbaa532fc),
	.w3(32'hbadfccaf),
	.w4(32'h3baabe9f),
	.w5(32'hbb92da8c),
	.w6(32'h3b30727a),
	.w7(32'h3c068e21),
	.w8(32'hbb4303c1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989c1b5),
	.w1(32'hbb439e1c),
	.w2(32'h3c1f6c20),
	.w3(32'hbae9ce13),
	.w4(32'h3c017e1c),
	.w5(32'h3b6d66ed),
	.w6(32'hbbbd8c6f),
	.w7(32'h3c000bf7),
	.w8(32'h3afbc594),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae69ed9),
	.w1(32'h3c110241),
	.w2(32'h3cc6e526),
	.w3(32'hbc012f88),
	.w4(32'hb8e8c68b),
	.w5(32'h3cdcdce2),
	.w6(32'hbb448ea3),
	.w7(32'h3a95c10e),
	.w8(32'hbb7ba4a1),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a7f43),
	.w1(32'hbae490de),
	.w2(32'h398798c1),
	.w3(32'h3b5c6440),
	.w4(32'h3c2158f3),
	.w5(32'h3ad8c146),
	.w6(32'h3b535cf3),
	.w7(32'hbc0c7162),
	.w8(32'hb9dbface),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05146a),
	.w1(32'hbbd97e6b),
	.w2(32'hbcc7477f),
	.w3(32'hba89044a),
	.w4(32'h3b0f6ff8),
	.w5(32'h3b6124a0),
	.w6(32'hbca65144),
	.w7(32'hbabfb220),
	.w8(32'h3ac06626),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1cf9a),
	.w1(32'hbb2b5960),
	.w2(32'h3b9ccdab),
	.w3(32'h3c5d5c99),
	.w4(32'hba6153cc),
	.w5(32'h39a4acb0),
	.w6(32'hbb9abbfe),
	.w7(32'hbc187ac4),
	.w8(32'hba93bfbb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06589a),
	.w1(32'hba9a21a6),
	.w2(32'h3a6b3ffc),
	.w3(32'hbba8060e),
	.w4(32'h39f4731f),
	.w5(32'h3c620656),
	.w6(32'h3bc8c4e8),
	.w7(32'h39a2a04d),
	.w8(32'h3b2853ba),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387fc7f2),
	.w1(32'hbc2aaded),
	.w2(32'h3cee3135),
	.w3(32'h3ca7e56b),
	.w4(32'h3ba8a262),
	.w5(32'hbc9d06b0),
	.w6(32'hb80e34c0),
	.w7(32'hbc12c97f),
	.w8(32'hbac1a54b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe091ca),
	.w1(32'hba8660ee),
	.w2(32'hba32b5d4),
	.w3(32'hbad80ca9),
	.w4(32'hba63c803),
	.w5(32'h3b67bb3e),
	.w6(32'h3aed6709),
	.w7(32'hbbb238bc),
	.w8(32'hbae9a35f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12230b),
	.w1(32'hbb0f4e8c),
	.w2(32'h3ab54d37),
	.w3(32'h3b4ed10a),
	.w4(32'hb820ca79),
	.w5(32'hbb8fcd14),
	.w6(32'h37811954),
	.w7(32'h3baff07c),
	.w8(32'h3ba135cc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ed7be),
	.w1(32'h3d1432ab),
	.w2(32'h3aaf1ef9),
	.w3(32'hbbcb7be2),
	.w4(32'h3bd4d0ed),
	.w5(32'h3b4affcd),
	.w6(32'hbb8d1530),
	.w7(32'hba853978),
	.w8(32'h3b3b46ce),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf7889),
	.w1(32'hbc7c69ab),
	.w2(32'h3b51173f),
	.w3(32'h3a905da6),
	.w4(32'hbba6c88a),
	.w5(32'hbba5c5eb),
	.w6(32'h3b034f7d),
	.w7(32'h3bf69f27),
	.w8(32'h3b4d0ea2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b4250),
	.w1(32'h3afee4d9),
	.w2(32'h3b6f2caa),
	.w3(32'h3c244e2d),
	.w4(32'h3cbe3617),
	.w5(32'hb8a4eaaf),
	.w6(32'hbbcda294),
	.w7(32'h3b5530cd),
	.w8(32'hbb79d219),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc63e48),
	.w1(32'hbc02b54e),
	.w2(32'hbbd7b4c3),
	.w3(32'h3b8a9cf0),
	.w4(32'h3be46372),
	.w5(32'h3b80176f),
	.w6(32'h3ca094ab),
	.w7(32'hbb16bc83),
	.w8(32'h3c9e053d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b493),
	.w1(32'hba61a788),
	.w2(32'h3bd43694),
	.w3(32'hb9111a44),
	.w4(32'hbb593ab4),
	.w5(32'h3b99168d),
	.w6(32'hbba82edd),
	.w7(32'hbbf89566),
	.w8(32'hbba052a3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8a1cf),
	.w1(32'hbbad8b4b),
	.w2(32'hba612f5e),
	.w3(32'hbb230fbf),
	.w4(32'h38d942ab),
	.w5(32'h3b956b6f),
	.w6(32'h39c06eb2),
	.w7(32'hba4c6f60),
	.w8(32'hbad50e37),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8437298),
	.w1(32'h3aa2d69c),
	.w2(32'hbb1ace18),
	.w3(32'hbc307625),
	.w4(32'hbb9a996c),
	.w5(32'h3c7127ab),
	.w6(32'hbbae994c),
	.w7(32'h3c7907b2),
	.w8(32'h3c15423c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81392c),
	.w1(32'hbb957c7c),
	.w2(32'hbc7ca90d),
	.w3(32'hbbf5e37c),
	.w4(32'hbb8853f7),
	.w5(32'hbaa814bc),
	.w6(32'hbb6f75fe),
	.w7(32'h3c0f8347),
	.w8(32'hb9563710),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb150f),
	.w1(32'h3913c252),
	.w2(32'hbb95e527),
	.w3(32'hbb0534ce),
	.w4(32'hbb8c768a),
	.w5(32'h3b53ee54),
	.w6(32'h3c44f994),
	.w7(32'h3c1ea52a),
	.w8(32'h3bb80e5f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd34834),
	.w1(32'h3c26ba2f),
	.w2(32'hba92f1a9),
	.w3(32'h3a031d59),
	.w4(32'hba7131e6),
	.w5(32'h3be7dd1d),
	.w6(32'hb98d7741),
	.w7(32'hbc4d5d3d),
	.w8(32'hba8d1b2e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c1c53),
	.w1(32'hbb37629b),
	.w2(32'hbae2bb76),
	.w3(32'h3b207eb6),
	.w4(32'h3c12a546),
	.w5(32'h3b30c7b9),
	.w6(32'h3bb5160a),
	.w7(32'h3c0c9619),
	.w8(32'hbb2a7909),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae9308),
	.w1(32'h3c5ee6e1),
	.w2(32'hbc3a9531),
	.w3(32'hbc734c21),
	.w4(32'h3b396687),
	.w5(32'hba213a0c),
	.w6(32'hbc01d553),
	.w7(32'h3c1ccc85),
	.w8(32'hb9b53b47),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ed2e8),
	.w1(32'hbaed6569),
	.w2(32'hbba93212),
	.w3(32'h3c911a84),
	.w4(32'h3b798143),
	.w5(32'h3b907f96),
	.w6(32'hbb416fa8),
	.w7(32'hba8c5ba4),
	.w8(32'hbb806d12),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20a95e),
	.w1(32'hbc957825),
	.w2(32'hbbf0469b),
	.w3(32'h3aaecb3a),
	.w4(32'hbbcf4998),
	.w5(32'hba9a6e43),
	.w6(32'hb99064c8),
	.w7(32'h3c6b3e2b),
	.w8(32'h3ca35fa7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202cb9),
	.w1(32'h3854a5e8),
	.w2(32'hbc345fea),
	.w3(32'h3b7a5494),
	.w4(32'h3be41988),
	.w5(32'hbb6d40c6),
	.w6(32'h3adffda7),
	.w7(32'h3c3547aa),
	.w8(32'h3b25888a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26e67f),
	.w1(32'h3c00805e),
	.w2(32'h3c289e9f),
	.w3(32'hbbd1ec78),
	.w4(32'h3c9491f3),
	.w5(32'h3bc691f9),
	.w6(32'hbc1dc8f4),
	.w7(32'h3b322bfd),
	.w8(32'h3ae15d07),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc03217),
	.w1(32'h3c6aa921),
	.w2(32'h3c4235c4),
	.w3(32'h3bc4ed6d),
	.w4(32'h3c648e90),
	.w5(32'hbbbfecdd),
	.w6(32'h3c04084c),
	.w7(32'h3b734945),
	.w8(32'h3bfb6746),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7eb54d),
	.w1(32'hbc3b0946),
	.w2(32'h3c31a7dd),
	.w3(32'hbc4abc82),
	.w4(32'hbc29abf9),
	.w5(32'hba58ea26),
	.w6(32'hbb710d32),
	.w7(32'hb9add10d),
	.w8(32'h3b771b80),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12562a),
	.w1(32'h3ce0d085),
	.w2(32'h3b14c27f),
	.w3(32'hbb242e0c),
	.w4(32'hbaae5ba3),
	.w5(32'hbc5773f3),
	.w6(32'h3b4fa656),
	.w7(32'hbc275cdc),
	.w8(32'h3abd21b4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fa5a5),
	.w1(32'h3b4f0e75),
	.w2(32'h3cb03e24),
	.w3(32'h39214b43),
	.w4(32'hbc150a4f),
	.w5(32'hbb8c1799),
	.w6(32'hbbbc1792),
	.w7(32'hbc44b8b4),
	.w8(32'hbc158a6e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc873291),
	.w1(32'h3bec469a),
	.w2(32'h3a6f07ca),
	.w3(32'hbc016533),
	.w4(32'h3ba76d5d),
	.w5(32'hbb40e2c2),
	.w6(32'hbba6f105),
	.w7(32'hb8d6451b),
	.w8(32'h3a0c007a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56a9c2),
	.w1(32'hbba28548),
	.w2(32'hbc0adb59),
	.w3(32'h3c056aac),
	.w4(32'hbc61a727),
	.w5(32'h3c3bd47e),
	.w6(32'hbb1ac386),
	.w7(32'hbaada1ff),
	.w8(32'h3c4942ae),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24d9aa),
	.w1(32'hbbcfca94),
	.w2(32'hba8898fb),
	.w3(32'h39800893),
	.w4(32'hba1b9ea2),
	.w5(32'hbb652b29),
	.w6(32'h3c5dde33),
	.w7(32'h3c0f7964),
	.w8(32'h3cb08a7f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c0029),
	.w1(32'hbc02f7a6),
	.w2(32'hbbac3aab),
	.w3(32'h3be06a51),
	.w4(32'h3b731b67),
	.w5(32'h3c16c636),
	.w6(32'hba9f65f2),
	.w7(32'h3a2f31dd),
	.w8(32'h3b692e7d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb84302),
	.w1(32'hbc3f4500),
	.w2(32'h3c33ea9e),
	.w3(32'hbbb9b942),
	.w4(32'h3bba2a03),
	.w5(32'h3ca7165f),
	.w6(32'h3c03be79),
	.w7(32'hbb65f321),
	.w8(32'hbb7f5d8e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a406),
	.w1(32'hbc3f3ac6),
	.w2(32'h3be0597f),
	.w3(32'hbc802eb6),
	.w4(32'hb8d98e44),
	.w5(32'hbc5cf8a0),
	.w6(32'h3c823395),
	.w7(32'hbb4fe63f),
	.w8(32'h3c2908eb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e1948),
	.w1(32'hbb47aa79),
	.w2(32'h3bda4fe4),
	.w3(32'hbc81d6c3),
	.w4(32'hb9bc3144),
	.w5(32'h3b394592),
	.w6(32'h3ba7da18),
	.w7(32'hbba6c40b),
	.w8(32'h3c1c87aa),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5dd30),
	.w1(32'h3b5fe78f),
	.w2(32'h34c8b74d),
	.w3(32'h39b48df7),
	.w4(32'hba2ce5c2),
	.w5(32'hbd00c580),
	.w6(32'h3b6efab9),
	.w7(32'h3c71f0b0),
	.w8(32'h3b190cd3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8674b),
	.w1(32'hba4bbf0d),
	.w2(32'hbb448101),
	.w3(32'h3c8aa971),
	.w4(32'h3ab0cd81),
	.w5(32'hbc3a5be0),
	.w6(32'h3a568fad),
	.w7(32'hba09900f),
	.w8(32'hbb1e91ab),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a13a9),
	.w1(32'h3b1c5c80),
	.w2(32'hbc323dc0),
	.w3(32'hbad5e864),
	.w4(32'hbc2ec2e9),
	.w5(32'h3b7f492e),
	.w6(32'hbc44fa8f),
	.w7(32'h3d06b412),
	.w8(32'h3c1f0e7d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1577da),
	.w1(32'h3a2b1e40),
	.w2(32'hbb3540a9),
	.w3(32'h3c209cbc),
	.w4(32'h3c0e80a5),
	.w5(32'h3bbca875),
	.w6(32'hbb3826b4),
	.w7(32'hbbbdaa4f),
	.w8(32'hbbe8b306),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aedfc3),
	.w1(32'hba539982),
	.w2(32'hbbf62757),
	.w3(32'hbbb0e472),
	.w4(32'hba727be6),
	.w5(32'h3c07b946),
	.w6(32'hb99b7118),
	.w7(32'h3a9c070f),
	.w8(32'h3bfcc456),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb876c11),
	.w1(32'h3bbf8653),
	.w2(32'h3b2065ac),
	.w3(32'h3b1b7138),
	.w4(32'hbb85a172),
	.w5(32'hbbbbeaec),
	.w6(32'h3a9a6b1f),
	.w7(32'h365b5c2d),
	.w8(32'h3b557856),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb194537),
	.w1(32'hbcabf1da),
	.w2(32'hbc9c226c),
	.w3(32'h3ab0c501),
	.w4(32'hbbf6d65d),
	.w5(32'h3c647134),
	.w6(32'hbb46f507),
	.w7(32'hba85c31e),
	.w8(32'h3a050ff3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbe1ac),
	.w1(32'hbc18d9d7),
	.w2(32'h3ab817f9),
	.w3(32'hbaa821b1),
	.w4(32'hbc5f30b9),
	.w5(32'h3ae68ec3),
	.w6(32'hbb2deec5),
	.w7(32'h3c71e15b),
	.w8(32'h3c64bdfb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0bf11),
	.w1(32'hbbad38cb),
	.w2(32'hbbc612a9),
	.w3(32'h3c3ea0c2),
	.w4(32'h3aaf5f16),
	.w5(32'hbbb0a54a),
	.w6(32'hbb96e685),
	.w7(32'h3d312002),
	.w8(32'hbba1fcce),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a156de3),
	.w1(32'hbc1c76d1),
	.w2(32'h3b4d7b54),
	.w3(32'hbc5ff639),
	.w4(32'h3bb2f639),
	.w5(32'h3cafd873),
	.w6(32'hbc4627a7),
	.w7(32'h3baddbcf),
	.w8(32'hbc099c5b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16577e),
	.w1(32'hbc9bd09c),
	.w2(32'h3779f3ed),
	.w3(32'hbbbf799b),
	.w4(32'h3b6f2e92),
	.w5(32'h3b893b4f),
	.w6(32'hb9db58b9),
	.w7(32'h3bce2a9d),
	.w8(32'hba016d1d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0b3b1),
	.w1(32'h3bea10a6),
	.w2(32'hbb1f1450),
	.w3(32'h39e6cdca),
	.w4(32'hba318c2c),
	.w5(32'h3b20dd80),
	.w6(32'hbba89333),
	.w7(32'h3b46f75f),
	.w8(32'h3c5df6b7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd65dad),
	.w1(32'h3ab801e6),
	.w2(32'hbc722380),
	.w3(32'hbb9af2c4),
	.w4(32'hbc9406fa),
	.w5(32'hbb86a4cc),
	.w6(32'h3b9f261f),
	.w7(32'hbaf638db),
	.w8(32'h3bf21b8a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b121a2b),
	.w1(32'hbc597695),
	.w2(32'h3c052960),
	.w3(32'hbb6df84a),
	.w4(32'h3c9a203f),
	.w5(32'h3c6d549a),
	.w6(32'h3c1c2954),
	.w7(32'h3c9a9a00),
	.w8(32'hbbaeb9f6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7be5f7),
	.w1(32'h3b1520ed),
	.w2(32'h3b8913ee),
	.w3(32'hba482dfe),
	.w4(32'hbb04529e),
	.w5(32'h3c7a1587),
	.w6(32'h385cafa3),
	.w7(32'h3c3047bd),
	.w8(32'hba4c3ab4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389bb298),
	.w1(32'hbafe3d9d),
	.w2(32'h3c1fcd6f),
	.w3(32'hbb6272f2),
	.w4(32'h3c2d5ead),
	.w5(32'h3b7f3b9e),
	.w6(32'h3c011006),
	.w7(32'h3af4c0ec),
	.w8(32'h3abdf8bc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdec518),
	.w1(32'h3995ec2f),
	.w2(32'hbb60ff9d),
	.w3(32'h3c823e2e),
	.w4(32'h3a5d2d0f),
	.w5(32'hbb52581c),
	.w6(32'h394bd3a4),
	.w7(32'h3bc20b6d),
	.w8(32'h3bb1340c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44dae4),
	.w1(32'h39555616),
	.w2(32'h38abe694),
	.w3(32'h3abf3874),
	.w4(32'h3bb0c4d5),
	.w5(32'h3bf0defd),
	.w6(32'hbc02c6fe),
	.w7(32'hbb8706cb),
	.w8(32'h3ab45c13),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d5ada),
	.w1(32'h3c959b4f),
	.w2(32'hbbd29780),
	.w3(32'h3c3baa6a),
	.w4(32'hbabf9db7),
	.w5(32'h3ba18aec),
	.w6(32'hbb416548),
	.w7(32'hbab1f5fa),
	.w8(32'h3c7278b5),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a40ab),
	.w1(32'h3b46b673),
	.w2(32'h3aba2e7c),
	.w3(32'h3c32d76d),
	.w4(32'hbaa21db2),
	.w5(32'h3bac9f09),
	.w6(32'hbbbdd9e7),
	.w7(32'h3c7362f8),
	.w8(32'hbb4ed638),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a430b1f),
	.w1(32'hbba59aaf),
	.w2(32'hbb7b4c3c),
	.w3(32'hbc424a18),
	.w4(32'h3ad7b3fe),
	.w5(32'hba3b82ec),
	.w6(32'hbac03186),
	.w7(32'h3ba45666),
	.w8(32'hbc015cc8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4ba6c),
	.w1(32'hbba9765d),
	.w2(32'h3c0b18c4),
	.w3(32'hb8fb196d),
	.w4(32'hbc75652a),
	.w5(32'hbc000226),
	.w6(32'h3c23a9bd),
	.w7(32'h3ba913d3),
	.w8(32'h389a92bc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c954f),
	.w1(32'hb9e114db),
	.w2(32'hbbe4f737),
	.w3(32'hbc087cee),
	.w4(32'hbaf7ecd1),
	.w5(32'h3b897d89),
	.w6(32'hbba1052f),
	.w7(32'h3c01f194),
	.w8(32'hbb98cdfd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb428be3),
	.w1(32'h3c1ce6bf),
	.w2(32'h3c43c4fd),
	.w3(32'hbc101714),
	.w4(32'hbb68c730),
	.w5(32'h3c592233),
	.w6(32'hbb7554dd),
	.w7(32'h38aba226),
	.w8(32'h3b13f0dc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd741e7),
	.w1(32'hbbff6a44),
	.w2(32'hbaf1667e),
	.w3(32'hbc1cc434),
	.w4(32'h39d50c5a),
	.w5(32'h3bb430ee),
	.w6(32'hbc3ba77f),
	.w7(32'hbd066af7),
	.w8(32'h3c6d54c0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c6968),
	.w1(32'h3a8ae262),
	.w2(32'h3a7d7a7b),
	.w3(32'h3b6cb54c),
	.w4(32'hbb38a6ce),
	.w5(32'h3c04105b),
	.w6(32'hbadc1943),
	.w7(32'hbac60ded),
	.w8(32'h3b1f798b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc688734),
	.w1(32'h3b1886b0),
	.w2(32'hba2a1932),
	.w3(32'hba889a4a),
	.w4(32'hbae325c0),
	.w5(32'h3c4c90d7),
	.w6(32'h3bc7aae4),
	.w7(32'h3bda259a),
	.w8(32'hb9b0a694),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9891e1),
	.w1(32'h3b9366ef),
	.w2(32'h3c1c852e),
	.w3(32'h3ad937cf),
	.w4(32'h3b5e7ef8),
	.w5(32'hbc677563),
	.w6(32'hbc2eaef2),
	.w7(32'h3b8be124),
	.w8(32'h396bfeb5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8e7f),
	.w1(32'h3b0be851),
	.w2(32'h3b159738),
	.w3(32'hbbcbc13a),
	.w4(32'h3c0d269a),
	.w5(32'hba3d7ad2),
	.w6(32'hbb0fe3d3),
	.w7(32'hbb2ba156),
	.w8(32'h3b411734),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944a85d),
	.w1(32'h3aed47fc),
	.w2(32'hbb83dab0),
	.w3(32'h36db93d9),
	.w4(32'hbbcf21fc),
	.w5(32'hb9492f87),
	.w6(32'h3aa13566),
	.w7(32'hbba6a2c6),
	.w8(32'h3c384205),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ab31a),
	.w1(32'h3ad513c0),
	.w2(32'h3bd0cc5f),
	.w3(32'h3a4b1c70),
	.w4(32'h3b1fb834),
	.w5(32'h3a4e47a4),
	.w6(32'hbbd4d6f0),
	.w7(32'hbb691631),
	.w8(32'hbb91902a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a01fe),
	.w1(32'h3b90768d),
	.w2(32'h3b80d15c),
	.w3(32'h3b1264db),
	.w4(32'hbabfbc52),
	.w5(32'hbc98b8df),
	.w6(32'hbbb5b712),
	.w7(32'hbc2631e5),
	.w8(32'hbcadb614),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21f50f),
	.w1(32'h3c5465de),
	.w2(32'h3bb75d01),
	.w3(32'h3c548b3d),
	.w4(32'h3b3bf9fd),
	.w5(32'hbc37b3ab),
	.w6(32'hba1df044),
	.w7(32'hba49d6d5),
	.w8(32'h3a8dfe85),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7cd25),
	.w1(32'h3b10d056),
	.w2(32'h3b34d793),
	.w3(32'h3b28d011),
	.w4(32'h3b3f0097),
	.w5(32'hbb2d4cf3),
	.w6(32'hbc4a189b),
	.w7(32'hbba9c054),
	.w8(32'h3bfd7e53),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f1993a),
	.w1(32'h3beb1612),
	.w2(32'h3b8e1d3f),
	.w3(32'h3a33e564),
	.w4(32'h3ca77726),
	.w5(32'hbb356c42),
	.w6(32'h3c2b6e56),
	.w7(32'h3c11f962),
	.w8(32'h3add24eb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fe834),
	.w1(32'h390cc0e8),
	.w2(32'hbc1f738d),
	.w3(32'h3bee6486),
	.w4(32'hbab409c3),
	.w5(32'h3c18ab70),
	.w6(32'h3b6e3ffd),
	.w7(32'hbb5b2558),
	.w8(32'hbc0e8510),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e68cd),
	.w1(32'hbb79d230),
	.w2(32'h3b01c517),
	.w3(32'h3c44b741),
	.w4(32'h3aa6b99f),
	.w5(32'h3a266d11),
	.w6(32'hbc235e8c),
	.w7(32'hbb0280ee),
	.w8(32'h3b53295c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2475f),
	.w1(32'h3ae69fe4),
	.w2(32'h3c0e8601),
	.w3(32'hbb899633),
	.w4(32'h3bcd0bfc),
	.w5(32'h3ba0bd57),
	.w6(32'h3cafafda),
	.w7(32'h3ad55cbd),
	.w8(32'hbbd4eef2),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927a7e9),
	.w1(32'hbc416653),
	.w2(32'hbaae8b47),
	.w3(32'h3c168c03),
	.w4(32'h3b2cc9a9),
	.w5(32'h3b20e0d1),
	.w6(32'h3c35784d),
	.w7(32'hbbeb5ae8),
	.w8(32'h3b94513e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32d1c5),
	.w1(32'hbabd1b76),
	.w2(32'hbb87a432),
	.w3(32'h391db642),
	.w4(32'hba8b1d1f),
	.w5(32'h3b9c8dec),
	.w6(32'hba33247f),
	.w7(32'h3b19984b),
	.w8(32'hb9640c78),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1707c8),
	.w1(32'hbb3ef6c4),
	.w2(32'hbc48e76e),
	.w3(32'hbb30a4fe),
	.w4(32'h3c993e2d),
	.w5(32'hbbae780a),
	.w6(32'hba11522a),
	.w7(32'h3bb38035),
	.w8(32'hbb9e1163),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a7410),
	.w1(32'hbb5bde68),
	.w2(32'h3bf72187),
	.w3(32'hbbcb2e44),
	.w4(32'hba9b46df),
	.w5(32'hbadc7a3a),
	.w6(32'h3c2824da),
	.w7(32'hbba1d5d8),
	.w8(32'hbc01dcba),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d7976),
	.w1(32'hbb338c0a),
	.w2(32'hbb3f619f),
	.w3(32'hbb83a18e),
	.w4(32'hbbaf0cf2),
	.w5(32'h3b2138e9),
	.w6(32'hb9fa98d6),
	.w7(32'hbb6f0db4),
	.w8(32'hbcb1509d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf11c72),
	.w1(32'h3ca795c3),
	.w2(32'h3bab55d0),
	.w3(32'hbc414f27),
	.w4(32'h3b16876e),
	.w5(32'h3cc1345d),
	.w6(32'hbba14631),
	.w7(32'hbc74391d),
	.w8(32'h3b4dc4fd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9620d0),
	.w1(32'hba0b5a16),
	.w2(32'hbc12c32b),
	.w3(32'h3b8420e4),
	.w4(32'h3a8137e3),
	.w5(32'h3a738512),
	.w6(32'hbc046ab5),
	.w7(32'hbc1f3510),
	.w8(32'hbb7cca81),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c166e65),
	.w1(32'hb9cac2be),
	.w2(32'hbab4d4d4),
	.w3(32'h3ca96564),
	.w4(32'h3b712861),
	.w5(32'hbbe3523d),
	.w6(32'hba9800bf),
	.w7(32'hbb447bb3),
	.w8(32'h3c016b20),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule