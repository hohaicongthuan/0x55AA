module layer_10_featuremap_151(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06c568),
	.w1(32'h395b552f),
	.w2(32'hba61ba90),
	.w3(32'h3a2af285),
	.w4(32'h3a665eb1),
	.w5(32'h3a4d9463),
	.w6(32'h39e6511b),
	.w7(32'h3a23c807),
	.w8(32'h3a1d80d4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a213050),
	.w1(32'h39d73b37),
	.w2(32'h39f39c4c),
	.w3(32'h3a8dcc1a),
	.w4(32'h39b1427f),
	.w5(32'h39b5ef1b),
	.w6(32'h383db095),
	.w7(32'h39486d0c),
	.w8(32'hb9b83a51),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987da87),
	.w1(32'h39dc7506),
	.w2(32'h3a35eec4),
	.w3(32'hb7690e3a),
	.w4(32'hb95de886),
	.w5(32'hb9c50840),
	.w6(32'hb928fff3),
	.w7(32'h39847a9b),
	.w8(32'hb897cc51),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6f175),
	.w1(32'hba327023),
	.w2(32'hba7ad0a7),
	.w3(32'hba1630f9),
	.w4(32'hbabafcff),
	.w5(32'hba8dd740),
	.w6(32'h3a523565),
	.w7(32'h3aa25c0e),
	.w8(32'h3a1d09a7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9552313),
	.w1(32'h397cb729),
	.w2(32'hb9b0d38b),
	.w3(32'hba78d1a9),
	.w4(32'h3941944e),
	.w5(32'hb98ba77a),
	.w6(32'h3928ebcd),
	.w7(32'h379835ad),
	.w8(32'h3a07ca5c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cd8149),
	.w1(32'h3a1bf647),
	.w2(32'h3a4295d5),
	.w3(32'hb96c5df5),
	.w4(32'h3a5b2868),
	.w5(32'h3a46aace),
	.w6(32'h39b2901d),
	.w7(32'h393f5158),
	.w8(32'h3973d664),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad522ab),
	.w1(32'h3a17e5b7),
	.w2(32'hba1f3cde),
	.w3(32'h3abec024),
	.w4(32'hb82d1397),
	.w5(32'hba7f148c),
	.w6(32'h398274d9),
	.w7(32'h38749e77),
	.w8(32'hba437be5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83cb22),
	.w1(32'hba5b30c5),
	.w2(32'hbacbb3cd),
	.w3(32'hbafd3a86),
	.w4(32'hbacdf006),
	.w5(32'hbad6230d),
	.w6(32'hba0d93cd),
	.w7(32'hbab9b762),
	.w8(32'hba9eb6ca),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a256ff5),
	.w1(32'h39f11e7b),
	.w2(32'hb9926b3b),
	.w3(32'h3a86a22e),
	.w4(32'h39979bcc),
	.w5(32'hba03bc9e),
	.w6(32'h3a341fec),
	.w7(32'hb9c29a2e),
	.w8(32'hba2a658b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bc4c3),
	.w1(32'hba376525),
	.w2(32'hbb555e81),
	.w3(32'hba835e10),
	.w4(32'hb9af9cb4),
	.w5(32'hbb3601eb),
	.w6(32'hbad91d8a),
	.w7(32'hba9ae40f),
	.w8(32'hbb5090ad),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d1a05a),
	.w1(32'h3a8ab8b3),
	.w2(32'h3a911521),
	.w3(32'hb87885d8),
	.w4(32'h3a1b7396),
	.w5(32'h3a4d9ad6),
	.w6(32'h3982e25f),
	.w7(32'h39e0f101),
	.w8(32'h39a4f667),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac41da2),
	.w1(32'h3adcd76a),
	.w2(32'h3881f376),
	.w3(32'h3ab79c65),
	.w4(32'h3b05957c),
	.w5(32'h3aa9fd9d),
	.w6(32'h3a2dac60),
	.w7(32'h3addf145),
	.w8(32'h38d50d53),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1450b3),
	.w1(32'hb9d4fc1e),
	.w2(32'hbb0ab2f9),
	.w3(32'hba3d3c53),
	.w4(32'hba882bbf),
	.w5(32'hbb18fcc1),
	.w6(32'hba46b641),
	.w7(32'hba97d33c),
	.w8(32'hbb0e6484),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab91145),
	.w1(32'h3ab592d4),
	.w2(32'h3a681812),
	.w3(32'h3aa5345e),
	.w4(32'h3aa6a9e6),
	.w5(32'h3a2ca6be),
	.w6(32'h3ac6b047),
	.w7(32'h3a4aff0a),
	.w8(32'h3a2e1dc9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34284d),
	.w1(32'hba22371d),
	.w2(32'hbb3ba2d6),
	.w3(32'h3a1ec27c),
	.w4(32'h3a4e7eb8),
	.w5(32'hba548476),
	.w6(32'h3a2c4971),
	.w7(32'h3ac67f31),
	.w8(32'h392a81a0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba217703),
	.w1(32'hb990f428),
	.w2(32'hbb03d99c),
	.w3(32'hba47dadf),
	.w4(32'hba431040),
	.w5(32'hbb059580),
	.w6(32'hba5e7863),
	.w7(32'hba9134db),
	.w8(32'hbb2cbb76),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b03b4),
	.w1(32'h3a72b607),
	.w2(32'h3a89e383),
	.w3(32'h38e2bd8e),
	.w4(32'h398bd072),
	.w5(32'hb99bd5f1),
	.w6(32'h39a5f89f),
	.w7(32'hb6c47442),
	.w8(32'hba2a55db),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f99e7d),
	.w1(32'hbac79758),
	.w2(32'hbb395c8e),
	.w3(32'hba1fbc61),
	.w4(32'hbb03c75f),
	.w5(32'hbb2de7ce),
	.w6(32'hba9a3840),
	.w7(32'hbade9726),
	.w8(32'hbb3fbd21),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a547a5d),
	.w1(32'hba8f43d4),
	.w2(32'hbb0524ca),
	.w3(32'hb8da9fd4),
	.w4(32'hbad7b43d),
	.w5(32'hbb26bd9b),
	.w6(32'hb995697d),
	.w7(32'hbab0c309),
	.w8(32'hbb154c84),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c37308),
	.w1(32'h3a1d416f),
	.w2(32'h398fe05b),
	.w3(32'hb9c5db6f),
	.w4(32'h39c20317),
	.w5(32'h39106ef8),
	.w6(32'h39f5d894),
	.w7(32'h391b547a),
	.w8(32'h38b344bf),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb716dbc5),
	.w1(32'h385fe1f5),
	.w2(32'hb917469d),
	.w3(32'h388a03e6),
	.w4(32'hb8862666),
	.w5(32'hb760d80f),
	.w6(32'hb940de76),
	.w7(32'hb9af9a98),
	.w8(32'hb9862917),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c9e3d7),
	.w1(32'h3abac384),
	.w2(32'h3a4324c5),
	.w3(32'h39d83812),
	.w4(32'h399e5998),
	.w5(32'hb9446b68),
	.w6(32'h3b3e0a73),
	.w7(32'h3b5d0c07),
	.w8(32'h3a8abe2f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b711a31),
	.w1(32'h3ae58e0c),
	.w2(32'hbb09ce3e),
	.w3(32'hb92dcb02),
	.w4(32'hb9fa3d82),
	.w5(32'hbb572959),
	.w6(32'hba6332d8),
	.w7(32'hba080202),
	.w8(32'hbb85ad23),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0ecf3),
	.w1(32'h3a0bd4fd),
	.w2(32'hbb01e0a9),
	.w3(32'h3a90da64),
	.w4(32'h3a8d510e),
	.w5(32'hbacc3c4f),
	.w6(32'h3a0a40aa),
	.w7(32'h3a6d9123),
	.w8(32'hbac0b384),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e29c5d),
	.w1(32'h38d38e62),
	.w2(32'hba9ffa4b),
	.w3(32'hba174aac),
	.w4(32'hb879accd),
	.w5(32'hba76bf69),
	.w6(32'hbaffbd50),
	.w7(32'hba405145),
	.w8(32'hbb0ba358),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9294583),
	.w1(32'h39e9c37a),
	.w2(32'h3a18fd55),
	.w3(32'h36a66b1c),
	.w4(32'h395c9675),
	.w5(32'h390fc2d4),
	.w6(32'h390dd11d),
	.w7(32'h38c64383),
	.w8(32'hb922581c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a704214),
	.w1(32'h39d9ead5),
	.w2(32'h399e0da8),
	.w3(32'h398f086a),
	.w4(32'h399939a0),
	.w5(32'h396d7c67),
	.w6(32'h39dd161a),
	.w7(32'h3986b107),
	.w8(32'h39a38ee5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6850fb),
	.w1(32'hba3537a2),
	.w2(32'hba6f91a3),
	.w3(32'h3a3d084f),
	.w4(32'hba420589),
	.w5(32'h3989c71e),
	.w6(32'h394899d6),
	.w7(32'hba54c5e2),
	.w8(32'hb9e11d4d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999615d),
	.w1(32'h392a903a),
	.w2(32'h39a3fc0b),
	.w3(32'h39813627),
	.w4(32'h3811f7ce),
	.w5(32'hb929bfe8),
	.w6(32'hba98bfba),
	.w7(32'h392e9722),
	.w8(32'h398e63c9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63d811),
	.w1(32'hba0b70a6),
	.w2(32'hbac18d8f),
	.w3(32'h396f7ac1),
	.w4(32'hba97f4b6),
	.w5(32'hbb261b77),
	.w6(32'hba8b11bf),
	.w7(32'hba6a1fda),
	.w8(32'hbb28ba6b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9861f0a),
	.w1(32'h39002bb7),
	.w2(32'h395a618d),
	.w3(32'hba27b848),
	.w4(32'h392bf0ee),
	.w5(32'h39375bd4),
	.w6(32'h38bb6a92),
	.w7(32'hb857c3ce),
	.w8(32'hb8ab5350),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386ecf37),
	.w1(32'h39ae8826),
	.w2(32'h3a01e90b),
	.w3(32'h3962c6c5),
	.w4(32'h39afc868),
	.w5(32'h39f48e38),
	.w6(32'h3a090f5c),
	.w7(32'h39cc4e45),
	.w8(32'h39c4d7e4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7edb3e),
	.w1(32'h3882a0ab),
	.w2(32'hbaa46495),
	.w3(32'h3a87e8eb),
	.w4(32'h398267da),
	.w5(32'hbad42b36),
	.w6(32'h39e72104),
	.w7(32'h3a066f20),
	.w8(32'hb9c3a654),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba595722),
	.w1(32'h3916aeab),
	.w2(32'hb9a12549),
	.w3(32'hbab26d64),
	.w4(32'h39e72490),
	.w5(32'h399ec032),
	.w6(32'hb9dd87a5),
	.w7(32'hb9ab28fa),
	.w8(32'hb969decd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08375f),
	.w1(32'hb917d4b9),
	.w2(32'hb9240650),
	.w3(32'hb886f9ad),
	.w4(32'hb6e91c33),
	.w5(32'h391352b2),
	.w6(32'hba1715a5),
	.w7(32'hba2e6d8e),
	.w8(32'hba6a9206),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b9cdf),
	.w1(32'h392677d2),
	.w2(32'hb98bdb97),
	.w3(32'h398ee9e5),
	.w4(32'h39153295),
	.w5(32'hb92415d1),
	.w6(32'h39a25676),
	.w7(32'h398f9eb6),
	.w8(32'hb9857a9e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f0ffa2),
	.w1(32'h3a71fc59),
	.w2(32'hbb086fca),
	.w3(32'h3a5e1a5f),
	.w4(32'h3aa2e136),
	.w5(32'hba9bddce),
	.w6(32'hba879338),
	.w7(32'h3aae2722),
	.w8(32'hbaad64db),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72595b),
	.w1(32'h3b1507e1),
	.w2(32'h3aae2d66),
	.w3(32'hb8c87277),
	.w4(32'h3b85de47),
	.w5(32'h3b09b866),
	.w6(32'hbb06ba27),
	.w7(32'h3b079d5c),
	.w8(32'h3a725d76),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c0048),
	.w1(32'h3af18491),
	.w2(32'h3ae418b1),
	.w3(32'hba780bcf),
	.w4(32'h3b005b50),
	.w5(32'h3adf2cad),
	.w6(32'hba9725ab),
	.w7(32'h39e2dba7),
	.w8(32'h39e5e994),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e51dcf),
	.w1(32'h3a2157d8),
	.w2(32'h38a7a61d),
	.w3(32'h3a2e9ec5),
	.w4(32'h3a828ffc),
	.w5(32'h39fb2732),
	.w6(32'hb9c14e9a),
	.w7(32'h39862636),
	.w8(32'h384b84d8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38660120),
	.w1(32'hb8c916f4),
	.w2(32'hb8617e1c),
	.w3(32'h389a2576),
	.w4(32'hba15499c),
	.w5(32'hb9fb9360),
	.w6(32'hb70165e3),
	.w7(32'hb8dfe68d),
	.w8(32'hb9690aea),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974b4c3),
	.w1(32'hb977dbcc),
	.w2(32'h3991d5ef),
	.w3(32'hb9fc720c),
	.w4(32'hb94ae4cc),
	.w5(32'h391cc509),
	.w6(32'hb8a1a935),
	.w7(32'h39029f0f),
	.w8(32'h383f5eb3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967ea49),
	.w1(32'h3a64c828),
	.w2(32'h3a15a082),
	.w3(32'h3923dc56),
	.w4(32'h3a9f8220),
	.w5(32'h3a0d20f7),
	.w6(32'h3a28c071),
	.w7(32'h3ab397fa),
	.w8(32'h38c5100f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70206d),
	.w1(32'hba839437),
	.w2(32'hbb586dac),
	.w3(32'hb926e2a2),
	.w4(32'hba18236c),
	.w5(32'hbb3d68aa),
	.w6(32'hbb175f24),
	.w7(32'hbb29166c),
	.w8(32'hbb938e04),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27db84),
	.w1(32'hb9ddfb37),
	.w2(32'hbb1b3d56),
	.w3(32'h397db661),
	.w4(32'h39e2de9e),
	.w5(32'hbaeed0df),
	.w6(32'hb9e2c463),
	.w7(32'h3a82db79),
	.w8(32'hbab344a4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecde21),
	.w1(32'hb931843b),
	.w2(32'hbb44258f),
	.w3(32'hba02a129),
	.w4(32'h383da3f6),
	.w5(32'hbb3f4373),
	.w6(32'hba46f7d3),
	.w7(32'h389d85f7),
	.w8(32'hbb3fc5af),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba014ee4),
	.w1(32'hb9f2c3e2),
	.w2(32'hbb26070a),
	.w3(32'hb94045b6),
	.w4(32'hb9264968),
	.w5(32'hb9e14921),
	.w6(32'h3a26123d),
	.w7(32'h3a5d8e67),
	.w8(32'hba36ab8f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a866220),
	.w1(32'hba3d3af9),
	.w2(32'hbb474f41),
	.w3(32'hbab0bd1a),
	.w4(32'hbb3beb2c),
	.w5(32'hbb83614f),
	.w6(32'hbb287c92),
	.w7(32'hbb9018e5),
	.w8(32'hbb991b53),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8aa11),
	.w1(32'h39f1d750),
	.w2(32'h39e08b6a),
	.w3(32'h399ec617),
	.w4(32'h39a224bd),
	.w5(32'h39238405),
	.w6(32'h3a2feb7c),
	.w7(32'h399f3858),
	.w8(32'h394b0361),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a72850),
	.w1(32'h37a18448),
	.w2(32'hb7685a30),
	.w3(32'h3921c430),
	.w4(32'h38d0217f),
	.w5(32'hb90e8340),
	.w6(32'h394c1a93),
	.w7(32'h390dd254),
	.w8(32'h38aa24fa),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14ab33),
	.w1(32'hb9831bcd),
	.w2(32'hb9ba8d30),
	.w3(32'h39fc5525),
	.w4(32'hb9b541dc),
	.w5(32'hba04c160),
	.w6(32'hba29f438),
	.w7(32'hba85471d),
	.w8(32'hba702cc0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8df238),
	.w1(32'hb7c251a4),
	.w2(32'hbaa53a35),
	.w3(32'hba987dac),
	.w4(32'hb9cab2d2),
	.w5(32'hb7963268),
	.w6(32'hb9ed13c2),
	.w7(32'hba35ff8f),
	.w8(32'hba91c5be),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bd9a3),
	.w1(32'h3a3b0828),
	.w2(32'h39d1b84e),
	.w3(32'hb9e8a951),
	.w4(32'h3a1ba54b),
	.w5(32'h39ba8fb5),
	.w6(32'h38f161d4),
	.w7(32'h37e17212),
	.w8(32'hb9ecf13e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c78d5),
	.w1(32'hbacc69cf),
	.w2(32'hbb871a05),
	.w3(32'h389dda3b),
	.w4(32'hba93e9a2),
	.w5(32'hbb7daec6),
	.w6(32'hba8545b2),
	.w7(32'hbaad5c2a),
	.w8(32'hbb28000e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb903d3c3),
	.w1(32'h37d65248),
	.w2(32'hb6057bce),
	.w3(32'hb98f11da),
	.w4(32'h39aba7d4),
	.w5(32'h390b10a9),
	.w6(32'hb997b4a0),
	.w7(32'hb9002080),
	.w8(32'hb9392135),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880a115),
	.w1(32'hb9c83d0e),
	.w2(32'h38814930),
	.w3(32'h38d7a6e0),
	.w4(32'hba48d9f2),
	.w5(32'hb9e2b7ae),
	.w6(32'hb86af67f),
	.w7(32'h3984a8c4),
	.w8(32'hb7fd5282),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b00cb7),
	.w1(32'hb9d0e83a),
	.w2(32'hb9c28618),
	.w3(32'hb9cddcb4),
	.w4(32'hba7da66d),
	.w5(32'hba9a97ab),
	.w6(32'hba162a16),
	.w7(32'hba33de73),
	.w8(32'hba3b143d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccbe3f),
	.w1(32'h3998c0f3),
	.w2(32'hb91a6a7c),
	.w3(32'hba33242d),
	.w4(32'h39ad8b1e),
	.w5(32'hb953a161),
	.w6(32'hb8881b7f),
	.w7(32'hb8e73d93),
	.w8(32'h38e0eb64),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba136db6),
	.w1(32'h38c79846),
	.w2(32'h39d561b4),
	.w3(32'hb9a901b2),
	.w4(32'h38089ea9),
	.w5(32'h370a415a),
	.w6(32'hb962a731),
	.w7(32'h39f32fc4),
	.w8(32'hb8885317),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dcc6b),
	.w1(32'h3a15e7c6),
	.w2(32'h39615141),
	.w3(32'hb91344ae),
	.w4(32'h3a1fd52c),
	.w5(32'h395f9c91),
	.w6(32'h3a23e0be),
	.w7(32'h39cdbb06),
	.w8(32'h38b558a6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa1f71),
	.w1(32'hb9f8d0ee),
	.w2(32'hba75915b),
	.w3(32'hb978ef21),
	.w4(32'hb9860de7),
	.w5(32'hba8bc6e3),
	.w6(32'hba91adc4),
	.w7(32'hb8157015),
	.w8(32'hba085e12),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56f5d2),
	.w1(32'hb9d3dd06),
	.w2(32'hba5e8d7e),
	.w3(32'hba8bd4aa),
	.w4(32'hb98e5629),
	.w5(32'hba6f3ff2),
	.w6(32'hba2d6bb4),
	.w7(32'hb98bca6b),
	.w8(32'hba41cc66),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984af5e),
	.w1(32'h38a0a773),
	.w2(32'hba30f001),
	.w3(32'hb861bea6),
	.w4(32'h39a0becf),
	.w5(32'hba23e387),
	.w6(32'h390500eb),
	.w7(32'hb9947348),
	.w8(32'h39b83621),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396721db),
	.w1(32'hb684a2a3),
	.w2(32'hb95bc065),
	.w3(32'hba3e6ac6),
	.w4(32'h39cdca9c),
	.w5(32'h393924bc),
	.w6(32'hb9f8ac43),
	.w7(32'hba07fabe),
	.w8(32'hba10d4f7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ecd780),
	.w1(32'hb9bb66d1),
	.w2(32'hb91c1b99),
	.w3(32'h3895614f),
	.w4(32'hb956f6d8),
	.w5(32'hb9bdd7d0),
	.w6(32'hb969d213),
	.w7(32'h39355894),
	.w8(32'h38943ec0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89dc220),
	.w1(32'h389980f6),
	.w2(32'hba0a12d1),
	.w3(32'hb980d6e8),
	.w4(32'h39340a02),
	.w5(32'hba70bbfe),
	.w6(32'hb8c6c384),
	.w7(32'hba2faf12),
	.w8(32'hba086bde),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8747c),
	.w1(32'hba473635),
	.w2(32'hbad94c73),
	.w3(32'hba7c8844),
	.w4(32'hbad1e560),
	.w5(32'hbb08821f),
	.w6(32'hba8429f3),
	.w7(32'hbaa91ee4),
	.w8(32'hbafb28a7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8a284),
	.w1(32'h39f903ad),
	.w2(32'hbb0458ea),
	.w3(32'hba1c91f0),
	.w4(32'h39031c62),
	.w5(32'hbb150ed3),
	.w6(32'h3a1d8c3e),
	.w7(32'h3a6f7cd5),
	.w8(32'hbac1c05f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f9602),
	.w1(32'h3a697f81),
	.w2(32'hb9610784),
	.w3(32'hb88cca52),
	.w4(32'h3ae9a900),
	.w5(32'h3a0d677b),
	.w6(32'hb9078af1),
	.w7(32'h3abbd776),
	.w8(32'h3916638e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83c78e),
	.w1(32'h3abe2f67),
	.w2(32'hbb1c0254),
	.w3(32'h3ada93f9),
	.w4(32'h3b0a9cb5),
	.w5(32'hba9e4bc0),
	.w6(32'hba158ac3),
	.w7(32'h3a1e1c97),
	.w8(32'hbb253240),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c5d70),
	.w1(32'h38112c2b),
	.w2(32'h39c74cc8),
	.w3(32'hba2a9e6d),
	.w4(32'hb9323022),
	.w5(32'h38818533),
	.w6(32'hb6df78ec),
	.w7(32'h380ae790),
	.w8(32'hb984e877),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38af1a8f),
	.w1(32'h39ba8b21),
	.w2(32'h3a06cc19),
	.w3(32'hb89ac06d),
	.w4(32'h399f07b1),
	.w5(32'h39d46287),
	.w6(32'h39d73139),
	.w7(32'h39eb6789),
	.w8(32'h39b39b03),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399745b5),
	.w1(32'h39f9ecc9),
	.w2(32'h39dc042a),
	.w3(32'h39eb99f7),
	.w4(32'h39d390e9),
	.w5(32'h39c258c3),
	.w6(32'h3a049801),
	.w7(32'h39a51e62),
	.w8(32'h3981c25c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad1961),
	.w1(32'h3a0e8dd5),
	.w2(32'h3997873c),
	.w3(32'h397468ab),
	.w4(32'h3a2e85f6),
	.w5(32'h39cea696),
	.w6(32'h391e02d0),
	.w7(32'h398a9d6c),
	.w8(32'h38964591),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2055fa),
	.w1(32'hb972a9a5),
	.w2(32'h388af11a),
	.w3(32'h3a5079ce),
	.w4(32'hb9ea1fd8),
	.w5(32'hb8669375),
	.w6(32'hb96e0f67),
	.w7(32'hb90b039a),
	.w8(32'hb955cc01),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393453af),
	.w1(32'hba4a38c8),
	.w2(32'hba07edeb),
	.w3(32'hb9b5bbd6),
	.w4(32'hba2bdd24),
	.w5(32'h3a8598b5),
	.w6(32'h3a059b23),
	.w7(32'h37836a57),
	.w8(32'hba04682f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e1305),
	.w1(32'hb9ec6854),
	.w2(32'hbaee0708),
	.w3(32'hba7b538f),
	.w4(32'hb9fae3bc),
	.w5(32'hbac31703),
	.w6(32'hba5a7cae),
	.w7(32'hb9b99fa4),
	.w8(32'hba9f68b1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba612bff),
	.w1(32'hbb0e8ded),
	.w2(32'hbb4317e4),
	.w3(32'hbac15a10),
	.w4(32'hbb365a3d),
	.w5(32'hbb495b52),
	.w6(32'hbb4833ff),
	.w7(32'hbb2bc487),
	.w8(32'hbb336c0e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba375b4a),
	.w1(32'h39bcb893),
	.w2(32'hba69c8c4),
	.w3(32'hba86fdbc),
	.w4(32'h3a179da6),
	.w5(32'hba8b6d0f),
	.w6(32'hb91ccd86),
	.w7(32'hba1b49da),
	.w8(32'hba005265),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab12146),
	.w1(32'h39fd9ac5),
	.w2(32'hba6f733f),
	.w3(32'h3a056ec2),
	.w4(32'hb8f004e6),
	.w5(32'hbaaf1005),
	.w6(32'h3989d588),
	.w7(32'hb9942dec),
	.w8(32'hba86c8f0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1650b3),
	.w1(32'hb9ab78ce),
	.w2(32'hba717b8f),
	.w3(32'hb900916d),
	.w4(32'hb876d407),
	.w5(32'hba1a2d0e),
	.w6(32'hb88a8847),
	.w7(32'h392f684a),
	.w8(32'hb9360697),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e53008),
	.w1(32'hba323b29),
	.w2(32'hbaca12d5),
	.w3(32'hb9fbe7aa),
	.w4(32'hba9ab0dc),
	.w5(32'hbafedb0f),
	.w6(32'hba9dc747),
	.w7(32'hba7fd905),
	.w8(32'hbadc6960),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdf56e),
	.w1(32'h39c29c14),
	.w2(32'h39e14273),
	.w3(32'hb96f6ab2),
	.w4(32'h385ceab6),
	.w5(32'h38b35ed7),
	.w6(32'h392133d2),
	.w7(32'h38715079),
	.w8(32'hb955d55f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a83ff),
	.w1(32'h36d4826c),
	.w2(32'h396e148a),
	.w3(32'h39260dd6),
	.w4(32'hb8a8562c),
	.w5(32'h39492e8f),
	.w6(32'hb86672ad),
	.w7(32'h39bb4d6a),
	.w8(32'h39357f33),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981274d),
	.w1(32'h3a295899),
	.w2(32'h3a2bac79),
	.w3(32'h3985fc9c),
	.w4(32'h39fe9443),
	.w5(32'h3a7b7394),
	.w6(32'h3a150bbe),
	.w7(32'hb91945c8),
	.w8(32'h39aaa553),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e055cd),
	.w1(32'hba4c7472),
	.w2(32'hb9d60843),
	.w3(32'h3a8171f9),
	.w4(32'hba95e64b),
	.w5(32'hba8060bd),
	.w6(32'hba4464cd),
	.w7(32'hba006337),
	.w8(32'hba5b3432),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4205b),
	.w1(32'h3a7bdb35),
	.w2(32'hb78f1c2c),
	.w3(32'hba98d21d),
	.w4(32'h3ae8f093),
	.w5(32'h3a94ea7f),
	.w6(32'hba5f2e59),
	.w7(32'h3a1c4f2a),
	.w8(32'h384ed401),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5d929),
	.w1(32'h39a10c50),
	.w2(32'h39752cba),
	.w3(32'hba2450ea),
	.w4(32'h395beb6d),
	.w5(32'h396101cd),
	.w6(32'hb90d5426),
	.w7(32'h35fe2390),
	.w8(32'hb9167ccc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20bb47),
	.w1(32'hb8c3792d),
	.w2(32'hbab44701),
	.w3(32'h3a0ac6e3),
	.w4(32'h3890f5c4),
	.w5(32'hba83902e),
	.w6(32'h385071f3),
	.w7(32'h38e25d3b),
	.w8(32'hba9997ae),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab46647),
	.w1(32'hbb0e4ac1),
	.w2(32'hbb11e6b4),
	.w3(32'hbb20d4bb),
	.w4(32'hbafefcb0),
	.w5(32'hbae40f05),
	.w6(32'hbb246146),
	.w7(32'hbb117e40),
	.w8(32'hbadd0d86),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381fefe4),
	.w1(32'h3a6e2417),
	.w2(32'h39f0f84c),
	.w3(32'h3949b931),
	.w4(32'h3ac7dd15),
	.w5(32'h3a4f7389),
	.w6(32'hb7f8866c),
	.w7(32'h3a3237cb),
	.w8(32'h3812f6e7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ae281),
	.w1(32'hb9a436be),
	.w2(32'hba8d4e66),
	.w3(32'hb9a1d4a2),
	.w4(32'hb6e24156),
	.w5(32'hba95d30f),
	.w6(32'hbaa1d110),
	.w7(32'hba7d8815),
	.w8(32'hbb0464fe),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f836e7),
	.w1(32'hb8fa3208),
	.w2(32'hba143f4c),
	.w3(32'h39a7aa57),
	.w4(32'h39cfc78e),
	.w5(32'hb9986983),
	.w6(32'hb7508561),
	.w7(32'h39a240a8),
	.w8(32'hb9c19cfd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb970f410),
	.w1(32'hb9dc9734),
	.w2(32'hbb271cce),
	.w3(32'h36b63462),
	.w4(32'hb8d6bdd6),
	.w5(32'hbabf9c8e),
	.w6(32'h3a084620),
	.w7(32'h3918b8f5),
	.w8(32'hbaabcb68),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8396cc),
	.w1(32'h3a75f345),
	.w2(32'h3928ac12),
	.w3(32'h3a31710a),
	.w4(32'h3a2e9d16),
	.w5(32'h392118cd),
	.w6(32'h39f3dbf0),
	.w7(32'h3a11eba8),
	.w8(32'h38940bcc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75ed4e),
	.w1(32'h3950ccbd),
	.w2(32'hb8daa493),
	.w3(32'h397aed99),
	.w4(32'h3ac94861),
	.w5(32'hb99a7744),
	.w6(32'hba37f68c),
	.w7(32'hb9acd4df),
	.w8(32'hba839d5b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3abab),
	.w1(32'hb8088956),
	.w2(32'hb8d74fe8),
	.w3(32'h3a1e6e46),
	.w4(32'hb8fbe1d4),
	.w5(32'h39aacc6f),
	.w6(32'hb8a6240a),
	.w7(32'h390ad8df),
	.w8(32'h3a1f403a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd027b),
	.w1(32'hba8e9a26),
	.w2(32'hbb6ebdfc),
	.w3(32'hb998d04f),
	.w4(32'hbab20a38),
	.w5(32'hbb311155),
	.w6(32'hba4b225d),
	.w7(32'hbaab0f61),
	.w8(32'hbb31bef0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9b941),
	.w1(32'h3ac5c0a2),
	.w2(32'hb9a7e01e),
	.w3(32'hb933f498),
	.w4(32'h3ab5ead2),
	.w5(32'hb8dea2ce),
	.w6(32'h3912edec),
	.w7(32'h3a323a24),
	.w8(32'hba5cd2e2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fe3cc),
	.w1(32'h38fb0b63),
	.w2(32'hbacf7889),
	.w3(32'hbb05063f),
	.w4(32'hbaa64178),
	.w5(32'hbae969ab),
	.w6(32'hbb474744),
	.w7(32'hba81a317),
	.w8(32'hbb364478),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b268e26),
	.w1(32'h3ba8ded5),
	.w2(32'h3a822ec1),
	.w3(32'h3aceb6a3),
	.w4(32'h3bc42333),
	.w5(32'h3ad2a9c6),
	.w6(32'hba160d95),
	.w7(32'h3b56ad68),
	.w8(32'h3ac4d388),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88327c),
	.w1(32'hba71993b),
	.w2(32'hbb29d11c),
	.w3(32'hbb027f22),
	.w4(32'hba2fa761),
	.w5(32'hbb1a3522),
	.w6(32'hba8595b1),
	.w7(32'hba555a37),
	.w8(32'hbb5dfe5b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbe516),
	.w1(32'h3b275c00),
	.w2(32'hb9dbc923),
	.w3(32'h3aa589fc),
	.w4(32'h3b397807),
	.w5(32'h399cc1d4),
	.w6(32'h3ae95648),
	.w7(32'h3af1b201),
	.w8(32'h39e71f64),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a746c15),
	.w1(32'h39cc69d1),
	.w2(32'h39c5c436),
	.w3(32'h3a95f4dc),
	.w4(32'h3925f3f7),
	.w5(32'h38d62946),
	.w6(32'h3a126303),
	.w7(32'h395517c4),
	.w8(32'h39cac7dd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba822362),
	.w1(32'hb99d2e73),
	.w2(32'hbb0a4f14),
	.w3(32'hba55ea5a),
	.w4(32'h38c6fb43),
	.w5(32'hbad11df3),
	.w6(32'hba0cfa7a),
	.w7(32'hb97b06dc),
	.w8(32'hba05113e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba017250),
	.w1(32'h3a605459),
	.w2(32'hb8c240fd),
	.w3(32'hb91da8a8),
	.w4(32'h3a130557),
	.w5(32'hba70fe0a),
	.w6(32'h39c3a1ef),
	.w7(32'h3a89a66b),
	.w8(32'hb9998e83),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37efe6eb),
	.w1(32'h399b0e7f),
	.w2(32'h3a29e5fb),
	.w3(32'hb834a90f),
	.w4(32'hb960b2c6),
	.w5(32'hb91361d1),
	.w6(32'hb7d5e03f),
	.w7(32'h39acf8cf),
	.w8(32'h37b8cca2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdb8b8),
	.w1(32'h387f4b5f),
	.w2(32'hb8977093),
	.w3(32'hb9949282),
	.w4(32'h39134b25),
	.w5(32'h36787c53),
	.w6(32'hb9a2ce3a),
	.w7(32'hb9b7c7e3),
	.w8(32'hb9d78346),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03200c),
	.w1(32'hba30b818),
	.w2(32'hbb308cf9),
	.w3(32'hb9a3cd3c),
	.w4(32'hba960d45),
	.w5(32'hbb2c092a),
	.w6(32'hbaa19a62),
	.w7(32'hbb008c5c),
	.w8(32'hbb333b92),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96823ac),
	.w1(32'hbaacfdf4),
	.w2(32'hbaf2a51e),
	.w3(32'hb93e7b42),
	.w4(32'hba97c9ba),
	.w5(32'hbad814ae),
	.w6(32'hbaabcf6d),
	.w7(32'hba072ea5),
	.w8(32'hbaf9d50c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96f2c7),
	.w1(32'h39107757),
	.w2(32'hba1e76e2),
	.w3(32'h39853f69),
	.w4(32'h38becb2c),
	.w5(32'hb855ce21),
	.w6(32'hb8b624c4),
	.w7(32'hba7f8786),
	.w8(32'hbae4ccc6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa31ac),
	.w1(32'h393f9170),
	.w2(32'hbaadfc8e),
	.w3(32'h3a883864),
	.w4(32'h398d601c),
	.w5(32'hb9358941),
	.w6(32'h37280a9d),
	.w7(32'hb9b5425c),
	.w8(32'hb97d919d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aa23d),
	.w1(32'h3ac95732),
	.w2(32'h3a3af8eb),
	.w3(32'h370318ec),
	.w4(32'h3ac636bb),
	.w5(32'h3a4cd70f),
	.w6(32'h3907daa6),
	.w7(32'h3a4eefc9),
	.w8(32'hb8e72c31),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee0b63),
	.w1(32'hba9d1575),
	.w2(32'hbae62b81),
	.w3(32'hb909102a),
	.w4(32'hba9212ee),
	.w5(32'hbafcf8aa),
	.w6(32'hba1b638f),
	.w7(32'hb9ce9709),
	.w8(32'hbae8db57),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d2e19e),
	.w1(32'hb99a2b6e),
	.w2(32'hba7947a9),
	.w3(32'hba281396),
	.w4(32'hb9be66ad),
	.w5(32'hba74637c),
	.w6(32'hb9a09ee1),
	.w7(32'hb9b8ccf5),
	.w8(32'hba9a9ee2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c39ae),
	.w1(32'h3a3bca91),
	.w2(32'h398277e1),
	.w3(32'h3983b275),
	.w4(32'h3a5d5c5a),
	.w5(32'h39842b72),
	.w6(32'h39f2f1ba),
	.w7(32'h39697fba),
	.w8(32'h3a0104ec),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da222b),
	.w1(32'h398c792a),
	.w2(32'h39a95676),
	.w3(32'h3a166565),
	.w4(32'h39a1a02c),
	.w5(32'h39999593),
	.w6(32'h395b18b0),
	.w7(32'h394b2439),
	.w8(32'h399fd1f5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cfc9c),
	.w1(32'h39fe19c9),
	.w2(32'h39abcf07),
	.w3(32'h3a1093b5),
	.w4(32'h39efcb70),
	.w5(32'h39b29f29),
	.w6(32'h39404af4),
	.w7(32'h3944a66d),
	.w8(32'h39b01b64),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3999a),
	.w1(32'h3a4c6c32),
	.w2(32'h37366ca8),
	.w3(32'h3a2364c9),
	.w4(32'h3a6623c3),
	.w5(32'h394c8010),
	.w6(32'h3a8cb191),
	.w7(32'h3abc159e),
	.w8(32'h3a72e185),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a406d0f),
	.w1(32'hb9172f61),
	.w2(32'hbacd5f96),
	.w3(32'h39e7630b),
	.w4(32'h39885d1f),
	.w5(32'hbafecb80),
	.w6(32'hb9baca91),
	.w7(32'hb901a210),
	.w8(32'hbababd3c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d0def),
	.w1(32'h3900bcff),
	.w2(32'h39d46a7f),
	.w3(32'hba556ece),
	.w4(32'h3a0fd273),
	.w5(32'h3a29bdda),
	.w6(32'h39c61c85),
	.w7(32'h3a15c1e8),
	.w8(32'h39a40b60),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a558a35),
	.w1(32'h39df4643),
	.w2(32'hba0dace8),
	.w3(32'h3a05249f),
	.w4(32'hb8e84bde),
	.w5(32'hba21c910),
	.w6(32'hb8033aeb),
	.w7(32'hb9e65312),
	.w8(32'hba49872a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e0201),
	.w1(32'h388b5992),
	.w2(32'hb9a8181a),
	.w3(32'hba6b3ca2),
	.w4(32'h3896c799),
	.w5(32'hb9a2b912),
	.w6(32'hbaa3b63b),
	.w7(32'hbaa89941),
	.w8(32'hbaba8c48),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13cb20),
	.w1(32'hb9ad794d),
	.w2(32'hba646a47),
	.w3(32'h3a1d2eac),
	.w4(32'h39ff5a19),
	.w5(32'hb9364ab3),
	.w6(32'h3a1bb1ad),
	.w7(32'h3ab2ffae),
	.w8(32'h38d3070d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39358f60),
	.w1(32'h3a1b83a4),
	.w2(32'h3a920325),
	.w3(32'h39d4e081),
	.w4(32'h3a754e62),
	.w5(32'h3a7f1b05),
	.w6(32'h393f8b10),
	.w7(32'hb7a2d3bb),
	.w8(32'h38b97692),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a4031),
	.w1(32'h39a94449),
	.w2(32'h3827eea2),
	.w3(32'h3a874951),
	.w4(32'h39d14d33),
	.w5(32'h3980a90e),
	.w6(32'h38bed17d),
	.w7(32'hb99ffb17),
	.w8(32'hb8d458c9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964cfe2),
	.w1(32'hb93587ec),
	.w2(32'hb9bf85b8),
	.w3(32'h394427bb),
	.w4(32'hb8fd2ed8),
	.w5(32'hb91d87a2),
	.w6(32'hba093205),
	.w7(32'hba0be785),
	.w8(32'hb9deeb37),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b115e),
	.w1(32'hb9ac7276),
	.w2(32'hbab77c48),
	.w3(32'h39c39bbc),
	.w4(32'h3943a0aa),
	.w5(32'hbaa2280c),
	.w6(32'h3a36a63b),
	.w7(32'h3a18a6cf),
	.w8(32'hba7b3e8f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b05002),
	.w1(32'hba539906),
	.w2(32'hbb1dfa7b),
	.w3(32'hb9717a33),
	.w4(32'hba5f3802),
	.w5(32'hbb0f09c8),
	.w6(32'h3915a2c2),
	.w7(32'h383795be),
	.w8(32'hbac9bfe3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378dd637),
	.w1(32'hb8068f85),
	.w2(32'hb8ac08a7),
	.w3(32'hb7e210da),
	.w4(32'hb83e059a),
	.w5(32'hb8564c39),
	.w6(32'hb7eb0c0b),
	.w7(32'hb78768e1),
	.w8(32'hb86dfbdf),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b635e0),
	.w1(32'hb93789a1),
	.w2(32'hba0705f3),
	.w3(32'hb9c560f2),
	.w4(32'hb92fe2ad),
	.w5(32'hba0b121a),
	.w6(32'hb9ffed5b),
	.w7(32'hb92d55f8),
	.w8(32'hb9e66b20),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e4f92c),
	.w1(32'h38c6e7ed),
	.w2(32'hb9763c29),
	.w3(32'hb9d3c6ff),
	.w4(32'hb9056b7f),
	.w5(32'hb9b36b34),
	.w6(32'hba19f041),
	.w7(32'hb9a31938),
	.w8(32'hba1fb67e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4e305),
	.w1(32'hba08ad40),
	.w2(32'hba59946c),
	.w3(32'hb9897325),
	.w4(32'hb9743a6e),
	.w5(32'hba3bf75d),
	.w6(32'hb96f00fd),
	.w7(32'hb911a3b9),
	.w8(32'hba35b2a6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e06508),
	.w1(32'h381ef55d),
	.w2(32'hba88ce7a),
	.w3(32'h3a1d973f),
	.w4(32'h38e0e07c),
	.w5(32'hba05ffdc),
	.w6(32'h393f3a57),
	.w7(32'hba0f4fc8),
	.w8(32'hba61315b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fb743),
	.w1(32'hb9156dc3),
	.w2(32'hbb012cf6),
	.w3(32'hb9a39376),
	.w4(32'hba3d967c),
	.w5(32'hbb2269a1),
	.w6(32'hba035a3f),
	.w7(32'hba498f48),
	.w8(32'hbb211673),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0b633),
	.w1(32'h3831a2b8),
	.w2(32'hba215d45),
	.w3(32'h392dfbd8),
	.w4(32'h3931b319),
	.w5(32'hb9f82bb8),
	.w6(32'hb9c324dd),
	.w7(32'hb902eeaf),
	.w8(32'hba707d72),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24ab9e),
	.w1(32'h3923a4ba),
	.w2(32'hbab47dcd),
	.w3(32'h39324b8c),
	.w4(32'h3a4004ad),
	.w5(32'hb9814c5a),
	.w6(32'h38dc1560),
	.w7(32'h39ec2361),
	.w8(32'hba08bfcd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8106b1c),
	.w1(32'hb94428eb),
	.w2(32'hba935d21),
	.w3(32'hb8d43c53),
	.w4(32'h380c0391),
	.w5(32'hba88965f),
	.w6(32'hb9d9524e),
	.w7(32'hb8db923f),
	.w8(32'hba965cb1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f23bf),
	.w1(32'h3873dcb4),
	.w2(32'hb8d2ca94),
	.w3(32'hb99a27cd),
	.w4(32'h398622d4),
	.w5(32'h38839db9),
	.w6(32'hb9cb91ba),
	.w7(32'h395133f3),
	.w8(32'hb97dd72e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ebbd2),
	.w1(32'h3918f99e),
	.w2(32'hbab67715),
	.w3(32'h39f6eef3),
	.w4(32'hb7407757),
	.w5(32'hba927bc7),
	.w6(32'h3a00003d),
	.w7(32'h38b5f1ab),
	.w8(32'hba8268fe),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84551fd),
	.w1(32'h37ac614a),
	.w2(32'hb9caafa9),
	.w3(32'hb89bee31),
	.w4(32'h37f9cc5b),
	.w5(32'hb9d712a7),
	.w6(32'hb94d0932),
	.w7(32'hb8748a50),
	.w8(32'hb9fc9721),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0c145),
	.w1(32'h3a630836),
	.w2(32'hba59ba7e),
	.w3(32'h3a8addaa),
	.w4(32'h3a8403d8),
	.w5(32'hb961d757),
	.w6(32'hb8960890),
	.w7(32'hb9a82fd1),
	.w8(32'hbae64df0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398445bc),
	.w1(32'h3aa27220),
	.w2(32'h3a506781),
	.w3(32'h37731fe3),
	.w4(32'h3a89f5a8),
	.w5(32'h3a19b59c),
	.w6(32'hb944eb08),
	.w7(32'h3a2487e3),
	.w8(32'h38c1fe81),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb721ab82),
	.w1(32'hb7871e56),
	.w2(32'hb789d95f),
	.w3(32'h36c67af8),
	.w4(32'hb61ee964),
	.w5(32'hb78ade8a),
	.w6(32'h376a823e),
	.w7(32'h3714177c),
	.w8(32'h361498fc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ad4226),
	.w1(32'h35281aa7),
	.w2(32'h369c48b5),
	.w3(32'hb4c0eef4),
	.w4(32'h34dfad62),
	.w5(32'hb6b307c9),
	.w6(32'h3739c44e),
	.w7(32'h3739429a),
	.w8(32'h37177787),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ed95b),
	.w1(32'hb7ceb597),
	.w2(32'hb9b5e643),
	.w3(32'hb9c86244),
	.w4(32'h386f3863),
	.w5(32'hb8a63b32),
	.w6(32'hb9b443b6),
	.w7(32'hb7c2cb62),
	.w8(32'hb92a6abd),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c8d876),
	.w1(32'h3928edae),
	.w2(32'hba3978fd),
	.w3(32'h398f640e),
	.w4(32'h3a858097),
	.w5(32'hb7bdcbb7),
	.w6(32'hb9153aae),
	.w7(32'h3a38d57f),
	.w8(32'hb9a39636),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0f2ee),
	.w1(32'hb95eb451),
	.w2(32'hbab373c0),
	.w3(32'hbb121f79),
	.w4(32'hbace27bb),
	.w5(32'hbb04c6d4),
	.w6(32'hbb02d48a),
	.w7(32'hbaee714c),
	.w8(32'hbb1760eb),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369e0535),
	.w1(32'h36427a44),
	.w2(32'h36cab575),
	.w3(32'h364111ed),
	.w4(32'hb484dfe7),
	.w5(32'h3626813f),
	.w6(32'h3690e619),
	.w7(32'h35bfed16),
	.w8(32'h369fe260),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38596ec8),
	.w1(32'hb9e8e980),
	.w2(32'hbb0ff8eb),
	.w3(32'hb9904bd3),
	.w4(32'hb9dd3164),
	.w5(32'hbb02cde3),
	.w6(32'hba3f5bbb),
	.w7(32'hba201ed2),
	.w8(32'hbaff9bdf),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9036b11),
	.w1(32'hba336fc8),
	.w2(32'hbadee392),
	.w3(32'hba0ffc22),
	.w4(32'hba43b340),
	.w5(32'hbab259f4),
	.w6(32'hba391c95),
	.w7(32'hba47597c),
	.w8(32'hbaaf3d2d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b2274),
	.w1(32'hbaa5a387),
	.w2(32'hbb3f7fa3),
	.w3(32'hba34ee6e),
	.w4(32'hbaa08e5d),
	.w5(32'hbb10e267),
	.w6(32'hba25a8d5),
	.w7(32'hbaa64779),
	.w8(32'hbaeb18c1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65d8d5),
	.w1(32'h38dbeb7c),
	.w2(32'hbab16f6c),
	.w3(32'h3a1afc77),
	.w4(32'h3a2ac9ca),
	.w5(32'hba9f6c8d),
	.w6(32'hb90647fb),
	.w7(32'hb902b418),
	.w8(32'hba892057),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e1e0e),
	.w1(32'h3a94af71),
	.w2(32'h3a5531fe),
	.w3(32'hb8d6a978),
	.w4(32'h3a4f42b4),
	.w5(32'h3a21ccf4),
	.w6(32'hb9e3aa47),
	.w7(32'h39c85d8a),
	.w8(32'h388aa1d0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7faa206),
	.w1(32'h37ccefa0),
	.w2(32'hb898c9a3),
	.w3(32'hb80370ba),
	.w4(32'hb876ee8e),
	.w5(32'hb91608cb),
	.w6(32'hb7cdf7dd),
	.w7(32'hb8b3ba0a),
	.w8(32'hb8d02b94),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c56371),
	.w1(32'h3a384dda),
	.w2(32'hb94e7176),
	.w3(32'h3a81eb83),
	.w4(32'h3acad009),
	.w5(32'h39be2b19),
	.w6(32'h3a2c010e),
	.w7(32'h3ac16db9),
	.w8(32'h39bdb68c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a864b03),
	.w1(32'h3b169545),
	.w2(32'h3b097965),
	.w3(32'h3aa7f670),
	.w4(32'h3b3f17bc),
	.w5(32'h3b3269a7),
	.w6(32'h3a605ff2),
	.w7(32'h3af9b60a),
	.w8(32'h3ab1cf51),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96354cc),
	.w1(32'h3a038c85),
	.w2(32'h39ec3735),
	.w3(32'h389284a7),
	.w4(32'h3a41d540),
	.w5(32'h3a1e423e),
	.w6(32'hb932d177),
	.w7(32'h3a02aacb),
	.w8(32'h39cfe2bd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370ab391),
	.w1(32'hb7bf052e),
	.w2(32'hb8ee8a17),
	.w3(32'hb8f09c65),
	.w4(32'hb9095365),
	.w5(32'hb966a297),
	.w6(32'hb8dbb553),
	.w7(32'hb807d8c8),
	.w8(32'hb926360b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc82d2),
	.w1(32'hb80ac2d7),
	.w2(32'hb87bea4d),
	.w3(32'hb694a778),
	.w4(32'hb81d3826),
	.w5(32'hb884df96),
	.w6(32'hb89d3d57),
	.w7(32'hb8d226a7),
	.w8(32'hb8fc02a2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0853db),
	.w1(32'hb95d108d),
	.w2(32'hbac1b7f5),
	.w3(32'h394ce3fd),
	.w4(32'hb9960dc1),
	.w5(32'hbaad1506),
	.w6(32'hb8549753),
	.w7(32'hb93cd01b),
	.w8(32'hba91b051),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d503f),
	.w1(32'h392dfc09),
	.w2(32'hb743986a),
	.w3(32'h398a688e),
	.w4(32'h3933217e),
	.w5(32'h384a9653),
	.w6(32'h391a9912),
	.w7(32'h38f80f1b),
	.w8(32'hb77c89de),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c0a94),
	.w1(32'h3953f730),
	.w2(32'hb9be9c47),
	.w3(32'h3a01c259),
	.w4(32'h39ec26ad),
	.w5(32'hb97a3c40),
	.w6(32'h3985ed36),
	.w7(32'h3a3636b1),
	.w8(32'h388b5e44),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378e4858),
	.w1(32'h375e9bac),
	.w2(32'h35e016f3),
	.w3(32'h36a16457),
	.w4(32'h3898a494),
	.w5(32'h380a2cbe),
	.w6(32'hb50a12a8),
	.w7(32'h38b24b3b),
	.w8(32'h37d59449),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba730d59),
	.w1(32'hb8d365f0),
	.w2(32'hb9d4e6e5),
	.w3(32'hbad0523e),
	.w4(32'hba7cc44e),
	.w5(32'hbaa9b7fb),
	.w6(32'hba189459),
	.w7(32'hb8fab657),
	.w8(32'hbaa0591c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3845c3a6),
	.w1(32'h37095d27),
	.w2(32'h35b14206),
	.w3(32'h38463e8d),
	.w4(32'h36610816),
	.w5(32'hb7ffbe95),
	.w6(32'h38225744),
	.w7(32'hb72be218),
	.w8(32'hb79f37df),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79a1366),
	.w1(32'hb7006151),
	.w2(32'hb78dad7c),
	.w3(32'hb80f3dd1),
	.w4(32'hb81bce00),
	.w5(32'h37ac8f05),
	.w6(32'h37e0eb38),
	.w7(32'hb5332435),
	.w8(32'hb7f9e117),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a482d50),
	.w1(32'h3a0380ff),
	.w2(32'hb9861925),
	.w3(32'h3a416446),
	.w4(32'h3a79912d),
	.w5(32'h396b8643),
	.w6(32'h39d4a500),
	.w7(32'h3a0d8fd6),
	.w8(32'hb8e22c1e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fca272),
	.w1(32'h38452dd1),
	.w2(32'hbb1bb8f4),
	.w3(32'hb93c5847),
	.w4(32'hb9950497),
	.w5(32'hbb2bb2aa),
	.w6(32'hb934e8a5),
	.w7(32'h3a01a6b5),
	.w8(32'hbaf6ecfe),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8e3da),
	.w1(32'h39a7c201),
	.w2(32'h3816b525),
	.w3(32'hb9edb224),
	.w4(32'h38faeb27),
	.w5(32'hb979740c),
	.w6(32'hba3bbebe),
	.w7(32'hb7514576),
	.w8(32'hb9040d92),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba092d30),
	.w1(32'hb9fd685d),
	.w2(32'hbad36079),
	.w3(32'hba579191),
	.w4(32'hb9af5614),
	.w5(32'hbac43a26),
	.w6(32'hbaa2571b),
	.w7(32'hba70e9fb),
	.w8(32'hbb0093e4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d7a1c),
	.w1(32'hb8158629),
	.w2(32'hb96ac39e),
	.w3(32'hb7e1edf0),
	.w4(32'hb8da5fe4),
	.w5(32'hb94e8049),
	.w6(32'hb8a2482e),
	.w7(32'hb976f5f3),
	.w8(32'hb9b04508),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaded0f5),
	.w1(32'hbaa731b4),
	.w2(32'hbb2de382),
	.w3(32'hba5934d2),
	.w4(32'hb9adfa23),
	.w5(32'hbae2a01c),
	.w6(32'hbaa8912f),
	.w7(32'hb9e34fa6),
	.w8(32'hbabd7e56),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba147a66),
	.w1(32'hb91ac18f),
	.w2(32'hbaa26558),
	.w3(32'hb9b4d9b2),
	.w4(32'h38cf98db),
	.w5(32'hba7e9a7f),
	.w6(32'hb9cfdefb),
	.w7(32'h3891f6d0),
	.w8(32'hba6d9155),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99faaac),
	.w1(32'hba6f0e00),
	.w2(32'hbb2dadd3),
	.w3(32'hba03173a),
	.w4(32'hba7ec43c),
	.w5(32'hbb2bbf7d),
	.w6(32'hb9ba6a10),
	.w7(32'hb98ddc47),
	.w8(32'hbb08c57d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3875860b),
	.w1(32'h37c5e25d),
	.w2(32'h379ab15a),
	.w3(32'h3864f8de),
	.w4(32'h388c1c4b),
	.w5(32'h37b16669),
	.w6(32'h3817b4f0),
	.w7(32'h37c94bcc),
	.w8(32'hb64eaf89),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0edc73),
	.w1(32'hb71ada4d),
	.w2(32'hba803b6b),
	.w3(32'h39e10fd2),
	.w4(32'h39733eef),
	.w5(32'hb9e934d0),
	.w6(32'h39c4a28a),
	.w7(32'h394fd1b0),
	.w8(32'hb96edbdf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374cbe9a),
	.w1(32'hb6d49f60),
	.w2(32'h36ea5614),
	.w3(32'h362c8fc0),
	.w4(32'hb7567359),
	.w5(32'h36c92515),
	.w6(32'h3716770a),
	.w7(32'hb6c3ba49),
	.w8(32'h3792844c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937afb0),
	.w1(32'hb95271e6),
	.w2(32'hba1ac5b3),
	.w3(32'hb954c648),
	.w4(32'hb9ace130),
	.w5(32'hba1db2b2),
	.w6(32'hb9e27be8),
	.w7(32'hba1827cf),
	.w8(32'hba6738bf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831b8f1),
	.w1(32'h381c8a8b),
	.w2(32'hb9119cba),
	.w3(32'hb814526c),
	.w4(32'hb791111f),
	.w5(32'hb92584e4),
	.w6(32'h3616a09f),
	.w7(32'hb9008e33),
	.w8(32'hb9804bc6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec11d2),
	.w1(32'hba495d3e),
	.w2(32'hbaf2aa34),
	.w3(32'hba7a4a9c),
	.w4(32'hba8e267d),
	.w5(32'hbab93db6),
	.w6(32'hbad31ed9),
	.w7(32'hbad898ba),
	.w8(32'hbb06d7e9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a3f87d),
	.w1(32'hb6426558),
	.w2(32'h3573cfb7),
	.w3(32'h36085318),
	.w4(32'hb6adca77),
	.w5(32'hb5261c66),
	.w6(32'h3656a663),
	.w7(32'hb5be7c8f),
	.w8(32'h364b2856),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365f86e8),
	.w1(32'hb76e75c5),
	.w2(32'hb7a8c13d),
	.w3(32'h35c7a1e8),
	.w4(32'hb75eec6c),
	.w5(32'hb7bceae3),
	.w6(32'hb5c40c63),
	.w7(32'hb4ca14ac),
	.w8(32'hb70a8afb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9beb648),
	.w1(32'hb84ede7e),
	.w2(32'hb8ad761d),
	.w3(32'hb97d6945),
	.w4(32'h36d228d1),
	.w5(32'hb8d016b0),
	.w6(32'hb91561a5),
	.w7(32'hb777cfa8),
	.w8(32'hb911ab29),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397606ad),
	.w1(32'h3a0bc580),
	.w2(32'hba9398ff),
	.w3(32'h390a9f93),
	.w4(32'h3a0e8f41),
	.w5(32'hba2152f7),
	.w6(32'hb9de726e),
	.w7(32'h39192738),
	.w8(32'hba0a33d1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b119e9),
	.w1(32'h390e766d),
	.w2(32'hb99cde2c),
	.w3(32'hb9885df6),
	.w4(32'h389394c2),
	.w5(32'hb8e78e4d),
	.w6(32'hb97023c5),
	.w7(32'h39a92488),
	.w8(32'hb5848840),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ee9df),
	.w1(32'hb82d7387),
	.w2(32'hb92efafd),
	.w3(32'hb96c7526),
	.w4(32'hb902998b),
	.w5(32'hb932e4b5),
	.w6(32'hb8fe8fb0),
	.w7(32'hb8595a40),
	.w8(32'hb930ec7e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2289c4),
	.w1(32'hbac994f5),
	.w2(32'hbbb8e496),
	.w3(32'hb9af2f1c),
	.w4(32'hb947acd9),
	.w5(32'hbb681035),
	.w6(32'h3a515965),
	.w7(32'h3af7d0c2),
	.w8(32'hba8c54f0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a382e12),
	.w1(32'h3af26467),
	.w2(32'hb8919da0),
	.w3(32'h39fbdf24),
	.w4(32'h3b3ae40e),
	.w5(32'h3ac4d06c),
	.w6(32'h39d1bbee),
	.w7(32'h3af0de1f),
	.w8(32'h39f7448b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393117f8),
	.w1(32'h3878ffc5),
	.w2(32'hb913f521),
	.w3(32'h39520be2),
	.w4(32'hb7b8cb65),
	.w5(32'hb91758ca),
	.w6(32'h38f6d63a),
	.w7(32'hb8592a13),
	.w8(32'hb900aab5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb668596a),
	.w1(32'hb61ac4d8),
	.w2(32'h361d347e),
	.w3(32'hb7d1c41c),
	.w4(32'hb71c2e31),
	.w5(32'hb7018f7c),
	.w6(32'hb7b51bab),
	.w7(32'hb7c01d65),
	.w8(32'hb626025e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8096fa9),
	.w1(32'hb82a360a),
	.w2(32'hb7a72199),
	.w3(32'hb7a3b164),
	.w4(32'hb79a939b),
	.w5(32'hb6cdb17a),
	.w6(32'hb723af2d),
	.w7(32'h37d68956),
	.w8(32'h37e4ad3b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b0817a),
	.w1(32'h344ecffd),
	.w2(32'h37313bf2),
	.w3(32'h35f8ef47),
	.w4(32'hb69a3de3),
	.w5(32'h37226a01),
	.w6(32'h3693ab02),
	.w7(32'hb46a3420),
	.w8(32'h37727c3a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a701b3e),
	.w1(32'h39d29bf0),
	.w2(32'hb9e74fed),
	.w3(32'h39d64afe),
	.w4(32'h395aff09),
	.w5(32'hb992edce),
	.w6(32'h39871d9a),
	.w7(32'hb7600113),
	.w8(32'hb9ea894d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f2af4),
	.w1(32'h3a6ffc5d),
	.w2(32'hb9621252),
	.w3(32'hb9f99b7e),
	.w4(32'hb888b4d1),
	.w5(32'hb9c29d38),
	.w6(32'hb9833fae),
	.w7(32'hb996e4e1),
	.w8(32'hba5a3293),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c0fc6),
	.w1(32'hbabaaa29),
	.w2(32'hbb111e20),
	.w3(32'hbad05701),
	.w4(32'hbaaf9a72),
	.w5(32'hbb0b5b4f),
	.w6(32'hbb0d6118),
	.w7(32'hbac188ed),
	.w8(32'hbb08e777),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9025c39),
	.w1(32'hb844ae98),
	.w2(32'hb94d35d5),
	.w3(32'hba09c450),
	.w4(32'hb971530a),
	.w5(32'hb9ac656e),
	.w6(32'hb9430cf6),
	.w7(32'hb89d8fd5),
	.w8(32'hb98f13ab),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba021941),
	.w1(32'hbaa49ebe),
	.w2(32'hbb3a4287),
	.w3(32'hba22eb81),
	.w4(32'hba9ab77e),
	.w5(32'hbb1e0a55),
	.w6(32'hbaca50b0),
	.w7(32'hbabac845),
	.w8(32'hbb203133),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4041fb),
	.w1(32'hb9d9f092),
	.w2(32'hba024d10),
	.w3(32'hba0f8082),
	.w4(32'hb9d058e6),
	.w5(32'hba0d99c5),
	.w6(32'hba13b5de),
	.w7(32'hb9b04813),
	.w8(32'hb9c7147c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3759c8c8),
	.w1(32'h36ef07e3),
	.w2(32'h37ae41c5),
	.w3(32'h3732280f),
	.w4(32'h369e61a7),
	.w5(32'h3790dbee),
	.w6(32'h379bcfcf),
	.w7(32'h375fe745),
	.w8(32'h37d62526),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6c5c3),
	.w1(32'hb9e2fea2),
	.w2(32'hb9f58f96),
	.w3(32'hb9a591d3),
	.w4(32'hb99c8096),
	.w5(32'hb959c48e),
	.w6(32'hb8bf9b1f),
	.w7(32'hb9125a14),
	.w8(32'hb93160b8),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377cc8cf),
	.w1(32'h35c30b8e),
	.w2(32'h383c4219),
	.w3(32'h3765678e),
	.w4(32'h362f12af),
	.w5(32'h384f504f),
	.w6(32'h3814d37e),
	.w7(32'h37c4a9d6),
	.w8(32'h388ea40a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d1bea),
	.w1(32'h368d62ee),
	.w2(32'hba0bbac3),
	.w3(32'hba602176),
	.w4(32'hb95a9425),
	.w5(32'hba6400c0),
	.w6(32'hba73e194),
	.w7(32'hba1b6a3f),
	.w8(32'hbab8fe87),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba818647),
	.w1(32'h3ac39b29),
	.w2(32'h3ac4c029),
	.w3(32'hb9e90022),
	.w4(32'h3b1cb9b9),
	.w5(32'h3b1eeb6e),
	.w6(32'hb9de7fc0),
	.w7(32'h3aef0316),
	.w8(32'h3ae77267),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911f240),
	.w1(32'h3724a74a),
	.w2(32'hba8a122a),
	.w3(32'h38768f3b),
	.w4(32'h39a0e6c7),
	.w5(32'hba2ba5b4),
	.w6(32'hb9d86787),
	.w7(32'h38353766),
	.w8(32'hba7ea263),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8928551),
	.w1(32'h39a3c31e),
	.w2(32'h395d9d87),
	.w3(32'hb874a08b),
	.w4(32'h398e0312),
	.w5(32'h392cede3),
	.w6(32'hb8b6efd4),
	.w7(32'h3981127c),
	.w8(32'h38c3c8d0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39082cf9),
	.w1(32'hb9546e41),
	.w2(32'hbaa5a5d8),
	.w3(32'hb882a539),
	.w4(32'hb89f2ca9),
	.w5(32'hba82e709),
	.w6(32'hba477741),
	.w7(32'hba3ff602),
	.w8(32'hbae538dd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14ad7b),
	.w1(32'hba09188d),
	.w2(32'hbab48cb1),
	.w3(32'hba479f32),
	.w4(32'hba13ec7d),
	.w5(32'hbaa251f6),
	.w6(32'hba4b5761),
	.w7(32'hb9f9c427),
	.w8(32'hbaa13213),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ba721),
	.w1(32'hbab8893e),
	.w2(32'hbb3c4f9b),
	.w3(32'hbb2b6a26),
	.w4(32'hbaeba19b),
	.w5(32'hbb30f74c),
	.w6(32'hbb4cd5a9),
	.w7(32'hbaf53d75),
	.w8(32'hbb3c2b94),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35292459),
	.w1(32'h368b8925),
	.w2(32'h374f479a),
	.w3(32'h36a8b4fa),
	.w4(32'h36cf2a41),
	.w5(32'h3749405a),
	.w6(32'h37438a5b),
	.w7(32'h37770572),
	.w8(32'h37c3acbb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4bccf),
	.w1(32'h37a0153f),
	.w2(32'h378a7f75),
	.w3(32'h37cba4d5),
	.w4(32'h36c46e59),
	.w5(32'hb70972ad),
	.w6(32'hb5078c36),
	.w7(32'h3729e7bf),
	.w8(32'h35dda914),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3feac),
	.w1(32'h3a3173b6),
	.w2(32'hba1f52de),
	.w3(32'hb7e518ec),
	.w4(32'h3a544585),
	.w5(32'hba193565),
	.w6(32'hb9d926cf),
	.w7(32'h3a65b0c8),
	.w8(32'hba0ca8cb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bca4a3),
	.w1(32'hb8e27f3b),
	.w2(32'hbb035288),
	.w3(32'hb7601f7f),
	.w4(32'hb8db9e5d),
	.w5(32'hbb0c854d),
	.w6(32'hb90aa2ca),
	.w7(32'h3a4b0042),
	.w8(32'hba958ecc),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b805a4),
	.w1(32'hb9b6f9e3),
	.w2(32'hbaec5830),
	.w3(32'hb950aac1),
	.w4(32'h3906f9ca),
	.w5(32'hbab3c67b),
	.w6(32'hba0cb605),
	.w7(32'hb8677c7b),
	.w8(32'hbabea2cc),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a326737),
	.w1(32'h3937c69a),
	.w2(32'hb930d73c),
	.w3(32'h3924a945),
	.w4(32'hb974bdee),
	.w5(32'hb9d48b7e),
	.w6(32'h39b3f0a7),
	.w7(32'h37de2d1c),
	.w8(32'hb98b3eb1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3810aad0),
	.w1(32'hb74f1837),
	.w2(32'hb80bb47c),
	.w3(32'h36ed336c),
	.w4(32'hb85c2ece),
	.w5(32'hb7f25513),
	.w6(32'h37277050),
	.w7(32'hb8103fab),
	.w8(32'hb76b90b9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c96e0),
	.w1(32'hb9201bc4),
	.w2(32'hb94976d2),
	.w3(32'hb83597cb),
	.w4(32'hb8d8d546),
	.w5(32'hb921bba3),
	.w6(32'hb77f0bbc),
	.w7(32'hb8803910),
	.w8(32'hb89d1058),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e6034),
	.w1(32'h3a33d898),
	.w2(32'hba361057),
	.w3(32'hb9973839),
	.w4(32'hb95fe2b3),
	.w5(32'hba96828f),
	.w6(32'hba0cc752),
	.w7(32'h39b3c8b8),
	.w8(32'hba42cf85),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42a893),
	.w1(32'hbadda34d),
	.w2(32'hbb495c15),
	.w3(32'hbb2124b3),
	.w4(32'hbac683f5),
	.w5(32'hbb544aa7),
	.w6(32'hbb1a1a30),
	.w7(32'hba54fe7c),
	.w8(32'hbb099858),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6cb64),
	.w1(32'h3a32f30d),
	.w2(32'hbaca2ac6),
	.w3(32'h3999e65f),
	.w4(32'h386b5fde),
	.w5(32'hba8f4b2f),
	.w6(32'hb97dbe8f),
	.w7(32'hba7b1255),
	.w8(32'hbab4e4e1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe428d),
	.w1(32'h3aa05209),
	.w2(32'h3a45bcc2),
	.w3(32'hb9231e63),
	.w4(32'h3aa4898a),
	.w5(32'h3a2a49ff),
	.w6(32'hb9f17e45),
	.w7(32'h3a38046b),
	.w8(32'h3967b95f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade047a),
	.w1(32'hba95947c),
	.w2(32'hbaf68d6f),
	.w3(32'hba7d9b83),
	.w4(32'hb9018047),
	.w5(32'hba8a569c),
	.w6(32'hba7b1859),
	.w7(32'hb90afd0a),
	.w8(32'hba4ec469),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ebc826),
	.w1(32'h36922d23),
	.w2(32'h37145a83),
	.w3(32'h36dae25b),
	.w4(32'h366ae0cb),
	.w5(32'h36e15403),
	.w6(32'h37089099),
	.w7(32'h36ef89be),
	.w8(32'h373f260e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3688f88d),
	.w1(32'h35ab1a56),
	.w2(32'h36ea00be),
	.w3(32'h371d1eb5),
	.w4(32'h367c234b),
	.w5(32'h3707ca27),
	.w6(32'h37a41f78),
	.w7(32'h3763dd97),
	.w8(32'h379805f4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e84b8),
	.w1(32'h391dcd63),
	.w2(32'hb7ce582e),
	.w3(32'h39190105),
	.w4(32'hb76acbbf),
	.w5(32'hb90db9e8),
	.w6(32'h39209cb3),
	.w7(32'h389088ca),
	.w8(32'hb6098a6b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3769890f),
	.w1(32'hb672cf31),
	.w2(32'hb4c96cb6),
	.w3(32'h37463730),
	.w4(32'hb6aa8ea8),
	.w5(32'h3584845a),
	.w6(32'h3761459c),
	.w7(32'h36ebcf60),
	.w8(32'h370567a6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39091d93),
	.w1(32'h38d65bca),
	.w2(32'hb9a96981),
	.w3(32'h3790a4e1),
	.w4(32'hb767f2dd),
	.w5(32'hb9aadc29),
	.w6(32'h37b06178),
	.w7(32'h38909150),
	.w8(32'hb95df263),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980d2cf),
	.w1(32'hb92cbe1f),
	.w2(32'hbaf68cda),
	.w3(32'h3909feb4),
	.w4(32'hb7aab0da),
	.w5(32'hbad540fd),
	.w6(32'h39603056),
	.w7(32'h3a1865ff),
	.w8(32'hba92e2e2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a663e0),
	.w1(32'hb8fc8000),
	.w2(32'hba944d71),
	.w3(32'hb87e0ce1),
	.w4(32'hb71ac226),
	.w5(32'hba51e57a),
	.w6(32'hb9423263),
	.w7(32'hb94a6bb0),
	.w8(32'hba9225c7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a91c1f),
	.w1(32'h3790741c),
	.w2(32'h379162ad),
	.w3(32'h3790e96e),
	.w4(32'h378b40af),
	.w5(32'h376891b9),
	.w6(32'h37b0bf3a),
	.w7(32'h37a2074f),
	.w8(32'h37bc1382),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380daa80),
	.w1(32'hb9136876),
	.w2(32'hbb152b42),
	.w3(32'hba1c86ee),
	.w4(32'hba12e959),
	.w5(32'hbb19aa7e),
	.w6(32'hba8d9ddb),
	.w7(32'hba0c7ebe),
	.w8(32'hbb088985),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849909f),
	.w1(32'hb9857724),
	.w2(32'hba539de8),
	.w3(32'hb8c79b30),
	.w4(32'hb9dc661c),
	.w5(32'hba60cde2),
	.w6(32'hb7cef2fa),
	.w7(32'hb988ffb0),
	.w8(32'hba35ff9f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9400ecf),
	.w1(32'hb8d0ab49),
	.w2(32'hb9273ea9),
	.w3(32'hb9387546),
	.w4(32'hb94040ee),
	.w5(32'hb9574e55),
	.w6(32'hb96d4c06),
	.w7(32'hb927e7a5),
	.w8(32'hb9674f7a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab6a5d),
	.w1(32'h3884d34c),
	.w2(32'hba16ffcf),
	.w3(32'hb787d118),
	.w4(32'hb8b31c31),
	.w5(32'hba210d4e),
	.w6(32'hb9b766ca),
	.w7(32'hb99522b6),
	.w8(32'hba365b3d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372d998f),
	.w1(32'h36f53b3a),
	.w2(32'h3736f3ad),
	.w3(32'h3713c61f),
	.w4(32'h3633e9ac),
	.w5(32'h3703398b),
	.w6(32'h37811858),
	.w7(32'h37312564),
	.w8(32'h3769b0db),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38679f4c),
	.w1(32'h38142b38),
	.w2(32'h37ef9f5e),
	.w3(32'h38114042),
	.w4(32'h38a5c128),
	.w5(32'h37866c86),
	.w6(32'h3874d5b6),
	.w7(32'h389c29ce),
	.w8(32'h38c50c22),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a7fd98),
	.w1(32'h37a0a468),
	.w2(32'hb74acfac),
	.w3(32'h37a56312),
	.w4(32'h3776b3f0),
	.w5(32'hb5dab3c6),
	.w6(32'h3800a758),
	.w7(32'h3792fe80),
	.w8(32'h37a35ae7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3624457a),
	.w1(32'hb408808e),
	.w2(32'h372cab78),
	.w3(32'h35d152bc),
	.w4(32'hb3fcf2af),
	.w5(32'h3752367e),
	.w6(32'h369a0202),
	.w7(32'h36959cff),
	.w8(32'h3774e867),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371c3c04),
	.w1(32'h3994970d),
	.w2(32'h39a535cb),
	.w3(32'h38e45878),
	.w4(32'h39262d98),
	.w5(32'h390df745),
	.w6(32'hb95003a4),
	.w7(32'h38f81fd9),
	.w8(32'h395a50af),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e249f),
	.w1(32'hba6864ae),
	.w2(32'hbb388b62),
	.w3(32'hb9261149),
	.w4(32'hba3c832f),
	.w5(32'hbb1ba71a),
	.w6(32'hb9ef8b3f),
	.w7(32'hba0d7364),
	.w8(32'hbb07f0db),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f3fdb2),
	.w1(32'hb98fe66b),
	.w2(32'hbad45d7a),
	.w3(32'h39db6820),
	.w4(32'h38e22ac6),
	.w5(32'hbaaeef9e),
	.w6(32'h3a0247bc),
	.w7(32'h39dd0dcf),
	.w8(32'hba8bc920),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa290f),
	.w1(32'hba8d28c6),
	.w2(32'hbb1d26c7),
	.w3(32'hb9a47cb0),
	.w4(32'hba510ec9),
	.w5(32'hbb008751),
	.w6(32'hba416d98),
	.w7(32'hba80ee93),
	.w8(32'hbaee9956),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dc43f5),
	.w1(32'hb4fcc4b3),
	.w2(32'hb5ce7086),
	.w3(32'hb80a39f0),
	.w4(32'hb7281193),
	.w5(32'hb7252df6),
	.w6(32'hb820a423),
	.w7(32'hb7a6b6cc),
	.w8(32'hb73079b1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb853cf35),
	.w1(32'hb8bf8198),
	.w2(32'hb8c4821b),
	.w3(32'hb85f536c),
	.w4(32'hb8903aa5),
	.w5(32'hb890c6fc),
	.w6(32'hb65b79bc),
	.w7(32'hb84e3991),
	.w8(32'hb8731c6b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6161772),
	.w1(32'hb65441cf),
	.w2(32'hb58f5963),
	.w3(32'hb69bd052),
	.w4(32'hb784704d),
	.w5(32'hb73c1bcd),
	.w6(32'hb74cfe3e),
	.w7(32'hb79fe3b0),
	.w8(32'hb6453af5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f0aee),
	.w1(32'h37e0c1cf),
	.w2(32'h37b6d1dc),
	.w3(32'h376f556f),
	.w4(32'h378c9029),
	.w5(32'h38022a79),
	.w6(32'h36fd3f32),
	.w7(32'h37a18f80),
	.w8(32'h37a909da),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9304758),
	.w1(32'hba5e8193),
	.w2(32'hbae14fd1),
	.w3(32'h38a84c35),
	.w4(32'hb911624b),
	.w5(32'hba792ccc),
	.w6(32'h38d8b2fb),
	.w7(32'h3837d147),
	.w8(32'hba3d74ec),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb745c2f6),
	.w1(32'hb8021097),
	.w2(32'hb7d2a2ee),
	.w3(32'hb72ae428),
	.w4(32'hb818dfc1),
	.w5(32'hb83c8847),
	.w6(32'hb64c65a3),
	.w7(32'hb7888479),
	.w8(32'hb79a90d4),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963300f),
	.w1(32'h39a03c04),
	.w2(32'h398e22b0),
	.w3(32'hb96d1363),
	.w4(32'h39712e7e),
	.w5(32'h391be701),
	.w6(32'hb954e1d7),
	.w7(32'h38d86016),
	.w8(32'hb72f4656),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06a0e3),
	.w1(32'hb98555e8),
	.w2(32'hb96df1da),
	.w3(32'hb9d17ea6),
	.w4(32'hb91c4032),
	.w5(32'hb8abc08e),
	.w6(32'hb98d8fff),
	.w7(32'h3662bdbb),
	.w8(32'hb83c5788),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370d2623),
	.w1(32'hb6e89735),
	.w2(32'hb7336fd5),
	.w3(32'hb67efea1),
	.w4(32'hb76c28d0),
	.w5(32'hb7459132),
	.w6(32'hb751ffa9),
	.w7(32'hb781538c),
	.w8(32'h35128660),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8430a35),
	.w1(32'hb94260bb),
	.w2(32'hb9dd4cee),
	.w3(32'hb98463f3),
	.w4(32'hb9a69b9b),
	.w5(32'hb9e66b3f),
	.w6(32'hba059294),
	.w7(32'hb9874db3),
	.w8(32'hba095405),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7edb203),
	.w1(32'hb82e42bd),
	.w2(32'hb81d1bd5),
	.w3(32'hb7bec692),
	.w4(32'hb7dceacf),
	.w5(32'hb7fde6d6),
	.w6(32'hb7b3041a),
	.w7(32'hb7e00d0f),
	.w8(32'hb805e710),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398805d6),
	.w1(32'hba853710),
	.w2(32'hbb298078),
	.w3(32'hb98d0209),
	.w4(32'hba3ead9a),
	.w5(32'hba9f3e2e),
	.w6(32'hba38213a),
	.w7(32'hba82a6da),
	.w8(32'hbac8c981),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377a1030),
	.w1(32'hb7acda6c),
	.w2(32'hb7db26cf),
	.w3(32'hb6270ccf),
	.w4(32'hb7ca9732),
	.w5(32'hb7d4da3f),
	.w6(32'h375f8674),
	.w7(32'hb712e7b5),
	.w8(32'hb581afd9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7e429),
	.w1(32'h3ae645fc),
	.w2(32'h3a9a7f8b),
	.w3(32'h3a2378d6),
	.w4(32'h3ac03cf3),
	.w5(32'h3a44a214),
	.w6(32'hba72adee),
	.w7(32'h3ad051ad),
	.w8(32'h3a9ef697),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule