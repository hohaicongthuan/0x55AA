module layer_10_featuremap_359(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a85b0),
	.w1(32'hba678448),
	.w2(32'hbc2fb4fa),
	.w3(32'hbbf30af6),
	.w4(32'hbc1bb154),
	.w5(32'h3b413346),
	.w6(32'h3a4ae266),
	.w7(32'hbc4ad2c4),
	.w8(32'h3c1600fe),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbfe3d),
	.w1(32'h3b42144f),
	.w2(32'h3b44e0a9),
	.w3(32'hbb85a8c4),
	.w4(32'hbb87bb1c),
	.w5(32'hbb9088ee),
	.w6(32'hbbc65191),
	.w7(32'hbbc9c2b0),
	.w8(32'hbc255380),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb73a2),
	.w1(32'hba84eca3),
	.w2(32'h3b0b489e),
	.w3(32'h3c050d34),
	.w4(32'h3c26b215),
	.w5(32'h3ab7c89b),
	.w6(32'h3b3dc93c),
	.w7(32'h3b4262bb),
	.w8(32'hbae56f52),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bc16a),
	.w1(32'hbb1ad9b0),
	.w2(32'h3b413ae3),
	.w3(32'h3b8d6745),
	.w4(32'h3c4eebad),
	.w5(32'h3bde4af6),
	.w6(32'hbb8ff1ee),
	.w7(32'h3c5e24af),
	.w8(32'h3c93c378),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b4577),
	.w1(32'hbc5cd3fd),
	.w2(32'hbb73afe1),
	.w3(32'hbca97154),
	.w4(32'h3c6f38da),
	.w5(32'hbbcefe12),
	.w6(32'hbcfc7fa1),
	.w7(32'h3966a4c2),
	.w8(32'hba2c0e53),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfb9b4),
	.w1(32'hb98a09a8),
	.w2(32'hbc252b94),
	.w3(32'hbbe12909),
	.w4(32'hbc194a77),
	.w5(32'hbb0a50dc),
	.w6(32'hbb5592ac),
	.w7(32'hbc3106f4),
	.w8(32'h3bb1b99c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba568c1),
	.w1(32'h3b3aef64),
	.w2(32'hbc052e48),
	.w3(32'hbbaa62fa),
	.w4(32'hbc4596f8),
	.w5(32'hbaa4224f),
	.w6(32'hbaac8c8e),
	.w7(32'hbc11d06f),
	.w8(32'h3b6574bd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4774d),
	.w1(32'h3b8e5a57),
	.w2(32'hbc0fb126),
	.w3(32'hbc13a76f),
	.w4(32'hbc9ba322),
	.w5(32'h3bda044e),
	.w6(32'hbb1c3ff8),
	.w7(32'hbbd44ca6),
	.w8(32'h3cdc5953),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca25b0d),
	.w1(32'h3c7e5bfa),
	.w2(32'hbc2c53f1),
	.w3(32'hbc591917),
	.w4(32'hbd0aebe2),
	.w5(32'hbb9540a3),
	.w6(32'h3bb8f43e),
	.w7(32'hbce6d33c),
	.w8(32'h3b00e91a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1536d9),
	.w1(32'hb81afa3b),
	.w2(32'hbbb77f66),
	.w3(32'hbbcaeb57),
	.w4(32'hba650ae0),
	.w5(32'h3a9b2f99),
	.w6(32'hbbab5eba),
	.w7(32'hbb9c561d),
	.w8(32'h3bf0f3d4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c8cbf),
	.w1(32'h3b67f7ff),
	.w2(32'hbbb5955a),
	.w3(32'h3a7cb428),
	.w4(32'hb9418968),
	.w5(32'h3be9f560),
	.w6(32'h3bbb8db1),
	.w7(32'h3a50eb0a),
	.w8(32'hbc5deb44),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92fe82),
	.w1(32'h3bc35fde),
	.w2(32'h3bd4002c),
	.w3(32'h3c5cfbe6),
	.w4(32'h3a3267de),
	.w5(32'h3bdb3712),
	.w6(32'hbb6caf56),
	.w7(32'h3c4d57f2),
	.w8(32'h3cdb5d86),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cce8ec9),
	.w1(32'h3c6301dc),
	.w2(32'hbbfe515d),
	.w3(32'hbcd3178e),
	.w4(32'hbcce19ae),
	.w5(32'h3ad27602),
	.w6(32'h3bbdd4fb),
	.w7(32'hbc9257b0),
	.w8(32'h3c0857da),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836803),
	.w1(32'hbb56e77c),
	.w2(32'hbb6594cd),
	.w3(32'hbb94cbd6),
	.w4(32'h3a6e3128),
	.w5(32'hbb800015),
	.w6(32'h3b98b36e),
	.w7(32'hba020f14),
	.w8(32'h3b62149d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58b1de),
	.w1(32'h3c583f25),
	.w2(32'hbb734e25),
	.w3(32'hbc028b10),
	.w4(32'hbc1e372a),
	.w5(32'h3bb7096a),
	.w6(32'h3b6f2592),
	.w7(32'hbc385796),
	.w8(32'h3cad496d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5019ae),
	.w1(32'h3bf207aa),
	.w2(32'hb7c96681),
	.w3(32'hbc9c8daf),
	.w4(32'hbb9b2550),
	.w5(32'h3c0e676e),
	.w6(32'hb828c2d3),
	.w7(32'hbc3513b4),
	.w8(32'h3c1ea6bc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7938a8),
	.w1(32'h3c21f433),
	.w2(32'h3a36685c),
	.w3(32'h395d6e74),
	.w4(32'hbc1a5b9d),
	.w5(32'hba853140),
	.w6(32'h3c86d1fd),
	.w7(32'hbb522104),
	.w8(32'hbb9c5945),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c0859),
	.w1(32'h3a2da977),
	.w2(32'h3b7855cd),
	.w3(32'h3c300e86),
	.w4(32'h3b20ddba),
	.w5(32'hbba1f0b3),
	.w6(32'h3c0470a4),
	.w7(32'h3c3d4a94),
	.w8(32'hbcad67ba),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9202e3),
	.w1(32'hbc719d95),
	.w2(32'h3bf674f5),
	.w3(32'h3c4714a1),
	.w4(32'h3c5bebb3),
	.w5(32'hbc210e30),
	.w6(32'hbc01bf0d),
	.w7(32'h3c74e4e3),
	.w8(32'h399d0039),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ecedd),
	.w1(32'h3b07775a),
	.w2(32'hbb652213),
	.w3(32'hbbcbae04),
	.w4(32'hbb81a69a),
	.w5(32'h3b5d119e),
	.w6(32'h3bec83a1),
	.w7(32'hbb76c1b9),
	.w8(32'h3bcb085e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e480c),
	.w1(32'h3c29b50b),
	.w2(32'hbb7f157e),
	.w3(32'hbc74f3de),
	.w4(32'hbbf0f70a),
	.w5(32'h3a714e82),
	.w6(32'hbad3db43),
	.w7(32'hbc89dc41),
	.w8(32'hbbefe3ff),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc538ef1),
	.w1(32'hbb571a3f),
	.w2(32'h3b67a685),
	.w3(32'h3b51e04c),
	.w4(32'h3b0374a1),
	.w5(32'h3809752e),
	.w6(32'hb9e9edf7),
	.w7(32'h3bb87e2f),
	.w8(32'hbbd2e0a6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89160),
	.w1(32'hbb863704),
	.w2(32'hbb1a61e0),
	.w3(32'hba9677f7),
	.w4(32'h3a6a97af),
	.w5(32'h39833009),
	.w6(32'hbae22dfa),
	.w7(32'hba2e5391),
	.w8(32'h3cd7e71b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe7c29),
	.w1(32'h3c545284),
	.w2(32'hbbd05771),
	.w3(32'hbc754e27),
	.w4(32'hbc074f9a),
	.w5(32'hba0cbe5d),
	.w6(32'hbb5cc2af),
	.w7(32'hbc27baa1),
	.w8(32'hbbc63eee),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4a328),
	.w1(32'hbbcd93e1),
	.w2(32'hbaad4945),
	.w3(32'hbbe6c39a),
	.w4(32'h3b903385),
	.w5(32'h3b1cc946),
	.w6(32'h3aa76855),
	.w7(32'h3a982e48),
	.w8(32'hb9a749d3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3e59e),
	.w1(32'h3b0f0de4),
	.w2(32'hbb002057),
	.w3(32'h3b4b3da0),
	.w4(32'hbb2a558b),
	.w5(32'hb9a26672),
	.w6(32'h3b9e78fb),
	.w7(32'hbb4217f5),
	.w8(32'hbbe4d582),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d25e2),
	.w1(32'hbc0a1b05),
	.w2(32'h3b872fbb),
	.w3(32'h3b17d963),
	.w4(32'h3c8294ec),
	.w5(32'hbb0977f2),
	.w6(32'hba98c014),
	.w7(32'h3c0a32a4),
	.w8(32'h3c2d8ee5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e371b),
	.w1(32'h3b03866f),
	.w2(32'hbc1af10c),
	.w3(32'hbc65c08f),
	.w4(32'hbc9ca660),
	.w5(32'hbc044b51),
	.w6(32'hbc18ca56),
	.w7(32'hbc932c7c),
	.w8(32'hbb63f5b4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8b8de),
	.w1(32'hbb0096b8),
	.w2(32'hbb35b2c7),
	.w3(32'h3813744a),
	.w4(32'h38d6588b),
	.w5(32'h3aa1880e),
	.w6(32'h3b9f39a7),
	.w7(32'h3b9594e5),
	.w8(32'h3c184e38),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16c9c7),
	.w1(32'h3b8c6f05),
	.w2(32'hbb8d505f),
	.w3(32'hbc748e70),
	.w4(32'hbbdeef67),
	.w5(32'hbb3e8bf9),
	.w6(32'h3a58f0f9),
	.w7(32'hbc0adbee),
	.w8(32'h3ba8fd94),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111b31),
	.w1(32'h3c7e5fc4),
	.w2(32'hbc133742),
	.w3(32'hbc0f2157),
	.w4(32'hbb857025),
	.w5(32'hbbc0dea4),
	.w6(32'hbb868244),
	.w7(32'hbb889521),
	.w8(32'hbc4602e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf02287),
	.w1(32'h3b1e8483),
	.w2(32'hbc1ae179),
	.w3(32'hbb120fb2),
	.w4(32'hba723503),
	.w5(32'h3c02b58f),
	.w6(32'hbc0fca51),
	.w7(32'h3aba4cf1),
	.w8(32'hbbe8f5e3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4deb7b),
	.w1(32'hbcbb40f6),
	.w2(32'h3c2735ed),
	.w3(32'h3c6fa004),
	.w4(32'h3c7939a8),
	.w5(32'hbbe74092),
	.w6(32'hbc48c670),
	.w7(32'h3c892aca),
	.w8(32'hbc249a19),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf8de8),
	.w1(32'hbc182030),
	.w2(32'h3bf4754b),
	.w3(32'h3bab10c0),
	.w4(32'h3c4a09ac),
	.w5(32'hbb9dbc42),
	.w6(32'hba785218),
	.w7(32'h3c7289f0),
	.w8(32'hbc6502a6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbada5fa),
	.w1(32'hbbeadf0c),
	.w2(32'hbb9bacc0),
	.w3(32'hbae2b4de),
	.w4(32'hbb3e22c9),
	.w5(32'hbbe76e52),
	.w6(32'h3c8a0867),
	.w7(32'hbb94c25e),
	.w8(32'hbc55515c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37c91),
	.w1(32'hbb8af7b6),
	.w2(32'h3bb5dfee),
	.w3(32'h3bafc7a8),
	.w4(32'h3befb94f),
	.w5(32'h3c42ad0b),
	.w6(32'h3b7bdb5e),
	.w7(32'h3a434423),
	.w8(32'hbc13d5b8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad818e5),
	.w1(32'hbbb989b5),
	.w2(32'h3be51c69),
	.w3(32'h3c02dee3),
	.w4(32'h3beb502c),
	.w5(32'h3c019313),
	.w6(32'hbacf7a99),
	.w7(32'h3be3d01a),
	.w8(32'h3b877a07),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41eb6b),
	.w1(32'hbb8e8bc6),
	.w2(32'hbb55071d),
	.w3(32'h3c4bc0e4),
	.w4(32'h3c3ca841),
	.w5(32'h3b078e0f),
	.w6(32'h3b79297c),
	.w7(32'h3b54f391),
	.w8(32'h3cc8be3e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2027d6),
	.w1(32'h3c65f6a3),
	.w2(32'hbbee90ba),
	.w3(32'hbc7eeea9),
	.w4(32'hbc32117c),
	.w5(32'h3bb8188f),
	.w6(32'h3c1f8c19),
	.w7(32'hbcc52a51),
	.w8(32'hbd120c31),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b9315),
	.w1(32'hbc881510),
	.w2(32'h3c5af8c5),
	.w3(32'h3cecb9a3),
	.w4(32'h3c9c5016),
	.w5(32'h3b431da0),
	.w6(32'hb9fe19e8),
	.w7(32'h3cf600c0),
	.w8(32'hbb839c99),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3ce9a),
	.w1(32'h3a52422c),
	.w2(32'hbad5b369),
	.w3(32'hba763c08),
	.w4(32'hbbcbb11c),
	.w5(32'h3c010d17),
	.w6(32'h3b563e57),
	.w7(32'h3b6ecdcb),
	.w8(32'hbbb065a7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24b125),
	.w1(32'h3af692e3),
	.w2(32'h3bec5b6e),
	.w3(32'h3c5a5e7e),
	.w4(32'h3c63364c),
	.w5(32'hbb903171),
	.w6(32'h3b97eaa3),
	.w7(32'h3c3231ba),
	.w8(32'hbc46f28b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb5d5d),
	.w1(32'hbba6f0fb),
	.w2(32'h3c364ba6),
	.w3(32'h3bc00dec),
	.w4(32'h3b7167cb),
	.w5(32'h3b86a36b),
	.w6(32'h3a80affc),
	.w7(32'h3c09692e),
	.w8(32'h3b9145cc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a252e3d),
	.w1(32'h3c004a99),
	.w2(32'h3befc231),
	.w3(32'hbbd3de96),
	.w4(32'hbc6b54fe),
	.w5(32'hbc642263),
	.w6(32'h3c61ba99),
	.w7(32'h3bc52063),
	.w8(32'hbd4b50ab),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2d44a0),
	.w1(32'hbd226a3a),
	.w2(32'h3bac2be0),
	.w3(32'h3c837616),
	.w4(32'h3cc3b7e4),
	.w5(32'hb8342bc0),
	.w6(32'hbcf28cbb),
	.w7(32'h3d00bfb2),
	.w8(32'hbc0bd40e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b5924),
	.w1(32'hbb81e41d),
	.w2(32'h3be8b0fa),
	.w3(32'hbb1b438e),
	.w4(32'h3b95a956),
	.w5(32'hbb7699e9),
	.w6(32'hbc0b21e4),
	.w7(32'h3b82634f),
	.w8(32'hbd0077d4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb56a1),
	.w1(32'hbc8fec09),
	.w2(32'h3c1b797d),
	.w3(32'h3c8fd84a),
	.w4(32'h3c9ead29),
	.w5(32'h3c445740),
	.w6(32'hbc7cd3f3),
	.w7(32'h3c90e6d6),
	.w8(32'h3d1d70cd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdaa234),
	.w1(32'h3c920735),
	.w2(32'hbc71d42a),
	.w3(32'hbcaf0ae1),
	.w4(32'hbcf65752),
	.w5(32'h3ada607c),
	.w6(32'h3bf14a33),
	.w7(32'hbd08102a),
	.w8(32'h3cd53572),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb48ec4),
	.w1(32'h3c8c4bd3),
	.w2(32'hbc555276),
	.w3(32'hbc51f8f5),
	.w4(32'hbc88c829),
	.w5(32'h3ba0a7a7),
	.w6(32'h3bba501c),
	.w7(32'hbc832bd4),
	.w8(32'h3a2a8846),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe025d5),
	.w1(32'hbadf5e82),
	.w2(32'h3bc160ac),
	.w3(32'h3aaeba32),
	.w4(32'h3b81670c),
	.w5(32'h3a7890cb),
	.w6(32'hb90a0046),
	.w7(32'h3b9b4e2e),
	.w8(32'h39931616),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba337057),
	.w1(32'hbc8a2301),
	.w2(32'hbbcd409c),
	.w3(32'h3b14376c),
	.w4(32'h3c28c40b),
	.w5(32'hba303d3e),
	.w6(32'hbc867a0a),
	.w7(32'h3c383754),
	.w8(32'hbc884ec4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf49a62),
	.w1(32'hbc5bf310),
	.w2(32'h3c2af134),
	.w3(32'h3befe6fd),
	.w4(32'h3b425ff7),
	.w5(32'h3b872220),
	.w6(32'hbbd77bdf),
	.w7(32'h3c85b797),
	.w8(32'hbba0a4c7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25a1f9),
	.w1(32'h3b89a6d5),
	.w2(32'h3a5c5044),
	.w3(32'hbb71319a),
	.w4(32'h3a41c888),
	.w5(32'h3b84915a),
	.w6(32'h3ae01ea8),
	.w7(32'h3be49026),
	.w8(32'h3b015966),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b351533),
	.w1(32'hbb0c19e0),
	.w2(32'h388bf4df),
	.w3(32'hbc0e10b1),
	.w4(32'hbb0d96d3),
	.w5(32'hbbffdd88),
	.w6(32'hbb38d814),
	.w7(32'h3a178359),
	.w8(32'hbb06f48e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea729),
	.w1(32'h3b303176),
	.w2(32'h3b8feb60),
	.w3(32'h3c421014),
	.w4(32'h3c1472af),
	.w5(32'h3b6b989d),
	.w6(32'h3b606914),
	.w7(32'h3c13552e),
	.w8(32'h3b9ee580),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d9a6f6),
	.w1(32'hbbbbda90),
	.w2(32'h395ffe8b),
	.w3(32'hbb2476aa),
	.w4(32'hba0b08ef),
	.w5(32'hbb6d3bb4),
	.w6(32'h3c323a50),
	.w7(32'h3c0ed064),
	.w8(32'h3b47c276),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04bbc6),
	.w1(32'hb9125a7d),
	.w2(32'hbae224fe),
	.w3(32'hbadb2291),
	.w4(32'hbbdc836c),
	.w5(32'hbb939ab7),
	.w6(32'h3be5ec4b),
	.w7(32'hbab441ac),
	.w8(32'hbac5113f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc4fd1),
	.w1(32'hbbacd85f),
	.w2(32'hbb3101c1),
	.w3(32'hbc009a59),
	.w4(32'hbb0e5f53),
	.w5(32'h3b886126),
	.w6(32'hbb31a656),
	.w7(32'hbabd23c5),
	.w8(32'h3bc4e6af),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ab284),
	.w1(32'h3ae81ad4),
	.w2(32'hba75edc4),
	.w3(32'h39547e12),
	.w4(32'hbb96f865),
	.w5(32'h3c6dee9f),
	.w6(32'h3afbf276),
	.w7(32'hbb71ed71),
	.w8(32'hb7242cda),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c330d),
	.w1(32'hbc23d7de),
	.w2(32'h3c561d60),
	.w3(32'h3c836465),
	.w4(32'h3c0dd961),
	.w5(32'hbb1946fe),
	.w6(32'hbba213a9),
	.w7(32'h3ca876a5),
	.w8(32'h3c88bfe6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3a3a6),
	.w1(32'h3c0c6e0a),
	.w2(32'hbc16b3fb),
	.w3(32'hbc5acc56),
	.w4(32'hbc219c60),
	.w5(32'hbaf230d4),
	.w6(32'h3b9fa6b5),
	.w7(32'hbc53090d),
	.w8(32'h3abfaee2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac14552),
	.w1(32'h3c1205f9),
	.w2(32'hbb927a7b),
	.w3(32'hbc109ea0),
	.w4(32'hbb95d668),
	.w5(32'h3a8dba8e),
	.w6(32'hbb3569c6),
	.w7(32'hbbf6b72e),
	.w8(32'h3a35bc18),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45fba9),
	.w1(32'hba00c532),
	.w2(32'h39a00e72),
	.w3(32'hbace39b5),
	.w4(32'hbb2ea38c),
	.w5(32'hba9814d7),
	.w6(32'h3c1ffc46),
	.w7(32'hbbd1d7d6),
	.w8(32'hbc036c7d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1dc08),
	.w1(32'hbc079921),
	.w2(32'h3b200959),
	.w3(32'h3aa25baa),
	.w4(32'hbaa74c9b),
	.w5(32'hbb90bae5),
	.w6(32'h3c4f11af),
	.w7(32'h3af7f49a),
	.w8(32'hbb3fd976),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ef650),
	.w1(32'hbc07ab97),
	.w2(32'hbb93dd00),
	.w3(32'hbada4935),
	.w4(32'h3a3c0462),
	.w5(32'hbb562961),
	.w6(32'h3bc8087a),
	.w7(32'h3aabf128),
	.w8(32'hbb880a89),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40d463),
	.w1(32'h3bf7af21),
	.w2(32'hba8f74c0),
	.w3(32'h3b9932fb),
	.w4(32'h3bb561fb),
	.w5(32'hbb5fd124),
	.w6(32'hbb8f6774),
	.w7(32'h3bf45121),
	.w8(32'h3bee8b0b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d46e0),
	.w1(32'h3c0e80b3),
	.w2(32'hbc6a7041),
	.w3(32'hbca789af),
	.w4(32'hbca1a957),
	.w5(32'hbaef37f9),
	.w6(32'h39833867),
	.w7(32'hbca92f65),
	.w8(32'h3ce28813),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47b6bd),
	.w1(32'h3ca50c0a),
	.w2(32'hbc4d4f8d),
	.w3(32'hbd005f8c),
	.w4(32'hbcfee97b),
	.w5(32'hbb84c12a),
	.w6(32'hbb36ef7e),
	.w7(32'hbd2aa436),
	.w8(32'h3b952f71),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91f18c),
	.w1(32'hbcc5b534),
	.w2(32'hbc37d636),
	.w3(32'hb953a740),
	.w4(32'h3bfe5b97),
	.w5(32'hbb744635),
	.w6(32'hbcb7940d),
	.w7(32'h3beac6d9),
	.w8(32'hbb9a3694),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac93f5c),
	.w1(32'hbad834b5),
	.w2(32'hb92a27cb),
	.w3(32'h3addb19b),
	.w4(32'h3aba3d90),
	.w5(32'h3bc281e6),
	.w6(32'h3babe554),
	.w7(32'h3c578ea4),
	.w8(32'hbc5878f2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc99b0b),
	.w1(32'hbb4b4a27),
	.w2(32'h3c3be9ee),
	.w3(32'h3c7485a1),
	.w4(32'h3c3bf993),
	.w5(32'h397d0663),
	.w6(32'h3b93d1e3),
	.w7(32'h3c84330d),
	.w8(32'h3c130571),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b002406),
	.w1(32'h3bea1eda),
	.w2(32'hbb287fd4),
	.w3(32'hbc1f5cfc),
	.w4(32'hbc7146d7),
	.w5(32'h3b05582c),
	.w6(32'h3b73b2c2),
	.w7(32'hbc6fd2e6),
	.w8(32'h3be0e92b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19a97e),
	.w1(32'h3c829ca7),
	.w2(32'hbbc0f00e),
	.w3(32'hbbde5e70),
	.w4(32'hbc012e78),
	.w5(32'h39bbf596),
	.w6(32'hbba5b25c),
	.w7(32'hbcb69988),
	.w8(32'hbb73b339),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf50ed),
	.w1(32'hbbede32e),
	.w2(32'h3ae82906),
	.w3(32'h3b184dfa),
	.w4(32'h3c20680b),
	.w5(32'h3920336d),
	.w6(32'hbbdb67a4),
	.w7(32'h3aae3254),
	.w8(32'h3c9bede3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f3e24),
	.w1(32'h3ac29b28),
	.w2(32'hbc231781),
	.w3(32'hbc89e343),
	.w4(32'hbc0b1f3f),
	.w5(32'hbb8ed5ad),
	.w6(32'h3b028772),
	.w7(32'hbc8195dd),
	.w8(32'h3b88a336),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbf53a),
	.w1(32'h3b25612c),
	.w2(32'hba44fb89),
	.w3(32'hbb7642cf),
	.w4(32'hbb840820),
	.w5(32'h3a8d61df),
	.w6(32'h39a25b78),
	.w7(32'h3a60bc66),
	.w8(32'hbb3e8d2f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4adbd),
	.w1(32'hbbb6cf0e),
	.w2(32'hbb8f5155),
	.w3(32'hbad67941),
	.w4(32'h3b67fc2d),
	.w5(32'hbc4e05ea),
	.w6(32'hbbf75c1e),
	.w7(32'h3b16e179),
	.w8(32'hbcdd4ea8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90d1e1),
	.w1(32'hbcb8e231),
	.w2(32'h3b84fdc9),
	.w3(32'h3bef04fc),
	.w4(32'h3c437c2f),
	.w5(32'h394bb42d),
	.w6(32'hbc9dcc85),
	.w7(32'h3c8b8591),
	.w8(32'hbbe81c3b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2c859),
	.w1(32'hbb9a36d8),
	.w2(32'hbb7eb7bd),
	.w3(32'h3c0670f8),
	.w4(32'h3b88482b),
	.w5(32'hbabd805b),
	.w6(32'hbbe3609e),
	.w7(32'h3c716c1b),
	.w8(32'h3ca4d4c2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c4430),
	.w1(32'h3ca34550),
	.w2(32'hbc27b5ab),
	.w3(32'hbc9d0d56),
	.w4(32'hbcde942d),
	.w5(32'h3ad1f328),
	.w6(32'h3a80cb88),
	.w7(32'hbce00afb),
	.w8(32'h3b9a3b38),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8157c8),
	.w1(32'h3c027a26),
	.w2(32'hbbfcf081),
	.w3(32'h3b9033c6),
	.w4(32'hbac7617f),
	.w5(32'h39057406),
	.w6(32'hbb765f02),
	.w7(32'h3a1da010),
	.w8(32'hbc133ae0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d74fe),
	.w1(32'hba69c0c6),
	.w2(32'hba4b1056),
	.w3(32'h3c144f17),
	.w4(32'h3bb8f9f0),
	.w5(32'h3b093c20),
	.w6(32'hb989e3d8),
	.w7(32'h3c0917e8),
	.w8(32'h3a16862b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acba20b),
	.w1(32'hbbc92dcc),
	.w2(32'h3ae7e57d),
	.w3(32'h3bb6701d),
	.w4(32'h3bbbc8d4),
	.w5(32'hbb69120a),
	.w6(32'hbb1f2f2e),
	.w7(32'h3a836b03),
	.w8(32'h3bd5286d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18dd79),
	.w1(32'h3bff7725),
	.w2(32'hbb917b3b),
	.w3(32'hbc837f7d),
	.w4(32'h3b9d6e64),
	.w5(32'hbb9ab070),
	.w6(32'hb999e204),
	.w7(32'hbbd465e3),
	.w8(32'hbc311c2d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac3b7a),
	.w1(32'hbbbddf5d),
	.w2(32'h39b36aa5),
	.w3(32'h3b4e36bb),
	.w4(32'h3a6cb0e3),
	.w5(32'hbb05e698),
	.w6(32'hbbc4288b),
	.w7(32'hbb735ec2),
	.w8(32'h3c31e777),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7ad53),
	.w1(32'h3c18304e),
	.w2(32'hbc384680),
	.w3(32'hba7d3954),
	.w4(32'h383b7e0c),
	.w5(32'h3bd764da),
	.w6(32'hb9e89ca6),
	.w7(32'hbbd945c2),
	.w8(32'hbb93a545),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd088cc),
	.w1(32'hba915c8a),
	.w2(32'h3bec34c0),
	.w3(32'h3b088ce3),
	.w4(32'h3bf2f86c),
	.w5(32'h3bb0d4a2),
	.w6(32'h3b84aff5),
	.w7(32'h3ba12979),
	.w8(32'h3bb34f75),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910410e),
	.w1(32'hba1c795a),
	.w2(32'hbb91aad1),
	.w3(32'h3aa0e945),
	.w4(32'h3b995e74),
	.w5(32'h3b1b4f17),
	.w6(32'h3c05559a),
	.w7(32'h3b60f060),
	.w8(32'h3c053578),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b810a66),
	.w1(32'h3c216cf6),
	.w2(32'hbb644254),
	.w3(32'hbb97cbd2),
	.w4(32'hbc47fb96),
	.w5(32'hbbbdecd4),
	.w6(32'h3bb617b2),
	.w7(32'hbc046754),
	.w8(32'h3c29486b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae3284),
	.w1(32'h3b3bb9b8),
	.w2(32'hbc10719a),
	.w3(32'hbbd929ba),
	.w4(32'hbae54349),
	.w5(32'h3a6124b1),
	.w6(32'hbb7d1e1a),
	.w7(32'hb9c7fd06),
	.w8(32'h3c54e1a3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c458582),
	.w1(32'h3c0f1bb3),
	.w2(32'hbb7a4131),
	.w3(32'hbbf838ff),
	.w4(32'hbbda872d),
	.w5(32'hbbace6a8),
	.w6(32'hbbcdb1bb),
	.w7(32'hbc05640e),
	.w8(32'hbbe6e4b3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc335e3f),
	.w1(32'hbbd86c77),
	.w2(32'hbb58c38b),
	.w3(32'h3b96b0f7),
	.w4(32'h3bb37dd0),
	.w5(32'h3b172634),
	.w6(32'hbbd18df8),
	.w7(32'h3bd5683d),
	.w8(32'h3b0053c2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11cee4),
	.w1(32'hbb8728e6),
	.w2(32'h3aa31afb),
	.w3(32'hbbd0c2bc),
	.w4(32'h3c48a66b),
	.w5(32'hbbc56cc7),
	.w6(32'h3b647298),
	.w7(32'h3b16af10),
	.w8(32'hbc49fbc5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b0040),
	.w1(32'hbc1ecb0a),
	.w2(32'hbc5f56f9),
	.w3(32'hbb647f1d),
	.w4(32'hbbeb81ae),
	.w5(32'h3ba9ecce),
	.w6(32'hbc3491ec),
	.w7(32'hbc899296),
	.w8(32'h3c02de3f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb320afa),
	.w1(32'h3b000f52),
	.w2(32'hba72e5f0),
	.w3(32'h3b641daa),
	.w4(32'h3bcdc759),
	.w5(32'hbbb76c51),
	.w6(32'h3bb381e0),
	.w7(32'h3b0ac4b8),
	.w8(32'hbc4367dd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f70c6),
	.w1(32'hbc28d3a9),
	.w2(32'hb9e0c857),
	.w3(32'h3b9e30a4),
	.w4(32'h3c687be1),
	.w5(32'hba050def),
	.w6(32'hbc40d247),
	.w7(32'h3bea87a5),
	.w8(32'hbc6798c2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c3b16),
	.w1(32'hbc9222ac),
	.w2(32'h3c2c8d72),
	.w3(32'h3c84dd58),
	.w4(32'h3cc77fbb),
	.w5(32'h39b5c53d),
	.w6(32'hbc9591d3),
	.w7(32'h3cf4599d),
	.w8(32'h393a5b2c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3a275),
	.w1(32'hbc902666),
	.w2(32'hb960f6d5),
	.w3(32'hbaf830ca),
	.w4(32'h3b801c06),
	.w5(32'hbbd21edc),
	.w6(32'hbc29477f),
	.w7(32'h3c07e884),
	.w8(32'hbbcb0adb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf802e9),
	.w1(32'hbbcbf635),
	.w2(32'hbbd36e7f),
	.w3(32'hbb801b58),
	.w4(32'hbb85cb59),
	.w5(32'h3c17fd8b),
	.w6(32'hb98b05d3),
	.w7(32'hbbf10558),
	.w8(32'h3c6c29bc),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1aff9e),
	.w1(32'hbac33f18),
	.w2(32'hbcbf1a74),
	.w3(32'hbb04b8b8),
	.w4(32'hbc25664b),
	.w5(32'h3bf48cae),
	.w6(32'hbba08c5f),
	.w7(32'hbca6cd7d),
	.w8(32'h3b9af521),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73c74e),
	.w1(32'hbc0d13d1),
	.w2(32'hbc2b1bac),
	.w3(32'hbc0477df),
	.w4(32'hbc046a43),
	.w5(32'h3b3b807b),
	.w6(32'h3bc7ccf1),
	.w7(32'hbc924fbd),
	.w8(32'h3afd6205),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49e906),
	.w1(32'h3b9bfeee),
	.w2(32'hbb89c28d),
	.w3(32'hbb8c4e9b),
	.w4(32'hbaa8309e),
	.w5(32'h3a4dbc74),
	.w6(32'hbb5e6512),
	.w7(32'h3b961fdb),
	.w8(32'h3adf7e8d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad2051),
	.w1(32'h3a011e18),
	.w2(32'h3939254b),
	.w3(32'h3979af85),
	.w4(32'hbba8fd93),
	.w5(32'h3c2d6fdb),
	.w6(32'hbafc5d13),
	.w7(32'hbaac0031),
	.w8(32'h3caae7a4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dbaf7),
	.w1(32'h3ba0b52e),
	.w2(32'hbc0cd059),
	.w3(32'h3bb3e711),
	.w4(32'hbc2db15b),
	.w5(32'h3bb54d97),
	.w6(32'hbb3e7f6f),
	.w7(32'hbbbb1b5f),
	.w8(32'h3bed1e93),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe28510),
	.w1(32'hbc411902),
	.w2(32'hbc206fae),
	.w3(32'hba82b4b6),
	.w4(32'hbaa7a87a),
	.w5(32'h3c03021d),
	.w6(32'h3c8fc517),
	.w7(32'hbbf40bf1),
	.w8(32'h3b841fde),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba566ed),
	.w1(32'h3b15dd99),
	.w2(32'h3b8063cd),
	.w3(32'h3bc84f8d),
	.w4(32'h3bf25c59),
	.w5(32'h3af69c57),
	.w6(32'hbc5f91c9),
	.w7(32'hbab3ee09),
	.w8(32'h3ccb822c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf822a2),
	.w1(32'hbbac21ed),
	.w2(32'hbc3e9c30),
	.w3(32'h3c33fb9c),
	.w4(32'h3a1306ea),
	.w5(32'h3ab9665f),
	.w6(32'hbc647d82),
	.w7(32'hbc47c499),
	.w8(32'hbb4499f4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a9fb6),
	.w1(32'h3bbef0c7),
	.w2(32'hbb4f3e89),
	.w3(32'h3bb76daf),
	.w4(32'hbb0da8aa),
	.w5(32'hbc0138c9),
	.w6(32'h3ba2849a),
	.w7(32'hbb2dbd4c),
	.w8(32'hbb7e090b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc018d18),
	.w1(32'hbc0d2cb3),
	.w2(32'hbc0b7be6),
	.w3(32'hbc061afa),
	.w4(32'hbbf8d160),
	.w5(32'hbbf791be),
	.w6(32'h39488dad),
	.w7(32'hbc265627),
	.w8(32'hbc96c174),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fddec),
	.w1(32'h3b926444),
	.w2(32'h3c82b812),
	.w3(32'hbb7ddc1c),
	.w4(32'h3c1bc725),
	.w5(32'h3bc4b1a9),
	.w6(32'hbc56d167),
	.w7(32'h3bff77af),
	.w8(32'h3ab5298e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd26853),
	.w1(32'h3b355869),
	.w2(32'h3b98b803),
	.w3(32'h3b3dd5ce),
	.w4(32'h3b5ea279),
	.w5(32'hb9f44eb8),
	.w6(32'h3b4ed3fa),
	.w7(32'hbba7c33d),
	.w8(32'hbb15c529),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b8968),
	.w1(32'h3abdd85b),
	.w2(32'hbc0b662f),
	.w3(32'h3b51e83b),
	.w4(32'hb98f9010),
	.w5(32'hbbb28f30),
	.w6(32'hb9c741fc),
	.w7(32'h3b04321b),
	.w8(32'hbc5c2129),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75f256),
	.w1(32'hbb469381),
	.w2(32'h3c1f2c91),
	.w3(32'h3bc0b397),
	.w4(32'h3c520dcc),
	.w5(32'h3b371125),
	.w6(32'hbbeafc81),
	.w7(32'h3c319170),
	.w8(32'h3b5fd728),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27b0be),
	.w1(32'hbbc0592b),
	.w2(32'hbb4d1f6b),
	.w3(32'h3b2f03b5),
	.w4(32'hbada1a24),
	.w5(32'h3c95e672),
	.w6(32'hba68a523),
	.w7(32'hbb743a7b),
	.w8(32'h3c1bc3a6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92fdc9),
	.w1(32'hbb4fec87),
	.w2(32'hbc338161),
	.w3(32'h3b0bb314),
	.w4(32'hbc211bda),
	.w5(32'hbb765604),
	.w6(32'h3be2036c),
	.w7(32'hbc417b60),
	.w8(32'hbb3ec463),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34b4b1),
	.w1(32'h3a86f503),
	.w2(32'hbc768e80),
	.w3(32'h3a9d2d35),
	.w4(32'hbb176976),
	.w5(32'hbc528de9),
	.w6(32'hbc030169),
	.w7(32'hbb99fafe),
	.w8(32'hbc148678),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c6f25),
	.w1(32'hbb908ff6),
	.w2(32'h3bc78dab),
	.w3(32'hb9af0869),
	.w4(32'h3bd41df8),
	.w5(32'h3c840559),
	.w6(32'h3c854851),
	.w7(32'h3c2ab876),
	.w8(32'h3c9104ba),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1afd17),
	.w1(32'hbbfa2b18),
	.w2(32'hbbb2398e),
	.w3(32'hbc608fcf),
	.w4(32'hbc0b29be),
	.w5(32'hbbb50613),
	.w6(32'hbb8dde74),
	.w7(32'hbc117e8c),
	.w8(32'hbb4aebd5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306434),
	.w1(32'hbb6a39eb),
	.w2(32'hbc190151),
	.w3(32'h3a69b3d4),
	.w4(32'hbbb1a752),
	.w5(32'h3a6f7a46),
	.w6(32'h3bc3a74c),
	.w7(32'hbc2d9cec),
	.w8(32'h3bbc1c97),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22a823),
	.w1(32'hbca67f44),
	.w2(32'hbcd3c068),
	.w3(32'hbc0dd54f),
	.w4(32'hbc928cb3),
	.w5(32'hbba0c323),
	.w6(32'hbcdc25b6),
	.w7(32'hbcedd19b),
	.w8(32'hbb56cf2f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16c6c6),
	.w1(32'hbb4b222f),
	.w2(32'hbbdd1c0f),
	.w3(32'hbba7e287),
	.w4(32'hbbd4ffc1),
	.w5(32'hbb46c0d8),
	.w6(32'hbc182c8a),
	.w7(32'hbbe013fb),
	.w8(32'h38ff6e20),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30ac2f),
	.w1(32'h3bc8c173),
	.w2(32'h3c707897),
	.w3(32'h3bd3c5bb),
	.w4(32'h3c020859),
	.w5(32'hbab50db2),
	.w6(32'hbc8b0d99),
	.w7(32'h3c8b292a),
	.w8(32'h3b8b43d4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfecc49),
	.w1(32'h3b9d3a9f),
	.w2(32'h3bb01a56),
	.w3(32'h3b3d6e30),
	.w4(32'h3bea72bc),
	.w5(32'h3b02861c),
	.w6(32'hbce2a6f5),
	.w7(32'h3b9118f3),
	.w8(32'hba73ebd1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafee343),
	.w1(32'h3bb1c35f),
	.w2(32'h3c57f030),
	.w3(32'h3bb3f452),
	.w4(32'h3bf725b9),
	.w5(32'hbc477573),
	.w6(32'hbc6cffb6),
	.w7(32'h3c7186f2),
	.w8(32'hbaa67697),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c118076),
	.w1(32'h3c0e9dad),
	.w2(32'h3c4d093d),
	.w3(32'hbbbdba83),
	.w4(32'h39b849fc),
	.w5(32'h3b36fced),
	.w6(32'hbc99c9ae),
	.w7(32'h3c7919ad),
	.w8(32'h39e87e9b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb765ea8),
	.w1(32'h3a877c5c),
	.w2(32'hbaf666ca),
	.w3(32'h3ae73193),
	.w4(32'hbb12a591),
	.w5(32'hbc021a37),
	.w6(32'hbbd144ba),
	.w7(32'hba281853),
	.w8(32'hbbfec454),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50c9d3),
	.w1(32'h3b5cf028),
	.w2(32'h3ba41cf9),
	.w3(32'hba93bfcb),
	.w4(32'hbbc81c20),
	.w5(32'h3c03f264),
	.w6(32'hb839ceed),
	.w7(32'hbb89e865),
	.w8(32'h3a58a380),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05764d),
	.w1(32'hbb7c462d),
	.w2(32'hbc23d0c0),
	.w3(32'h3bcc8bd8),
	.w4(32'hbb603c99),
	.w5(32'hbbffb60d),
	.w6(32'h3bafc509),
	.w7(32'hbbdba757),
	.w8(32'hbc594a93),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d08e2),
	.w1(32'hbb5b7009),
	.w2(32'h3c319af5),
	.w3(32'h3b4cd455),
	.w4(32'h3c1a3cd4),
	.w5(32'h3c0b9c4c),
	.w6(32'hbd139f94),
	.w7(32'h3b93fda1),
	.w8(32'h3bf1ec48),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b490010),
	.w1(32'h39b8b21c),
	.w2(32'h3bffdf14),
	.w3(32'h3b4d6513),
	.w4(32'h39f3ff98),
	.w5(32'hb91ec9a1),
	.w6(32'hbbbd3213),
	.w7(32'h3bec811a),
	.w8(32'h3c350a56),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1a878),
	.w1(32'hbb8455a0),
	.w2(32'hbc0f324f),
	.w3(32'h3aabe486),
	.w4(32'hbbde104a),
	.w5(32'hbc2a21bd),
	.w6(32'hbae34704),
	.w7(32'hbaff45eb),
	.w8(32'hbb3c9d16),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ff189),
	.w1(32'hbb92126f),
	.w2(32'hbbed2a25),
	.w3(32'hbba610d1),
	.w4(32'hbc18b91d),
	.w5(32'hbad5dd72),
	.w6(32'h3c144a31),
	.w7(32'hbbe9a361),
	.w8(32'h3c4b8874),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1da769),
	.w1(32'h3b1938a0),
	.w2(32'hbc466956),
	.w3(32'h3b9fdb0e),
	.w4(32'hbbaced64),
	.w5(32'hbc278d94),
	.w6(32'h3ba285c6),
	.w7(32'h3c34d901),
	.w8(32'hbc3088b1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26c535),
	.w1(32'h3b5958fc),
	.w2(32'h3bfbb688),
	.w3(32'hbb1e6e1a),
	.w4(32'h3ac8378d),
	.w5(32'hbc2473e9),
	.w6(32'hb840448f),
	.w7(32'h3be9ef2b),
	.w8(32'hbbe5c168),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc318945),
	.w1(32'hbb9275fb),
	.w2(32'h3be23a6a),
	.w3(32'hbb99c2f1),
	.w4(32'hba854500),
	.w5(32'hbc954864),
	.w6(32'h3aeb5353),
	.w7(32'h3c035831),
	.w8(32'hbc032696),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb78e79),
	.w1(32'h3b0c5170),
	.w2(32'hbbfe6e24),
	.w3(32'h3b64a276),
	.w4(32'h3c2ba6d2),
	.w5(32'hbc1f89af),
	.w6(32'h3c9367e2),
	.w7(32'h3ab1ecf8),
	.w8(32'hbc8e07d8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6618),
	.w1(32'hb94eefe8),
	.w2(32'h3c867bf5),
	.w3(32'hbb47a08f),
	.w4(32'h3c4ff650),
	.w5(32'hbc306a9c),
	.w6(32'hbb9feb6c),
	.w7(32'h3c895b15),
	.w8(32'hbc3ae6ef),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc561843),
	.w1(32'h3ad4870e),
	.w2(32'h3b3a94c8),
	.w3(32'hbb69ec5a),
	.w4(32'hbb00cfae),
	.w5(32'hbc308cd3),
	.w6(32'hb8865472),
	.w7(32'h3bd5a073),
	.w8(32'hbaa5b3be),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2430e3),
	.w1(32'h399b8eaa),
	.w2(32'hbb8719fd),
	.w3(32'hb8fcfca7),
	.w4(32'hbb819a12),
	.w5(32'hbb64a010),
	.w6(32'h3b8b3a69),
	.w7(32'h3b60b531),
	.w8(32'h3bf6780f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace808e),
	.w1(32'h3b37fdac),
	.w2(32'h3b2f8c4a),
	.w3(32'hb8dbbc56),
	.w4(32'hba20795f),
	.w5(32'h3c2f79b1),
	.w6(32'h3ba1636e),
	.w7(32'hbbdc32df),
	.w8(32'h3bd6d427),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf04a24),
	.w1(32'h3c1a9e6c),
	.w2(32'h3c3ae0bf),
	.w3(32'h3c86bb91),
	.w4(32'h3c6fb28c),
	.w5(32'hbaf10e78),
	.w6(32'hbc711538),
	.w7(32'h3c1438f0),
	.w8(32'h3b2556a4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5e7dd),
	.w1(32'h3bd4292a),
	.w2(32'hbbeefcb3),
	.w3(32'h3b893f6b),
	.w4(32'hbc1bed50),
	.w5(32'h3bc9c267),
	.w6(32'hbb3f21eb),
	.w7(32'hb8b0fadd),
	.w8(32'h3adeed19),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14cef0),
	.w1(32'h3bb2ec92),
	.w2(32'h3b1778b5),
	.w3(32'h3ada87f8),
	.w4(32'hb9860428),
	.w5(32'h3b88397a),
	.w6(32'h3bf4becc),
	.w7(32'h39f74e52),
	.w8(32'h3bd59ec5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f7db2),
	.w1(32'hbb163151),
	.w2(32'hb924a44a),
	.w3(32'h3ba2d182),
	.w4(32'hbbd32f45),
	.w5(32'h3b3d00f4),
	.w6(32'hbc5ec249),
	.w7(32'h394367ac),
	.w8(32'hbbca72ee),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0803f5),
	.w1(32'hbbb07d75),
	.w2(32'h3c2c63c8),
	.w3(32'h3c1e8d91),
	.w4(32'h3c1ba278),
	.w5(32'h3b8d8649),
	.w6(32'hbaabdb9a),
	.w7(32'h3bab7860),
	.w8(32'h3b9a48aa),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce9c22),
	.w1(32'h3b7b7c33),
	.w2(32'hbb65e375),
	.w3(32'hb944b128),
	.w4(32'hba675267),
	.w5(32'h3a1642a6),
	.w6(32'hbbd0a4c6),
	.w7(32'hbb0e54cf),
	.w8(32'h3c2ecba2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15dd22),
	.w1(32'hbac58810),
	.w2(32'hbc051840),
	.w3(32'hbbc6145d),
	.w4(32'hbbb211b5),
	.w5(32'h3b8db7ef),
	.w6(32'hba40902a),
	.w7(32'hbc34786e),
	.w8(32'h3beab119),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3f583),
	.w1(32'hbc139a10),
	.w2(32'hbb8d4ce7),
	.w3(32'h399e44e6),
	.w4(32'hbbda3322),
	.w5(32'h3baf3a96),
	.w6(32'hbc21911f),
	.w7(32'h3aacccf2),
	.w8(32'h3ba92d79),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7b7a9),
	.w1(32'h3a3829b9),
	.w2(32'h3c0f41ca),
	.w3(32'hbb838b34),
	.w4(32'h3b84772b),
	.w5(32'hbc4dd974),
	.w6(32'hbce69a0a),
	.w7(32'h3bcf7e15),
	.w8(32'hbc032a45),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bcf8f),
	.w1(32'hbb90f5b5),
	.w2(32'hbb994f89),
	.w3(32'hbb91b61a),
	.w4(32'hbb59cc6b),
	.w5(32'h3b1a55e3),
	.w6(32'h3c508f7b),
	.w7(32'hbb8d614f),
	.w8(32'h3b8048b8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3203c4),
	.w1(32'hbb2b1f09),
	.w2(32'hba180752),
	.w3(32'h3b8de477),
	.w4(32'hbb78ad16),
	.w5(32'h3becc23b),
	.w6(32'hbbae16f7),
	.w7(32'hbbf3f23e),
	.w8(32'h3b6e4925),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb366f),
	.w1(32'h3c1f18ba),
	.w2(32'h3b8e6384),
	.w3(32'h39a912dd),
	.w4(32'h3b97a6a7),
	.w5(32'h3b63e98c),
	.w6(32'hbc6908c4),
	.w7(32'h3ca68a60),
	.w8(32'h3bda3c30),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b763c5c),
	.w1(32'h3bcb53f5),
	.w2(32'hbc3ebd7a),
	.w3(32'hbb6b325b),
	.w4(32'hbb2c3990),
	.w5(32'hbbf9cf09),
	.w6(32'hbc24d3f0),
	.w7(32'h399f121a),
	.w8(32'hbc6012d6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ac472),
	.w1(32'hbbaea69f),
	.w2(32'hbb5109ae),
	.w3(32'hbc28f5a3),
	.w4(32'hbb3800ad),
	.w5(32'hbc168904),
	.w6(32'h3ad4449c),
	.w7(32'hbc0f2af1),
	.w8(32'hbbf6aeb6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccb402),
	.w1(32'hbc3f8862),
	.w2(32'hbc3c5009),
	.w3(32'hbc1ab800),
	.w4(32'hbc2d6147),
	.w5(32'hbba3c3dd),
	.w6(32'h3b29e750),
	.w7(32'hbc63e58c),
	.w8(32'hbca0ace5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0e094),
	.w1(32'h3b493c45),
	.w2(32'h3cb2b41b),
	.w3(32'hbb5fd4b0),
	.w4(32'h3c69221f),
	.w5(32'h3be185ed),
	.w6(32'hbce0f0ab),
	.w7(32'h3c6713fe),
	.w8(32'h3c829aeb),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba585dc5),
	.w1(32'h3bc3f3e2),
	.w2(32'h3ba44f5a),
	.w3(32'hbbc63ba2),
	.w4(32'hbc0dc59e),
	.w5(32'hbafd4068),
	.w6(32'hbbb2802e),
	.w7(32'h3b6f8c2e),
	.w8(32'hba8c3d82),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9b38),
	.w1(32'h3bf44332),
	.w2(32'h3aee857a),
	.w3(32'h3b65f1ec),
	.w4(32'hba43e27a),
	.w5(32'hbae08e2c),
	.w6(32'hbc12f30b),
	.w7(32'h3c0d3480),
	.w8(32'hbb042e42),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56dbe8),
	.w1(32'h3a0eb4e6),
	.w2(32'h3a284a13),
	.w3(32'hbb9c735e),
	.w4(32'h3c031070),
	.w5(32'h3bb98370),
	.w6(32'hbbbe41e7),
	.w7(32'hbb971c7d),
	.w8(32'h3c10b505),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a064),
	.w1(32'hbbb430b5),
	.w2(32'h3b82a65e),
	.w3(32'h3c4f4c4a),
	.w4(32'hbaa13af2),
	.w5(32'h3ba7d529),
	.w6(32'h3bd5aa08),
	.w7(32'h3b9b1c0d),
	.w8(32'hbba2f4d2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be904e7),
	.w1(32'h3886ea7d),
	.w2(32'hbc45e2b6),
	.w3(32'hbbfdce79),
	.w4(32'hbb2bfbcf),
	.w5(32'h3c5481af),
	.w6(32'h3b38c689),
	.w7(32'hbc57918f),
	.w8(32'h3c39696d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c0f1b),
	.w1(32'h3968773d),
	.w2(32'h3b962871),
	.w3(32'h3b7786b9),
	.w4(32'h3bde87b9),
	.w5(32'h3af96c70),
	.w6(32'hbc4384ac),
	.w7(32'h3c1d8082),
	.w8(32'h3b9fa19e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb714ceb),
	.w1(32'h3ab370a1),
	.w2(32'hbbe1223d),
	.w3(32'hbb99047e),
	.w4(32'hbbfefa78),
	.w5(32'h3bbcb04a),
	.w6(32'hbbe0c248),
	.w7(32'hbb263e03),
	.w8(32'h3c3939b1),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74be90),
	.w1(32'h3b38aaef),
	.w2(32'h3b96b300),
	.w3(32'h3b358f47),
	.w4(32'h3b27350a),
	.w5(32'h3c861ea9),
	.w6(32'hbc90cb0b),
	.w7(32'h3b73b87e),
	.w8(32'h3c8b37cd),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b960da4),
	.w1(32'hbb12bf6c),
	.w2(32'hbbeb942e),
	.w3(32'h3b8fb01c),
	.w4(32'h3bb81b6d),
	.w5(32'hbc07f804),
	.w6(32'hbb3489d9),
	.w7(32'hbb98ea90),
	.w8(32'hbc33ae1e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc00fad),
	.w1(32'hbb279050),
	.w2(32'h3bad64d8),
	.w3(32'hbbee4895),
	.w4(32'hbb3d72ad),
	.w5(32'hb9c957be),
	.w6(32'h3b356552),
	.w7(32'h3b8e5214),
	.w8(32'hba23dd77),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcab4bb),
	.w1(32'h3b0acfb8),
	.w2(32'h3b81bccc),
	.w3(32'h399cb74f),
	.w4(32'h3baa328d),
	.w5(32'hbc1c23fc),
	.w6(32'hbc8a16ca),
	.w7(32'h3c501350),
	.w8(32'hbc7e0380),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3cb81),
	.w1(32'hbbc3b8a2),
	.w2(32'hbb946d3c),
	.w3(32'hbc27d1dc),
	.w4(32'hbbe6a225),
	.w5(32'h3b285d58),
	.w6(32'hbaed4e87),
	.w7(32'hbb771a8e),
	.w8(32'h3b68669b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2f7d0),
	.w1(32'hbb994737),
	.w2(32'h3bc54e27),
	.w3(32'h3ba03d94),
	.w4(32'h3b876073),
	.w5(32'hbb93fe74),
	.w6(32'hbbc78f4d),
	.w7(32'h3b3c0edd),
	.w8(32'hbc0897f6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfab08),
	.w1(32'hbbd0aead),
	.w2(32'hbc0252dc),
	.w3(32'hbba59563),
	.w4(32'hbc02b4f4),
	.w5(32'h3b7a5559),
	.w6(32'h3bbe7459),
	.w7(32'hbc570a60),
	.w8(32'h3bcd67b8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba4073),
	.w1(32'hbb8e6c78),
	.w2(32'hbb764155),
	.w3(32'hb8ed5d1c),
	.w4(32'hbb8aac04),
	.w5(32'hbacf5ae5),
	.w6(32'hb9ff6543),
	.w7(32'hbb3f3fe3),
	.w8(32'h3c66ac4a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85712b),
	.w1(32'h3b3662fb),
	.w2(32'hbbf86fff),
	.w3(32'hbbd2171f),
	.w4(32'hbc84f6b7),
	.w5(32'h3adeed52),
	.w6(32'h3cab1b90),
	.w7(32'hbc207eb9),
	.w8(32'h3b188e74),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b319ba2),
	.w1(32'hbc0aa007),
	.w2(32'hbc929045),
	.w3(32'hbc567b57),
	.w4(32'hbc4052eb),
	.w5(32'h3be27b48),
	.w6(32'hbb51f432),
	.w7(32'hbca8a20d),
	.w8(32'h3a9bde67),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be43202),
	.w1(32'hb87b1339),
	.w2(32'h3bb146e9),
	.w3(32'h3b28827c),
	.w4(32'h3c1242a7),
	.w5(32'h3c06e057),
	.w6(32'hbc02d0c5),
	.w7(32'hbbeb1a7e),
	.w8(32'h3c840c7b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13df7d),
	.w1(32'hbc4f5b9e),
	.w2(32'hbc950143),
	.w3(32'hbc07cea2),
	.w4(32'hbc359584),
	.w5(32'hbc482c97),
	.w6(32'hbc629dec),
	.w7(32'hbca10afc),
	.w8(32'hbc97fa03),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50e51a),
	.w1(32'hba267e7d),
	.w2(32'h3c4ec438),
	.w3(32'h3b41efff),
	.w4(32'h3c2e227d),
	.w5(32'h3b884aa6),
	.w6(32'h3c146ed3),
	.w7(32'h3c838891),
	.w8(32'hbb824fdb),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c124eb1),
	.w1(32'h3c8c411e),
	.w2(32'h3c93453e),
	.w3(32'h3bc8d1a6),
	.w4(32'h3c82cb35),
	.w5(32'hbc6cc49f),
	.w6(32'hbc9c8381),
	.w7(32'h3c7ef8a9),
	.w8(32'hbc523d58),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70b75f),
	.w1(32'hbbd834d4),
	.w2(32'hbb9490be),
	.w3(32'hb5f611ac),
	.w4(32'hbadd0d80),
	.w5(32'hbae9661f),
	.w6(32'h3c5b07c9),
	.w7(32'hbb1d5352),
	.w8(32'hbb8859e4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc053e47),
	.w1(32'hbbad3dfa),
	.w2(32'hbb45d06e),
	.w3(32'hbb9294b5),
	.w4(32'h3c31856b),
	.w5(32'h3ba90845),
	.w6(32'hbbcfd950),
	.w7(32'h3ab8c0ac),
	.w8(32'h3b8c122f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08dd2d),
	.w1(32'hbb2e37da),
	.w2(32'hbc0614c3),
	.w3(32'hbc376f4f),
	.w4(32'hbc73933c),
	.w5(32'hbb6980df),
	.w6(32'h39a265b4),
	.w7(32'hbc09a358),
	.w8(32'h3bf4a66b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4b80),
	.w1(32'hbc017f30),
	.w2(32'hbc14f18d),
	.w3(32'h39ce9a2e),
	.w4(32'h3b1317a5),
	.w5(32'h3c2a4e69),
	.w6(32'hbbec1195),
	.w7(32'hbb7d8ec4),
	.w8(32'hbb060906),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb684c6f),
	.w1(32'h393ac650),
	.w2(32'h3be811e0),
	.w3(32'h3c40ad5a),
	.w4(32'h3bf5e3d4),
	.w5(32'h3bc664c4),
	.w6(32'hbbe42b3f),
	.w7(32'hbaff46cd),
	.w8(32'h3c1af365),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e5cf3),
	.w1(32'hbba17825),
	.w2(32'hbb0d6711),
	.w3(32'hb9a67e13),
	.w4(32'hbc6d1656),
	.w5(32'h3c05ed6f),
	.w6(32'hbb6e3b60),
	.w7(32'h3ab0440a),
	.w8(32'h3ba28ac1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4643c7),
	.w1(32'h3b57cf2b),
	.w2(32'hbbba1ae3),
	.w3(32'h3bd01e6a),
	.w4(32'hbb8418dd),
	.w5(32'h3bac736d),
	.w6(32'hbc15932e),
	.w7(32'hbb3c7bf0),
	.w8(32'hbb5ff5c1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcd434),
	.w1(32'hba2e9021),
	.w2(32'h3b8005f8),
	.w3(32'h3ac19a63),
	.w4(32'h3b5a5b9e),
	.w5(32'h3bd83673),
	.w6(32'hbb16d86e),
	.w7(32'h3bd69795),
	.w8(32'h3c5ce46e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb5482),
	.w1(32'h3bac6e01),
	.w2(32'h3b21d3c1),
	.w3(32'h3c67b524),
	.w4(32'h3a466f4b),
	.w5(32'hbc3ee615),
	.w6(32'h3bc77624),
	.w7(32'hba13ed89),
	.w8(32'hbc5fcf34),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f359c),
	.w1(32'hbbd82e19),
	.w2(32'hbab1e7d6),
	.w3(32'h3933aa90),
	.w4(32'h3aff61e1),
	.w5(32'hbc059b01),
	.w6(32'h3c44928e),
	.w7(32'h3b31816b),
	.w8(32'h3bcc2b6e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7893c),
	.w1(32'hbba782c4),
	.w2(32'hbc4e14e5),
	.w3(32'hbb80dfb2),
	.w4(32'hbb5a4615),
	.w5(32'hbb0f0db4),
	.w6(32'h3cc6a07e),
	.w7(32'hbafd1432),
	.w8(32'hbb7b5362),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16d7be),
	.w1(32'h3bb2cc97),
	.w2(32'h3a76c067),
	.w3(32'h3b3a5f69),
	.w4(32'h3bce45e6),
	.w5(32'hbb3428f8),
	.w6(32'hbbe97c75),
	.w7(32'h3bddd026),
	.w8(32'hbb205edc),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc166655),
	.w1(32'hbbc1a896),
	.w2(32'hbbb8b53d),
	.w3(32'hba85ca2e),
	.w4(32'hbb81aebd),
	.w5(32'hbb1d4c15),
	.w6(32'hbb8c0b6d),
	.w7(32'hbbd0fa04),
	.w8(32'h3b5e90ce),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978f87),
	.w1(32'hbb31465b),
	.w2(32'hbc63e95b),
	.w3(32'h3956a768),
	.w4(32'hbb0d84b5),
	.w5(32'h3c28b7fc),
	.w6(32'hbbd6a8e9),
	.w7(32'h3a9c11d2),
	.w8(32'h3c2997fa),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8efbc3),
	.w1(32'h3b487414),
	.w2(32'hbbcb4afa),
	.w3(32'h3b8738ae),
	.w4(32'hbbe7c669),
	.w5(32'h3ae79ea5),
	.w6(32'hbbdc58d4),
	.w7(32'hbaf355d5),
	.w8(32'h3c006303),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb883def),
	.w1(32'h3b09e1b5),
	.w2(32'h3b726010),
	.w3(32'hb94d96f7),
	.w4(32'hbc6c69c9),
	.w5(32'hba9097fb),
	.w6(32'hbbe40bb3),
	.w7(32'h3b9ba961),
	.w8(32'h3beb1784),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffad18),
	.w1(32'hbb42f1f3),
	.w2(32'hbb9f0ba5),
	.w3(32'hb9ca88e6),
	.w4(32'hbc0f00b9),
	.w5(32'hbbff1c4d),
	.w6(32'hbbacf554),
	.w7(32'hbb51ab89),
	.w8(32'h3b155a41),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb675b88),
	.w1(32'h3ad8d9d5),
	.w2(32'hba864bc5),
	.w3(32'h3c20ba27),
	.w4(32'h3a2d3f08),
	.w5(32'h3c42ceba),
	.w6(32'h3b0606e5),
	.w7(32'hbb6cfc4c),
	.w8(32'h3b6f58eb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d1e27),
	.w1(32'h3cae99df),
	.w2(32'h3c93fddd),
	.w3(32'h3b041926),
	.w4(32'h3c31980f),
	.w5(32'hbbbfca08),
	.w6(32'h3be33abc),
	.w7(32'h3c96eabf),
	.w8(32'hbc1e5da5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37207a3d),
	.w1(32'hba22e1c1),
	.w2(32'hb822b0fa),
	.w3(32'hbb08b158),
	.w4(32'hbb8a927e),
	.w5(32'h3b685b88),
	.w6(32'hba119b6e),
	.w7(32'h3c3e88b5),
	.w8(32'h3bc1bfff),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88dd10),
	.w1(32'hbb55a292),
	.w2(32'hbb062aca),
	.w3(32'h3c12b7db),
	.w4(32'h3a5e0e06),
	.w5(32'h3b082bd2),
	.w6(32'h3c9c63cf),
	.w7(32'hbc589958),
	.w8(32'h3b86f429),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fc7f3),
	.w1(32'hbb9d125b),
	.w2(32'hbc1a5866),
	.w3(32'hbbbcbe09),
	.w4(32'hbc0ab8fb),
	.w5(32'h3ab8822f),
	.w6(32'h3bca6d0f),
	.w7(32'hbc475408),
	.w8(32'h3b8bd02f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1528a8),
	.w1(32'h3c1cdb4d),
	.w2(32'h3bac261a),
	.w3(32'hba2c0c5f),
	.w4(32'h3c1349e4),
	.w5(32'hbb5fe706),
	.w6(32'hbc42b25d),
	.w7(32'h3b808672),
	.w8(32'hbb589dac),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b0f7),
	.w1(32'h3bb70b9a),
	.w2(32'h3c9da570),
	.w3(32'hbbbf757c),
	.w4(32'h3a0d0a02),
	.w5(32'h3bcddccf),
	.w6(32'hbca89c70),
	.w7(32'h3c0cfb9d),
	.w8(32'h3bfa00fc),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4aaea8),
	.w1(32'h3bb06b3e),
	.w2(32'h3c389320),
	.w3(32'h3bc1d7ba),
	.w4(32'h3c0aea4d),
	.w5(32'hbadc7add),
	.w6(32'hbc0ed5a2),
	.w7(32'h3c36172a),
	.w8(32'h3ad6944f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6f28c),
	.w1(32'hbb3c2d85),
	.w2(32'h3be843a3),
	.w3(32'h3c21ac47),
	.w4(32'h3b89c2f4),
	.w5(32'h3c28399a),
	.w6(32'hbbd9c878),
	.w7(32'h3ba693e3),
	.w8(32'h3c254b50),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33e0e4),
	.w1(32'h3c80098c),
	.w2(32'h3c30298a),
	.w3(32'h3c0c7953),
	.w4(32'h3c203c94),
	.w5(32'hb8e46c35),
	.w6(32'hbc55338a),
	.w7(32'h3c50bfa8),
	.w8(32'h3b6a991b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f821c),
	.w1(32'hbbf61d4d),
	.w2(32'hbb1aeb07),
	.w3(32'h3badbcf5),
	.w4(32'hbb1723a3),
	.w5(32'h3c43829d),
	.w6(32'hba161910),
	.w7(32'hbbdbe204),
	.w8(32'h3c915dd7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72428),
	.w1(32'hbbe108d2),
	.w2(32'hbc7ea993),
	.w3(32'hb79f367a),
	.w4(32'hbc46e2c4),
	.w5(32'hbbe2c207),
	.w6(32'h3b8fd26c),
	.w7(32'hbc614162),
	.w8(32'hbbf99bc2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb19bd),
	.w1(32'h3bea53d3),
	.w2(32'h3bff0ba3),
	.w3(32'hba0c4956),
	.w4(32'h3b2972e8),
	.w5(32'hb8b9a3dd),
	.w6(32'hbc0ba7c8),
	.w7(32'h3b92827a),
	.w8(32'hbbeb4b20),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9839f01),
	.w1(32'h3c2bd3cb),
	.w2(32'h3c934b4c),
	.w3(32'hbac24497),
	.w4(32'h3c3b97f8),
	.w5(32'hbbab84f9),
	.w6(32'hbc4148d6),
	.w7(32'h3c38762e),
	.w8(32'h3b1a1751),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d1233),
	.w1(32'h3c4df0bc),
	.w2(32'h3bc7ac38),
	.w3(32'h3c082df6),
	.w4(32'h3c2cfc22),
	.w5(32'h3b3e702e),
	.w6(32'h3c1a7c38),
	.w7(32'h3c00da32),
	.w8(32'hba723814),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c02f00),
	.w1(32'h3b8579c3),
	.w2(32'h3b8f6162),
	.w3(32'h3ba16e62),
	.w4(32'h3bd45a4c),
	.w5(32'hbb836d5f),
	.w6(32'hbc52ce17),
	.w7(32'h3b214c9c),
	.w8(32'h38d6d3d8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64fae5),
	.w1(32'h38501e6d),
	.w2(32'hbb2dbb6d),
	.w3(32'hbb484755),
	.w4(32'hba92487d),
	.w5(32'hba1f4359),
	.w6(32'hbbf8ec07),
	.w7(32'h38f42c82),
	.w8(32'h3ba8f6fd),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f4e5d),
	.w1(32'h3ca28423),
	.w2(32'h3c10b309),
	.w3(32'h3b82b17a),
	.w4(32'hb9ca978e),
	.w5(32'h3a22a479),
	.w6(32'h3c7de5fc),
	.w7(32'h3c108fa9),
	.w8(32'h3af04a73),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca4d6),
	.w1(32'hbc032768),
	.w2(32'hbbbc5427),
	.w3(32'hbb2714c6),
	.w4(32'hbb4cde59),
	.w5(32'hbb403bec),
	.w6(32'hbc06f0af),
	.w7(32'hbbe06f16),
	.w8(32'hb9b2ad72),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce4434),
	.w1(32'h3c4bcd78),
	.w2(32'h3b3b9aa1),
	.w3(32'h3b52fde4),
	.w4(32'h3add54f5),
	.w5(32'hbbe43cf0),
	.w6(32'hbb856079),
	.w7(32'h3ba8e7fc),
	.w8(32'h3b957902),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88f57d),
	.w1(32'hbb9b4370),
	.w2(32'hbc10f1b5),
	.w3(32'h39dad44f),
	.w4(32'hbb64e3b4),
	.w5(32'h3aef8e57),
	.w6(32'h3bb6a35b),
	.w7(32'hbc07fa02),
	.w8(32'h3ba944f1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ce426),
	.w1(32'h3b8deac7),
	.w2(32'hbacc1ff3),
	.w3(32'hb9d584df),
	.w4(32'h3af7d024),
	.w5(32'h3ae230f7),
	.w6(32'hbbcdb1cd),
	.w7(32'h3a8fba3b),
	.w8(32'hbb941cb6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0b701),
	.w1(32'hbad30adc),
	.w2(32'h3c3904eb),
	.w3(32'h3be72c9b),
	.w4(32'h3c1f57cb),
	.w5(32'h39a26190),
	.w6(32'h3c14c4a9),
	.w7(32'h3c2ec6ba),
	.w8(32'hbb90fea5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae54cbb),
	.w1(32'hbb44563e),
	.w2(32'h3be0632c),
	.w3(32'hb9bdc68d),
	.w4(32'h3bc35ddd),
	.w5(32'hb8bfab86),
	.w6(32'hbc1fdea5),
	.w7(32'h3c7a2dfd),
	.w8(32'hbbaa7774),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f9c98),
	.w1(32'hbbbe998d),
	.w2(32'h3c6ef7c0),
	.w3(32'hba5819b0),
	.w4(32'h3bf91369),
	.w5(32'hbb0668b6),
	.w6(32'hbc654381),
	.w7(32'h3c9135fe),
	.w8(32'hbb2c854d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe43a8e),
	.w1(32'hba3ae362),
	.w2(32'hbc20265c),
	.w3(32'hbb773a7e),
	.w4(32'hbc4437a5),
	.w5(32'h3bf348bf),
	.w6(32'hba40d9c2),
	.w7(32'hbba8f8be),
	.w8(32'h3c07f0f3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb79a77),
	.w1(32'hbbf4031d),
	.w2(32'hbc64504f),
	.w3(32'h39c62c5f),
	.w4(32'hbc385b7d),
	.w5(32'hbc00d75c),
	.w6(32'h3ba615f2),
	.w7(32'hbbf07182),
	.w8(32'hbb3204bf),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb77aae),
	.w1(32'h3b885e0b),
	.w2(32'hbb8f87da),
	.w3(32'h3b845f95),
	.w4(32'hbb9741d8),
	.w5(32'hbbd174e6),
	.w6(32'h3b9f8c91),
	.w7(32'hbb155c4b),
	.w8(32'hbbca8ec2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb529c0d),
	.w1(32'h3b464462),
	.w2(32'h3be8bcf9),
	.w3(32'hbaf024f1),
	.w4(32'h3bdcdccb),
	.w5(32'h3afe0be4),
	.w6(32'hba79f505),
	.w7(32'h3c500961),
	.w8(32'h3c56859a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b885c6c),
	.w1(32'hbc3901d9),
	.w2(32'hbab56e49),
	.w3(32'h3b5a27ae),
	.w4(32'hbbf870d0),
	.w5(32'hbbc9574a),
	.w6(32'h3b974ae2),
	.w7(32'hbb9fe4a7),
	.w8(32'hbc10655d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa89a4),
	.w1(32'h3c281e08),
	.w2(32'h3ba58606),
	.w3(32'h3a577161),
	.w4(32'hb9b3729d),
	.w5(32'h3b81403e),
	.w6(32'hb957396b),
	.w7(32'h3beb9512),
	.w8(32'hbb8e3d84),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6f6fe),
	.w1(32'h3b36c48b),
	.w2(32'hbb459138),
	.w3(32'hbb755b44),
	.w4(32'h3b8d916b),
	.w5(32'hba30ddd6),
	.w6(32'h3c1262fd),
	.w7(32'h3b8b563d),
	.w8(32'hba317384),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6a547),
	.w1(32'hbacfa7e9),
	.w2(32'hba67ca40),
	.w3(32'hbaaf89ec),
	.w4(32'hba5a19d3),
	.w5(32'hba0a08b7),
	.w6(32'hbb001f8b),
	.w7(32'hbad5283d),
	.w8(32'h3b34d343),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b3dd6),
	.w1(32'hbb92f8d8),
	.w2(32'hbb88753e),
	.w3(32'h3ab27701),
	.w4(32'hb9a51e36),
	.w5(32'hba533b1a),
	.w6(32'hbb2a747f),
	.w7(32'hb9e08057),
	.w8(32'hba998862),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac26bff),
	.w1(32'h39ba22d1),
	.w2(32'hb9f45b0a),
	.w3(32'h39f3b76a),
	.w4(32'h3ab3b84f),
	.w5(32'h3990b48d),
	.w6(32'hbb018f43),
	.w7(32'hbae4368c),
	.w8(32'h3b4dd363),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820f46),
	.w1(32'hbb31f64b),
	.w2(32'hba5cb2bd),
	.w3(32'hbb351b4a),
	.w4(32'h3b45e5f1),
	.w5(32'h3a368a93),
	.w6(32'h3a09c018),
	.w7(32'hba22c5d1),
	.w8(32'hb93b6e30),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19147e),
	.w1(32'hbb32712d),
	.w2(32'hbb3141f7),
	.w3(32'hbb20f1c4),
	.w4(32'hb9b979b3),
	.w5(32'hbbc1b7c5),
	.w6(32'h389b4071),
	.w7(32'hb9b79d0f),
	.w8(32'hbaadb890),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7402a6),
	.w1(32'h3b037bb6),
	.w2(32'hbaf9b532),
	.w3(32'hbb30b092),
	.w4(32'hbb328c97),
	.w5(32'hb93aeca8),
	.w6(32'hba31ec71),
	.w7(32'hb963bd9c),
	.w8(32'hbb01e167),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec477b),
	.w1(32'hbb17b5f6),
	.w2(32'hb96ac8d3),
	.w3(32'h3a64f274),
	.w4(32'h3a78ca3a),
	.w5(32'h3b02b12f),
	.w6(32'hba63c0dc),
	.w7(32'hb7eea5f3),
	.w8(32'h3ba1a040),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccf9c1),
	.w1(32'h39091fdb),
	.w2(32'h39ff351f),
	.w3(32'h3bb63d3d),
	.w4(32'h3b8ba306),
	.w5(32'h3afa67a9),
	.w6(32'h3a826c5b),
	.w7(32'h3acb7ee5),
	.w8(32'h3afd0c4d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac759fe),
	.w1(32'hbaa2f6bb),
	.w2(32'hbb100949),
	.w3(32'h3b3c2b05),
	.w4(32'h3b419313),
	.w5(32'hba71c7a4),
	.w6(32'h3b060e84),
	.w7(32'hbad92b7a),
	.w8(32'hba7bbe0a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ed5b9),
	.w1(32'hb7365732),
	.w2(32'h38cc6963),
	.w3(32'hb8d8e110),
	.w4(32'h39af5606),
	.w5(32'h37e42928),
	.w6(32'h39a7f657),
	.w7(32'h3a80c038),
	.w8(32'hba96fb4d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fdaae),
	.w1(32'hbab805a6),
	.w2(32'hbad3f2b1),
	.w3(32'hba954b58),
	.w4(32'hbaac43d8),
	.w5(32'hba1248c1),
	.w6(32'hbb2db043),
	.w7(32'hbb4dcee5),
	.w8(32'hb89ccc98),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35161d),
	.w1(32'hba43a5e3),
	.w2(32'hba3f1c79),
	.w3(32'hba17cb00),
	.w4(32'hb9f2700b),
	.w5(32'hbaac5d4b),
	.w6(32'hba7d2c26),
	.w7(32'hbaf111b3),
	.w8(32'hbab02443),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e34eff),
	.w1(32'hbac6586d),
	.w2(32'hbac57fcf),
	.w3(32'hba7741e7),
	.w4(32'h3a9aefd7),
	.w5(32'hbacecc12),
	.w6(32'hbb353e3c),
	.w7(32'hba5625c4),
	.w8(32'h3ab48f45),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd3f06),
	.w1(32'hbadcfcb7),
	.w2(32'hba99cfeb),
	.w3(32'hbad035f7),
	.w4(32'h3ae7505a),
	.w5(32'hbb14e462),
	.w6(32'h3b028c45),
	.w7(32'h3a6d0b15),
	.w8(32'h398b51ac),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba361d4a),
	.w1(32'hbaa216e1),
	.w2(32'hba4817f3),
	.w3(32'h3a090325),
	.w4(32'h3aed038e),
	.w5(32'hb99b871d),
	.w6(32'h3a8a03c4),
	.w7(32'hbac6f6e6),
	.w8(32'h3a31f399),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d6776),
	.w1(32'h3a297897),
	.w2(32'h3b0dcb24),
	.w3(32'hba0779cf),
	.w4(32'h3a0f0f95),
	.w5(32'hbaef8657),
	.w6(32'hba31e493),
	.w7(32'h3b049aa4),
	.w8(32'hbaab2e93),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35b66a),
	.w1(32'hbb1f11af),
	.w2(32'h3ab970d4),
	.w3(32'hba4ac4cd),
	.w4(32'hbacaecdc),
	.w5(32'hbaa5083e),
	.w6(32'h381eb3e9),
	.w7(32'h39870630),
	.w8(32'h3b802713),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add019b),
	.w1(32'hba45ef3f),
	.w2(32'hb89bd9d7),
	.w3(32'hba2447dd),
	.w4(32'h3b81fdb0),
	.w5(32'hb90959ab),
	.w6(32'h3bb2b410),
	.w7(32'h3b3b8b97),
	.w8(32'hb9b52f7d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7be38a),
	.w1(32'hb9c3d641),
	.w2(32'hba458ace),
	.w3(32'hb9eba536),
	.w4(32'hb9f357ee),
	.w5(32'h3a5a09c8),
	.w6(32'hb9c373d8),
	.w7(32'hba4b8680),
	.w8(32'hba8936f1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5b5c9),
	.w1(32'hbb7a0295),
	.w2(32'hbaf66fd6),
	.w3(32'h3950212d),
	.w4(32'h39c154f2),
	.w5(32'h3b14657f),
	.w6(32'hbb4eefff),
	.w7(32'h38aa4b57),
	.w8(32'h3b01a069),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18ec6d),
	.w1(32'hb9959df7),
	.w2(32'hb9410242),
	.w3(32'hb9f61fad),
	.w4(32'h392fe518),
	.w5(32'hbbcbe63b),
	.w6(32'hba766259),
	.w7(32'hb9006e1b),
	.w8(32'hbbb56773),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d1170),
	.w1(32'hbb0dbd32),
	.w2(32'hbb8ad273),
	.w3(32'hbbe24f96),
	.w4(32'hbb3e7b9f),
	.w5(32'hbb960c33),
	.w6(32'hbbf8b8b1),
	.w7(32'hbbb50d70),
	.w8(32'hbad4b45f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc508c),
	.w1(32'h3ade61ff),
	.w2(32'h3a80ef6e),
	.w3(32'hbb87c01f),
	.w4(32'hbb790c4b),
	.w5(32'hbac44d7a),
	.w6(32'hba0a964b),
	.w7(32'h3942521e),
	.w8(32'hb95b1df7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaa7d0),
	.w1(32'h3aadcee5),
	.w2(32'h3adfef83),
	.w3(32'hba0b32e8),
	.w4(32'hbac16804),
	.w5(32'hbae95ed5),
	.w6(32'h3b00eea3),
	.w7(32'h3afc7737),
	.w8(32'h3b735fbb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909cd3),
	.w1(32'hbbbe0ace),
	.w2(32'hbba92da0),
	.w3(32'hb9a43cee),
	.w4(32'h3af08947),
	.w5(32'h3a140235),
	.w6(32'h38b18978),
	.w7(32'hba37bd29),
	.w8(32'h395d85ab),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b097adf),
	.w1(32'h3aa2c63d),
	.w2(32'h3aa37242),
	.w3(32'h3b072dc5),
	.w4(32'h3a55dbac),
	.w5(32'h3908138d),
	.w6(32'h3a797a1c),
	.w7(32'hba2628a3),
	.w8(32'h3aab2b92),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbe2f8),
	.w1(32'hbb4803ff),
	.w2(32'hbb0eb1e6),
	.w3(32'hbb2ae59e),
	.w4(32'h39a99e00),
	.w5(32'hb9255910),
	.w6(32'h3b621630),
	.w7(32'h3b162e6b),
	.w8(32'hbb1da58c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0e7a8),
	.w1(32'hbab80be8),
	.w2(32'h3af9f05d),
	.w3(32'h39629d9d),
	.w4(32'h3a40c068),
	.w5(32'hba7bdc20),
	.w6(32'hba94a9f1),
	.w7(32'h3b1edcad),
	.w8(32'hbaaec652),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41484a),
	.w1(32'hb932fd08),
	.w2(32'hb975f6d6),
	.w3(32'h384ec7f2),
	.w4(32'hbae8383e),
	.w5(32'hb76aa4c1),
	.w6(32'h39d23b75),
	.w7(32'h3a26f503),
	.w8(32'hbb04f831),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6af5100),
	.w1(32'h395d9d4e),
	.w2(32'h38a4d825),
	.w3(32'h39b1a864),
	.w4(32'h3a38f20e),
	.w5(32'h394fef20),
	.w6(32'hbb28db0a),
	.w7(32'hba832d85),
	.w8(32'h3b21c7e3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule