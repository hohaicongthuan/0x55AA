module layer_10_featuremap_210(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90abd8f),
	.w1(32'hba101a31),
	.w2(32'hbaf55fa9),
	.w3(32'hb9584f3c),
	.w4(32'hb9c61176),
	.w5(32'hbac79c93),
	.w6(32'hb9be5ec5),
	.w7(32'hb9a93149),
	.w8(32'hb8b57a71),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28a177),
	.w1(32'h3a6a0264),
	.w2(32'hba1b0579),
	.w3(32'hbb49606f),
	.w4(32'h3a8e46a6),
	.w5(32'h38821705),
	.w6(32'hb98fbdd7),
	.w7(32'h38dfc086),
	.w8(32'h3a23c662),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea8a65),
	.w1(32'hb9ea333d),
	.w2(32'hba7543e9),
	.w3(32'h39fef5ca),
	.w4(32'hb99618bd),
	.w5(32'hb9c5504f),
	.w6(32'hba1ca407),
	.w7(32'hba4474e1),
	.w8(32'hb9dd01b8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba551140),
	.w1(32'hbaa3404b),
	.w2(32'hba057529),
	.w3(32'hb97c38a7),
	.w4(32'h3916595b),
	.w5(32'h3aa12f69),
	.w6(32'hb8a37808),
	.w7(32'hb937cae0),
	.w8(32'h3a77e911),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ad891),
	.w1(32'h39994d3c),
	.w2(32'hb9c27228),
	.w3(32'h3a7d5eb9),
	.w4(32'h39bad821),
	.w5(32'hb9adab5c),
	.w6(32'h39e7b90f),
	.w7(32'hb9bb5681),
	.w8(32'hb86eeec3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ab297),
	.w1(32'hba543a79),
	.w2(32'hba314cd1),
	.w3(32'hb9b99dd9),
	.w4(32'hba507819),
	.w5(32'hba25df0b),
	.w6(32'hba22c3ba),
	.w7(32'hba3d1051),
	.w8(32'hba280a5f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10469a),
	.w1(32'h3a24dd7d),
	.w2(32'h3b683015),
	.w3(32'hb9e49d3a),
	.w4(32'h3b1d77e4),
	.w5(32'h3ab788df),
	.w6(32'h3ac64db1),
	.w7(32'h3b4bf801),
	.w8(32'h3adaed9e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd25dc),
	.w1(32'hbbc5441c),
	.w2(32'hbb92125e),
	.w3(32'h3b61538e),
	.w4(32'hbbaca669),
	.w5(32'hbbff1187),
	.w6(32'h3a45f938),
	.w7(32'hba80a971),
	.w8(32'hbbbe6e47),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacac468),
	.w1(32'hba670ca5),
	.w2(32'hba59d37b),
	.w3(32'hba53427e),
	.w4(32'hb928f54f),
	.w5(32'hb999dd1d),
	.w6(32'hb940d427),
	.w7(32'h376bd6d2),
	.w8(32'hb9d28607),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba519407),
	.w1(32'h3ac4aa24),
	.w2(32'h3a7b3912),
	.w3(32'h3a269d5b),
	.w4(32'h399d1917),
	.w5(32'hbb17637e),
	.w6(32'h3b96fc8f),
	.w7(32'h3b35377e),
	.w8(32'hba4bae5b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ccca7),
	.w1(32'hb8dde2fe),
	.w2(32'h395ce297),
	.w3(32'h3a8fb0af),
	.w4(32'h3953011d),
	.w5(32'h3a026dda),
	.w6(32'hba3f2013),
	.w7(32'hba2c91d6),
	.w8(32'hba18f553),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7f5dd),
	.w1(32'hb9a57380),
	.w2(32'h3bba9155),
	.w3(32'h3b8b6357),
	.w4(32'h3b1fd5fe),
	.w5(32'h3ba4de86),
	.w6(32'h3b37dba2),
	.w7(32'h3b30c3e3),
	.w8(32'h3b3af09e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e773e3),
	.w1(32'h389c32cb),
	.w2(32'h3af3aa24),
	.w3(32'h3a13c248),
	.w4(32'hbacf139b),
	.w5(32'hbb5ae796),
	.w6(32'h3b0c7fe2),
	.w7(32'h3a9810f3),
	.w8(32'hbb4bf89f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c9139),
	.w1(32'h398b4840),
	.w2(32'hbb090bd1),
	.w3(32'h3b535ea0),
	.w4(32'hb9bbf5e5),
	.w5(32'hbb50d56f),
	.w6(32'h3afcdd42),
	.w7(32'hb9df5536),
	.w8(32'hbb4fc8d4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90add4),
	.w1(32'hba3d773d),
	.w2(32'hbb0a52d3),
	.w3(32'hbb43cadd),
	.w4(32'h3b0739f6),
	.w5(32'h39acdc3e),
	.w6(32'hba0dabda),
	.w7(32'h3a788c87),
	.w8(32'h3aa00b71),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb032be9),
	.w1(32'h3b5f4a29),
	.w2(32'hb9968bac),
	.w3(32'h39ae6f02),
	.w4(32'hbb4636db),
	.w5(32'hbb65d0c3),
	.w6(32'h3ac157d4),
	.w7(32'hbb4867c4),
	.w8(32'hbbc8e71e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399de133),
	.w1(32'h39829f49),
	.w2(32'h38d593cf),
	.w3(32'h39ab771a),
	.w4(32'h38151044),
	.w5(32'hb8d7084e),
	.w6(32'h39a40c9c),
	.w7(32'h388a612c),
	.w8(32'h39830a1c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58faf3),
	.w1(32'hbb1b99fd),
	.w2(32'h3b10d9a8),
	.w3(32'h3b573607),
	.w4(32'hbb2724d6),
	.w5(32'hbb38a4ae),
	.w6(32'h3b8dce10),
	.w7(32'hb99632a5),
	.w8(32'hbb9e2559),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8784b60),
	.w1(32'hbaad1059),
	.w2(32'h3a5b9acb),
	.w3(32'h3ad38565),
	.w4(32'hbacd65b6),
	.w5(32'hba97f679),
	.w6(32'h3ae533d2),
	.w7(32'h38925ba0),
	.w8(32'hbb00e705),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd6fef),
	.w1(32'h36f107f8),
	.w2(32'h39346ac4),
	.w3(32'h393d630d),
	.w4(32'h38f82875),
	.w5(32'h3941d77c),
	.w6(32'hb906384f),
	.w7(32'h38282471),
	.w8(32'hb8dcc44e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391741f5),
	.w1(32'hba443ae7),
	.w2(32'hba45d4d1),
	.w3(32'h39012390),
	.w4(32'hba1b90de),
	.w5(32'hba2b2ab6),
	.w6(32'hba1f4f2c),
	.w7(32'hba47eb4f),
	.w8(32'hb9cb2d94),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0061f1),
	.w1(32'h3a30944d),
	.w2(32'hb8df394c),
	.w3(32'hba337e32),
	.w4(32'h3a368fed),
	.w5(32'h391ab6e1),
	.w6(32'hba98adac),
	.w7(32'hba11ff1d),
	.w8(32'h393eae1d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c30a7),
	.w1(32'hbb22dfd1),
	.w2(32'hbb0c2dd4),
	.w3(32'h39e4fd19),
	.w4(32'h3aeab85a),
	.w5(32'hb88d2518),
	.w6(32'hbac110ad),
	.w7(32'h3b026859),
	.w8(32'h3b12fe51),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf98e8a),
	.w1(32'hba7b08a1),
	.w2(32'hba8589c0),
	.w3(32'hb9b42b4c),
	.w4(32'hba668eb6),
	.w5(32'hbaddfcd5),
	.w6(32'hb9025775),
	.w7(32'h3ace0584),
	.w8(32'h391ab1ca),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d2747),
	.w1(32'h3acef73d),
	.w2(32'hb993689c),
	.w3(32'hbbe6f490),
	.w4(32'hba55a2b5),
	.w5(32'h394fadf7),
	.w6(32'hbb623b82),
	.w7(32'hba04edcc),
	.w8(32'h3a9a97ae),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7749f),
	.w1(32'hb9838c52),
	.w2(32'h39da40ba),
	.w3(32'hb61587d0),
	.w4(32'hba18f472),
	.w5(32'hba510d70),
	.w6(32'hb95c7ad2),
	.w7(32'h391a3d03),
	.w8(32'h386bb165),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c83806),
	.w1(32'hb95a35a2),
	.w2(32'h39696f2b),
	.w3(32'hb9b0e809),
	.w4(32'hb95016cc),
	.w5(32'h390863d2),
	.w6(32'hb97c293b),
	.w7(32'hb934985c),
	.w8(32'hb90f18d3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9d1b7),
	.w1(32'hbb5e0d3c),
	.w2(32'h3881e4fc),
	.w3(32'hbbe80c56),
	.w4(32'hbc1d70e6),
	.w5(32'h3b849285),
	.w6(32'hbaaa90d8),
	.w7(32'hbc074012),
	.w8(32'h3a9d936e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7ede5),
	.w1(32'h399a5d41),
	.w2(32'hb995fdfa),
	.w3(32'h3addd513),
	.w4(32'h3a112823),
	.w5(32'h38eb0088),
	.w6(32'hb91a2bb0),
	.w7(32'hb9a41aaa),
	.w8(32'h38e61fbc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b4ccb),
	.w1(32'h3ae9987c),
	.w2(32'hbb0ab923),
	.w3(32'hbbacc3b9),
	.w4(32'hbb889a39),
	.w5(32'hbb58ee16),
	.w6(32'hbae153f5),
	.w7(32'hba28d8b6),
	.w8(32'h3a812afe),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df52fa),
	.w1(32'hb9e94450),
	.w2(32'hb9d3d970),
	.w3(32'hba5329dc),
	.w4(32'hb9e6d646),
	.w5(32'hb9884c90),
	.w6(32'hb9fc5ab7),
	.w7(32'hb9edaa2e),
	.w8(32'hb9526b1e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909efc4),
	.w1(32'hb9e75679),
	.w2(32'hb9195bb8),
	.w3(32'hb970a2e9),
	.w4(32'hb9f42615),
	.w5(32'hb955de47),
	.w6(32'hb9fb349d),
	.w7(32'hb9c1c81f),
	.w8(32'hb985998a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2bd8a),
	.w1(32'h3900b432),
	.w2(32'hb9c4c525),
	.w3(32'h3a96761b),
	.w4(32'h37563eab),
	.w5(32'hbab59954),
	.w6(32'h3a5d1ecc),
	.w7(32'h3a4e26e0),
	.w8(32'hba90d2f4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6b58),
	.w1(32'hba2c343f),
	.w2(32'hb884ee5f),
	.w3(32'hbb13d2b8),
	.w4(32'hb97cdeac),
	.w5(32'h38b4bd42),
	.w6(32'hbac10bbb),
	.w7(32'h39a31975),
	.w8(32'h399c4e8d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39862bed),
	.w1(32'h397c3a9e),
	.w2(32'h3a10851f),
	.w3(32'h3a04ef24),
	.w4(32'h3995c07d),
	.w5(32'h3a19ccd8),
	.w6(32'h3a779c3c),
	.w7(32'hb7ce7b49),
	.w8(32'h3a344274),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d1bf6),
	.w1(32'hb9e2e91d),
	.w2(32'h3a7c85ad),
	.w3(32'h3aa7ba7e),
	.w4(32'h3a004a96),
	.w5(32'hba54a75e),
	.w6(32'h38a75342),
	.w7(32'h3ad9f577),
	.w8(32'h397eda88),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5df23),
	.w1(32'hbc2bca3e),
	.w2(32'h3b473e3d),
	.w3(32'h3a803e55),
	.w4(32'h3bb7592f),
	.w5(32'h3c2973e2),
	.w6(32'h3b830b07),
	.w7(32'h3c169552),
	.w8(32'h3c5b4835),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1aa48),
	.w1(32'h39ae228c),
	.w2(32'hb9a6484c),
	.w3(32'hbc0c7ef0),
	.w4(32'h3b015f94),
	.w5(32'h3bace978),
	.w6(32'hbbc90cf7),
	.w7(32'hba4562ef),
	.w8(32'h3b76a2f8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ab78e),
	.w1(32'h38aec06b),
	.w2(32'hb523e820),
	.w3(32'hba99cb5a),
	.w4(32'hbb21d60b),
	.w5(32'h3a6bd3d9),
	.w6(32'hba439c27),
	.w7(32'hbb36f9c9),
	.w8(32'h3902d040),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98b478),
	.w1(32'h3936c436),
	.w2(32'h38b09500),
	.w3(32'hbb077711),
	.w4(32'h38ffc1e2),
	.w5(32'h3a0d43d9),
	.w6(32'hba7eb8d0),
	.w7(32'hb7d044a9),
	.w8(32'h3a0204af),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9240cad),
	.w1(32'h3849c1d4),
	.w2(32'hb9a32df7),
	.w3(32'hb8274c1c),
	.w4(32'hb51217df),
	.w5(32'hb9ed9c8a),
	.w6(32'h3922a0fb),
	.w7(32'hb95b75e1),
	.w8(32'h3934aa2d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b90064),
	.w1(32'hba390e94),
	.w2(32'hb9f2b288),
	.w3(32'hba336ba2),
	.w4(32'hb98300a0),
	.w5(32'h38d7cd64),
	.w6(32'h383c2eb3),
	.w7(32'hb99d8e13),
	.w8(32'h3902bff8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f8cbf),
	.w1(32'h39bcbba1),
	.w2(32'h3a97ed33),
	.w3(32'hb9b1c809),
	.w4(32'h39d4a738),
	.w5(32'h399a284f),
	.w6(32'hb9e0aaf1),
	.w7(32'h3914464c),
	.w8(32'hb977a655),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0cb25),
	.w1(32'hb9f66da3),
	.w2(32'h39c8ca83),
	.w3(32'hbb38540a),
	.w4(32'hbb582c5a),
	.w5(32'hb9923e32),
	.w6(32'h3b7cb669),
	.w7(32'h39f4f6b2),
	.w8(32'hba3a0307),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65926f),
	.w1(32'hb9db3b0e),
	.w2(32'hb8c6b998),
	.w3(32'hbb52313d),
	.w4(32'hb9f6de70),
	.w5(32'h3a6dca72),
	.w6(32'hba93f9fb),
	.w7(32'h3ab83081),
	.w8(32'h3b3bf54e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64b755),
	.w1(32'hbad21050),
	.w2(32'hba2e063c),
	.w3(32'hbb57576a),
	.w4(32'hb88908ca),
	.w5(32'hba212124),
	.w6(32'hbac21b4f),
	.w7(32'h3b3386f4),
	.w8(32'h3b827b8f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe4e8),
	.w1(32'hbb07a824),
	.w2(32'h3a9264eb),
	.w3(32'hbb2bda56),
	.w4(32'hbad4626b),
	.w5(32'h3a702fd2),
	.w6(32'hb836c698),
	.w7(32'hb966a367),
	.w8(32'h38fdff99),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c0f2),
	.w1(32'h3a7cdd4d),
	.w2(32'h3b910f9b),
	.w3(32'h3bd8c577),
	.w4(32'h3961fe5b),
	.w5(32'hbade0426),
	.w6(32'h3ba2afd3),
	.w7(32'h3b388e58),
	.w8(32'hbb58bc3c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2dda2b),
	.w1(32'hba4345a2),
	.w2(32'hb95ed3df),
	.w3(32'hba05cb69),
	.w4(32'hba2e8ec2),
	.w5(32'hb9b44769),
	.w6(32'hba2211e3),
	.w7(32'hb9e44639),
	.w8(32'hba1663a3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf998ca),
	.w1(32'hbae59e1d),
	.w2(32'hbaae8c39),
	.w3(32'hba6674bb),
	.w4(32'hbae456d0),
	.w5(32'hbaf5c024),
	.w6(32'hba781907),
	.w7(32'hba43ffe5),
	.w8(32'hba9b5c21),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cc299),
	.w1(32'h3946d97d),
	.w2(32'hb965c8c9),
	.w3(32'hba264bba),
	.w4(32'h39a5fc66),
	.w5(32'hb9768253),
	.w6(32'h3a480cc8),
	.w7(32'h3a2378f9),
	.w8(32'h396c386c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd1a09),
	.w1(32'hbb01cc0f),
	.w2(32'hba6e1ec3),
	.w3(32'hba833e66),
	.w4(32'hba817c97),
	.w5(32'hb73d6768),
	.w6(32'hbab5b2c2),
	.w7(32'hba8e6357),
	.w8(32'h3a2de1b6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f503d),
	.w1(32'hba3e3dc1),
	.w2(32'hbaafcc26),
	.w3(32'h39f98e73),
	.w4(32'hba4fff57),
	.w5(32'hbab31eb6),
	.w6(32'h38de0063),
	.w7(32'hba03f811),
	.w8(32'hba3359f4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb453245),
	.w1(32'hbb646fa2),
	.w2(32'h3ae5166e),
	.w3(32'h3acc1d38),
	.w4(32'hbb47ad68),
	.w5(32'hba8c9295),
	.w6(32'h3bb2c7fa),
	.w7(32'hb86b2595),
	.w8(32'hbb121e48),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade6d83),
	.w1(32'hbaf00510),
	.w2(32'hb9824696),
	.w3(32'hbab9d903),
	.w4(32'hbacd0d6a),
	.w5(32'hba2feb8a),
	.w6(32'hba29d130),
	.w7(32'hb990d175),
	.w8(32'hba010d48),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba509bb6),
	.w1(32'hb91fb784),
	.w2(32'hba3d34b9),
	.w3(32'hba76f781),
	.w4(32'h38b3748f),
	.w5(32'hb9a8787b),
	.w6(32'hb9eb7952),
	.w7(32'hb9d35b7b),
	.w8(32'hb9892b64),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d27f00),
	.w1(32'hb9b47237),
	.w2(32'hb96eb183),
	.w3(32'hb904068e),
	.w4(32'hba06a069),
	.w5(32'hb9bd31a6),
	.w6(32'hba00c796),
	.w7(32'hb985bee1),
	.w8(32'hb8f58ebe),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b71a50),
	.w1(32'hba30da93),
	.w2(32'hba2734fb),
	.w3(32'hb8442f86),
	.w4(32'hba6132a5),
	.w5(32'hba60137a),
	.w6(32'h38f998aa),
	.w7(32'hba25b4fd),
	.w8(32'h39f17265),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a242cd6),
	.w1(32'h3a92e32f),
	.w2(32'h3a498583),
	.w3(32'h396318f0),
	.w4(32'h3a8e464f),
	.w5(32'h3a874071),
	.w6(32'h3a155f5c),
	.w7(32'h3a18ac8b),
	.w8(32'h3a84dffb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972e15e),
	.w1(32'hba24ddf5),
	.w2(32'h3a026caa),
	.w3(32'hb90e49e3),
	.w4(32'hba8c5869),
	.w5(32'h398d471c),
	.w6(32'hba7d775e),
	.w7(32'hba56870f),
	.w8(32'hb8eabfb0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39571940),
	.w1(32'hb9d2542c),
	.w2(32'hba525284),
	.w3(32'h3aa1467e),
	.w4(32'hbabff27c),
	.w5(32'hbad9790a),
	.w6(32'h3afed8f3),
	.w7(32'hba2c4cea),
	.w8(32'hbb32b5fa),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2cb63),
	.w1(32'hbb992a47),
	.w2(32'hba99bf1d),
	.w3(32'hbacf2309),
	.w4(32'hbc115552),
	.w5(32'hb8f7c041),
	.w6(32'hbb07458a),
	.w7(32'hbbd3323a),
	.w8(32'hbb027714),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba723d4d),
	.w1(32'hb94c7f0d),
	.w2(32'hba301e9f),
	.w3(32'hba4afa97),
	.w4(32'hb929b8c7),
	.w5(32'h3884965f),
	.w6(32'hb9fe331a),
	.w7(32'hba51d982),
	.w8(32'hba3486e7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab00316),
	.w1(32'h3abe2c0f),
	.w2(32'h3a5552c0),
	.w3(32'hbaab21fc),
	.w4(32'h3adfd097),
	.w5(32'h3a8af377),
	.w6(32'h3aec552c),
	.w7(32'h3ab16028),
	.w8(32'h3ad0c096),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a758117),
	.w1(32'hb947484c),
	.w2(32'hb9ae8bc5),
	.w3(32'h3a8c90ed),
	.w4(32'hb90e6d73),
	.w5(32'hb980a996),
	.w6(32'hb9b39f44),
	.w7(32'hb9d5b3a6),
	.w8(32'hb9ddc68f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3cc71),
	.w1(32'hba1901a6),
	.w2(32'h39303391),
	.w3(32'h38390214),
	.w4(32'hb9ff04d2),
	.w5(32'hb9f381ad),
	.w6(32'hb9dcfcf8),
	.w7(32'hb9e93ff1),
	.w8(32'h39ca7eba),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891a64),
	.w1(32'hbbe85a64),
	.w2(32'h3a31b25f),
	.w3(32'h3b6ec721),
	.w4(32'hbbe7013f),
	.w5(32'h39d78816),
	.w6(32'h3bbbed4d),
	.w7(32'hbbf69620),
	.w8(32'hbbf1abb3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc74b37),
	.w1(32'hba8f82de),
	.w2(32'hbb812d65),
	.w3(32'h3ba5e98e),
	.w4(32'hba53bf7b),
	.w5(32'hbbcdf8b9),
	.w6(32'h3996de55),
	.w7(32'h3b81fe97),
	.w8(32'h3b254915),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b9d33),
	.w1(32'hbb585901),
	.w2(32'hbb6432e0),
	.w3(32'hb9a4cde3),
	.w4(32'hbb3ed85d),
	.w5(32'hbb443889),
	.w6(32'hba2ecaaf),
	.w7(32'hbac3c347),
	.w8(32'hba715bcb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7c73e),
	.w1(32'h3976895a),
	.w2(32'h3ae07181),
	.w3(32'hbc2f8d24),
	.w4(32'hba22e2d2),
	.w5(32'h3b608ef4),
	.w6(32'hbbd51509),
	.w7(32'hbad0bd23),
	.w8(32'h3ba82d8c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcc9e7),
	.w1(32'h3a1bcf1e),
	.w2(32'h395f8e56),
	.w3(32'h3ab41dcf),
	.w4(32'h3a3dfbc2),
	.w5(32'h39e54b5f),
	.w6(32'h3a09b792),
	.w7(32'h39d85cf3),
	.w8(32'h3a21bb28),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd710d),
	.w1(32'hba204170),
	.w2(32'hb9a47056),
	.w3(32'h3a01c553),
	.w4(32'hba085d5c),
	.w5(32'hb94d19b2),
	.w6(32'hba236176),
	.w7(32'hba18d472),
	.w8(32'hb9a16e03),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab3665),
	.w1(32'hba049e11),
	.w2(32'hb9a09e42),
	.w3(32'hb994600a),
	.w4(32'hba06b93d),
	.w5(32'hb9941368),
	.w6(32'hba0f40f8),
	.w7(32'hb9edc861),
	.w8(32'hb9a1a8ad),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb833f1e1),
	.w1(32'hba799452),
	.w2(32'h39f3eb09),
	.w3(32'h3a0d88f5),
	.w4(32'hba9d1ad7),
	.w5(32'hba142537),
	.w6(32'h3a1d8d5d),
	.w7(32'hba750e08),
	.w8(32'hbac6d6f2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6ded2),
	.w1(32'hb980644c),
	.w2(32'hb9650f48),
	.w3(32'hb967ab94),
	.w4(32'h397ade3e),
	.w5(32'h3924e0fb),
	.w6(32'h3997819c),
	.w7(32'hb856228f),
	.w8(32'h39836c68),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5da399),
	.w1(32'hbadf4645),
	.w2(32'h3add419f),
	.w3(32'h3b248fbb),
	.w4(32'h39504608),
	.w5(32'h3a88b7a1),
	.w6(32'h3b3575fd),
	.w7(32'h3a98870d),
	.w8(32'h38fb0898),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0f6d),
	.w1(32'hbb4341f2),
	.w2(32'hbb8b8d94),
	.w3(32'h3bb4a5ff),
	.w4(32'hba066ccc),
	.w5(32'hbbc145bd),
	.w6(32'h3b8d1cf6),
	.w7(32'h3b0a862f),
	.w8(32'hbb976bd8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f749d),
	.w1(32'h3abdd482),
	.w2(32'h3a219175),
	.w3(32'hbb79af0a),
	.w4(32'h3a4348a8),
	.w5(32'h3a663ec2),
	.w6(32'hba3c1f40),
	.w7(32'h3a051e27),
	.w8(32'h3a84e68d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ec3387),
	.w1(32'hbb0c535b),
	.w2(32'hba9954f4),
	.w3(32'h3ad573da),
	.w4(32'hbaf55e8c),
	.w5(32'hbb2e43d1),
	.w6(32'h3b23bb6e),
	.w7(32'hb9c82ab6),
	.w8(32'hbb326b17),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2efa7),
	.w1(32'hbb28ec11),
	.w2(32'h3ad8705a),
	.w3(32'h3ace3308),
	.w4(32'hba8f6140),
	.w5(32'hb9cd82b6),
	.w6(32'h3b0d4df7),
	.w7(32'hbac1ffe7),
	.w8(32'hbb1e61f9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaefe5),
	.w1(32'h394de9d2),
	.w2(32'hba2cf856),
	.w3(32'hbad53e75),
	.w4(32'hb9ec2742),
	.w5(32'hb92f8d44),
	.w6(32'hb9bbd516),
	.w7(32'hb9123cc7),
	.w8(32'h396804da),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92c9c8),
	.w1(32'hb9253cff),
	.w2(32'h3a85c72f),
	.w3(32'h3a7efff3),
	.w4(32'hb9d36eba),
	.w5(32'hba1be68a),
	.w6(32'h3a4ce446),
	.w7(32'h39125351),
	.w8(32'hbad667ab),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d635ad),
	.w1(32'hb897c955),
	.w2(32'hb9b5691f),
	.w3(32'hba1ed438),
	.w4(32'h39469fe0),
	.w5(32'h37817f20),
	.w6(32'h3896d4c3),
	.w7(32'hb89cb96b),
	.w8(32'h37f0199d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985e0a9),
	.w1(32'h3894dc9a),
	.w2(32'hb987128c),
	.w3(32'hb84abb04),
	.w4(32'h39366b80),
	.w5(32'hb8aab229),
	.w6(32'hb86c5771),
	.w7(32'hb97a3e74),
	.w8(32'hb9b3d82e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98aa34c),
	.w1(32'h39d30806),
	.w2(32'hb7818789),
	.w3(32'hb92309a0),
	.w4(32'h3989fe87),
	.w5(32'h393fe1c1),
	.w6(32'h388fd7bd),
	.w7(32'hb88f9c11),
	.w8(32'h38f6de6a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee2b5f),
	.w1(32'h38a419b7),
	.w2(32'h39eb5442),
	.w3(32'h39187485),
	.w4(32'h39db251c),
	.w5(32'h3a07212d),
	.w6(32'h39618fb0),
	.w7(32'h3a341630),
	.w8(32'h3a472cae),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb837e16),
	.w1(32'hbab7f4c5),
	.w2(32'h39878201),
	.w3(32'hbb8f4dd4),
	.w4(32'hb992d89d),
	.w5(32'h3abf1300),
	.w6(32'hbb3d4e99),
	.w7(32'hb91ecf77),
	.w8(32'h3ac720e0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8f038),
	.w1(32'h390fe21c),
	.w2(32'h39eca544),
	.w3(32'hb839522a),
	.w4(32'h39582309),
	.w5(32'h3a0ffbbb),
	.w6(32'hb9de5b47),
	.w7(32'hb8c90cb0),
	.w8(32'h39a3a055),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e5bc1),
	.w1(32'hbafada10),
	.w2(32'hbaa98009),
	.w3(32'hbb545c46),
	.w4(32'hba853b0b),
	.w5(32'hbae744b4),
	.w6(32'hbac3f18b),
	.w7(32'h3a87586d),
	.w8(32'h3a6d5671),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ca8a4),
	.w1(32'hba721474),
	.w2(32'h3a17fd07),
	.w3(32'h3aec1e39),
	.w4(32'hba1830da),
	.w5(32'hba638987),
	.w6(32'h3ac0a7e1),
	.w7(32'h3a120070),
	.w8(32'hba35bd8f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299568),
	.w1(32'hb8820584),
	.w2(32'h3aafe57f),
	.w3(32'hbb8ab5a2),
	.w4(32'hb97bff5a),
	.w5(32'h3b48cf5c),
	.w6(32'hbb1041e7),
	.w7(32'hb9e8ab72),
	.w8(32'h3b24fd39),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb91f2b),
	.w1(32'hbad06796),
	.w2(32'h38990ef3),
	.w3(32'h3b1b9d11),
	.w4(32'h3a4fabde),
	.w5(32'h39eb76c0),
	.w6(32'h3b5485a5),
	.w7(32'h3a86dcfa),
	.w8(32'hbb5f7ff6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985065c),
	.w1(32'hb929eb32),
	.w2(32'h3b1eeb46),
	.w3(32'hba8f3d7a),
	.w4(32'h3a84a899),
	.w5(32'h3b0a6544),
	.w6(32'hbabbe4bd),
	.w7(32'hb9581bac),
	.w8(32'h3b665082),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1751a1),
	.w1(32'hbb93e247),
	.w2(32'hbb3c69be),
	.w3(32'h3b79887c),
	.w4(32'hbbaf9654),
	.w5(32'hbba3639b),
	.w6(32'h3b76e77f),
	.w7(32'hbb74737e),
	.w8(32'hbbd93b3f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f3512),
	.w1(32'hb8b1db10),
	.w2(32'hba41bb0d),
	.w3(32'hbac75728),
	.w4(32'h39a7a055),
	.w5(32'hb8a06328),
	.w6(32'h3a7c8ecd),
	.w7(32'h3913a313),
	.w8(32'hbaf5f998),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88cb9d),
	.w1(32'h38e27ecc),
	.w2(32'hb9bcf44c),
	.w3(32'hbba7f15d),
	.w4(32'hb849917f),
	.w5(32'h3aa9ff00),
	.w6(32'hbaeef96a),
	.w7(32'hba34617e),
	.w8(32'h3abcb371),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45f9b3),
	.w1(32'hb8604c9a),
	.w2(32'hba288879),
	.w3(32'hb960817f),
	.w4(32'h397b7e4c),
	.w5(32'hba103383),
	.w6(32'h39f528fc),
	.w7(32'h38862e44),
	.w8(32'hb9997c27),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6292b),
	.w1(32'hbb3da43d),
	.w2(32'hbb28bc41),
	.w3(32'h3ae215f9),
	.w4(32'hbafe9ca5),
	.w5(32'hbb7290b9),
	.w6(32'h3b23840d),
	.w7(32'h39e283ca),
	.w8(32'hbb1c8467),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf25e4e),
	.w1(32'hbbb9641e),
	.w2(32'h3b8f7810),
	.w3(32'hba763d51),
	.w4(32'hbb23a3d7),
	.w5(32'h3b8a899e),
	.w6(32'h3b1c177b),
	.w7(32'hba7ec636),
	.w8(32'h3940208c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad09552),
	.w1(32'hbb05329b),
	.w2(32'h3a00b655),
	.w3(32'hb8e2b616),
	.w4(32'h3b1b664a),
	.w5(32'h3c0ba797),
	.w6(32'h3a365f2c),
	.w7(32'h3b4aaadb),
	.w8(32'h3c1e4197),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ed507),
	.w1(32'hbb7546e7),
	.w2(32'h39dd0ee7),
	.w3(32'hbc314c19),
	.w4(32'hbb334001),
	.w5(32'h3a5411f3),
	.w6(32'hbbcc2513),
	.w7(32'h3a3081c8),
	.w8(32'h3b3625a6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5165d6),
	.w1(32'h38a1ae7b),
	.w2(32'h3a25a3f6),
	.w3(32'hbb81e8f0),
	.w4(32'h39a313cb),
	.w5(32'hba93e1f0),
	.w6(32'hbaee0106),
	.w7(32'h3a9b539c),
	.w8(32'h3afac97e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b3899),
	.w1(32'hbbe80a15),
	.w2(32'h3b26fe89),
	.w3(32'h3ae90c9f),
	.w4(32'h3b0b55c3),
	.w5(32'h3b2aa0ad),
	.w6(32'h3a294147),
	.w7(32'h3b85b0a4),
	.w8(32'hb97971ab),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf69506),
	.w1(32'hbab196bb),
	.w2(32'hba85ab01),
	.w3(32'hba75f9c3),
	.w4(32'hba135005),
	.w5(32'h391a216e),
	.w6(32'hb95da26f),
	.w7(32'h39f075df),
	.w8(32'h3a03b331),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc246a12),
	.w1(32'hbc1ecbe6),
	.w2(32'hbb3eaab0),
	.w3(32'hbb9c760a),
	.w4(32'hb9afcabc),
	.w5(32'h3b9672e5),
	.w6(32'h3aa2fe1b),
	.w7(32'h3b74c7ef),
	.w8(32'h3bb661b2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b138e),
	.w1(32'hbb9e1786),
	.w2(32'hba6c8839),
	.w3(32'hba2591f9),
	.w4(32'hbac51f17),
	.w5(32'h39dd2aa2),
	.w6(32'hb9c95a7d),
	.w7(32'h39b08629),
	.w8(32'h3b150020),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926e252),
	.w1(32'hba2ddac9),
	.w2(32'hba7b588c),
	.w3(32'hb99557be),
	.w4(32'hb9feb742),
	.w5(32'hb9db8bb1),
	.w6(32'hb9d8bdb8),
	.w7(32'hba65d4d8),
	.w8(32'hba4f0237),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1024f0),
	.w1(32'h3a20b9db),
	.w2(32'hba88bedb),
	.w3(32'hba2a15f9),
	.w4(32'hb963d70d),
	.w5(32'hb9ce35b6),
	.w6(32'hba8691b1),
	.w7(32'hba5ea7f6),
	.w8(32'hba2d29f0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bedcc),
	.w1(32'hb92db479),
	.w2(32'hb95bd5b1),
	.w3(32'h3b164768),
	.w4(32'hb9181577),
	.w5(32'hbb16d07e),
	.w6(32'h3b385b45),
	.w7(32'h3ab3c969),
	.w8(32'hbb0076b0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5929ed),
	.w1(32'hba470d12),
	.w2(32'hbb01321c),
	.w3(32'hbb5faf3b),
	.w4(32'hba2f182f),
	.w5(32'hbadd5df7),
	.w6(32'hba96eb18),
	.w7(32'h392d088c),
	.w8(32'h38820ecb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4ae14),
	.w1(32'hbb4dd2e5),
	.w2(32'hbb24f2d6),
	.w3(32'hbbcc52a0),
	.w4(32'hbb796e41),
	.w5(32'h39d5814b),
	.w6(32'hbb2ef63d),
	.w7(32'hbb0d4065),
	.w8(32'h3ac3f45c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba402ff),
	.w1(32'hbb0b6c33),
	.w2(32'hba40e40e),
	.w3(32'hbb9ca5bf),
	.w4(32'hba860cdc),
	.w5(32'h3a547e42),
	.w6(32'hbb324f3e),
	.w7(32'hbaa6f682),
	.w8(32'h39c109ef),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadec120),
	.w1(32'h3abf247f),
	.w2(32'h3a998c20),
	.w3(32'hbb9e22b9),
	.w4(32'hb837361a),
	.w5(32'h3a9e6a8a),
	.w6(32'hbb3c499c),
	.w7(32'h3aa0b12c),
	.w8(32'h3a7f3bfd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac02058),
	.w1(32'h3b39798c),
	.w2(32'hba98e621),
	.w3(32'h3a54c3ab),
	.w4(32'hbad3eeae),
	.w5(32'hbaff8b2b),
	.w6(32'h39cf625a),
	.w7(32'hbb164830),
	.w8(32'hbb9571da),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcbbab),
	.w1(32'hb969e0f3),
	.w2(32'h38582e47),
	.w3(32'hba7bb17a),
	.w4(32'hba3dfa76),
	.w5(32'hba43e4d1),
	.w6(32'h37e4d900),
	.w7(32'h3a7a3b40),
	.w8(32'h3a280658),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba643efa),
	.w1(32'hbaa8c9cd),
	.w2(32'hba981b2c),
	.w3(32'hba4ee040),
	.w4(32'hba983fca),
	.w5(32'hba778ab0),
	.w6(32'hba6caaee),
	.w7(32'hba765e6c),
	.w8(32'hba231358),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cdaec),
	.w1(32'hba80d22d),
	.w2(32'hba7b2973),
	.w3(32'hba610f43),
	.w4(32'hba67f743),
	.w5(32'hba26f2cc),
	.w6(32'hba43f371),
	.w7(32'hba465874),
	.w8(32'hba238b9f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba002329),
	.w1(32'hba526e4d),
	.w2(32'hba24077c),
	.w3(32'hb9ff53c9),
	.w4(32'hba3af60d),
	.w5(32'hb9fcaf78),
	.w6(32'hba13223b),
	.w7(32'hba313965),
	.w8(32'hb9ec4abf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391edc0a),
	.w1(32'hba4fcd21),
	.w2(32'hb96a5f6a),
	.w3(32'h3844fa41),
	.w4(32'h39b92f7a),
	.w5(32'hb78a1250),
	.w6(32'hb9ee0f01),
	.w7(32'hba3e4d98),
	.w8(32'hba21c882),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07a1a5),
	.w1(32'hb9b813fc),
	.w2(32'hba85f109),
	.w3(32'hbadec670),
	.w4(32'hba2ff486),
	.w5(32'hba9ef8e9),
	.w6(32'hb90a437c),
	.w7(32'h3a90f468),
	.w8(32'h3a8828b9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804d26),
	.w1(32'hba1f8757),
	.w2(32'h39d70b4c),
	.w3(32'hb987f835),
	.w4(32'hb8a4ef5a),
	.w5(32'h3a7af75a),
	.w6(32'hb927cad1),
	.w7(32'hb96c8858),
	.w8(32'hb8e1b5cd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39988176),
	.w1(32'hb9c4c3f6),
	.w2(32'h3b3247ed),
	.w3(32'h3aea6eb2),
	.w4(32'h383dc048),
	.w5(32'h3a9bd8d4),
	.w6(32'h3aafca98),
	.w7(32'h39d1695b),
	.w8(32'h37b725bc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2243d8),
	.w1(32'hba394714),
	.w2(32'hbaa75900),
	.w3(32'hbb8c9423),
	.w4(32'hbac58cec),
	.w5(32'h3a3c9ef3),
	.w6(32'hbb43f234),
	.w7(32'hbad36d74),
	.w8(32'h3915d852),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e3d8a),
	.w1(32'hba2ee14c),
	.w2(32'hb9fed65f),
	.w3(32'hba2cead4),
	.w4(32'h395f5e27),
	.w5(32'hb9bf709c),
	.w6(32'hba1e6447),
	.w7(32'hba179607),
	.w8(32'h393e9294),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0f4af),
	.w1(32'hb7b22e35),
	.w2(32'hb85112d5),
	.w3(32'hba57ade9),
	.w4(32'hb8509214),
	.w5(32'hb9c90ec0),
	.w6(32'hb716ed4d),
	.w7(32'hb92881cf),
	.w8(32'hb9ad9514),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03b2e7),
	.w1(32'hba03e2a9),
	.w2(32'hb997fff3),
	.w3(32'hba3e1474),
	.w4(32'hb9baab75),
	.w5(32'hb900030e),
	.w6(32'hba0b6e57),
	.w7(32'hb9e94c4c),
	.w8(32'hb93c7edf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9650b5b),
	.w1(32'h39967066),
	.w2(32'hb913019a),
	.w3(32'h38819237),
	.w4(32'h39ca6ada),
	.w5(32'h389e7f54),
	.w6(32'h39cb0e85),
	.w7(32'h3a09e4ce),
	.w8(32'h39e73644),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ea0ea),
	.w1(32'h3b3ff18a),
	.w2(32'hba857be9),
	.w3(32'h3bbeddb9),
	.w4(32'h3809fce8),
	.w5(32'hbbb0e98c),
	.w6(32'hba506f82),
	.w7(32'h3b8ec866),
	.w8(32'hb9d889f2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8602332),
	.w1(32'hb7ac039d),
	.w2(32'h3a4b1f48),
	.w3(32'h3ac79f87),
	.w4(32'hbb438819),
	.w5(32'hbb3ae920),
	.w6(32'h3b17869f),
	.w7(32'hbb01657d),
	.w8(32'hbb498394),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d93fd),
	.w1(32'hb92bf9a4),
	.w2(32'h392a9887),
	.w3(32'h3a300808),
	.w4(32'h39153808),
	.w5(32'h38ff68aa),
	.w6(32'h39df5294),
	.w7(32'h39b3ea11),
	.w8(32'hb9a68eee),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90451ca),
	.w1(32'hbab16dd0),
	.w2(32'hba29f114),
	.w3(32'h3a11c91c),
	.w4(32'h39497cbd),
	.w5(32'hbafefcf1),
	.w6(32'h39274e52),
	.w7(32'h3a8cef87),
	.w8(32'hb9db48ba),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f0a23),
	.w1(32'h392742cb),
	.w2(32'h38b174bf),
	.w3(32'hba941f03),
	.w4(32'hbaa58c7d),
	.w5(32'hb767ae9b),
	.w6(32'hb8951a7e),
	.w7(32'h38b2d57c),
	.w8(32'h3aad034c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d11078),
	.w1(32'hbaeccad1),
	.w2(32'h39086bab),
	.w3(32'h3a8f261c),
	.w4(32'hbacebecd),
	.w5(32'hbb1a5073),
	.w6(32'h3ad13e88),
	.w7(32'hba3b40a1),
	.w8(32'hbabf3fb9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a1c94),
	.w1(32'h395e8cb4),
	.w2(32'hba99ed5c),
	.w3(32'hb9bbf96e),
	.w4(32'hb9598528),
	.w5(32'h3ad03e1f),
	.w6(32'h3b17e978),
	.w7(32'hb96319b1),
	.w8(32'h36be1472),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9628fae),
	.w1(32'hbabcdca2),
	.w2(32'h3b925b9b),
	.w3(32'h3b43e1b3),
	.w4(32'hba57a7f0),
	.w5(32'h3aaf8a10),
	.w6(32'h3ad18110),
	.w7(32'hb959618c),
	.w8(32'hbb76fdee),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb531202),
	.w1(32'h39703305),
	.w2(32'h3998507d),
	.w3(32'hbb99616d),
	.w4(32'hb8a9a89a),
	.w5(32'h38654acd),
	.w6(32'hbad943bd),
	.w7(32'h3992ed54),
	.w8(32'h3a009e94),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c9085),
	.w1(32'h3aa246a8),
	.w2(32'h39800eae),
	.w3(32'hb9a2459b),
	.w4(32'h3a4ad44d),
	.w5(32'h39587774),
	.w6(32'hb9494f0c),
	.w7(32'h3a864079),
	.w8(32'hb8b2182e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f79fc),
	.w1(32'hba96a63c),
	.w2(32'h3ab02d5b),
	.w3(32'h3a19e4ec),
	.w4(32'h3a1e22db),
	.w5(32'h3b02fe73),
	.w6(32'h3aa66980),
	.w7(32'h3b273391),
	.w8(32'hba6da094),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0e0a2),
	.w1(32'hb9f1f421),
	.w2(32'hbaa43e70),
	.w3(32'hbb07cca0),
	.w4(32'h38cf6fd9),
	.w5(32'h38887deb),
	.w6(32'hbb227637),
	.w7(32'hb9f32121),
	.w8(32'h3acd02ea),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33499d),
	.w1(32'h38b5ae68),
	.w2(32'h3972a72b),
	.w3(32'h3a9d29a1),
	.w4(32'h39c74f7f),
	.w5(32'hbb0d251a),
	.w6(32'h3b3742cb),
	.w7(32'h3aa4c993),
	.w8(32'hbb11b9ef),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1914b0),
	.w1(32'hb87759f3),
	.w2(32'hb94ee6ba),
	.w3(32'h398c9ddd),
	.w4(32'hb90e4346),
	.w5(32'hb98b287d),
	.w6(32'h39a0928b),
	.w7(32'h3a28f46a),
	.w8(32'h3986c06b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4461),
	.w1(32'hb9198256),
	.w2(32'h3ab10628),
	.w3(32'hbba34748),
	.w4(32'hbb6dfe85),
	.w5(32'h39e4c2db),
	.w6(32'hbae99fe1),
	.w7(32'hbaf80aeb),
	.w8(32'h3aca49ba),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb199605),
	.w1(32'hbafefbc0),
	.w2(32'hbabbcfd7),
	.w3(32'hbb15d155),
	.w4(32'hbad2d866),
	.w5(32'hba69eb1a),
	.w6(32'hbab03655),
	.w7(32'h3a85c3ef),
	.w8(32'h39712225),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47a55e),
	.w1(32'h39737014),
	.w2(32'h39e8db6c),
	.w3(32'hba49c3f4),
	.w4(32'h38d2ca36),
	.w5(32'hb8f1b952),
	.w6(32'h3950afc4),
	.w7(32'h39920e25),
	.w8(32'h3813cc69),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8001df1),
	.w1(32'hb9f7b550),
	.w2(32'hba3ff8cf),
	.w3(32'hb8d295f6),
	.w4(32'h39752c83),
	.w5(32'hb81d3e5d),
	.w6(32'h39a50f4d),
	.w7(32'hb99bb53c),
	.w8(32'h399456a4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad08a85),
	.w1(32'hbb01d787),
	.w2(32'hba4b9b2f),
	.w3(32'h3a098791),
	.w4(32'hbaad3827),
	.w5(32'hb9871468),
	.w6(32'hb7b2d048),
	.w7(32'hba1344bd),
	.w8(32'hba914510),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbde87),
	.w1(32'hbae787c2),
	.w2(32'hb9f5ac3f),
	.w3(32'hbc01117a),
	.w4(32'hbaa9ea04),
	.w5(32'h3a808049),
	.w6(32'hbbb0d320),
	.w7(32'hbad87ed8),
	.w8(32'h3aa1e274),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efc96a),
	.w1(32'hb9d26914),
	.w2(32'h3aac659d),
	.w3(32'h3a46e823),
	.w4(32'hb9a746e6),
	.w5(32'hbab19050),
	.w6(32'h3b418529),
	.w7(32'h3acd8546),
	.w8(32'hb92eee0b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916a6c1),
	.w1(32'hb96c39eb),
	.w2(32'h38dc3245),
	.w3(32'hb955e548),
	.w4(32'hb995ec37),
	.w5(32'hb9a0768d),
	.w6(32'hb86324da),
	.w7(32'hb91ec0ec),
	.w8(32'hb84dade3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf9e3f),
	.w1(32'hbafd2260),
	.w2(32'h3abd8b7f),
	.w3(32'h3a82e6eb),
	.w4(32'hbb21ee0b),
	.w5(32'hbb250db7),
	.w6(32'h3b16efe2),
	.w7(32'hba875313),
	.w8(32'hbb65b712),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ae705),
	.w1(32'h3a7d6f52),
	.w2(32'h3ab655e1),
	.w3(32'h39f163df),
	.w4(32'h3a938df1),
	.w5(32'hb983842d),
	.w6(32'h3a52e66c),
	.w7(32'h3ab0ffc7),
	.w8(32'hb98e02e8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf4029),
	.w1(32'hba566fde),
	.w2(32'h3b062c1d),
	.w3(32'h3ba2a2fe),
	.w4(32'h3b1891c6),
	.w5(32'h39d7d290),
	.w6(32'h3b5c0b71),
	.w7(32'h3b2f9e9d),
	.w8(32'hbaa1c07f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf430d2),
	.w1(32'hbb8bd99d),
	.w2(32'hbb0c766a),
	.w3(32'hbc05cb61),
	.w4(32'hbb9a5aea),
	.w5(32'h3b68fa76),
	.w6(32'hbba50efd),
	.w7(32'hbb1c0e19),
	.w8(32'h3ae33a01),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8f69c),
	.w1(32'h38d00e10),
	.w2(32'hba5cd02b),
	.w3(32'hbac46753),
	.w4(32'h38b87f37),
	.w5(32'h39dbccee),
	.w6(32'h39b41ba2),
	.w7(32'h398dec4e),
	.w8(32'h3a0286b4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e4030),
	.w1(32'hb993e9bb),
	.w2(32'h3a5002d9),
	.w3(32'h3a3d333c),
	.w4(32'h3a727c6e),
	.w5(32'h3a5d0fbc),
	.w6(32'h3a502755),
	.w7(32'h3a8bede0),
	.w8(32'h3ac8ae64),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09f943),
	.w1(32'hb9cc1baa),
	.w2(32'h3aac12c1),
	.w3(32'hbb4c3567),
	.w4(32'hba8ec60c),
	.w5(32'hba00f3dd),
	.w6(32'hbab86cc7),
	.w7(32'h3a31ac03),
	.w8(32'h3aa28b8b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb957b4a),
	.w1(32'hbb65a002),
	.w2(32'hba9b330a),
	.w3(32'hbb264731),
	.w4(32'hba9f4d29),
	.w5(32'h3a5b7a3e),
	.w6(32'hbad50bdf),
	.w7(32'hbb2d3641),
	.w8(32'h38c2732d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74397a),
	.w1(32'h3a45e62c),
	.w2(32'h3988e35c),
	.w3(32'hb99efbc4),
	.w4(32'h3a756da7),
	.w5(32'h3a107ade),
	.w6(32'hba3f7372),
	.w7(32'h39186532),
	.w8(32'h3a330c03),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba932ae2),
	.w1(32'hba905a84),
	.w2(32'h3a04d8d8),
	.w3(32'h39de05dd),
	.w4(32'h38296230),
	.w5(32'h3994c389),
	.w6(32'h39e23b22),
	.w7(32'hb7dcfa9d),
	.w8(32'hb9b1f065),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8392382),
	.w1(32'h39333e24),
	.w2(32'h39771d92),
	.w3(32'hb825ebea),
	.w4(32'h390dc677),
	.w5(32'hb71d4a9d),
	.w6(32'h393273ca),
	.w7(32'h39c54290),
	.w8(32'h38eb3e77),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cafad2),
	.w1(32'hba733417),
	.w2(32'h3aacb4c0),
	.w3(32'h3b0aca69),
	.w4(32'hba571089),
	.w5(32'h3a087ee1),
	.w6(32'h3b08d532),
	.w7(32'h3ab18dc4),
	.w8(32'h3984ed1a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ca0b77),
	.w1(32'hbaa2552d),
	.w2(32'h39e3d165),
	.w3(32'h3a1bce70),
	.w4(32'hba42df4c),
	.w5(32'h3a06b4b5),
	.w6(32'hb9cca8b3),
	.w7(32'h38d2211d),
	.w8(32'h39e8a7e2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c1756),
	.w1(32'hb9fc423e),
	.w2(32'hba9d98b8),
	.w3(32'hbb4a5458),
	.w4(32'hbb3236db),
	.w5(32'hba18895d),
	.w6(32'hbad8c6c2),
	.w7(32'hb9d62e13),
	.w8(32'h39945261),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba262aef),
	.w1(32'h3a203697),
	.w2(32'h3a4b7f7c),
	.w3(32'hba60d432),
	.w4(32'h39e88abb),
	.w5(32'h3941881f),
	.w6(32'h3937d1fc),
	.w7(32'h39399e4c),
	.w8(32'h39763c40),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc948fd),
	.w1(32'h3ad17975),
	.w2(32'h3a632ff3),
	.w3(32'h3ba096e2),
	.w4(32'h39c563ba),
	.w5(32'hb9c1e285),
	.w6(32'h3b539552),
	.w7(32'h3ab8847f),
	.w8(32'hbab5fc91),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a13bf),
	.w1(32'hb9ece66e),
	.w2(32'h39c6f353),
	.w3(32'hba48c602),
	.w4(32'hb9bd023a),
	.w5(32'hb7e76ba7),
	.w6(32'hba306934),
	.w7(32'hb94acf41),
	.w8(32'hb9d3e532),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07fda3),
	.w1(32'hb85a3ca1),
	.w2(32'h39863725),
	.w3(32'hb9eb82b6),
	.w4(32'hb910501e),
	.w5(32'hb93f8b14),
	.w6(32'h39bde407),
	.w7(32'h381ab637),
	.w8(32'hb9b6541c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bd05a),
	.w1(32'hba84d77f),
	.w2(32'hb9c39f97),
	.w3(32'hbb1a7ca5),
	.w4(32'h39f1e300),
	.w5(32'h39a55336),
	.w6(32'hba8eaddd),
	.w7(32'h3a6325e2),
	.w8(32'h3ad520f5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b179fa),
	.w1(32'hba0526e6),
	.w2(32'h3b079c91),
	.w3(32'h3a7ee93e),
	.w4(32'hba872b52),
	.w5(32'hbb5b57fa),
	.w6(32'hba4f709c),
	.w7(32'h3b60ae15),
	.w8(32'hba47ee3d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fec8c),
	.w1(32'h3a908592),
	.w2(32'h3a5147bf),
	.w3(32'h39a5ca0a),
	.w4(32'h39b568b5),
	.w5(32'h38f89b40),
	.w6(32'h3a26a546),
	.w7(32'h3a0f2e2a),
	.w8(32'h38d4b035),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe0edb),
	.w1(32'h3b20d0dc),
	.w2(32'h3a02b8a0),
	.w3(32'hbb453d21),
	.w4(32'h39f00f84),
	.w5(32'hba7bc4d5),
	.w6(32'h3a5b07ef),
	.w7(32'h3b3023c0),
	.w8(32'h39dc2177),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca2fe4),
	.w1(32'hbb04a876),
	.w2(32'hb98fbdc7),
	.w3(32'hba87ffeb),
	.w4(32'hbb232be0),
	.w5(32'h3a0dc31e),
	.w6(32'hb9d334e0),
	.w7(32'hbb10be88),
	.w8(32'hb9f4f3dc),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ff0a6),
	.w1(32'hbb81c4e7),
	.w2(32'hba684d0e),
	.w3(32'hbb38f466),
	.w4(32'hbb9cb4fe),
	.w5(32'hbaadba9c),
	.w6(32'hba89cb40),
	.w7(32'hbb8185fc),
	.w8(32'hbb2786f9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5faf7f),
	.w1(32'hbad57a2c),
	.w2(32'hba228de5),
	.w3(32'h379dab09),
	.w4(32'hb9c68773),
	.w5(32'hba8fa8e1),
	.w6(32'h3a5dd7b4),
	.w7(32'h39c3a905),
	.w8(32'hba7bb9b8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43518f),
	.w1(32'hba812445),
	.w2(32'hbae38fdc),
	.w3(32'hba27992e),
	.w4(32'hbae52f84),
	.w5(32'hbb5cbfda),
	.w6(32'h3b30fadf),
	.w7(32'h3b0659df),
	.w8(32'hbb182eba),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9875cac),
	.w1(32'h397b8d6d),
	.w2(32'hb90fece2),
	.w3(32'h3a9ee669),
	.w4(32'h39fed5c7),
	.w5(32'hb944b67a),
	.w6(32'h3901cf06),
	.w7(32'h38565f6a),
	.w8(32'h39bb6984),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae610a0),
	.w1(32'hbb082088),
	.w2(32'h39959727),
	.w3(32'h3a17ee0f),
	.w4(32'hbb363994),
	.w5(32'hba221d20),
	.w6(32'h3b2fe740),
	.w7(32'hbabdbefc),
	.w8(32'hbb080031),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382c148a),
	.w1(32'hb89ee31d),
	.w2(32'h396c292b),
	.w3(32'hb93b8952),
	.w4(32'hb8538ef0),
	.w5(32'hb79b29a4),
	.w6(32'h3917e3e5),
	.w7(32'h3808c837),
	.w8(32'h38c40b25),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e6aa8),
	.w1(32'hba8cba2b),
	.w2(32'h39cafe12),
	.w3(32'hba95be2e),
	.w4(32'hba5fb423),
	.w5(32'h3a24e79c),
	.w6(32'hba74e413),
	.w7(32'hb9ae4cbb),
	.w8(32'hb8a40d98),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85bc7d),
	.w1(32'hb9d0454c),
	.w2(32'h39be3b63),
	.w3(32'hbaa93676),
	.w4(32'hb921d9a4),
	.w5(32'hba66b8a5),
	.w6(32'h38c6feee),
	.w7(32'h3a0a6a56),
	.w8(32'h39c5475c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab9ff2),
	.w1(32'h3ad0c2d7),
	.w2(32'h3ab8abb6),
	.w3(32'h3b2c8011),
	.w4(32'hba8e7ec3),
	.w5(32'hba153e16),
	.w6(32'h3b057543),
	.w7(32'hbaa0021a),
	.w8(32'hbb38f638),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a924cb),
	.w1(32'h394e8254),
	.w2(32'h3916499b),
	.w3(32'hb9e5bef7),
	.w4(32'h39be79a0),
	.w5(32'hb8245dcd),
	.w6(32'h39dcba9e),
	.w7(32'h392b7759),
	.w8(32'h39db05d6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e3646),
	.w1(32'hb99d0259),
	.w2(32'hba0c3275),
	.w3(32'hba12c99c),
	.w4(32'hb9ad1599),
	.w5(32'hb99bf6a2),
	.w6(32'h397d3968),
	.w7(32'hb889a3f3),
	.w8(32'hb8636c27),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de795f),
	.w1(32'h39b23622),
	.w2(32'h390cf7a7),
	.w3(32'hbabf670a),
	.w4(32'hba2aa79b),
	.w5(32'h3a20fbe4),
	.w6(32'h38367f2b),
	.w7(32'h39488c7d),
	.w8(32'h39bc7786),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb417889),
	.w1(32'hbada1003),
	.w2(32'hba226202),
	.w3(32'h3a60bf3d),
	.w4(32'h3ab75027),
	.w5(32'hba07443f),
	.w6(32'h39a40acd),
	.w7(32'h3b0575a6),
	.w8(32'h3a328bb6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb185b19),
	.w1(32'hbbd26fd7),
	.w2(32'h39be08c2),
	.w3(32'hb96b152a),
	.w4(32'hbae9f961),
	.w5(32'h3b784867),
	.w6(32'h3accf3b5),
	.w7(32'h3a9c8ffe),
	.w8(32'h3b9b8e6d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53df7c),
	.w1(32'hba2c5bd7),
	.w2(32'hba1b3f6c),
	.w3(32'h38ff5daf),
	.w4(32'hba83908b),
	.w5(32'hba963166),
	.w6(32'hba6af822),
	.w7(32'hba239670),
	.w8(32'hbab90553),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09c002),
	.w1(32'h39fdc9f2),
	.w2(32'hba0755e2),
	.w3(32'h3b8f974d),
	.w4(32'hba9438e8),
	.w5(32'hbbe16291),
	.w6(32'h3bbac30e),
	.w7(32'h3ae62113),
	.w8(32'hbbd767c8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc279342),
	.w1(32'hbbac0b87),
	.w2(32'h3a4f7f28),
	.w3(32'hbc1864e6),
	.w4(32'hbbb5f359),
	.w5(32'h3bad85a8),
	.w6(32'hbb2034da),
	.w7(32'hbb834dbb),
	.w8(32'h3a005547),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba291542),
	.w1(32'hbabb9884),
	.w2(32'h3ab34557),
	.w3(32'h39a66cd8),
	.w4(32'hba107f33),
	.w5(32'h3a4e1b0a),
	.w6(32'h3a5091e0),
	.w7(32'hb821d87c),
	.w8(32'h38ab0ecd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380fe742),
	.w1(32'hba02ced8),
	.w2(32'hb9f19a31),
	.w3(32'hb89087ba),
	.w4(32'hb9e380a7),
	.w5(32'hba807c5e),
	.w6(32'h3a112cda),
	.w7(32'hb8ecef97),
	.w8(32'h38d214d5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d26130),
	.w1(32'hba2ef0d7),
	.w2(32'hba1a5677),
	.w3(32'h399446de),
	.w4(32'hb999fc9d),
	.w5(32'hb9e34db0),
	.w6(32'hb9abb707),
	.w7(32'hb9a00f22),
	.w8(32'hba038612),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f4400),
	.w1(32'hb84669e0),
	.w2(32'h38c829f3),
	.w3(32'hb9c51103),
	.w4(32'hb953a1ca),
	.w5(32'h3996f972),
	.w6(32'hb95d5225),
	.w7(32'h39418a3a),
	.w8(32'h37a168a1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba3274),
	.w1(32'h388d2aeb),
	.w2(32'h3b37bf86),
	.w3(32'h3ab1a099),
	.w4(32'h39f1e839),
	.w5(32'h3a5d76d4),
	.w6(32'h3a87a47d),
	.w7(32'h3b0e892d),
	.w8(32'h3a5cd2df),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a14df),
	.w1(32'hbb0ff1b3),
	.w2(32'hb9c396b0),
	.w3(32'h39a0595f),
	.w4(32'hba97cf63),
	.w5(32'h39e23f94),
	.w6(32'hbab8dd13),
	.w7(32'hba6dcba8),
	.w8(32'hba701227),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb340b18),
	.w1(32'hba1927b5),
	.w2(32'hb92902ef),
	.w3(32'hbb8bbef6),
	.w4(32'hb9c9756f),
	.w5(32'h387df789),
	.w6(32'hba973b77),
	.w7(32'h3a9ddc14),
	.w8(32'h3a28e391),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb804bff6),
	.w1(32'hba047d25),
	.w2(32'h3a010212),
	.w3(32'hba1a3cfb),
	.w4(32'hb9b7ce92),
	.w5(32'hb9467535),
	.w6(32'h38a3dbf1),
	.w7(32'h39bb005c),
	.w8(32'h3a0b8853),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecc831),
	.w1(32'h392fdfef),
	.w2(32'h3ab900cf),
	.w3(32'h3ae4e0c5),
	.w4(32'h3aa7c6a0),
	.w5(32'hba00a7c8),
	.w6(32'h3aa9de16),
	.w7(32'h3b185f77),
	.w8(32'hbab2bd4e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3cff1),
	.w1(32'hbb0ebf4d),
	.w2(32'hbac74b7d),
	.w3(32'hbae95635),
	.w4(32'hba6a37b4),
	.w5(32'hba79097c),
	.w6(32'hbab172ea),
	.w7(32'h37312783),
	.w8(32'h39bce05c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e4253),
	.w1(32'hb8acfbca),
	.w2(32'h392ab12f),
	.w3(32'hba26c95a),
	.w4(32'hb9299338),
	.w5(32'hb96a923a),
	.w6(32'h390425f5),
	.w7(32'hb8f7913e),
	.w8(32'h385e3305),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a0177),
	.w1(32'h39b875ec),
	.w2(32'hba998207),
	.w3(32'h3918590f),
	.w4(32'hbacccabc),
	.w5(32'hbb05bf12),
	.w6(32'h3a001487),
	.w7(32'hba0e00b3),
	.w8(32'hbad27774),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6850c35),
	.w1(32'h39c3fe95),
	.w2(32'h3a2177fd),
	.w3(32'hb9457e3e),
	.w4(32'h39280cad),
	.w5(32'hb854351b),
	.w6(32'h393608db),
	.w7(32'h391e60ac),
	.w8(32'h38a9d748),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba245570),
	.w1(32'hb9ba8c48),
	.w2(32'hb8753f20),
	.w3(32'hb8cb6764),
	.w4(32'hb8caadf7),
	.w5(32'h39dd318b),
	.w6(32'hb8426089),
	.w7(32'h3a4b82d3),
	.w8(32'h38506881),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb473fc4),
	.w1(32'hb99017d6),
	.w2(32'hbb1a0ab1),
	.w3(32'hbb84d5bd),
	.w4(32'hb9d2f669),
	.w5(32'h3b06fadd),
	.w6(32'hb91f2caf),
	.w7(32'h3a08522d),
	.w8(32'h3b14b3c5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285e56),
	.w1(32'h38c24da8),
	.w2(32'h3a0aa988),
	.w3(32'hb9f28bf3),
	.w4(32'h3978a541),
	.w5(32'h3a505eb7),
	.w6(32'hb9ce9c78),
	.w7(32'h39f926d7),
	.w8(32'h3abea676),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b4e45),
	.w1(32'h39901e7c),
	.w2(32'hb8951f24),
	.w3(32'h3a0f3eae),
	.w4(32'hb928de86),
	.w5(32'hb9ac601a),
	.w6(32'h39ba2f1c),
	.w7(32'hb9c40741),
	.w8(32'hb950a42f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a136d),
	.w1(32'h390ca134),
	.w2(32'hba3b4039),
	.w3(32'hbb490499),
	.w4(32'hbb03534e),
	.w5(32'h3aa029fe),
	.w6(32'h3a234557),
	.w7(32'hba5030aa),
	.w8(32'h3a32ebf9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85f66e),
	.w1(32'hb9aa2410),
	.w2(32'hba6e6d21),
	.w3(32'h3b032ff6),
	.w4(32'hbaabf072),
	.w5(32'hbb4bc164),
	.w6(32'h3affff22),
	.w7(32'hb9b1a1bd),
	.w8(32'hbaf8be79),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab37318),
	.w1(32'h3a27ea64),
	.w2(32'h3af45623),
	.w3(32'h3ae4403c),
	.w4(32'hb97107a8),
	.w5(32'hb9ad39ac),
	.w6(32'h3b06a656),
	.w7(32'h3aec772a),
	.w8(32'hba70a3cf),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964cb32),
	.w1(32'hba4a05de),
	.w2(32'hb9264e00),
	.w3(32'hb99165c5),
	.w4(32'hb9fe0a2b),
	.w5(32'hb9ed2fb2),
	.w6(32'hb979ef24),
	.w7(32'hb9a9be0a),
	.w8(32'hb9d3e447),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b8fd8),
	.w1(32'hb93703c4),
	.w2(32'hb885d2a9),
	.w3(32'hb94fb8ae),
	.w4(32'hb9ad6e96),
	.w5(32'hb9c82502),
	.w6(32'h39ca6e1c),
	.w7(32'hb99e9d9b),
	.w8(32'hb994f2bf),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87bbdc),
	.w1(32'hbb4ed83c),
	.w2(32'hb8d174bf),
	.w3(32'h3aaa536e),
	.w4(32'h396be7d0),
	.w5(32'hba8322e8),
	.w6(32'hba88f8ed),
	.w7(32'h3af49431),
	.w8(32'h3b52e881),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998e263),
	.w1(32'hba10a725),
	.w2(32'hba9f8897),
	.w3(32'h395eabdf),
	.w4(32'hba612fa6),
	.w5(32'hbb63a221),
	.w6(32'h391d0a12),
	.w7(32'h3b20db16),
	.w8(32'hb9dd5e8f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb0a9b),
	.w1(32'hba885d76),
	.w2(32'hb9d9d2bd),
	.w3(32'hbb1aa8a6),
	.w4(32'hba10c119),
	.w5(32'hb9125f02),
	.w6(32'hba700625),
	.w7(32'h3aa58165),
	.w8(32'h3a90d4cb),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d8ed),
	.w1(32'hbb4e8d5c),
	.w2(32'h3af3a9d8),
	.w3(32'h3b0f334c),
	.w4(32'h396f7f2f),
	.w5(32'h3b21a39b),
	.w6(32'h3b837374),
	.w7(32'hb9927d73),
	.w8(32'hbb22e5e4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ff117),
	.w1(32'h3a52c19c),
	.w2(32'hba070196),
	.w3(32'h39342152),
	.w4(32'h386c0a0d),
	.w5(32'hba69825e),
	.w6(32'hb952e8bb),
	.w7(32'hb9dea91e),
	.w8(32'hba77012d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a18cb),
	.w1(32'hb9dcdd67),
	.w2(32'hb9ec9f13),
	.w3(32'h39d02ad5),
	.w4(32'hba2e103f),
	.w5(32'hbaa72c31),
	.w6(32'h39e4dd1f),
	.w7(32'h3946b477),
	.w8(32'hb9d388f8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801aa0),
	.w1(32'hbb487fb5),
	.w2(32'h3bb9c536),
	.w3(32'hbb55b8f1),
	.w4(32'h3ac7cac3),
	.w5(32'h3beb1e42),
	.w6(32'hbb9fae05),
	.w7(32'h3b77b47e),
	.w8(32'h3c0975e2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b019d59),
	.w1(32'hbaaaf7b2),
	.w2(32'h3b0f138b),
	.w3(32'h3b31c815),
	.w4(32'hbb448680),
	.w5(32'hbae1a87a),
	.w6(32'h3b4882d1),
	.w7(32'hb96e4f81),
	.w8(32'hbb546430),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5f603),
	.w1(32'hbade438c),
	.w2(32'h3aa1b85e),
	.w3(32'h3b4a9634),
	.w4(32'h3a849b39),
	.w5(32'h3b10bc18),
	.w6(32'h3a8a8eb1),
	.w7(32'h3b2dc633),
	.w8(32'h392a7460),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5c491),
	.w1(32'hb8734ac2),
	.w2(32'hba0d1210),
	.w3(32'hbb6b33e4),
	.w4(32'hba6bab79),
	.w5(32'h398f970c),
	.w6(32'hbb250149),
	.w7(32'hba8011de),
	.w8(32'h3a6bafd8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb829465),
	.w1(32'h39e73af8),
	.w2(32'hb8bc26be),
	.w3(32'hbb8957a7),
	.w4(32'hb9ccc3a7),
	.w5(32'h3ab40ad5),
	.w6(32'hbabd67fe),
	.w7(32'hb9de1bf9),
	.w8(32'h398e3955),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd5beb),
	.w1(32'h39bf752a),
	.w2(32'h39ee389c),
	.w3(32'h3908d9a5),
	.w4(32'h39286ee3),
	.w5(32'hb81078b7),
	.w6(32'h39c0ed0e),
	.w7(32'h398911a6),
	.w8(32'h38185bf8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378bd256),
	.w1(32'h39a225f7),
	.w2(32'h39b587db),
	.w3(32'h36e89018),
	.w4(32'h399d85bd),
	.w5(32'h3a10d79b),
	.w6(32'h39c7d6c8),
	.w7(32'h39841d09),
	.w8(32'h38f7e96d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfb487),
	.w1(32'h3a25e73e),
	.w2(32'h3afd7650),
	.w3(32'hb9d7c825),
	.w4(32'hba64018e),
	.w5(32'h3a8a69c9),
	.w6(32'h399fe7a4),
	.w7(32'h390473d7),
	.w8(32'h3acb1d07),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae336ea),
	.w1(32'h38ba06a8),
	.w2(32'h39eb2927),
	.w3(32'h3aeebe95),
	.w4(32'hb8e0c73a),
	.w5(32'hb90c4b48),
	.w6(32'h38a05d64),
	.w7(32'h39ca7150),
	.w8(32'h399a925e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76e69f),
	.w1(32'hba28bdc7),
	.w2(32'h3a70c3b7),
	.w3(32'h3a945b83),
	.w4(32'hb9109427),
	.w5(32'hb8c7e04a),
	.w6(32'h39e6f89c),
	.w7(32'h3a1429ca),
	.w8(32'hb8c94d50),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8f90e),
	.w1(32'h3a8d1ced),
	.w2(32'hba9be130),
	.w3(32'h3b6f3518),
	.w4(32'h3aa70d07),
	.w5(32'hbb0377b7),
	.w6(32'h3ada60cb),
	.w7(32'h3b369ee7),
	.w8(32'h3af5f2c0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba681f4b),
	.w1(32'hb99019c3),
	.w2(32'h3aa2d0b7),
	.w3(32'hbafca660),
	.w4(32'hb9bde619),
	.w5(32'h3a04ba3d),
	.w6(32'hba2400a1),
	.w7(32'h3adb6b80),
	.w8(32'h3af5ce58),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e3c15),
	.w1(32'hba77f197),
	.w2(32'hb7af6bab),
	.w3(32'h3a4cf844),
	.w4(32'hb7e3f3a1),
	.w5(32'h38ffce76),
	.w6(32'hba941e16),
	.w7(32'hba979aec),
	.w8(32'hb8ea3ed8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f9552),
	.w1(32'hba50447f),
	.w2(32'h3b815f35),
	.w3(32'h3b5b51d4),
	.w4(32'h3b096cc5),
	.w5(32'h3a9a5c61),
	.w6(32'h3aa9a50f),
	.w7(32'h3bc12db4),
	.w8(32'hba1b213f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a704a8c),
	.w1(32'hb943f593),
	.w2(32'h3a1a3b60),
	.w3(32'h3ac36029),
	.w4(32'hb998eb3c),
	.w5(32'hba0ec572),
	.w6(32'h3ab4bdd5),
	.w7(32'h3a6df8d0),
	.w8(32'hbab1fe64),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973fc46),
	.w1(32'h3919ef25),
	.w2(32'h39da9976),
	.w3(32'h38933746),
	.w4(32'h3983fe9e),
	.w5(32'h39dd82e3),
	.w6(32'h39d237d1),
	.w7(32'h3981603d),
	.w8(32'h39bd01ff),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cf281),
	.w1(32'h3991c14f),
	.w2(32'h3b1a46b3),
	.w3(32'h3ae47e49),
	.w4(32'h39c7ed34),
	.w5(32'h3a27ab37),
	.w6(32'h3aa78300),
	.w7(32'h388a86be),
	.w8(32'hba29c746),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380c8015),
	.w1(32'h38cdcd13),
	.w2(32'h36d54729),
	.w3(32'hb8eee7e2),
	.w4(32'hb90e5011),
	.w5(32'hb9dfc291),
	.w6(32'hb7d56bf8),
	.w7(32'hb966bef8),
	.w8(32'hb9acf1dc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c07080),
	.w1(32'h3987fe92),
	.w2(32'h38e8e1f3),
	.w3(32'hb94e7732),
	.w4(32'hb87e59a7),
	.w5(32'hba02676c),
	.w6(32'h39b96313),
	.w7(32'h3a30173c),
	.w8(32'h397df92f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d00363),
	.w1(32'h39197e91),
	.w2(32'h39e263a3),
	.w3(32'hb98e884a),
	.w4(32'h3989c917),
	.w5(32'h39b9f86c),
	.w6(32'h39c36c0e),
	.w7(32'h396b40ab),
	.w8(32'h39c30ff6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ffbcd6),
	.w1(32'hb9073d84),
	.w2(32'hba531380),
	.w3(32'h3993e955),
	.w4(32'hb99d2f1e),
	.w5(32'hb9de410d),
	.w6(32'h398cd608),
	.w7(32'hb9a485df),
	.w8(32'h392777cd),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d0378),
	.w1(32'h3a5e3e66),
	.w2(32'h3b18fb83),
	.w3(32'hbb1788d1),
	.w4(32'h3a13d727),
	.w5(32'h3aab4ba4),
	.w6(32'hbae76316),
	.w7(32'h3a09066f),
	.w8(32'h3abbdd26),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87a0b4),
	.w1(32'h3a34f80b),
	.w2(32'h38fdd668),
	.w3(32'hba0dfda0),
	.w4(32'hbb52744e),
	.w5(32'hbb01a44b),
	.w6(32'h3b690648),
	.w7(32'hba9a583a),
	.w8(32'hbb340e78),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d67c5b),
	.w1(32'hbaeb99a1),
	.w2(32'h3abf29e6),
	.w3(32'h3b12fec6),
	.w4(32'hba71cd05),
	.w5(32'hba5efda1),
	.w6(32'h3aeb2e1a),
	.w7(32'h3a742b30),
	.w8(32'hba01c94d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb177da7),
	.w1(32'hba075172),
	.w2(32'h3ac7c7e2),
	.w3(32'hba3147a4),
	.w4(32'hbb219590),
	.w5(32'h39e621c8),
	.w6(32'h3b013aca),
	.w7(32'hb9ff6aec),
	.w8(32'hbaec05a8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ab28c),
	.w1(32'h39c26b86),
	.w2(32'h39e31236),
	.w3(32'hba250ba1),
	.w4(32'hb75ee67f),
	.w5(32'h392b2b5c),
	.w6(32'h33a69d0f),
	.w7(32'h39c784f3),
	.w8(32'h39a3fc37),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34794f),
	.w1(32'h3a0fd231),
	.w2(32'h397e6aa7),
	.w3(32'h3a1a0997),
	.w4(32'h39ea5f14),
	.w5(32'h39c2bb7f),
	.w6(32'h3a9361e3),
	.w7(32'h39d5d3d4),
	.w8(32'h38fedeef),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f546a7),
	.w1(32'h3927e7f7),
	.w2(32'h39866590),
	.w3(32'h39919d2a),
	.w4(32'h399cd05b),
	.w5(32'h3979e2f1),
	.w6(32'h3a01c686),
	.w7(32'h39604116),
	.w8(32'h39292e44),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39290a72),
	.w1(32'h3992a149),
	.w2(32'h3993ee2a),
	.w3(32'h38c4149f),
	.w4(32'h39aad7ed),
	.w5(32'h392bd500),
	.w6(32'h3a1e1391),
	.w7(32'h39a05608),
	.w8(32'h39775e69),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e7322),
	.w1(32'hbaed5a9d),
	.w2(32'hba94aa6e),
	.w3(32'h3aae61c7),
	.w4(32'hbb8525be),
	.w5(32'hbb309051),
	.w6(32'h3b27c3c4),
	.w7(32'hbb1b10f1),
	.w8(32'hbb3341b2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba442b51),
	.w1(32'hb9db627e),
	.w2(32'h3a83ca4f),
	.w3(32'hb942f717),
	.w4(32'hba084e21),
	.w5(32'h3981fefb),
	.w6(32'hb8fdfdf3),
	.w7(32'h3a2a83d2),
	.w8(32'h38d6cdf5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa17a28),
	.w1(32'h3a7fcb16),
	.w2(32'h3a9347c0),
	.w3(32'h3a649a53),
	.w4(32'h39d59f58),
	.w5(32'h39d4a469),
	.w6(32'h3aa8e574),
	.w7(32'h3a573bcc),
	.w8(32'h3a26c173),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b34fa0),
	.w1(32'hb9872882),
	.w2(32'hba96bf5d),
	.w3(32'hbac23e38),
	.w4(32'hbaa91afa),
	.w5(32'hbaafad86),
	.w6(32'h39a3770c),
	.w7(32'hba49eb8d),
	.w8(32'h366fab96),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3879c1ed),
	.w1(32'h39742164),
	.w2(32'h39b73ef8),
	.w3(32'hb987c999),
	.w4(32'h3931d600),
	.w5(32'h37c9cfbc),
	.w6(32'h398cb742),
	.w7(32'h395c5a53),
	.w8(32'h393907b3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41047e),
	.w1(32'h3a71137a),
	.w2(32'h3b0613cd),
	.w3(32'h3aa78dd3),
	.w4(32'h3a839955),
	.w5(32'h3aa93bd2),
	.w6(32'h38f1ac8d),
	.w7(32'hb9f1245c),
	.w8(32'hb74dd872),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f144f4),
	.w1(32'h39972291),
	.w2(32'hb8d9ff30),
	.w3(32'h3a1dd99e),
	.w4(32'h3a10ae2f),
	.w5(32'hba108ad5),
	.w6(32'h3a81d7ed),
	.w7(32'h38f854f0),
	.w8(32'hba7ec52b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf0a66),
	.w1(32'hbac4fc71),
	.w2(32'h3abac132),
	.w3(32'hba766fcc),
	.w4(32'hbc09d52b),
	.w5(32'hb97cad83),
	.w6(32'h3acf8a7d),
	.w7(32'hbbfd1ec3),
	.w8(32'hbbbc1e39),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d34308),
	.w1(32'h38bcde46),
	.w2(32'h38f68cf4),
	.w3(32'hb9b0eac2),
	.w4(32'h38db4e9b),
	.w5(32'h38c582f3),
	.w6(32'h37c81ace),
	.w7(32'h380e7c9e),
	.w8(32'hb6d0996b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93e03c),
	.w1(32'hbb141f9d),
	.w2(32'h37490249),
	.w3(32'hbb921fb0),
	.w4(32'hba88d80c),
	.w5(32'h3a30eda5),
	.w6(32'hbb3ec353),
	.w7(32'h3aac43cb),
	.w8(32'h3b2dda78),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule