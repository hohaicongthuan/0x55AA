module layer_8_featuremap_40(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4f4f3),
	.w1(32'hb8c7c1ea),
	.w2(32'h3924fa46),
	.w3(32'h3985387c),
	.w4(32'h37b7bd9c),
	.w5(32'h38873b51),
	.w6(32'hb6200ee3),
	.w7(32'h39a38497),
	.w8(32'hb96064d0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b80ab6),
	.w1(32'hb92a49c8),
	.w2(32'hb9503ed0),
	.w3(32'h3859c987),
	.w4(32'hb8c5af96),
	.w5(32'hb953e969),
	.w6(32'hb97ca71c),
	.w7(32'hb88b2dfe),
	.w8(32'hb9386fc9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b52b64),
	.w1(32'hb92c417d),
	.w2(32'hb937cb73),
	.w3(32'h3877123b),
	.w4(32'hb919b7a9),
	.w5(32'hb964cb58),
	.w6(32'hb970998c),
	.w7(32'hb8cf6bf2),
	.w8(32'h39aafa88),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ab30f0),
	.w1(32'h3a961032),
	.w2(32'h394746db),
	.w3(32'h39f631e0),
	.w4(32'h3ac0f19b),
	.w5(32'h3a848d13),
	.w6(32'hb6a60535),
	.w7(32'hba3ca279),
	.w8(32'h39e7d51a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efd87f),
	.w1(32'h387583f4),
	.w2(32'h39a369ab),
	.w3(32'h39d95450),
	.w4(32'h38882495),
	.w5(32'h390d244c),
	.w6(32'h3863811a),
	.w7(32'h39fffdf3),
	.w8(32'h3ad2a281),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4be23),
	.w1(32'h39f33b90),
	.w2(32'h3a843b02),
	.w3(32'h39825a53),
	.w4(32'h3a1daf9b),
	.w5(32'h3a5c5294),
	.w6(32'h3b0c15ee),
	.w7(32'h3b32907d),
	.w8(32'hb8fc5ae4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e35e5d),
	.w1(32'hb92e29d6),
	.w2(32'h37c3a2ab),
	.w3(32'h39530a88),
	.w4(32'hb8cef49e),
	.w5(32'hb948017e),
	.w6(32'hb889d487),
	.w7(32'h39a180f3),
	.w8(32'h3a1a5d8a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a293fa2),
	.w1(32'h38fe6378),
	.w2(32'h39e09ae8),
	.w3(32'h3a449f34),
	.w4(32'h39c9c388),
	.w5(32'h39d00a16),
	.w6(32'hb76df1b4),
	.w7(32'h39dfaf5c),
	.w8(32'hb92052ba),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c9797),
	.w1(32'hb926c71d),
	.w2(32'hb8a2caab),
	.w3(32'h3982f534),
	.w4(32'hb95f8df3),
	.w5(32'hb9a1ae48),
	.w6(32'hb95b114e),
	.w7(32'h3946eb65),
	.w8(32'hb8ab5ee1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab40e52),
	.w1(32'hbad61c82),
	.w2(32'hba7d3185),
	.w3(32'hba94f44d),
	.w4(32'hb99a624f),
	.w5(32'hb9d70192),
	.w6(32'hba2128bd),
	.w7(32'hbaab6a85),
	.w8(32'h39d268da),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20d963),
	.w1(32'h392f98ad),
	.w2(32'h39a1807b),
	.w3(32'h3a06c3f4),
	.w4(32'h3868625d),
	.w5(32'h377f634b),
	.w6(32'h38a11709),
	.w7(32'h398dff3e),
	.w8(32'hb9a6877a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88df934),
	.w1(32'hb9a18330),
	.w2(32'hb959ff0f),
	.w3(32'h38fe3ae7),
	.w4(32'hb89a5f7a),
	.w5(32'hb91eba7a),
	.w6(32'hb9c8274b),
	.w7(32'hb8d27223),
	.w8(32'h38e38a03),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39383ebb),
	.w1(32'hb8c8154a),
	.w2(32'h3850dff7),
	.w3(32'h39716118),
	.w4(32'hb917c0ad),
	.w5(32'hb9307562),
	.w6(32'hb8e3cfbb),
	.w7(32'h39af4809),
	.w8(32'h3af506f4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d28bf),
	.w1(32'h39cc789c),
	.w2(32'h3a97d946),
	.w3(32'h39150917),
	.w4(32'h3a1b6289),
	.w5(32'h3a75faed),
	.w6(32'h3b2e616c),
	.w7(32'h3b615822),
	.w8(32'h3a0c1f9b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80466ac),
	.w1(32'h395d6a4b),
	.w2(32'h39cb9a63),
	.w3(32'h3985d273),
	.w4(32'h399ecc95),
	.w5(32'h39a88f46),
	.w6(32'h3a5caa80),
	.w7(32'h3a9cf85a),
	.w8(32'hb888c5c8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9322f48),
	.w1(32'h382b459a),
	.w2(32'h390a81d4),
	.w3(32'hb925bb09),
	.w4(32'hb9438fdd),
	.w5(32'hb9007891),
	.w6(32'h37e25572),
	.w7(32'h38251359),
	.w8(32'h39c81f08),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac367b8),
	.w1(32'h3a734671),
	.w2(32'hb9464a0e),
	.w3(32'h3aafa5e2),
	.w4(32'h3b7d6f51),
	.w5(32'h3b236db4),
	.w6(32'h3ada582f),
	.w7(32'h3a8a62fb),
	.w8(32'h3995a525),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39add3f2),
	.w1(32'h37275784),
	.w2(32'h3994d2ee),
	.w3(32'h3a49ca59),
	.w4(32'h38ac437e),
	.w5(32'h39979a79),
	.w6(32'hb8b436a7),
	.w7(32'h39d058e1),
	.w8(32'h3915c445),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f0b75),
	.w1(32'hba2dfe59),
	.w2(32'hb8f39e55),
	.w3(32'h39d5461a),
	.w4(32'hba37a83b),
	.w5(32'hb98a3977),
	.w6(32'hba1b1fe3),
	.w7(32'h390bef8a),
	.w8(32'h3ae67633),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4de841),
	.w1(32'hba6338c3),
	.w2(32'hbb0a5adc),
	.w3(32'h3a608be6),
	.w4(32'h3a479297),
	.w5(32'h3a9be65d),
	.w6(32'h3a0819cb),
	.w7(32'h3963b848),
	.w8(32'hb8d36353),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd67cc),
	.w1(32'hb9b8b6b4),
	.w2(32'h3743adae),
	.w3(32'h394844c5),
	.w4(32'hb9592a2c),
	.w5(32'h38d29d94),
	.w6(32'hb820e1fb),
	.w7(32'h39d8a816),
	.w8(32'h395f38aa),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b22aa5),
	.w1(32'hba416b51),
	.w2(32'hba22f175),
	.w3(32'hb7eea006),
	.w4(32'hba2887b7),
	.w5(32'hba2f9bdf),
	.w6(32'hb960b648),
	.w7(32'hb9b1367a),
	.w8(32'h38bb9758),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8871a30),
	.w1(32'hb99520a5),
	.w2(32'h3a0a69f2),
	.w3(32'hba8bdf7f),
	.w4(32'hba391bb4),
	.w5(32'h3951a445),
	.w6(32'h3a43d172),
	.w7(32'h3adcd68e),
	.w8(32'h3a119eb5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370c9682),
	.w1(32'hba125968),
	.w2(32'h399ba3d2),
	.w3(32'h3988afcb),
	.w4(32'hb90a3c4c),
	.w5(32'h3a0ce7d5),
	.w6(32'hb9959725),
	.w7(32'h399d8ca0),
	.w8(32'hbadcd67b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16bc96),
	.w1(32'hbb0c966e),
	.w2(32'hbad9d894),
	.w3(32'hbb03e9c6),
	.w4(32'hbb0d4e9e),
	.w5(32'hbac97dca),
	.w6(32'hbb117e4e),
	.w7(32'hbb19a102),
	.w8(32'h3a1653b6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f90734),
	.w1(32'hba381351),
	.w2(32'h38cb44a8),
	.w3(32'hba8938ec),
	.w4(32'hba5ab062),
	.w5(32'hb80db353),
	.w6(32'h3a0e424e),
	.w7(32'h3aaf7c16),
	.w8(32'h3a0048f1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d87aaf),
	.w1(32'hba20aa95),
	.w2(32'h39004799),
	.w3(32'hba79581c),
	.w4(32'hba4a4db9),
	.w5(32'hb8357479),
	.w6(32'h39f35983),
	.w7(32'h3a92b883),
	.w8(32'hb946d2ac),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391400aa),
	.w1(32'h39203eb5),
	.w2(32'h396faa74),
	.w3(32'hb9ade003),
	.w4(32'hb99ae94e),
	.w5(32'hb7584a39),
	.w6(32'hb99d05db),
	.w7(32'h3a0a73c0),
	.w8(32'hb9a7395b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf46345),
	.w1(32'hba988b59),
	.w2(32'h3adc7930),
	.w3(32'hba2aa25e),
	.w4(32'hba7914fe),
	.w5(32'hba432cec),
	.w6(32'h3abca134),
	.w7(32'h3a209d12),
	.w8(32'hb8f7f5ef),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388415e4),
	.w1(32'h37ec7add),
	.w2(32'hb8b4fee5),
	.w3(32'h38bf9259),
	.w4(32'hb767c191),
	.w5(32'hb951fec5),
	.w6(32'hb94c0bdf),
	.w7(32'hb9484f04),
	.w8(32'hba8a8e0d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62fac6),
	.w1(32'hbab4d004),
	.w2(32'hbba664cd),
	.w3(32'hba2c4dbf),
	.w4(32'h3a699698),
	.w5(32'h3a38e167),
	.w6(32'hba6f1191),
	.w7(32'hbafd0126),
	.w8(32'hb9b9ec9a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddaffa),
	.w1(32'hba812243),
	.w2(32'hb918be87),
	.w3(32'hb94a8987),
	.w4(32'hbaa55d72),
	.w5(32'hba1ff15e),
	.w6(32'hb9e0001b),
	.w7(32'h39d966b3),
	.w8(32'hb54775a6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5d481),
	.w1(32'hba0062ff),
	.w2(32'hbab92ffb),
	.w3(32'h3a1f5eb2),
	.w4(32'h3a3eb988),
	.w5(32'h3a13d5fb),
	.w6(32'hb92029a0),
	.w7(32'hba8eb3d6),
	.w8(32'hbabb4364),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb6a89),
	.w1(32'h39dc5af2),
	.w2(32'hbae1a994),
	.w3(32'hbaa954f3),
	.w4(32'hb9ef1e41),
	.w5(32'hba1ac4fd),
	.w6(32'hbaa2786e),
	.w7(32'hbaeefe85),
	.w8(32'h3ae086a2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94323fa),
	.w1(32'h39a5f3f2),
	.w2(32'h3a75fe4c),
	.w3(32'h390d3c4a),
	.w4(32'h3a015276),
	.w5(32'h3a477058),
	.w6(32'h3b164aab),
	.w7(32'h3b41a9fd),
	.w8(32'hb728595d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378d1a31),
	.w1(32'hba30add3),
	.w2(32'hb90f77f1),
	.w3(32'h389bceaa),
	.w4(32'hba24c6c6),
	.w5(32'hb8f13406),
	.w6(32'hb9fc231c),
	.w7(32'h38be8f51),
	.w8(32'hba5d64fc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e563f),
	.w1(32'hbabd5418),
	.w2(32'hbabf1ee8),
	.w3(32'hba6239d2),
	.w4(32'hba6f235f),
	.w5(32'hba53b4ea),
	.w6(32'hba9b80c1),
	.w7(32'hbacd7527),
	.w8(32'hb93dc0a6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f9d6d),
	.w1(32'hb9b47c3b),
	.w2(32'hb9a9021c),
	.w3(32'h385db0fc),
	.w4(32'hb994310a),
	.w5(32'hb9ce6807),
	.w6(32'hb9d32876),
	.w7(32'hb9906aec),
	.w8(32'h3a1153e3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af16c3),
	.w1(32'h377456a0),
	.w2(32'h39abff12),
	.w3(32'h39af00e1),
	.w4(32'h39801914),
	.w5(32'h39919e87),
	.w6(32'h3a62d316),
	.w7(32'h3ad5cf83),
	.w8(32'hb9d16119),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f03b52),
	.w1(32'hb9b4e251),
	.w2(32'hb9b6839f),
	.w3(32'hb9ed6efd),
	.w4(32'hba33826e),
	.w5(32'hba166d8c),
	.w6(32'hb8c0787f),
	.w7(32'hb90b6169),
	.w8(32'h396de436),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9818f47),
	.w1(32'hb9860f43),
	.w2(32'h38d7aec9),
	.w3(32'hba01a739),
	.w4(32'hb99f5c63),
	.w5(32'h37095b05),
	.w6(32'h38d21dcb),
	.w7(32'h39eab737),
	.w8(32'hb9633be5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7114279),
	.w1(32'hbb172b54),
	.w2(32'hbb5b63f2),
	.w3(32'hb98ff9ce),
	.w4(32'h38ef74bf),
	.w5(32'hbab25aba),
	.w6(32'hbb1f7055),
	.w7(32'hbb580277),
	.w8(32'hba4acd17),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5effa),
	.w1(32'hbb8b91b8),
	.w2(32'hbb074725),
	.w3(32'hbc29e69d),
	.w4(32'hbc07db44),
	.w5(32'h3ab66cfa),
	.w6(32'hbaa4a258),
	.w7(32'hbc1af04b),
	.w8(32'hba9b0b7f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab52350),
	.w1(32'hbb2c2dd7),
	.w2(32'hbbcb70c0),
	.w3(32'h3b93a1a0),
	.w4(32'h3b397c09),
	.w5(32'hba77a98b),
	.w6(32'hbbc00b66),
	.w7(32'hbbec4bf0),
	.w8(32'hbb172e2f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b9316),
	.w1(32'hbb059d2d),
	.w2(32'hbb984b64),
	.w3(32'h3b126011),
	.w4(32'h3ae26a08),
	.w5(32'hbaaa1678),
	.w6(32'hbbb7b4e5),
	.w7(32'hbbd3acc0),
	.w8(32'h3ae41cdf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08a44d),
	.w1(32'hbaadee99),
	.w2(32'hbb0919e4),
	.w3(32'hbba76e59),
	.w4(32'hbb9f3ef3),
	.w5(32'hb9edf7d7),
	.w6(32'hb93285b4),
	.w7(32'hba52d7fc),
	.w8(32'hbb696221),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fedd2),
	.w1(32'h3be49513),
	.w2(32'h3b50c610),
	.w3(32'hbb8946a4),
	.w4(32'h3b895f32),
	.w5(32'h3bcc4eec),
	.w6(32'hbbbe6bd8),
	.w7(32'hbb241a30),
	.w8(32'hbbb6ea76),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc560f9a),
	.w1(32'hbb27b0a5),
	.w2(32'h3bf82958),
	.w3(32'hbc3410a9),
	.w4(32'hbba8b8e8),
	.w5(32'h3b8fec12),
	.w6(32'h3ac236cb),
	.w7(32'h3b510056),
	.w8(32'hbb1d7256),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8340e8),
	.w1(32'h3a8996e9),
	.w2(32'h3c9138b5),
	.w3(32'hbcd1c85a),
	.w4(32'hbc8391f3),
	.w5(32'hb51fcc88),
	.w6(32'h3c8a537a),
	.w7(32'h3cf1a09e),
	.w8(32'hbaeb5069),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d1c37),
	.w1(32'hbae00582),
	.w2(32'hbb92544e),
	.w3(32'h39337a6a),
	.w4(32'h3a097932),
	.w5(32'hba982b4d),
	.w6(32'hbb8a17b2),
	.w7(32'hbbc08a4b),
	.w8(32'h39559e01),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b069f20),
	.w1(32'hba8adc12),
	.w2(32'hbb86bbcd),
	.w3(32'h3b7e5044),
	.w4(32'h3b0effa0),
	.w5(32'hba16f739),
	.w6(32'hbb6758e7),
	.w7(32'hbba35d61),
	.w8(32'h3a328da0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ac7b),
	.w1(32'hbb795845),
	.w2(32'hbc18ae22),
	.w3(32'h3c093b49),
	.w4(32'h3b883849),
	.w5(32'hbaf45e3b),
	.w6(32'hbc0ff57f),
	.w7(32'hbc3c3bbb),
	.w8(32'hbc221e1a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7989f1),
	.w1(32'hbc3f6b7a),
	.w2(32'hbc8387f4),
	.w3(32'hba609c31),
	.w4(32'hbba62686),
	.w5(32'hbbe8d7c4),
	.w6(32'hbca9cece),
	.w7(32'hbc81a353),
	.w8(32'hbbd862b2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72c67b),
	.w1(32'h3a8a321e),
	.w2(32'h3c506894),
	.w3(32'hbcaa6f06),
	.w4(32'hbc1fc144),
	.w5(32'h3a9b4a58),
	.w6(32'h3c25ab77),
	.w7(32'h3cb2b8eb),
	.w8(32'hbb6356f7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a02593),
	.w1(32'h3af23e64),
	.w2(32'h3c37e269),
	.w3(32'hbc1877bb),
	.w4(32'h3ba796e0),
	.w5(32'h3c62aa82),
	.w6(32'hbb596565),
	.w7(32'hbb9f4351),
	.w8(32'h3b269cba),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc84bc8),
	.w1(32'h3bee7298),
	.w2(32'hba4ddc56),
	.w3(32'hba81ac8b),
	.w4(32'h3c286416),
	.w5(32'h3b57c0a1),
	.w6(32'h3a776807),
	.w7(32'hbae99e07),
	.w8(32'hbb3bffef),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fad68),
	.w1(32'h3b065431),
	.w2(32'hbb9eab7b),
	.w3(32'hbb3d0b22),
	.w4(32'hbb43447e),
	.w5(32'hbb661e3d),
	.w6(32'hb9718010),
	.w7(32'hbb9bdec4),
	.w8(32'h3c103637),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba72f07),
	.w1(32'hba60eca8),
	.w2(32'h3c236a00),
	.w3(32'hbc1e51e7),
	.w4(32'h39007e30),
	.w5(32'h3bdfed88),
	.w6(32'h3c468ff2),
	.w7(32'h3b916b79),
	.w8(32'h3b0dfe9d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e85fb),
	.w1(32'h3a4184f5),
	.w2(32'hbb8c5da9),
	.w3(32'h3bb8fdda),
	.w4(32'h3b03b52c),
	.w5(32'hbb3b76df),
	.w6(32'hbacdaf87),
	.w7(32'hbb9a4696),
	.w8(32'h3a0628f7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05bad0),
	.w1(32'hbba57df2),
	.w2(32'hbaba5a9b),
	.w3(32'hbb98f974),
	.w4(32'hbba2a6ae),
	.w5(32'hba9536e2),
	.w6(32'hbb1663ee),
	.w7(32'h3a5e73b6),
	.w8(32'h3a790ed4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb22373),
	.w1(32'h3be993dd),
	.w2(32'hbb50265a),
	.w3(32'hbaf1a5ed),
	.w4(32'hbb72cc4b),
	.w5(32'h3a178ca9),
	.w6(32'h3ada79b1),
	.w7(32'h3a28c719),
	.w8(32'h3ba17a49),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb415642),
	.w1(32'hba0caa66),
	.w2(32'h39f80289),
	.w3(32'hbbd1ed8c),
	.w4(32'hbb5b5eda),
	.w5(32'h3adc1870),
	.w6(32'h3b8bd14c),
	.w7(32'h3a925d7c),
	.w8(32'hbb36db65),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70b891),
	.w1(32'h3adb3fd7),
	.w2(32'hbbd638a7),
	.w3(32'h3bc79018),
	.w4(32'h3b80ca7a),
	.w5(32'hbb57b64d),
	.w6(32'hbbb37f5a),
	.w7(32'hbc21628d),
	.w8(32'h3bd2cdaf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d20f6),
	.w1(32'hb85c2ad2),
	.w2(32'hbb45e72f),
	.w3(32'hbae165e1),
	.w4(32'hbab56889),
	.w5(32'hb971c6fa),
	.w6(32'h3bc3066d),
	.w7(32'h3be821ba),
	.w8(32'hbb4432c4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86b85b),
	.w1(32'hbaea57e2),
	.w2(32'hbb77b02d),
	.w3(32'h3a959450),
	.w4(32'h3a28abe2),
	.w5(32'hbaa9a38f),
	.w6(32'hbb87f4f8),
	.w7(32'hbb92b5f9),
	.w8(32'h3a5ac1fe),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2af0f9),
	.w1(32'hb9fb922f),
	.w2(32'hbb17bcc9),
	.w3(32'h3b84c1b3),
	.w4(32'h3b22d572),
	.w5(32'h390f754b),
	.w6(32'hbb51ef5c),
	.w7(32'hbb6a33e7),
	.w8(32'hb8a77202),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a583d16),
	.w1(32'hbac3e259),
	.w2(32'hbb5194e0),
	.w3(32'h3b148aef),
	.w4(32'h3a839e69),
	.w5(32'hba4e4d16),
	.w6(32'hbb36cb36),
	.w7(32'hbb5eb6d8),
	.w8(32'h3aadc42f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6002cb),
	.w1(32'h3998700a),
	.w2(32'hbb3ca9ed),
	.w3(32'hbbc9331b),
	.w4(32'hbbe979ae),
	.w5(32'hbbf0be2d),
	.w6(32'hba945e08),
	.w7(32'h3af7d288),
	.w8(32'hbaf1e704),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10a892),
	.w1(32'hbb0d09c1),
	.w2(32'hbb86adaf),
	.w3(32'h38a0f3b6),
	.w4(32'h39315d78),
	.w5(32'hbaae43b2),
	.w6(32'hbb89c8d4),
	.w7(32'hbba45e2f),
	.w8(32'h3bca79df),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6b419),
	.w1(32'h3a0da002),
	.w2(32'hbcd5676a),
	.w3(32'h3d16341b),
	.w4(32'h3cac352e),
	.w5(32'hbb8b2fab),
	.w6(32'hbca91469),
	.w7(32'hbd2340fb),
	.w8(32'hba930fbb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efe574),
	.w1(32'hbb3b7bd4),
	.w2(32'hbb82a527),
	.w3(32'h3a883d41),
	.w4(32'h3943d958),
	.w5(32'hbaf5f833),
	.w6(32'hbb5fa7eb),
	.w7(32'hbb70e261),
	.w8(32'hbb1468e6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf512b0),
	.w1(32'hbb636ac8),
	.w2(32'hbb92903a),
	.w3(32'hbb1b1aa6),
	.w4(32'hbad9738a),
	.w5(32'hbad6607a),
	.w6(32'hbb8fef53),
	.w7(32'hbbb4f6e5),
	.w8(32'hba2a89cc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8140c7),
	.w1(32'hbb4d5b7a),
	.w2(32'hbb725725),
	.w3(32'h3b3268d6),
	.w4(32'h3a9e06ec),
	.w5(32'hba234bc6),
	.w6(32'hbbaff4db),
	.w7(32'hbb943633),
	.w8(32'hb9d5fd8a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf23f5b),
	.w1(32'hbbee57b3),
	.w2(32'hbc1606b1),
	.w3(32'hbc6be68a),
	.w4(32'hbc4af6ef),
	.w5(32'hbc190db1),
	.w6(32'hbbab37d3),
	.w7(32'hbc019923),
	.w8(32'hbb078e0c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43acb6),
	.w1(32'hbbb4d509),
	.w2(32'hbba981d0),
	.w3(32'hbb502173),
	.w4(32'hbb5be7f0),
	.w5(32'hbb20cf3e),
	.w6(32'hbba75397),
	.w7(32'hbba9d7a3),
	.w8(32'hba47c39e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a154909),
	.w1(32'hbb068872),
	.w2(32'hbb98124e),
	.w3(32'h3b2fc73e),
	.w4(32'h3ad871de),
	.w5(32'hbaa7101f),
	.w6(32'hbb734828),
	.w7(32'hbb9cfab0),
	.w8(32'hba90dd44),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8c7a0),
	.w1(32'hbb6ca37e),
	.w2(32'hbb86306a),
	.w3(32'hba994a51),
	.w4(32'hba938aa1),
	.w5(32'hbafefb76),
	.w6(32'hbb7506ec),
	.w7(32'hbb81cc4c),
	.w8(32'h3be8424f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc9023),
	.w1(32'h3a08488b),
	.w2(32'hbcef3cd0),
	.w3(32'h3d26e1b8),
	.w4(32'h3cbc8e04),
	.w5(32'hbbad35e9),
	.w6(32'hbcb90ec6),
	.w7(32'hbd35a2b4),
	.w8(32'h3b0794d7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52f79e),
	.w1(32'h3a3a1413),
	.w2(32'hbc6da2d0),
	.w3(32'h3ca75b63),
	.w4(32'h3c4cd6fd),
	.w5(32'hbb159433),
	.w6(32'hbc4bc40d),
	.w7(32'hbcc61eea),
	.w8(32'hba59cdcf),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7762ef),
	.w1(32'hbb0b8da3),
	.w2(32'hbaee126a),
	.w3(32'h3a833fe9),
	.w4(32'h3a591083),
	.w5(32'hb8fa6be3),
	.w6(32'hbb658cf2),
	.w7(32'hbb5623e9),
	.w8(32'hb7ac61b1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5544eb),
	.w1(32'hbbbdb282),
	.w2(32'hbc85b499),
	.w3(32'hbb633254),
	.w4(32'hbb90f4fa),
	.w5(32'hbbdc1398),
	.w6(32'hbb71d720),
	.w7(32'hb94d77c5),
	.w8(32'h3987e5db),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e22d1),
	.w1(32'hbb255670),
	.w2(32'hbb1d3d12),
	.w3(32'hba8b8e95),
	.w4(32'hb9db4fd3),
	.w5(32'h3986f77d),
	.w6(32'hba9f2402),
	.w7(32'hbab0fbd3),
	.w8(32'hbb2fcc17),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52922),
	.w1(32'hbbd15de7),
	.w2(32'hbb9a909b),
	.w3(32'hbbba87ae),
	.w4(32'hbb51dd73),
	.w5(32'h39d4e52e),
	.w6(32'hbbd33d4a),
	.w7(32'hbbd02363),
	.w8(32'h3be01d20),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe6f9b),
	.w1(32'h3bb87e75),
	.w2(32'h3b81920b),
	.w3(32'h3bc2f5b3),
	.w4(32'h3c2b749e),
	.w5(32'h3c29a6af),
	.w6(32'h39e674bb),
	.w7(32'hbbe7a823),
	.w8(32'hbb785355),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc526bb0),
	.w1(32'hba43b654),
	.w2(32'h3c00a641),
	.w3(32'hbca04428),
	.w4(32'hbc31ace1),
	.w5(32'hbb148c38),
	.w6(32'h3bf04ce6),
	.w7(32'h3c63f28b),
	.w8(32'hbac3f0fc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2404e),
	.w1(32'hba3370f1),
	.w2(32'hbba125a6),
	.w3(32'h3b3674e2),
	.w4(32'h3b073b90),
	.w5(32'hbb0ce9f5),
	.w6(32'hbba662f1),
	.w7(32'hbbee2213),
	.w8(32'hbb393e71),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadd464),
	.w1(32'h3ab3448c),
	.w2(32'h3cc025f3),
	.w3(32'hbd0ad448),
	.w4(32'hbcae333a),
	.w5(32'h35dc6ac9),
	.w6(32'h3cb73ef6),
	.w7(32'h3d1fedbe),
	.w8(32'hbb996286),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86d527),
	.w1(32'hbaf24eee),
	.w2(32'hbad0b0c4),
	.w3(32'hbb013b3c),
	.w4(32'h396d3bcf),
	.w5(32'h3a521022),
	.w6(32'hbb9bdbf9),
	.w7(32'hbaed36e5),
	.w8(32'h3b026aff),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaadf60),
	.w1(32'hbbd59ab8),
	.w2(32'h3abbf76b),
	.w3(32'hbc139a00),
	.w4(32'hbc365606),
	.w5(32'hbab16387),
	.w6(32'h3b2e1966),
	.w7(32'h3bd30358),
	.w8(32'hbb37d596),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca25730),
	.w1(32'h3aa9b93d),
	.w2(32'h3cb44321),
	.w3(32'hbd01d88a),
	.w4(32'hbca305a1),
	.w5(32'h37bb6897),
	.w6(32'h3cab1203),
	.w7(32'h3d15a8bc),
	.w8(32'hbb186298),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ac7a1),
	.w1(32'h3a93c1da),
	.w2(32'h3c9a0a25),
	.w3(32'hbcdddaa1),
	.w4(32'hbc8b2d95),
	.w5(32'h37ba53d1),
	.w6(32'h3c9305fd),
	.w7(32'h3d002522),
	.w8(32'hbb621fcd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5011bf),
	.w1(32'h39259280),
	.w2(32'h3c4a9f0f),
	.w3(32'hbc91d0c6),
	.w4(32'hbc10b897),
	.w5(32'h3b0081a2),
	.w6(32'h3c1ce910),
	.w7(32'h3ca12aac),
	.w8(32'hbc91f57f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b378b),
	.w1(32'hbbfdaa71),
	.w2(32'hbafc79c4),
	.w3(32'hbc50546b),
	.w4(32'hbc1b4dda),
	.w5(32'hbb5a8f99),
	.w6(32'hbc5802de),
	.w7(32'hbc17fbb4),
	.w8(32'h39ccbd9b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9e43b),
	.w1(32'hba6af7eb),
	.w2(32'hbb582d02),
	.w3(32'h3b52fa8c),
	.w4(32'h3b01d6d1),
	.w5(32'hb9ffc774),
	.w6(32'hbb2359b6),
	.w7(32'hbb758be3),
	.w8(32'h3c608c9c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0365b5),
	.w1(32'hb9f97812),
	.w2(32'hbbaaa704),
	.w3(32'hbbd4bf24),
	.w4(32'h3c123a61),
	.w5(32'h3c13d422),
	.w6(32'h3c331b5e),
	.w7(32'h3a767708),
	.w8(32'hbc1d4cab),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb76e09),
	.w1(32'hbc00cad5),
	.w2(32'h3b9ef029),
	.w3(32'hbd000dd4),
	.w4(32'hbcaecbbd),
	.w5(32'hbc0d2724),
	.w6(32'h3bca7f2c),
	.w7(32'h3c8797ec),
	.w8(32'h3bac6d5e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2a604),
	.w1(32'h3af0a061),
	.w2(32'hb99b43ed),
	.w3(32'hbb39cc5c),
	.w4(32'h3ad3bc14),
	.w5(32'h3b5b1885),
	.w6(32'h3bc8e6b2),
	.w7(32'h3bb423e6),
	.w8(32'hbb5cd12b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc99605),
	.w1(32'h3a1e8653),
	.w2(32'h3b396f3a),
	.w3(32'hba8f31c6),
	.w4(32'h3b7746fe),
	.w5(32'hb99dd261),
	.w6(32'hba1e16eb),
	.w7(32'h3a671846),
	.w8(32'h3bcb6e27),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc11a50),
	.w1(32'h39dd7f04),
	.w2(32'hbcd20adf),
	.w3(32'h3d12896d),
	.w4(32'h3ca59909),
	.w5(32'hbb96b1fa),
	.w6(32'hbca23bb4),
	.w7(32'hbd1f5b66),
	.w8(32'hbb2b8478),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79196),
	.w1(32'hbb16e99f),
	.w2(32'hbb0ea76b),
	.w3(32'hb91683cd),
	.w4(32'h3ab8e658),
	.w5(32'h3a9b4e39),
	.w6(32'hbbc0a72a),
	.w7(32'hbb86640f),
	.w8(32'hbb342331),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde9eea),
	.w1(32'hbba13732),
	.w2(32'h3b50b5cc),
	.w3(32'hbc79a085),
	.w4(32'hbc159c5e),
	.w5(32'hbac33eb7),
	.w6(32'h3afe01c5),
	.w7(32'h3c29a9cd),
	.w8(32'h38b9c08c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb53b5),
	.w1(32'hbab2d651),
	.w2(32'hbb987d77),
	.w3(32'h3b799bc4),
	.w4(32'h3ae79cad),
	.w5(32'hba888457),
	.w6(32'hbb7f61e5),
	.w7(32'hbbb0976f),
	.w8(32'h3b15e40b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca84752),
	.w1(32'h3b135ed8),
	.w2(32'hbcba25b5),
	.w3(32'h3cfed8b3),
	.w4(32'h3ca79a3f),
	.w5(32'hbb89deed),
	.w6(32'hbc9f86d4),
	.w7(32'hbd2129b0),
	.w8(32'hbba86bda),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74c13e),
	.w1(32'hbb759888),
	.w2(32'h3c0e2b1e),
	.w3(32'hbca8bfac),
	.w4(32'hbc4ece5d),
	.w5(32'hba65f3fc),
	.w6(32'h3be41a2b),
	.w7(32'h3c8495f0),
	.w8(32'hbab610ae),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08f220),
	.w1(32'h39f06bb4),
	.w2(32'h3c171544),
	.w3(32'hbc59ceec),
	.w4(32'hbc06f9ff),
	.w5(32'h39380bf0),
	.w6(32'h3c0e679d),
	.w7(32'h3c7afbef),
	.w8(32'hbafc45c2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb325559),
	.w1(32'hbb088f46),
	.w2(32'hb9d0dfdd),
	.w3(32'hbb618b72),
	.w4(32'hbb1667af),
	.w5(32'hb85cb39b),
	.w6(32'hbaa35da0),
	.w7(32'h3a3b7ad9),
	.w8(32'hbb43af1e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c5e8),
	.w1(32'h391a77e9),
	.w2(32'hb93a4077),
	.w3(32'h3ac8d490),
	.w4(32'h3b175cd8),
	.w5(32'hba8c6d5c),
	.w6(32'h3a6488cc),
	.w7(32'h3b8f506a),
	.w8(32'hbba9ea4e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f010d),
	.w1(32'hbb433216),
	.w2(32'hbb1658e8),
	.w3(32'hbb9d5083),
	.w4(32'hbb2536bf),
	.w5(32'hba188b09),
	.w6(32'hbb6d4587),
	.w7(32'hbb6aeab2),
	.w8(32'h3bbf76a5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f81c),
	.w1(32'h3b94a26c),
	.w2(32'h3b8d3f31),
	.w3(32'h3b91e36c),
	.w4(32'h3b8a1b83),
	.w5(32'h3bbbc1fc),
	.w6(32'h3b91aab9),
	.w7(32'h3b6c217a),
	.w8(32'hbae99f9e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07170c),
	.w1(32'hbbee6adb),
	.w2(32'hbb7e2597),
	.w3(32'h3a1c3fec),
	.w4(32'hbb561e45),
	.w5(32'hbb256be8),
	.w6(32'hbb5fde30),
	.w7(32'h3a1fa875),
	.w8(32'hbaf4e7a3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11d225),
	.w1(32'hba7b5f06),
	.w2(32'h3a68d6bd),
	.w3(32'h39d361fb),
	.w4(32'hbb20c1aa),
	.w5(32'h3b22c3ac),
	.w6(32'hb9aa6fe6),
	.w7(32'h3bccdc37),
	.w8(32'h39c5ae90),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecb20e),
	.w1(32'hbb950050),
	.w2(32'hbb747d11),
	.w3(32'h3b4f363e),
	.w4(32'hbb23afac),
	.w5(32'hbaea0c69),
	.w6(32'hbb0668e5),
	.w7(32'hba74874a),
	.w8(32'h3ca86d28),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e1eb8),
	.w1(32'h3c28e901),
	.w2(32'h3c70cdbc),
	.w3(32'h3c921ee0),
	.w4(32'h3c4c2fae),
	.w5(32'h3c6676d6),
	.w6(32'h3c693821),
	.w7(32'h3c9965dc),
	.w8(32'h3b3ab267),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25179f),
	.w1(32'h39b9b342),
	.w2(32'h39f18a02),
	.w3(32'h3a83bc1c),
	.w4(32'h39805f7a),
	.w5(32'h3abbb2b4),
	.w6(32'h3a94edc5),
	.w7(32'h3982cb40),
	.w8(32'hba9e7248),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c26e9),
	.w1(32'hbab24a43),
	.w2(32'hbaab9836),
	.w3(32'hbaaab268),
	.w4(32'hba7fd468),
	.w5(32'hba07156b),
	.w6(32'hbaa14e33),
	.w7(32'hbac492dd),
	.w8(32'hbb567165),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37cfc2),
	.w1(32'hbb14252b),
	.w2(32'hbb1a8b55),
	.w3(32'hbb77687f),
	.w4(32'hbb1c55f6),
	.w5(32'hba8ec61f),
	.w6(32'hbb367646),
	.w7(32'hbb6228b8),
	.w8(32'hbbad3e92),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcae7c5),
	.w1(32'h3b435afd),
	.w2(32'hba055ce4),
	.w3(32'hbbaed360),
	.w4(32'h3b0393bd),
	.w5(32'hbb14fd1e),
	.w6(32'h3aab38a7),
	.w7(32'h3b851857),
	.w8(32'h3c40d5ad),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c595425),
	.w1(32'h3ca3c310),
	.w2(32'h3c8f0aa9),
	.w3(32'h3c5c3037),
	.w4(32'h3c98bb96),
	.w5(32'h3c6d7239),
	.w6(32'h3c9141a5),
	.w7(32'h3c843c81),
	.w8(32'h3c12ac95),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f1197),
	.w1(32'hbb80f2f5),
	.w2(32'h3a2d8f95),
	.w3(32'h3a447cf6),
	.w4(32'hbbb3452e),
	.w5(32'h3aa331d2),
	.w6(32'hb6b245a4),
	.w7(32'h3b8d24be),
	.w8(32'hbbfba7fa),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf03ae7),
	.w1(32'hbbb28f11),
	.w2(32'hbb42d497),
	.w3(32'hbb6a619d),
	.w4(32'hb98d1f48),
	.w5(32'hbb3fab62),
	.w6(32'hbbfa65b2),
	.w7(32'hbb7d4940),
	.w8(32'hbb4197fb),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09748a),
	.w1(32'hbba7e2bf),
	.w2(32'hba03c2c4),
	.w3(32'hbbd6994b),
	.w4(32'hbba2331b),
	.w5(32'hbb39f9c1),
	.w6(32'hbb732099),
	.w7(32'h3abf3a9e),
	.w8(32'h3b84f8c0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0e4b1),
	.w1(32'hbb84d4c6),
	.w2(32'hbaa69fe7),
	.w3(32'hbabe0a8b),
	.w4(32'hbbd439cd),
	.w5(32'hb993ddaa),
	.w6(32'hba8a8d54),
	.w7(32'h3adaec7e),
	.w8(32'h3c431509),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1641dc),
	.w1(32'hbb9b5c54),
	.w2(32'hbaa9d3eb),
	.w3(32'h3b90b451),
	.w4(32'hbb4e9381),
	.w5(32'h38982fff),
	.w6(32'h3a92b99a),
	.w7(32'h3b841033),
	.w8(32'hbc81d34c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca23fc),
	.w1(32'hbd112fe0),
	.w2(32'hbcb0ca75),
	.w3(32'hbc807e75),
	.w4(32'hbce0a1be),
	.w5(32'hbc90b6e3),
	.w6(32'hbcc55fed),
	.w7(32'hbc1082c2),
	.w8(32'h3b7d1c5f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae4fcf),
	.w1(32'hbb81a4d4),
	.w2(32'hba211022),
	.w3(32'hbb97c4d0),
	.w4(32'hbb018f58),
	.w5(32'hbbd2bd56),
	.w6(32'h3a4cb93e),
	.w7(32'h3b7d363f),
	.w8(32'hbb958808),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77f87),
	.w1(32'hbbf002f3),
	.w2(32'hbb8c6a81),
	.w3(32'hbb31769d),
	.w4(32'hbaa5ba96),
	.w5(32'hb8159d5a),
	.w6(32'hbba85077),
	.w7(32'hbad890d6),
	.w8(32'h3bd9b5d9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3e91b),
	.w1(32'h3af456d2),
	.w2(32'h39ea9c15),
	.w3(32'h3ba030f2),
	.w4(32'h3af1b771),
	.w5(32'h3ab36654),
	.w6(32'h3b307ca2),
	.w7(32'h389c2b50),
	.w8(32'h39a231cb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda0cbc),
	.w1(32'h3bbcb43f),
	.w2(32'hba714eae),
	.w3(32'h3b1b398c),
	.w4(32'hbba2ecd0),
	.w5(32'hbb9eb3e7),
	.w6(32'hba4b637b),
	.w7(32'hbaa474b4),
	.w8(32'hbb75b2d0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule