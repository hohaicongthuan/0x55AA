module layer_8_featuremap_255(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8e3c0),
	.w1(32'h3c7b144f),
	.w2(32'h3bd7c93d),
	.w3(32'hbba01d3c),
	.w4(32'h3c2e53b5),
	.w5(32'h3bf3754e),
	.w6(32'hbaf1ab14),
	.w7(32'h3abeb10c),
	.w8(32'hbab29d17),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e0d3a),
	.w1(32'hbcb43aaa),
	.w2(32'hbc884deb),
	.w3(32'h3aa86c16),
	.w4(32'hbd5f58a1),
	.w5(32'hbdd97ec8),
	.w6(32'h3cf03fdf),
	.w7(32'h3db7def0),
	.w8(32'h3d8b4476),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb58079),
	.w1(32'hb916924d),
	.w2(32'hbb01945d),
	.w3(32'hbd6c9b2b),
	.w4(32'hbb129452),
	.w5(32'hbbc89cbf),
	.w6(32'h3a4ae13b),
	.w7(32'hbbe7e7c4),
	.w8(32'hbc304c06),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc2a6a),
	.w1(32'hbc1946fc),
	.w2(32'hbc85bebd),
	.w3(32'hbba5cad0),
	.w4(32'hbafa2e0c),
	.w5(32'hbc0786a4),
	.w6(32'hbb9a67dd),
	.w7(32'hbc0eea3b),
	.w8(32'hbb8ba682),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb350a0),
	.w1(32'h3b840328),
	.w2(32'h39964118),
	.w3(32'hbb84cd8c),
	.w4(32'hbd8136eb),
	.w5(32'hbe114c89),
	.w6(32'h3d8842eb),
	.w7(32'h3e0db6e3),
	.w8(32'h3dbfe82f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21bc97),
	.w1(32'h3b98f747),
	.w2(32'h3ba1c2cd),
	.w3(32'hbda19abe),
	.w4(32'h3c5fb945),
	.w5(32'h3c767b9f),
	.w6(32'h3b464ca3),
	.w7(32'hbb0e96e2),
	.w8(32'h3c4d3889),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3f605),
	.w1(32'h3c1a7261),
	.w2(32'h3bbaa40d),
	.w3(32'hba960a00),
	.w4(32'h3cd1b7e2),
	.w5(32'h3d68a44a),
	.w6(32'hbcb584fc),
	.w7(32'hbd55b3df),
	.w8(32'hbd1df670),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaafc38),
	.w1(32'h3c235fa1),
	.w2(32'h3c2bee5f),
	.w3(32'h3d246ec6),
	.w4(32'h3c46519c),
	.w5(32'h3c36fea3),
	.w6(32'h3c2f6202),
	.w7(32'h3c9814bc),
	.w8(32'h3c503a83),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cd9e6),
	.w1(32'hbba0e23d),
	.w2(32'hbc1b5b53),
	.w3(32'hb8971ef3),
	.w4(32'hbd5823b2),
	.w5(32'hbe00b0e5),
	.w6(32'h3d7c1efa),
	.w7(32'h3e06cd26),
	.w8(32'h3da8e6ab),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c862444),
	.w1(32'hb9acde95),
	.w2(32'h3c1f49b0),
	.w3(32'hbd767eba),
	.w4(32'hbb30d325),
	.w5(32'h3c1155d8),
	.w6(32'hba8138e5),
	.w7(32'hba9ceca9),
	.w8(32'hbb9b375c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c685fde),
	.w1(32'h3c08ccab),
	.w2(32'hbad4d4c7),
	.w3(32'h3be98441),
	.w4(32'h3be8e5dd),
	.w5(32'h3b350b4d),
	.w6(32'hbb69d992),
	.w7(32'h3a162078),
	.w8(32'hbc371151),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c7ba),
	.w1(32'h3c041465),
	.w2(32'h3b3dfe2a),
	.w3(32'hbba69968),
	.w4(32'h3c3c3d9d),
	.w5(32'h3c183e51),
	.w6(32'hbb7a5738),
	.w7(32'hbb4f53b0),
	.w8(32'h3b750332),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904ad8e),
	.w1(32'hbc42e9aa),
	.w2(32'hbc5cc45a),
	.w3(32'h3c09e7a4),
	.w4(32'hbbf80a76),
	.w5(32'hbbaa5c43),
	.w6(32'hbc272ee3),
	.w7(32'hbb98402f),
	.w8(32'hb94f7747),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb194cf2),
	.w1(32'hbb80f04d),
	.w2(32'hbb25cd9d),
	.w3(32'hbbd3cf60),
	.w4(32'h3b41d736),
	.w5(32'hbbd313ad),
	.w6(32'h3b9ff038),
	.w7(32'hbac332dc),
	.w8(32'h39c90d24),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76c74e),
	.w1(32'hba085ab7),
	.w2(32'h3b8139f7),
	.w3(32'hba86fbf1),
	.w4(32'h3d36590f),
	.w5(32'h3dccf94c),
	.w6(32'hbd46e637),
	.w7(32'hbdc185ec),
	.w8(32'hbd7aad34),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3824d0),
	.w1(32'h3b04afc2),
	.w2(32'h3c151827),
	.w3(32'h3d49367a),
	.w4(32'h3bd90f2f),
	.w5(32'h3b625e32),
	.w6(32'h3b5633dc),
	.w7(32'h3c166bba),
	.w8(32'h3be2fa70),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c672ef1),
	.w1(32'h3b1e639d),
	.w2(32'h3b912102),
	.w3(32'h3afa4a2a),
	.w4(32'hbab24ad0),
	.w5(32'h3b1d6e1a),
	.w6(32'hbb7e692f),
	.w7(32'hbad652b5),
	.w8(32'h3a7221c4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd3c9c),
	.w1(32'h3adf329c),
	.w2(32'hbbb9501d),
	.w3(32'h3ab4354c),
	.w4(32'h3ba7ac03),
	.w5(32'h3aa8386b),
	.w6(32'h3ad279a7),
	.w7(32'hbb99f757),
	.w8(32'hbbacfee3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e9bfc),
	.w1(32'h3c877338),
	.w2(32'hbbdbe83e),
	.w3(32'hbad093c0),
	.w4(32'h3c9b2a0d),
	.w5(32'h3c032f01),
	.w6(32'hbcb6a89f),
	.w7(32'hbc6b4029),
	.w8(32'hbca062a2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce56d37),
	.w1(32'h3d1fe616),
	.w2(32'h3cca4b68),
	.w3(32'h3c269284),
	.w4(32'h3d893f28),
	.w5(32'h3e0088b6),
	.w6(32'hbd33a085),
	.w7(32'hbddf4033),
	.w8(32'hbdb466be),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0762fe),
	.w1(32'hb8623df5),
	.w2(32'h3bb9eb7b),
	.w3(32'h3d7dae22),
	.w4(32'hba36fe04),
	.w5(32'h3ba09eef),
	.w6(32'hbaf57cb4),
	.w7(32'hbab937da),
	.w8(32'h3ba55ea9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901ef4),
	.w1(32'hbb73f63e),
	.w2(32'hbc3af32d),
	.w3(32'hbbc5d807),
	.w4(32'hbba9f060),
	.w5(32'hbbc29c0f),
	.w6(32'hbbafbb3d),
	.w7(32'h3b56ed63),
	.w8(32'hbb2b5a1b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc459a2),
	.w1(32'h3d127f47),
	.w2(32'h3c90d694),
	.w3(32'h3c3a82a1),
	.w4(32'h3c8c88bc),
	.w5(32'h3bd744d9),
	.w6(32'hb9e106ff),
	.w7(32'h3b8f6044),
	.w8(32'hbbc23af6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21473c),
	.w1(32'h3c3df0c7),
	.w2(32'h3c503c57),
	.w3(32'h3ba7c933),
	.w4(32'h3c18d634),
	.w5(32'h3acf590c),
	.w6(32'h3abd2040),
	.w7(32'h3c1ecdba),
	.w8(32'hba96313f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe79c3b),
	.w1(32'hbaa99bf8),
	.w2(32'hbce5d27d),
	.w3(32'h3b9135fa),
	.w4(32'h3b5b5427),
	.w5(32'h3b20d14d),
	.w6(32'hb8f80a3c),
	.w7(32'hbbf5990f),
	.w8(32'hbbd95061),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb421888),
	.w1(32'h3c76520a),
	.w2(32'h3b4f6f45),
	.w3(32'h3c35a981),
	.w4(32'h3c803b54),
	.w5(32'h3c1f3ed0),
	.w6(32'hbc436e1b),
	.w7(32'hbbac91e9),
	.w8(32'hbc2fdc50),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ed6e7),
	.w1(32'hba322b87),
	.w2(32'h3b4a1ef1),
	.w3(32'hbc153544),
	.w4(32'hbb1a9ab7),
	.w5(32'h3c026fd7),
	.w6(32'hb9c45b3e),
	.w7(32'hbc19fbfc),
	.w8(32'hbb834e7e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fcde4),
	.w1(32'h3d0a8014),
	.w2(32'h3d26da16),
	.w3(32'h3c228457),
	.w4(32'h3cdd6f79),
	.w5(32'h3cf4e020),
	.w6(32'hbd945cd3),
	.w7(32'hbd4dc767),
	.w8(32'hbd1683e5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc76449),
	.w1(32'h3b45a749),
	.w2(32'h38a2c68d),
	.w3(32'hbc0dd3fd),
	.w4(32'hbaf7c775),
	.w5(32'h3915fbbc),
	.w6(32'h3bd61c26),
	.w7(32'h3b94c68b),
	.w8(32'hbb0ec37d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26ef18),
	.w1(32'hbb05f93a),
	.w2(32'hbba7081b),
	.w3(32'hbb4bd578),
	.w4(32'h3c6c1c52),
	.w5(32'h3c1a4d20),
	.w6(32'h384410af),
	.w7(32'h3c075ad1),
	.w8(32'hbb4682b1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4016b2),
	.w1(32'hbc7516c0),
	.w2(32'hbcb30346),
	.w3(32'h3b77efda),
	.w4(32'hbc46f4a2),
	.w5(32'hbb068ccc),
	.w6(32'hbbe746c0),
	.w7(32'hbbdc0cea),
	.w8(32'hbb5e0fa8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71282b),
	.w1(32'h3a8a1965),
	.w2(32'h3c37d837),
	.w3(32'h3b06e90f),
	.w4(32'h3b7cbf2c),
	.w5(32'h3c244aaa),
	.w6(32'h3bbc27dc),
	.w7(32'h3c5b73fe),
	.w8(32'h3cb403ae),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e9058),
	.w1(32'hbab05ca6),
	.w2(32'h3b103b42),
	.w3(32'hbab5e038),
	.w4(32'h3af8e50c),
	.w5(32'h3bcb28cf),
	.w6(32'h3bb76ef2),
	.w7(32'hbb907716),
	.w8(32'h3c1df8fc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390700d6),
	.w1(32'h3b175573),
	.w2(32'h3bbfc90c),
	.w3(32'h3bf46aef),
	.w4(32'hbbf9c244),
	.w5(32'hba7d2ea5),
	.w6(32'h3b4fab2c),
	.w7(32'hba13a331),
	.w8(32'hba8b662b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25c7d0),
	.w1(32'hbafe5d41),
	.w2(32'hbb240f45),
	.w3(32'h3bc06056),
	.w4(32'h3b4bff7f),
	.w5(32'h3ba0c6d4),
	.w6(32'hba84b4f1),
	.w7(32'h3b23534c),
	.w8(32'hba763e29),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52f73d),
	.w1(32'hb7dbe1c4),
	.w2(32'hbb4101e1),
	.w3(32'h3c4e93c7),
	.w4(32'hbb2a9345),
	.w5(32'hbbf33101),
	.w6(32'hbb1ac7c2),
	.w7(32'hbbbefc18),
	.w8(32'hbb09f022),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60e142),
	.w1(32'hbc053244),
	.w2(32'hbc2c221f),
	.w3(32'h3a68e219),
	.w4(32'hbbf102aa),
	.w5(32'hbba91949),
	.w6(32'hbad1cb2f),
	.w7(32'hbb6cebaf),
	.w8(32'hbb261040),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e73e5),
	.w1(32'hbbd68ed1),
	.w2(32'hbae3e6d5),
	.w3(32'hbbcac13e),
	.w4(32'hbbcf0c25),
	.w5(32'hbc65b92e),
	.w6(32'h3bbdbd7d),
	.w7(32'h3cca9e86),
	.w8(32'h3cedaa97),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026023),
	.w1(32'hba29ee18),
	.w2(32'hbb40fb97),
	.w3(32'hbbf1bb63),
	.w4(32'h3ba450a1),
	.w5(32'h3c097001),
	.w6(32'h3bebd799),
	.w7(32'h3bcb02bc),
	.w8(32'h3af88cd1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2c4dc),
	.w1(32'hbb873036),
	.w2(32'hbb1716b1),
	.w3(32'h3b914d2f),
	.w4(32'hb9fd566c),
	.w5(32'h3abf18f0),
	.w6(32'h38ea4f64),
	.w7(32'h3aadb69c),
	.w8(32'hbb055ea5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ced6e),
	.w1(32'h3b9c1df9),
	.w2(32'h3bf9bcf7),
	.w3(32'hbc2f8e3b),
	.w4(32'h3be8367e),
	.w5(32'h3c6584f1),
	.w6(32'hbc216615),
	.w7(32'hbbaae8ed),
	.w8(32'hb9f9e644),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c3df3),
	.w1(32'h3a8985e9),
	.w2(32'h3bb78378),
	.w3(32'h3b65420a),
	.w4(32'hbb7bbc3a),
	.w5(32'h3c04f46f),
	.w6(32'hba52fcce),
	.w7(32'h3b5e1cbd),
	.w8(32'h3c1d47cb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e22ae),
	.w1(32'h3a907d0c),
	.w2(32'hbbff144d),
	.w3(32'h3c21e0dc),
	.w4(32'h3bf09e8d),
	.w5(32'h39213af4),
	.w6(32'hbb3514a6),
	.w7(32'hbbf9a11b),
	.w8(32'h3b7165b9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba724ca),
	.w1(32'h3b9fa199),
	.w2(32'h3b19e93b),
	.w3(32'h3b5d7506),
	.w4(32'h3b1cee61),
	.w5(32'h3b31c788),
	.w6(32'hba81bc8d),
	.w7(32'h3b768b32),
	.w8(32'h3b62f40a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc591de),
	.w1(32'h3b884743),
	.w2(32'hbb8377e4),
	.w3(32'h3a3e1b37),
	.w4(32'h3b47dceb),
	.w5(32'hbb6ec158),
	.w6(32'hbca1e10d),
	.w7(32'hbc004354),
	.w8(32'hbc607ad4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc058),
	.w1(32'h3ac5e484),
	.w2(32'h3b9c7796),
	.w3(32'h3b04d1d6),
	.w4(32'h3d32d2da),
	.w5(32'h3dc33986),
	.w6(32'hbd35d787),
	.w7(32'hbdb8da97),
	.w8(32'hbd926f5a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15660a),
	.w1(32'hbb43fb4f),
	.w2(32'hbad998ba),
	.w3(32'h3d6ba1c6),
	.w4(32'h3b77c204),
	.w5(32'hba2f9da3),
	.w6(32'h3b642f6f),
	.w7(32'h3b2fa1fb),
	.w8(32'h3c3a4189),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbcb4e),
	.w1(32'h3cca3325),
	.w2(32'h3bbec1b0),
	.w3(32'h3c7380b1),
	.w4(32'h3c45f23f),
	.w5(32'h3bc90b2a),
	.w6(32'h3bd03996),
	.w7(32'h3c27a175),
	.w8(32'hbbb5df16),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd5725),
	.w1(32'h3c0f2752),
	.w2(32'h3b6b7b01),
	.w3(32'h3b4f6ee7),
	.w4(32'hba4ecece),
	.w5(32'h394aedc2),
	.w6(32'h3a519d58),
	.w7(32'h3bdf4ae9),
	.w8(32'h3bae4ccf),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c7e42),
	.w1(32'h3c1e74b5),
	.w2(32'hbbbdcb4e),
	.w3(32'h3b82041d),
	.w4(32'h3c57503e),
	.w5(32'hbb0c39f2),
	.w6(32'h3695c138),
	.w7(32'hbb58f798),
	.w8(32'hbb9eb1d5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55133b),
	.w1(32'hbb266511),
	.w2(32'hbaea07b8),
	.w3(32'hbc1eac46),
	.w4(32'h3b9ec62c),
	.w5(32'h3c830b02),
	.w6(32'h3b4efb75),
	.w7(32'h3c0d8251),
	.w8(32'h3c685697),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f027b0),
	.w1(32'h3c5fda18),
	.w2(32'hbbe73cae),
	.w3(32'h3c91bc09),
	.w4(32'h3ce99b47),
	.w5(32'h3c26cb1d),
	.w6(32'h3baf257a),
	.w7(32'h3bc2aadb),
	.w8(32'hbbb30e4a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d5706),
	.w1(32'hbb973476),
	.w2(32'hbb629e83),
	.w3(32'h3c908d4c),
	.w4(32'hbc84b729),
	.w5(32'hbd591838),
	.w6(32'h3c332e62),
	.w7(32'h3d67b7bc),
	.w8(32'h3d15dd00),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73b67e),
	.w1(32'h3bd357c5),
	.w2(32'h3c615024),
	.w3(32'hbcbe739f),
	.w4(32'h3bdc6f9b),
	.w5(32'hbb85febc),
	.w6(32'h3be369ac),
	.w7(32'h3c2c26e0),
	.w8(32'h3be4fbeb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c205225),
	.w1(32'h3aca0988),
	.w2(32'hbb54b2cc),
	.w3(32'h3c3cbe5e),
	.w4(32'h3b4f6d82),
	.w5(32'h3bd4e613),
	.w6(32'hba083c3b),
	.w7(32'hbb281f1c),
	.w8(32'hbb99f069),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b654a40),
	.w1(32'h3cc54eb3),
	.w2(32'h3bf9fe56),
	.w3(32'h3be9ec5c),
	.w4(32'h3a98d5cb),
	.w5(32'h3be30153),
	.w6(32'h3b5b20a1),
	.w7(32'hbb22ad5a),
	.w8(32'hbc8c28e6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcef46a),
	.w1(32'hbabfa9cd),
	.w2(32'h3bc431c2),
	.w3(32'hbad58109),
	.w4(32'h3c5fcd84),
	.w5(32'h3c2dca08),
	.w6(32'h3c13786e),
	.w7(32'hbaeef3c1),
	.w8(32'h3b6ba41d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94fd5e),
	.w1(32'h3bccea3e),
	.w2(32'hbba69d1a),
	.w3(32'h3c608911),
	.w4(32'h3c127903),
	.w5(32'hbb94981a),
	.w6(32'hba1364dc),
	.w7(32'h3918b859),
	.w8(32'hbbb100e2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5ee6),
	.w1(32'h3a22aef2),
	.w2(32'hbbba9675),
	.w3(32'hbb5c6a04),
	.w4(32'h3bdfe5a2),
	.w5(32'h3c2af2e5),
	.w6(32'hbc11d1ef),
	.w7(32'hbc9f5918),
	.w8(32'hbc2d6b4f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c3788),
	.w1(32'h3bc312bf),
	.w2(32'hba24f498),
	.w3(32'h3c9ca5ca),
	.w4(32'h3b79a044),
	.w5(32'h3b877a51),
	.w6(32'h3ac9c990),
	.w7(32'h3b0e4582),
	.w8(32'hbb9434e2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8bf99),
	.w1(32'hbc31635d),
	.w2(32'hbbde073e),
	.w3(32'hbadf8101),
	.w4(32'hbaa2a7e9),
	.w5(32'h3bd627aa),
	.w6(32'hbb818835),
	.w7(32'h3b78910f),
	.w8(32'h3b5d84c7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d443e),
	.w1(32'hbc90bb3a),
	.w2(32'hbce101ea),
	.w3(32'h3b0252a1),
	.w4(32'hbc9f6456),
	.w5(32'hbc9ceb19),
	.w6(32'hbb8a930c),
	.w7(32'hbaaa4924),
	.w8(32'hbb90b910),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd614de),
	.w1(32'h3c5fba2b),
	.w2(32'h3caf46fe),
	.w3(32'hbc44a8de),
	.w4(32'h3c2ecbc6),
	.w5(32'h3ca7e9a1),
	.w6(32'h3b1839bb),
	.w7(32'h3c9d2966),
	.w8(32'h3c51102f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cb6c9),
	.w1(32'hba990b4a),
	.w2(32'hbbe6560e),
	.w3(32'hbae38874),
	.w4(32'h3c263598),
	.w5(32'h3b7b65b8),
	.w6(32'hbc1f30fd),
	.w7(32'hbc343b3d),
	.w8(32'hbbd955de),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f4112),
	.w1(32'hbbb8e51b),
	.w2(32'h3b825e9b),
	.w3(32'h3c2d0804),
	.w4(32'h3c93fc46),
	.w5(32'h3d2d9416),
	.w6(32'hbcd2eefd),
	.w7(32'hbd096b9c),
	.w8(32'hbc84c768),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf76023),
	.w1(32'h3c1123bf),
	.w2(32'h3c06c442),
	.w3(32'h3ce6014d),
	.w4(32'h3bc43540),
	.w5(32'hba4bec6b),
	.w6(32'h3bb2e26d),
	.w7(32'h3bff9660),
	.w8(32'hba2ae74a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924e81d),
	.w1(32'h3be58955),
	.w2(32'h3c3a9b90),
	.w3(32'hbb7eec2b),
	.w4(32'hba429d89),
	.w5(32'hbaca03d3),
	.w6(32'h3a3c4345),
	.w7(32'h3bcc628a),
	.w8(32'h3b781159),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3aa72f),
	.w1(32'hba8ec518),
	.w2(32'hbb31badd),
	.w3(32'hbb7a17e9),
	.w4(32'hb9fcd408),
	.w5(32'hbb820aa3),
	.w6(32'h3ab3ff05),
	.w7(32'h3a05bd1e),
	.w8(32'hbb812913),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd19bf),
	.w1(32'h3c1742ff),
	.w2(32'h3a5a5532),
	.w3(32'hbb86e75c),
	.w4(32'hbabeceb8),
	.w5(32'h3b29d6a4),
	.w6(32'h3becd7e2),
	.w7(32'h3b8349cb),
	.w8(32'h3a9c069a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf19a1),
	.w1(32'h3c87f31f),
	.w2(32'hb9b46eec),
	.w3(32'h39983d86),
	.w4(32'h3c978535),
	.w5(32'h3ba7404f),
	.w6(32'hbc481eee),
	.w7(32'hbc283786),
	.w8(32'hbc3e8a71),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc574c8b),
	.w1(32'h3bbbf0c7),
	.w2(32'h3bb4582e),
	.w3(32'hbbd0b06c),
	.w4(32'hbba88a9d),
	.w5(32'hba09b02f),
	.w6(32'h3c02c259),
	.w7(32'h3b61bc65),
	.w8(32'hbc352ba3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eeeed),
	.w1(32'h3bd93eb9),
	.w2(32'h3bb77eb6),
	.w3(32'h3bece6e2),
	.w4(32'h3b94ecd0),
	.w5(32'hbad6976b),
	.w6(32'h3b05e90c),
	.w7(32'hba720914),
	.w8(32'hbac896da),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d519d5),
	.w1(32'hbbdcb46d),
	.w2(32'hbbbbbff6),
	.w3(32'hbbd0e65e),
	.w4(32'hbb122f08),
	.w5(32'h3b3857f4),
	.w6(32'h39f67614),
	.w7(32'h38f219e7),
	.w8(32'h3b3da13d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b119949),
	.w1(32'h3be8bf66),
	.w2(32'h36e3fc14),
	.w3(32'hbb3aa381),
	.w4(32'h3b359d73),
	.w5(32'h3ae31ace),
	.w6(32'h3b84590f),
	.w7(32'hbaf181de),
	.w8(32'hbbaf295c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6276ef),
	.w1(32'hbb8242a9),
	.w2(32'hbcce8cdc),
	.w3(32'h3b8e2327),
	.w4(32'hbb98b70e),
	.w5(32'hbc7d2768),
	.w6(32'h3bd1d5b5),
	.w7(32'hbc31fc21),
	.w8(32'hbc43e3fd),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc901af2),
	.w1(32'h3c022118),
	.w2(32'hbbcd79d2),
	.w3(32'hbbaef402),
	.w4(32'h3c032f12),
	.w5(32'h3bd7018f),
	.w6(32'h3be3c45e),
	.w7(32'h3b9d18a3),
	.w8(32'h3bd3d2a0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71128e),
	.w1(32'h3a14eb5e),
	.w2(32'h39382982),
	.w3(32'hbb283889),
	.w4(32'h3bedcf10),
	.w5(32'h3b2ca3dd),
	.w6(32'h3b0bc2f1),
	.w7(32'hbb893cf6),
	.w8(32'hbba991a7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803bc9),
	.w1(32'h3c39e206),
	.w2(32'h3b936bb6),
	.w3(32'h3ba6c09e),
	.w4(32'h3c7f53fe),
	.w5(32'h3c3f26ac),
	.w6(32'hbc108249),
	.w7(32'hbc002160),
	.w8(32'hbc2056a7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025902),
	.w1(32'h3c2ff728),
	.w2(32'h3c20b8a3),
	.w3(32'h3ba3344a),
	.w4(32'h3bfd1dd8),
	.w5(32'h3c878af2),
	.w6(32'hbb94b840),
	.w7(32'hbba011e3),
	.w8(32'hbb8be5c1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b112cc0),
	.w1(32'h3a630737),
	.w2(32'hbb3f4075),
	.w3(32'h3c5da827),
	.w4(32'h3938b482),
	.w5(32'hbb486a48),
	.w6(32'hb771ec68),
	.w7(32'h3c137726),
	.w8(32'hb9413a15),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9a7cd),
	.w1(32'h3adc02c5),
	.w2(32'hbb77aa10),
	.w3(32'hbb986788),
	.w4(32'h3b4fde11),
	.w5(32'hbb10d89a),
	.w6(32'h3b109b66),
	.w7(32'h3ba36c49),
	.w8(32'hbc018315),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9712e),
	.w1(32'h3bfff24a),
	.w2(32'h3b9058da),
	.w3(32'hbb44a73e),
	.w4(32'hba4314e6),
	.w5(32'h39d9bd0c),
	.w6(32'h3b1e8008),
	.w7(32'h3c670fec),
	.w8(32'h3c049193),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b567e20),
	.w1(32'h3bc2abc3),
	.w2(32'h3bcd4e4c),
	.w3(32'h3b400598),
	.w4(32'h3c6700cf),
	.w5(32'h3b3dde4f),
	.w6(32'hbbf65624),
	.w7(32'hbb569362),
	.w8(32'hbb63c3b0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0a6ea),
	.w1(32'h3c4d8749),
	.w2(32'h3c02124e),
	.w3(32'h3c0f1406),
	.w4(32'h3c473476),
	.w5(32'h3c128b1b),
	.w6(32'h3c147308),
	.w7(32'h3c77a6e3),
	.w8(32'h3c38ec12),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c751542),
	.w1(32'h3ce80a0e),
	.w2(32'h3c073337),
	.w3(32'h3c1824e2),
	.w4(32'h3c57a636),
	.w5(32'hb9334674),
	.w6(32'hbc83f52a),
	.w7(32'hbbb5289d),
	.w8(32'hbc814c2b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc792b3),
	.w1(32'h3c5f0934),
	.w2(32'h3b1b78a7),
	.w3(32'h3a3180c8),
	.w4(32'h3c5a7b50),
	.w5(32'h3bac3b96),
	.w6(32'hbb6fee3b),
	.w7(32'hbac91759),
	.w8(32'hbb47cd5c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc143880),
	.w1(32'h3c7e8204),
	.w2(32'h3c8acaee),
	.w3(32'hbb75b657),
	.w4(32'h3c3d756d),
	.w5(32'h3c5934b5),
	.w6(32'h3ba57ef9),
	.w7(32'h3c2b750b),
	.w8(32'h3b71ca47),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3371b5),
	.w1(32'hbb2c75d7),
	.w2(32'hbbc387c5),
	.w3(32'h3baedc04),
	.w4(32'h3c53fb8a),
	.w5(32'h3c12299a),
	.w6(32'hbb7916d5),
	.w7(32'hb8f590e3),
	.w8(32'h3bf4fa46),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6a3b6),
	.w1(32'h3b8c87f0),
	.w2(32'h3b3dd351),
	.w3(32'h3bf5c28e),
	.w4(32'h3bf090cd),
	.w5(32'h3c7ae35c),
	.w6(32'hba2962a7),
	.w7(32'h3b125a6b),
	.w8(32'h3b43bd43),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5231c),
	.w1(32'h3ba281f5),
	.w2(32'hbc30e224),
	.w3(32'h3c6bfd2d),
	.w4(32'h3a662335),
	.w5(32'hbbbb3e3d),
	.w6(32'h3b867e74),
	.w7(32'h392b27ea),
	.w8(32'h3b6011bf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3289f),
	.w1(32'h3ade3c26),
	.w2(32'hbb5b46d5),
	.w3(32'hbb0f1bc0),
	.w4(32'h39c08ec4),
	.w5(32'hbbf214de),
	.w6(32'hbbaaddf9),
	.w7(32'hb8b1c88c),
	.w8(32'hbb0cca59),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994eebd),
	.w1(32'hbb64d495),
	.w2(32'h3b54bbe3),
	.w3(32'hbbcfb0f5),
	.w4(32'hbb053c21),
	.w5(32'h3bbfb5e8),
	.w6(32'hbbcf5d4b),
	.w7(32'hbb5af4c1),
	.w8(32'h38bb3098),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba730546),
	.w1(32'h3a99ced9),
	.w2(32'h3bbd5be8),
	.w3(32'hbb20a8b6),
	.w4(32'hbb620d21),
	.w5(32'hbc5d9cca),
	.w6(32'h3c3344e7),
	.w7(32'h3c9a8552),
	.w8(32'h3caed287),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2355b6),
	.w1(32'hbae31d76),
	.w2(32'hbb8b0fde),
	.w3(32'hbb55867e),
	.w4(32'hbcad6eb2),
	.w5(32'hbd38fc33),
	.w6(32'h3c0b7285),
	.w7(32'h3cfd16fb),
	.w8(32'h3cb2b3c1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cdee8),
	.w1(32'h3b630e70),
	.w2(32'hbb337b89),
	.w3(32'hbcae7ede),
	.w4(32'h3b04c701),
	.w5(32'h3b88a895),
	.w6(32'h3c016d56),
	.w7(32'hbba23f67),
	.w8(32'hbb42d717),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28480f),
	.w1(32'h3c274adb),
	.w2(32'h3c6590f7),
	.w3(32'hb662a490),
	.w4(32'h3b9a0009),
	.w5(32'h3bb30d90),
	.w6(32'h3b850eb5),
	.w7(32'h3c0a0fd5),
	.w8(32'hba84fa4d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c310932),
	.w1(32'h3cd16c2e),
	.w2(32'h3bd13d88),
	.w3(32'hbab46a39),
	.w4(32'h3c348419),
	.w5(32'h3c4e5bdc),
	.w6(32'hbaac64f9),
	.w7(32'h395cce87),
	.w8(32'hbbbb4c71),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9067c6),
	.w1(32'h3a557a68),
	.w2(32'h3b521843),
	.w3(32'hba8f6e8d),
	.w4(32'h399898c3),
	.w5(32'h3a7df347),
	.w6(32'h3b83a0bf),
	.w7(32'h3b949f38),
	.w8(32'hb92e6b38),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be29ae4),
	.w1(32'hbb867282),
	.w2(32'hbb4df44f),
	.w3(32'h3aa57e86),
	.w4(32'h3b8a4804),
	.w5(32'h3bba6644),
	.w6(32'hba0a0ba8),
	.w7(32'h395b0721),
	.w8(32'h3b290f0a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f1f0c),
	.w1(32'h3c0d7cd2),
	.w2(32'hba3a2c89),
	.w3(32'h3bedc159),
	.w4(32'h3a9119e7),
	.w5(32'h3bab79e4),
	.w6(32'h3ab77186),
	.w7(32'hbbb49310),
	.w8(32'h393d372e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1ed0),
	.w1(32'h3c00b8c6),
	.w2(32'hbad9b695),
	.w3(32'h3bf4b2b3),
	.w4(32'h3b992c12),
	.w5(32'h3bd5d32d),
	.w6(32'hbb73bfe0),
	.w7(32'hbb081cd9),
	.w8(32'hbbb4de89),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b272fde),
	.w1(32'h3907ff65),
	.w2(32'h3baa9ebf),
	.w3(32'hbb226cb4),
	.w4(32'hba15e9bb),
	.w5(32'h3bed1027),
	.w6(32'hbc2171fc),
	.w7(32'hba7abbd3),
	.w8(32'hbbb5a5cf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c037d44),
	.w1(32'h3b726d05),
	.w2(32'h3bcc7890),
	.w3(32'h3b88817e),
	.w4(32'h39f0903e),
	.w5(32'hb99a9c37),
	.w6(32'h3ad54eb9),
	.w7(32'h3c15779b),
	.w8(32'h3c13c26e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d76bc),
	.w1(32'h3bb3be80),
	.w2(32'h3a4b4909),
	.w3(32'hbac1a2e4),
	.w4(32'hbb8ff718),
	.w5(32'hbc2237b5),
	.w6(32'h3b4558fc),
	.w7(32'h3b7434d6),
	.w8(32'hbb55a4f7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb630454),
	.w1(32'hb90c6990),
	.w2(32'hbb4a6af8),
	.w3(32'hbbdce0b7),
	.w4(32'hb6aec929),
	.w5(32'h3aaa2ce3),
	.w6(32'h3c1a0c75),
	.w7(32'hbc11c188),
	.w8(32'hbad3c300),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba19dec),
	.w1(32'h3ba611fb),
	.w2(32'h3c2a4322),
	.w3(32'h3b37cc4a),
	.w4(32'h3d30c6a5),
	.w5(32'h3dc0fead),
	.w6(32'hbd680278),
	.w7(32'hbdaf94a3),
	.w8(32'hbd7b37fb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2951b),
	.w1(32'h3c2914e7),
	.w2(32'h3c2d24e0),
	.w3(32'h3d54b609),
	.w4(32'h3c44ed9b),
	.w5(32'h3c713de0),
	.w6(32'h3882c789),
	.w7(32'hbb94b51b),
	.w8(32'hbb9ef7cb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92e42d),
	.w1(32'hbc30340a),
	.w2(32'hbc8c4eb0),
	.w3(32'h3c01ee74),
	.w4(32'hbb13cafb),
	.w5(32'hbb660e89),
	.w6(32'hbb751a85),
	.w7(32'hbbe57523),
	.w8(32'h3a96c9af),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95fdfb),
	.w1(32'hba89141c),
	.w2(32'h3b030609),
	.w3(32'h3b2f4955),
	.w4(32'h3a9eb9a7),
	.w5(32'h3a8475c2),
	.w6(32'h3a9328f7),
	.w7(32'h3b77491d),
	.w8(32'h3b128a5b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76310c),
	.w1(32'hbbde4808),
	.w2(32'hbbbeda8f),
	.w3(32'hbb1da9de),
	.w4(32'hbcecd696),
	.w5(32'hbd7d670a),
	.w6(32'h3c9b4c50),
	.w7(32'h3d73fd1a),
	.w8(32'h3d312ff3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf263c),
	.w1(32'hbaa93cc0),
	.w2(32'h3b60a7b2),
	.w3(32'hbd03fcdf),
	.w4(32'h3b1d0cc1),
	.w5(32'hb9da474d),
	.w6(32'h3c076ed5),
	.w7(32'h3b868f9a),
	.w8(32'h3b887d0a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33552f),
	.w1(32'h3b9ad93a),
	.w2(32'h3b5b9d31),
	.w3(32'hbb3ceeee),
	.w4(32'h3ca5a8f9),
	.w5(32'h3d32718a),
	.w6(32'hbc911443),
	.w7(32'hbd0c1d2d),
	.w8(32'hbcd89b36),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f8489),
	.w1(32'hbc2028ba),
	.w2(32'hbc043b28),
	.w3(32'h3cfb114e),
	.w4(32'hbc081842),
	.w5(32'hbbd7ab7d),
	.w6(32'h3c03d77d),
	.w7(32'hbb97e399),
	.w8(32'hba0d063c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5a1a2),
	.w1(32'hbb7e70ed),
	.w2(32'hbbe134c1),
	.w3(32'hbb5252d8),
	.w4(32'hba988201),
	.w5(32'hbc08d9af),
	.w6(32'hbb8d3418),
	.w7(32'hbbb4f38d),
	.w8(32'hbb9cadd9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5aaf53),
	.w1(32'h3b64b809),
	.w2(32'h3b10325e),
	.w3(32'hbbc01463),
	.w4(32'h3b173f95),
	.w5(32'h3c2aa0a7),
	.w6(32'h3b0ab154),
	.w7(32'h3b87c2f2),
	.w8(32'h3b788432),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd68726),
	.w1(32'hbc6a5a34),
	.w2(32'hbc014f73),
	.w3(32'hbb045236),
	.w4(32'hbcbb0e76),
	.w5(32'hbd1dd0cc),
	.w6(32'hbb108733),
	.w7(32'h3cd1f744),
	.w8(32'h3cb69f9d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beeb593),
	.w1(32'h3c2dded0),
	.w2(32'h3bd3c52e),
	.w3(32'hbc831b44),
	.w4(32'h3c60138c),
	.w5(32'h3bdfc2e8),
	.w6(32'h3c1fdbbc),
	.w7(32'h3bbd3a6f),
	.w8(32'h3c301928),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7547ac),
	.w1(32'h3b1365fe),
	.w2(32'hbb27ca2d),
	.w3(32'h3b055e8a),
	.w4(32'hbae46e48),
	.w5(32'hbb21154b),
	.w6(32'hbb95efee),
	.w7(32'hbbdf4526),
	.w8(32'hbbe33343),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08c981),
	.w1(32'hbafd5e00),
	.w2(32'hbc500ae5),
	.w3(32'hbc29a29f),
	.w4(32'hbb9c6995),
	.w5(32'hbad42122),
	.w6(32'hbbee3f23),
	.w7(32'hbacacaf3),
	.w8(32'h3b9cc3e0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef253c),
	.w1(32'h3ae52fb7),
	.w2(32'hbbe96daa),
	.w3(32'hbb875853),
	.w4(32'h39bc5e88),
	.w5(32'hbbb5c2c0),
	.w6(32'h3bac8774),
	.w7(32'hbb9986cd),
	.w8(32'hbbb847b3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d1bb0),
	.w1(32'h3c04d345),
	.w2(32'h3c3bcbdc),
	.w3(32'hbb266bda),
	.w4(32'h3bd88650),
	.w5(32'h3a6a783b),
	.w6(32'h3c4242fa),
	.w7(32'h3c35c703),
	.w8(32'hba81efd4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb047a96),
	.w1(32'h3b12e1a9),
	.w2(32'h3ba7fcbe),
	.w3(32'h3ba308de),
	.w4(32'hbbb60718),
	.w5(32'h3ba2e5a9),
	.w6(32'h3b43cc62),
	.w7(32'hba84d1f0),
	.w8(32'h3c254173),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c669b20),
	.w1(32'hbc3a7c86),
	.w2(32'hbc286111),
	.w3(32'h3b9f2fb5),
	.w4(32'hbcd81eea),
	.w5(32'hbd5d53e5),
	.w6(32'h3c22676c),
	.w7(32'h3d395c7d),
	.w8(32'h3cde8db3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa2f5a),
	.w1(32'hbb667f91),
	.w2(32'hbbf55248),
	.w3(32'hbca211ab),
	.w4(32'hbb1f545d),
	.w5(32'h3a5dddef),
	.w6(32'h3bb54b6d),
	.w7(32'hbb37acc2),
	.w8(32'h3be162dc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7fedc),
	.w1(32'h3ab130a0),
	.w2(32'h3ad188bb),
	.w3(32'hbbcee01d),
	.w4(32'hbad1bf6d),
	.w5(32'hbc1282e9),
	.w6(32'h3b32904c),
	.w7(32'hbb6334af),
	.w8(32'hbb346109),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b6acd),
	.w1(32'h3b1b0b05),
	.w2(32'h3c129443),
	.w3(32'hbc1eeac4),
	.w4(32'h3a1b2bf3),
	.w5(32'h3ab28c46),
	.w6(32'hba44af60),
	.w7(32'h3b8e26af),
	.w8(32'h3b14a164),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05bc05),
	.w1(32'h3b812449),
	.w2(32'h3b914dff),
	.w3(32'hba260bb4),
	.w4(32'hbacf5709),
	.w5(32'h38c3eaa5),
	.w6(32'h3a94fb1a),
	.w7(32'h3b2c4d5f),
	.w8(32'h3b280c42),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0ec27),
	.w1(32'hbb71dd86),
	.w2(32'hbc03e931),
	.w3(32'h3b416577),
	.w4(32'h3a35ed83),
	.w5(32'hbb19ff32),
	.w6(32'hbb4f511f),
	.w7(32'hbbd34b25),
	.w8(32'hbaf44365),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule