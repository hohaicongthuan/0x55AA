module layer_8_featuremap_96(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd76163),
	.w1(32'hbb7b7df9),
	.w2(32'hbbe43a85),
	.w3(32'h3bc87f33),
	.w4(32'hbc77c136),
	.w5(32'hbbf8320c),
	.w6(32'hbc84ab33),
	.w7(32'hb943e50f),
	.w8(32'h3be1d7f5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e89211),
	.w1(32'hbc146ac7),
	.w2(32'h3b327944),
	.w3(32'hbc82c8d8),
	.w4(32'hbbfe71ee),
	.w5(32'hbcd860b4),
	.w6(32'hbc078d0a),
	.w7(32'h3c31b620),
	.w8(32'h3cb7b078),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c7234),
	.w1(32'h3c9c7e0f),
	.w2(32'h3c90623f),
	.w3(32'hbce1d2c8),
	.w4(32'hbc758c24),
	.w5(32'hbc8e04d4),
	.w6(32'h3bfb0a7c),
	.w7(32'h3a2c3ce8),
	.w8(32'h3c0ff6c9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c109a1b),
	.w1(32'hbc24b1df),
	.w2(32'hbcb23d7a),
	.w3(32'hbbc85d5a),
	.w4(32'h3b768e88),
	.w5(32'h3b82dff5),
	.w6(32'h39c4fefb),
	.w7(32'h3af73405),
	.w8(32'h3cb13417),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af50f9),
	.w1(32'hbb3d1b97),
	.w2(32'hbc30aaf1),
	.w3(32'hbb09c000),
	.w4(32'hbbf12602),
	.w5(32'hbbe4bd36),
	.w6(32'hbc5f3139),
	.w7(32'hbc9d98dd),
	.w8(32'hbcc38631),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03437e),
	.w1(32'hbc6855eb),
	.w2(32'h3b4124b2),
	.w3(32'h3c524139),
	.w4(32'h3bf51675),
	.w5(32'hbb642dc5),
	.w6(32'hbc59873d),
	.w7(32'h3b9e0383),
	.w8(32'h3c8d6453),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fa698),
	.w1(32'h3bea2052),
	.w2(32'h3c03a09a),
	.w3(32'hbc0c0117),
	.w4(32'h3b3f7a02),
	.w5(32'hba0a2bec),
	.w6(32'h3be0cdfb),
	.w7(32'h3c0a2b16),
	.w8(32'h3bb8e687),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6626a),
	.w1(32'h3c04c49c),
	.w2(32'hbbd68dda),
	.w3(32'h3bc3e9d8),
	.w4(32'h3b0e9233),
	.w5(32'h3bf31691),
	.w6(32'hba231297),
	.w7(32'hbc217e25),
	.w8(32'hbbd005bd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e2ab2),
	.w1(32'h3be57bdf),
	.w2(32'hbc0b491e),
	.w3(32'hbc57fd1d),
	.w4(32'h3c5f4234),
	.w5(32'h3ca90a12),
	.w6(32'hbc35583f),
	.w7(32'hbc582c88),
	.w8(32'hbcacfb9a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc77c11),
	.w1(32'hbc1c319c),
	.w2(32'hbaa1a737),
	.w3(32'h3b4cb30d),
	.w4(32'h3bc0a7c5),
	.w5(32'hbc54b24c),
	.w6(32'hbc97a5d6),
	.w7(32'h3c524cbd),
	.w8(32'h3d1423a5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb47e35),
	.w1(32'h3c6757ee),
	.w2(32'hbbde4b70),
	.w3(32'hbcc82b06),
	.w4(32'h3c072f47),
	.w5(32'h3d44fbaf),
	.w6(32'h3b0f9d3e),
	.w7(32'hbcd263e5),
	.w8(32'hbcff9e19),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc867159),
	.w1(32'hbbbb8fca),
	.w2(32'hbb9c4e8d),
	.w3(32'h3c75afe5),
	.w4(32'h3bd3edae),
	.w5(32'hbb5aa496),
	.w6(32'hbb7a5a1a),
	.w7(32'h3adc1b09),
	.w8(32'h3b297be7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d60cc1),
	.w1(32'h39ab8546),
	.w2(32'h3a86ad6e),
	.w3(32'hbb2e7c39),
	.w4(32'h3ab006ce),
	.w5(32'h3ae66870),
	.w6(32'hbb32b175),
	.w7(32'h3a26e9fa),
	.w8(32'h3a33a86a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdf0a3),
	.w1(32'h3ae6d34a),
	.w2(32'h3b11ca67),
	.w3(32'h3aa155a9),
	.w4(32'h3aa58f72),
	.w5(32'h3ae9a05b),
	.w6(32'hb9a8bb76),
	.w7(32'h3824cb77),
	.w8(32'h3a80f097),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bbe011),
	.w1(32'hb89cc697),
	.w2(32'h381f8bcc),
	.w3(32'hb8901455),
	.w4(32'h3821318b),
	.w5(32'h390781af),
	.w6(32'hb8a4c404),
	.w7(32'h3877889d),
	.w8(32'h390ac44a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23155e),
	.w1(32'h3950200c),
	.w2(32'h39db977f),
	.w3(32'h3a19d667),
	.w4(32'h3969cc2c),
	.w5(32'h39cada76),
	.w6(32'h3a8c7862),
	.w7(32'h3a433d3b),
	.w8(32'h395cc247),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a607765),
	.w1(32'hb9800de4),
	.w2(32'hb89336b1),
	.w3(32'h3a25112d),
	.w4(32'hb9cfce3d),
	.w5(32'h3a93c883),
	.w6(32'h3afd7405),
	.w7(32'h3a772a93),
	.w8(32'h3a97988b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb346120),
	.w1(32'hbb2c73e2),
	.w2(32'hb87e422f),
	.w3(32'hbb3da660),
	.w4(32'hba848513),
	.w5(32'hba851812),
	.w6(32'hbb478931),
	.w7(32'hbaa0538c),
	.w8(32'hb953346f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39852475),
	.w1(32'h3a9e4fe7),
	.w2(32'h3a5d9151),
	.w3(32'hb968c17b),
	.w4(32'h39990a4a),
	.w5(32'h37b7b63a),
	.w6(32'hbac55fd7),
	.w7(32'h3991cf2c),
	.w8(32'h39da8969),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d09c9),
	.w1(32'hba8c028d),
	.w2(32'hb9540d45),
	.w3(32'hba466a7e),
	.w4(32'hb8a135b6),
	.w5(32'hba27b360),
	.w6(32'hbb26c867),
	.w7(32'hba1a5f1a),
	.w8(32'hbb0d477b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba21bf),
	.w1(32'hb9d9f192),
	.w2(32'h3adf9641),
	.w3(32'h3b055eea),
	.w4(32'h3af789ed),
	.w5(32'hb74d3cf9),
	.w6(32'hba59514a),
	.w7(32'hbb033f97),
	.w8(32'h3842bc75),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf43c5),
	.w1(32'h3b437a27),
	.w2(32'h3ba69bfc),
	.w3(32'h3b062166),
	.w4(32'h3b7979d6),
	.w5(32'h3b6f77af),
	.w6(32'hbb6ddea5),
	.w7(32'hb723d64f),
	.w8(32'h3b1662e3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9e87f),
	.w1(32'hba99d844),
	.w2(32'hbb335708),
	.w3(32'h3b07e92d),
	.w4(32'h39c10952),
	.w5(32'hb9ad6245),
	.w6(32'h3bb685ee),
	.w7(32'h3b8f985e),
	.w8(32'h3b5757ca),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b7ec1),
	.w1(32'hbb18b7e9),
	.w2(32'hba5b55f0),
	.w3(32'hba6ba007),
	.w4(32'hba857008),
	.w5(32'hb901b910),
	.w6(32'hbb30b466),
	.w7(32'hbb16f5ea),
	.w8(32'hba2024ef),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf762cf),
	.w1(32'h3b5f8b91),
	.w2(32'h3b4dee31),
	.w3(32'h3bf54f8e),
	.w4(32'h3b31d18a),
	.w5(32'h3aeef3de),
	.w6(32'h3c39571d),
	.w7(32'h3bb6b43d),
	.w8(32'h3b91ae41),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e0daf),
	.w1(32'hbad84852),
	.w2(32'hbacbdb01),
	.w3(32'hb99474d5),
	.w4(32'hba9f0f66),
	.w5(32'hbaff5fa7),
	.w6(32'hbadfcf6e),
	.w7(32'hba74bd77),
	.w8(32'hb96f91ec),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04b141),
	.w1(32'hbb024724),
	.w2(32'hbacacf16),
	.w3(32'hbb19af7f),
	.w4(32'hbb00d8de),
	.w5(32'hbaa28cb5),
	.w6(32'hbb06e844),
	.w7(32'hbb087f4a),
	.w8(32'hbaaa5a86),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d1717),
	.w1(32'h39ff419d),
	.w2(32'h3ab6baee),
	.w3(32'h3b4651eb),
	.w4(32'h3b11c89c),
	.w5(32'hb9eca9a2),
	.w6(32'h3bea83de),
	.w7(32'h3b876bef),
	.w8(32'h3b64b4d1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13b8aa),
	.w1(32'hba30b665),
	.w2(32'hba4cee19),
	.w3(32'hba0cde8e),
	.w4(32'hb9f28eb1),
	.w5(32'hba18e946),
	.w6(32'hb9ce4c63),
	.w7(32'hb9c24fd4),
	.w8(32'hba18a592),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e963f),
	.w1(32'hb9ce7a0e),
	.w2(32'h3a23b53b),
	.w3(32'h3a0d4dde),
	.w4(32'h3a0cebfd),
	.w5(32'h3aa023ed),
	.w6(32'h39b768c4),
	.w7(32'h39d2e014),
	.w8(32'h3978e3f6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce6f64),
	.w1(32'hbb91d778),
	.w2(32'hbb46f3e1),
	.w3(32'hbbe6925b),
	.w4(32'hbb911e79),
	.w5(32'hbb6042b3),
	.w6(32'hbc097fc0),
	.w7(32'hbbebed06),
	.w8(32'hbbb21626),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a90e8),
	.w1(32'hba473f9d),
	.w2(32'hbacdd24e),
	.w3(32'hba441068),
	.w4(32'hbabe1ab9),
	.w5(32'hbad8442a),
	.w6(32'hb9a16ccd),
	.w7(32'hb99b3b41),
	.w8(32'hb9bae646),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994caa1),
	.w1(32'h39b858f7),
	.w2(32'h3907b564),
	.w3(32'h39d5fb19),
	.w4(32'h392dc6f4),
	.w5(32'h389748e5),
	.w6(32'h38d7ae5b),
	.w7(32'h3956e085),
	.w8(32'h3829b87e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3859dbac),
	.w1(32'hb7eb8171),
	.w2(32'hb88b136b),
	.w3(32'hb8cd8e20),
	.w4(32'h388e0529),
	.w5(32'hb8960155),
	.w6(32'h37ae3e74),
	.w7(32'h382a3a02),
	.w8(32'h385b703a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0be60),
	.w1(32'hbad4977e),
	.w2(32'hba4f795b),
	.w3(32'hba680c16),
	.w4(32'hba5c6ba7),
	.w5(32'hba0b5356),
	.w6(32'hbac67d98),
	.w7(32'hba85698a),
	.w8(32'hba5971a6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33be4c),
	.w1(32'hba03288e),
	.w2(32'hba636b84),
	.w3(32'hb9c724ef),
	.w4(32'hba0e69a0),
	.w5(32'hba258660),
	.w6(32'hb9d97fcd),
	.w7(32'hb98155d3),
	.w8(32'hb8616c84),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92857ed),
	.w1(32'hba01ae07),
	.w2(32'hb97ac54b),
	.w3(32'hb881c19b),
	.w4(32'hb82d32e4),
	.w5(32'h39fcb907),
	.w6(32'h39b50f4f),
	.w7(32'h39bef5f0),
	.w8(32'h398ab927),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5b427),
	.w1(32'hbad0944f),
	.w2(32'hbac751b7),
	.w3(32'hbb085405),
	.w4(32'hbab011b3),
	.w5(32'hba2fd126),
	.w6(32'hbb2abea1),
	.w7(32'hba969483),
	.w8(32'hba366005),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb892d666),
	.w1(32'h37ffacce),
	.w2(32'hb90f5d78),
	.w3(32'hb87e675e),
	.w4(32'hb8cdb2b9),
	.w5(32'hb8db42f8),
	.w6(32'h38b1965e),
	.w7(32'h39532273),
	.w8(32'h38e85f40),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36b87d),
	.w1(32'h3a0d1ba6),
	.w2(32'h3a0058fd),
	.w3(32'h3a3456e2),
	.w4(32'h3981ec4c),
	.w5(32'h3a08dec7),
	.w6(32'hb985bc97),
	.w7(32'hb9a9cd94),
	.w8(32'h3946fe6f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3863a3ec),
	.w1(32'hb89fc016),
	.w2(32'hb9654cb3),
	.w3(32'h385feff8),
	.w4(32'hb8bf5e89),
	.w5(32'h390324f0),
	.w6(32'hb7e31a06),
	.w7(32'h39a2d81d),
	.w8(32'h39139f48),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f2e61),
	.w1(32'hba5b00d8),
	.w2(32'hba52cd03),
	.w3(32'hbabdabc5),
	.w4(32'hba819c23),
	.w5(32'hba5fc16a),
	.w6(32'hbabd7463),
	.w7(32'hbabadbe7),
	.w8(32'hb9dd2c56),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980bf03),
	.w1(32'h3790faac),
	.w2(32'h37a188c4),
	.w3(32'h38634a0f),
	.w4(32'hb995abe7),
	.w5(32'h39d498dd),
	.w6(32'h3946f699),
	.w7(32'hb84f28bb),
	.w8(32'h388666b5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f5375),
	.w1(32'h39aaf5e1),
	.w2(32'hb7b9a0ff),
	.w3(32'h3ace0e94),
	.w4(32'h3a4e6c1f),
	.w5(32'h3a57809c),
	.w6(32'h3abe9b75),
	.w7(32'h3a8ecbc7),
	.w8(32'h3a659fef),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144845),
	.w1(32'hba833aad),
	.w2(32'hb980d810),
	.w3(32'hbaedcd93),
	.w4(32'hba37f44f),
	.w5(32'hba53ce2a),
	.w6(32'hbb85020f),
	.w7(32'hbb5af8e4),
	.w8(32'hbb1568ef),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933f85),
	.w1(32'hb9f89c74),
	.w2(32'hb9d90f78),
	.w3(32'hbadc8712),
	.w4(32'hbaab70a2),
	.w5(32'hba38e2a0),
	.w6(32'hbb342e82),
	.w7(32'hbb0df4fa),
	.w8(32'hbabe9a21),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39042c40),
	.w1(32'h3866e43a),
	.w2(32'hb7f0e396),
	.w3(32'hb8c0937e),
	.w4(32'hb81f9a31),
	.w5(32'hb870da2a),
	.w6(32'hb8d50444),
	.w7(32'hb895f5da),
	.w8(32'hb73ef044),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956a88d),
	.w1(32'hb9f174e9),
	.w2(32'h3ad63941),
	.w3(32'h3a3f30ba),
	.w4(32'h3aeefb02),
	.w5(32'h3b53f45b),
	.w6(32'hba6f324b),
	.w7(32'h38832230),
	.w8(32'h39736c8d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a27c59),
	.w1(32'hb9997439),
	.w2(32'h3715ca38),
	.w3(32'hb95306de),
	.w4(32'h3954168b),
	.w5(32'h3921b87e),
	.w6(32'hb8ac4bc3),
	.w7(32'hb9d2e7a6),
	.w8(32'hb91942c3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaef194),
	.w1(32'hbbb1c179),
	.w2(32'hbb35d925),
	.w3(32'hbb93eda8),
	.w4(32'hbb339708),
	.w5(32'hba4a473e),
	.w6(32'hbb97d9a8),
	.w7(32'hbb5cd2d9),
	.w8(32'hbae7baeb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14762a),
	.w1(32'hbac06d01),
	.w2(32'hbb18c9e0),
	.w3(32'hbb381df9),
	.w4(32'hbb155b2f),
	.w5(32'hbb357941),
	.w6(32'hbb367488),
	.w7(32'hbb480c55),
	.w8(32'hbb483074),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b880bae),
	.w1(32'h3b8ec932),
	.w2(32'h3ba48efb),
	.w3(32'h3b2850c1),
	.w4(32'h3b613178),
	.w5(32'h3aff502d),
	.w6(32'h3a21afb0),
	.w7(32'h3a702cfd),
	.w8(32'h3a8cf55c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a409422),
	.w1(32'hb96859b3),
	.w2(32'h3a956d68),
	.w3(32'h39ce6386),
	.w4(32'hb9bf4dd2),
	.w5(32'h3b0f6e1e),
	.w6(32'h3b2a8036),
	.w7(32'h3b227c5c),
	.w8(32'h3b35b04b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b8ec7),
	.w1(32'hb92be37e),
	.w2(32'hb94ef4b0),
	.w3(32'h3a01caec),
	.w4(32'hb858df08),
	.w5(32'h39203d72),
	.w6(32'hb9b1b0e2),
	.w7(32'h399371b1),
	.w8(32'h39cc8863),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36165fcf),
	.w1(32'hb76becce),
	.w2(32'hb718f95f),
	.w3(32'h371713cd),
	.w4(32'hb84113f3),
	.w5(32'h387831a2),
	.w6(32'h384419c8),
	.w7(32'h38aa3005),
	.w8(32'hb888afe4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f692),
	.w1(32'hbb38480c),
	.w2(32'hbb09ff18),
	.w3(32'hbb580a0c),
	.w4(32'hbb35f2c2),
	.w5(32'hbb0415cf),
	.w6(32'hbb83086e),
	.w7(32'hbaa32144),
	.w8(32'hb9ed2e80),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95badf),
	.w1(32'h3a41a885),
	.w2(32'h3a39a95a),
	.w3(32'h3a45a67e),
	.w4(32'h39a0bfb9),
	.w5(32'h39d7c05a),
	.w6(32'h3a9eaa13),
	.w7(32'h3a104ffd),
	.w8(32'h3a2a645e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab12f92),
	.w1(32'hbabf32b4),
	.w2(32'hba08e41c),
	.w3(32'hb91b3278),
	.w4(32'hba0b7b36),
	.w5(32'h39ae099c),
	.w6(32'h3b0a8c77),
	.w7(32'h39ecfb85),
	.w8(32'h38fe864e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984a85e),
	.w1(32'h391ec9a5),
	.w2(32'hb81727c8),
	.w3(32'h39c8df81),
	.w4(32'h38d00d18),
	.w5(32'h391dec90),
	.w6(32'h39968dd1),
	.w7(32'h39847344),
	.w8(32'h399fd98d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cde20),
	.w1(32'hb9f54c1c),
	.w2(32'h38c07089),
	.w3(32'h3811bab3),
	.w4(32'hb8b6e96a),
	.w5(32'h39e65bef),
	.w6(32'h3ab23fa2),
	.w7(32'h3a918620),
	.w8(32'h3a8ff1dd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe49f0),
	.w1(32'h398edefb),
	.w2(32'h3a82861c),
	.w3(32'h3b1976ef),
	.w4(32'h3a82ed0b),
	.w5(32'h3b1c0801),
	.w6(32'h3b8c56ab),
	.w7(32'h3b553020),
	.w8(32'h3b5dadf0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17027d),
	.w1(32'hb984b226),
	.w2(32'hb991a1f0),
	.w3(32'hb9872c3d),
	.w4(32'hb96f2202),
	.w5(32'hb8e8b512),
	.w6(32'hb9bdceb2),
	.w7(32'hb9c0cf50),
	.w8(32'hb91d3d71),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96424c),
	.w1(32'hba96e82d),
	.w2(32'hba9d885c),
	.w3(32'hbaae5c25),
	.w4(32'hba96b887),
	.w5(32'hba62b91b),
	.w6(32'hbacc7ddb),
	.w7(32'hbab4ed88),
	.w8(32'hba6fc99e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a50d3),
	.w1(32'h3a586b5a),
	.w2(32'h3a541303),
	.w3(32'h39be2327),
	.w4(32'h3a14a8ba),
	.w5(32'h399c80e0),
	.w6(32'hb90752e6),
	.w7(32'h3906040b),
	.w8(32'h390f92ed),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93342b3),
	.w1(32'hb9044abd),
	.w2(32'hb9169647),
	.w3(32'hb9b529bd),
	.w4(32'hb90a3a41),
	.w5(32'hb90a579d),
	.w6(32'hb9d623f3),
	.w7(32'hb888c37d),
	.w8(32'h3715e4f1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9231e17),
	.w1(32'hba8294f5),
	.w2(32'hba7b3cf3),
	.w3(32'h38b8794c),
	.w4(32'hba35d596),
	.w5(32'h38e2f17e),
	.w6(32'h3ab89ff1),
	.w7(32'h3a06a18f),
	.w8(32'h3a2ec491),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3826f2),
	.w1(32'h3b2f07ac),
	.w2(32'h3b4cba6c),
	.w3(32'h3b661479),
	.w4(32'h3b6fe7bc),
	.w5(32'h3b5faec5),
	.w6(32'h3b8793c3),
	.w7(32'h3b92af4f),
	.w8(32'h3b685b83),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c800c),
	.w1(32'hbb56fed6),
	.w2(32'hbad35f8a),
	.w3(32'hba972ede),
	.w4(32'hbac2fef7),
	.w5(32'h3a1f1ecf),
	.w6(32'h3aa09c7a),
	.w7(32'h3a7d3a8f),
	.w8(32'h3a746f63),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43b4c2),
	.w1(32'hbb151712),
	.w2(32'hbb196196),
	.w3(32'hbaafb10a),
	.w4(32'hbb0aec41),
	.w5(32'hba98c883),
	.w6(32'hba553162),
	.w7(32'hba7a6db2),
	.w8(32'hba706678),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aee9cb),
	.w1(32'hba236cb7),
	.w2(32'hba69e4e8),
	.w3(32'h3a5e14e3),
	.w4(32'h398a5afe),
	.w5(32'h3a7ee320),
	.w6(32'h3a654d6d),
	.w7(32'h3aebc330),
	.w8(32'h3ac3b8e7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fabbe),
	.w1(32'hb9e126c1),
	.w2(32'hb9d84f4c),
	.w3(32'hbaa43099),
	.w4(32'hba6fbdfe),
	.w5(32'hba385671),
	.w6(32'hba8e1d21),
	.w7(32'hba934c6c),
	.w8(32'hba85e19b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90b5a0),
	.w1(32'hbab28904),
	.w2(32'hbafa3904),
	.w3(32'hba5dc618),
	.w4(32'hba9c0f79),
	.w5(32'hba309962),
	.w6(32'hb99d29ad),
	.w7(32'h37148249),
	.w8(32'h39c7f1c5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23c9ab),
	.w1(32'hbb37b6a0),
	.w2(32'hbac689c6),
	.w3(32'hbb2140cd),
	.w4(32'hbaf168e1),
	.w5(32'hba5ec2f9),
	.w6(32'hbb1f8bae),
	.w7(32'hbaba05bb),
	.w8(32'hba21aee7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d8d98),
	.w1(32'hba5652f0),
	.w2(32'hbaa315d2),
	.w3(32'h3b8764ec),
	.w4(32'h398d265d),
	.w5(32'h3aff08ff),
	.w6(32'h3b6dea41),
	.w7(32'h3b3cc417),
	.w8(32'h3b47671c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39003cb1),
	.w1(32'hb8311031),
	.w2(32'h38ff4bf8),
	.w3(32'hb888cca8),
	.w4(32'hb6da5395),
	.w5(32'hb81ec93b),
	.w6(32'h378a5232),
	.w7(32'hb8099365),
	.w8(32'h3711575c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d28450),
	.w1(32'hba912e07),
	.w2(32'hba1f1ea3),
	.w3(32'h3a971e93),
	.w4(32'h3926cc61),
	.w5(32'h3a3ec36b),
	.w6(32'h3b67884c),
	.w7(32'h3b0b3b25),
	.w8(32'h3af84ed1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912ffee),
	.w1(32'hb9a4dcc9),
	.w2(32'hbb6f8517),
	.w3(32'hb9ef2bc4),
	.w4(32'h3bab0a89),
	.w5(32'hbb0d3aee),
	.w6(32'hba0ddd77),
	.w7(32'h3923ea36),
	.w8(32'hbc1ca1e8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7c71f),
	.w1(32'hbb53e9e1),
	.w2(32'h3b8ac16a),
	.w3(32'h3ad1029b),
	.w4(32'hbb8696ce),
	.w5(32'h3a35bc67),
	.w6(32'hbb1036fb),
	.w7(32'h3bd48e21),
	.w8(32'h3bd48d3f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82d5a8),
	.w1(32'hbc1b9710),
	.w2(32'hba9d42bb),
	.w3(32'h3b04ac6a),
	.w4(32'hbbc4e76e),
	.w5(32'hbb915c7b),
	.w6(32'h3b584b13),
	.w7(32'hba864be4),
	.w8(32'h3a678ccd),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fd27d),
	.w1(32'hbbd33ba6),
	.w2(32'hba89f834),
	.w3(32'h3b1b9462),
	.w4(32'h3c43fd75),
	.w5(32'hba4ba2db),
	.w6(32'hbb22fb6d),
	.w7(32'hba08985b),
	.w8(32'h3b045a87),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34e430),
	.w1(32'h3a07ea15),
	.w2(32'h3c1934b5),
	.w3(32'hbbdc4bc2),
	.w4(32'hb9b57a43),
	.w5(32'hbbca6c4a),
	.w6(32'hbb6889d2),
	.w7(32'h3b83abc2),
	.w8(32'h3b29c45a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab6c99),
	.w1(32'hbc4e038a),
	.w2(32'h3ac3079d),
	.w3(32'hbc802f2d),
	.w4(32'h3c2d3b65),
	.w5(32'h3c21e32f),
	.w6(32'hbc26df0b),
	.w7(32'h3c6a58b5),
	.w8(32'hbcb68600),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb73b44),
	.w1(32'h3b9a6d7a),
	.w2(32'h3ce2aea6),
	.w3(32'hbb7ebefc),
	.w4(32'h391a4e50),
	.w5(32'h3cd4edb1),
	.w6(32'hbbd45566),
	.w7(32'h3bda37a4),
	.w8(32'hbb238563),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc159cbd),
	.w1(32'h3c48d43e),
	.w2(32'hbbf969b7),
	.w3(32'hbbaa8851),
	.w4(32'h3ca84fa1),
	.w5(32'h3c2167df),
	.w6(32'h3bfebe37),
	.w7(32'hbbe357fd),
	.w8(32'h3c2e7514),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b860106),
	.w1(32'hbcc892ce),
	.w2(32'hbc3de64a),
	.w3(32'h396de672),
	.w4(32'h39dfdaac),
	.w5(32'hba05e0c5),
	.w6(32'h3d05d8e9),
	.w7(32'hbc326c18),
	.w8(32'h3d51f2d9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92b56d),
	.w1(32'hbd016275),
	.w2(32'h3ba9a52a),
	.w3(32'h3c9b8e19),
	.w4(32'hbb149cb6),
	.w5(32'hbacd740c),
	.w6(32'hbc8addd6),
	.w7(32'h3cb45094),
	.w8(32'h3ca8c3d7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca41628),
	.w1(32'hbb71e455),
	.w2(32'h3bff00c5),
	.w3(32'h3c003551),
	.w4(32'h3c88a704),
	.w5(32'hbcce0a2f),
	.w6(32'hbb0c81b2),
	.w7(32'hbc277285),
	.w8(32'h3c279585),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1841e),
	.w1(32'hbc2f5285),
	.w2(32'hbbc5d7c0),
	.w3(32'h3b64fa6b),
	.w4(32'h3c99836a),
	.w5(32'h3c38cffb),
	.w6(32'h3b8a50a5),
	.w7(32'h3b7f3aff),
	.w8(32'h3bac518a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9ab46),
	.w1(32'hbbe94584),
	.w2(32'h3b822919),
	.w3(32'hbb3d04f3),
	.w4(32'hbbca8fa6),
	.w5(32'hbc3c5a9d),
	.w6(32'hbac88dfe),
	.w7(32'hbc2d737a),
	.w8(32'h3b67996a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d6478),
	.w1(32'hbba31b43),
	.w2(32'h3c023bf5),
	.w3(32'hbabd264e),
	.w4(32'hbb903a80),
	.w5(32'hbb6afac7),
	.w6(32'h3b8fbed6),
	.w7(32'hbc0f2ef1),
	.w8(32'h3d4460d9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c44ce9),
	.w1(32'hbca38a45),
	.w2(32'hbc8786fd),
	.w3(32'h3bcbbe75),
	.w4(32'h3c8c34f5),
	.w5(32'h3a7b8e72),
	.w6(32'h3a81ad75),
	.w7(32'hb8f25c33),
	.w8(32'hbca671df),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf76211),
	.w1(32'h3bcfad5f),
	.w2(32'hb8e19868),
	.w3(32'hbc48d7e2),
	.w4(32'h39b0efd0),
	.w5(32'h3c3b8711),
	.w6(32'h3c208fe1),
	.w7(32'hbc015cfe),
	.w8(32'hbc37beb2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20a833),
	.w1(32'h3c47c0f7),
	.w2(32'hba1242c8),
	.w3(32'h3b75c878),
	.w4(32'hbc0cbcc5),
	.w5(32'h3b63b640),
	.w6(32'hbb91e9e7),
	.w7(32'hbcc3f553),
	.w8(32'h3cb35ba1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01d880),
	.w1(32'hbb3d4db6),
	.w2(32'h399c1277),
	.w3(32'hba4066f8),
	.w4(32'h3bc9a6d7),
	.w5(32'hbc3868df),
	.w6(32'h3b45dc2f),
	.w7(32'hbcf6a725),
	.w8(32'h3d2810d3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a6694),
	.w1(32'hbae09ea7),
	.w2(32'h3b3cfd6b),
	.w3(32'h3bc40760),
	.w4(32'h3b09acb0),
	.w5(32'h3b2fcf11),
	.w6(32'hbb76e291),
	.w7(32'h3aacd6f1),
	.w8(32'h3aca6ac4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed0e83),
	.w1(32'h3bcb1399),
	.w2(32'hbc909732),
	.w3(32'h3bed847a),
	.w4(32'h3c99de63),
	.w5(32'h3c537ff7),
	.w6(32'h3b933e3a),
	.w7(32'h3c9b4daa),
	.w8(32'hbd13d683),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e7270),
	.w1(32'hbbcf8ed3),
	.w2(32'hbb337c08),
	.w3(32'hbc078213),
	.w4(32'h3baa39c6),
	.w5(32'hbcb35a07),
	.w6(32'hbca604be),
	.w7(32'hbca0ea92),
	.w8(32'hbc74f716),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8a5b0),
	.w1(32'h3b917740),
	.w2(32'hbafec060),
	.w3(32'hbbdee842),
	.w4(32'h3ba3ad1c),
	.w5(32'h3c77686d),
	.w6(32'h3bad3499),
	.w7(32'h3c728da6),
	.w8(32'hbb8fd802),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca36a3a),
	.w1(32'hbbd2c1c9),
	.w2(32'hbbfe2b64),
	.w3(32'hbc8df117),
	.w4(32'hbcbf1e0c),
	.w5(32'hbc5c8594),
	.w6(32'h3c1abb26),
	.w7(32'hbcbc3be4),
	.w8(32'h3b0b3b5e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e66ea),
	.w1(32'hbc05f26f),
	.w2(32'hbc2cfa7d),
	.w3(32'h3b01ea7b),
	.w4(32'h3c03a6ce),
	.w5(32'hbd0450a7),
	.w6(32'hba41da9d),
	.w7(32'hbc92c17d),
	.w8(32'hbc168fe1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a72b0),
	.w1(32'h3c72d126),
	.w2(32'h3bda17aa),
	.w3(32'h3ba123d1),
	.w4(32'h3bb90966),
	.w5(32'h3c2a5a63),
	.w6(32'h3c6ab909),
	.w7(32'hbc48221f),
	.w8(32'h3adc23f8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78418b),
	.w1(32'h3978aaff),
	.w2(32'hbb82d1ac),
	.w3(32'hba9ee9c9),
	.w4(32'h3c099a63),
	.w5(32'hbc419be3),
	.w6(32'h39aa830b),
	.w7(32'h3bdfe014),
	.w8(32'hbce916a0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9129cc),
	.w1(32'hbb56e838),
	.w2(32'hbbd89c36),
	.w3(32'hbc0fc324),
	.w4(32'h3b6a393c),
	.w5(32'h3bb2182f),
	.w6(32'h3bcb7d97),
	.w7(32'h3bc2541b),
	.w8(32'hbbd81ac9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba80fe),
	.w1(32'hbc1fa73b),
	.w2(32'hba2b442d),
	.w3(32'hbafe0412),
	.w4(32'h3c565939),
	.w5(32'h3aa9fe13),
	.w6(32'hbafa68c0),
	.w7(32'hbb8844ca),
	.w8(32'hb8e5dd07),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce151),
	.w1(32'hbbe35b16),
	.w2(32'hbb287167),
	.w3(32'h3b32a66a),
	.w4(32'h3afa2d06),
	.w5(32'h3bde88e5),
	.w6(32'h3c161905),
	.w7(32'h3ca20df2),
	.w8(32'hbc063eec),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19791a),
	.w1(32'hbbfabde4),
	.w2(32'hbbc2acdc),
	.w3(32'hbc3cbd9c),
	.w4(32'hbc8789e1),
	.w5(32'h3a07145b),
	.w6(32'h3d0ec8ac),
	.w7(32'hbc6320b5),
	.w8(32'hbb98e47a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03f40c),
	.w1(32'h3be2d4ce),
	.w2(32'hbb226965),
	.w3(32'h3bfbed35),
	.w4(32'h3c51c4d8),
	.w5(32'hbcbf55dd),
	.w6(32'hbcb35be0),
	.w7(32'hbd07a00e),
	.w8(32'hbbf577a3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f45f),
	.w1(32'h3cbf6822),
	.w2(32'hba018b4f),
	.w3(32'hba801b6f),
	.w4(32'h3b97646e),
	.w5(32'hbb9e9e3f),
	.w6(32'hbc133d2b),
	.w7(32'hbaf7d7b2),
	.w8(32'hbc3ea5d7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc384bde),
	.w1(32'hbbe593c2),
	.w2(32'hbc8ba9fb),
	.w3(32'hbc008070),
	.w4(32'hbce14a6f),
	.w5(32'hbb949f6c),
	.w6(32'hbc0db75c),
	.w7(32'hbcf745f5),
	.w8(32'h3b46d3e0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20c9f7),
	.w1(32'h3bb76ea6),
	.w2(32'hbc106c2d),
	.w3(32'h3b99f5cb),
	.w4(32'hbbd86876),
	.w5(32'hbce29f09),
	.w6(32'h3b9123a2),
	.w7(32'hbcc71070),
	.w8(32'hbc0694d5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf6083),
	.w1(32'h3c850f27),
	.w2(32'hbad3ec76),
	.w3(32'h3c221549),
	.w4(32'hbc811786),
	.w5(32'hbc562321),
	.w6(32'hbb5d4024),
	.w7(32'hbcddd7a9),
	.w8(32'h3c792167),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87de66),
	.w1(32'h392d8930),
	.w2(32'h3ba9b0f5),
	.w3(32'hba7a0a60),
	.w4(32'h3c28992b),
	.w5(32'hbc335d5f),
	.w6(32'h3bf938cf),
	.w7(32'hbb782711),
	.w8(32'h3c2948fc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf4a09),
	.w1(32'h3a2dc9bc),
	.w2(32'hbc3dc7f1),
	.w3(32'h3bf9590a),
	.w4(32'h3c119867),
	.w5(32'h3c44f99a),
	.w6(32'h3ca444cc),
	.w7(32'h3cfefe0f),
	.w8(32'hbcb60776),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1cfd5),
	.w1(32'hbb12facf),
	.w2(32'hbc958a99),
	.w3(32'hbbc88528),
	.w4(32'h3cbbe3ec),
	.w5(32'h3bc834ac),
	.w6(32'hbd124bbb),
	.w7(32'h3d189dfe),
	.w8(32'hbd1e6da2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2f62c0),
	.w1(32'hbd060c01),
	.w2(32'hbbe2da0d),
	.w3(32'hbd0afdd6),
	.w4(32'h3b91101e),
	.w5(32'h3c81adb4),
	.w6(32'hbd0d38dc),
	.w7(32'hbc7adb8b),
	.w8(32'h3c963e38),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba8c7a),
	.w1(32'hbc2f7900),
	.w2(32'hbb9b9e20),
	.w3(32'hbb212dee),
	.w4(32'hbcfc0131),
	.w5(32'hbc3d73fb),
	.w6(32'h3a9bce9f),
	.w7(32'hbcd236a0),
	.w8(32'h3d30372e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd5ab36),
	.w1(32'hbc33dad2),
	.w2(32'h3c9dcaf2),
	.w3(32'h3ca8372b),
	.w4(32'hbc6176d3),
	.w5(32'h3d3e2c0e),
	.w6(32'h3cac9c34),
	.w7(32'h3d53afe7),
	.w8(32'hbd015667),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34e9f),
	.w1(32'h3b793b99),
	.w2(32'hb9fe8fca),
	.w3(32'h3c210e3c),
	.w4(32'hbaf57fbe),
	.w5(32'hbac82165),
	.w6(32'h3c752772),
	.w7(32'h3a6a1d21),
	.w8(32'hbb6a0b8b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5144a5),
	.w1(32'hbb1ab067),
	.w2(32'h3c618b9c),
	.w3(32'hb82a7d65),
	.w4(32'hbc9a178d),
	.w5(32'hbb3730d2),
	.w6(32'hb907c569),
	.w7(32'hbd03935f),
	.w8(32'h3d53d1f2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb321abe),
	.w1(32'hbc8778d0),
	.w2(32'hbb0db703),
	.w3(32'h3bec19f8),
	.w4(32'h3caa1490),
	.w5(32'h3b7df405),
	.w6(32'hbb16c979),
	.w7(32'h3ce6912f),
	.w8(32'hbd1cb3b0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad68ff),
	.w1(32'hbc6b8b93),
	.w2(32'hb84272cc),
	.w3(32'hbcc37a47),
	.w4(32'h3c277d50),
	.w5(32'h3bbb282b),
	.w6(32'hbc666e44),
	.w7(32'h3ba63a6a),
	.w8(32'h3b546874),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6d1bd),
	.w1(32'hbc2339b8),
	.w2(32'h3c106dd3),
	.w3(32'hbb2de212),
	.w4(32'hbc13f2a6),
	.w5(32'h3ba8cad1),
	.w6(32'hbae43cd0),
	.w7(32'hbc952682),
	.w8(32'h3d04c60d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce2c24),
	.w1(32'hbbc462f9),
	.w2(32'hbb42809d),
	.w3(32'hbc744cba),
	.w4(32'hb95605e9),
	.w5(32'hbb877492),
	.w6(32'hbb367ff2),
	.w7(32'h39849c91),
	.w8(32'hbc0c6773),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886725),
	.w1(32'hbb764d3b),
	.w2(32'hbb1fc5b6),
	.w3(32'hbb55eb77),
	.w4(32'h3c9d41f5),
	.w5(32'h3b15f87f),
	.w6(32'hbad46c38),
	.w7(32'h3c449d03),
	.w8(32'hbd0ab179),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f0c80),
	.w1(32'hbc2ff31b),
	.w2(32'hbbd12bce),
	.w3(32'hbc011641),
	.w4(32'h3d033572),
	.w5(32'h3ca22824),
	.w6(32'hbca2946e),
	.w7(32'h3cddcb20),
	.w8(32'hbd22fd25),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e3936),
	.w1(32'hbcaa87c2),
	.w2(32'h3b361480),
	.w3(32'hbc89fd98),
	.w4(32'h3bb8fb3d),
	.w5(32'h3c30f623),
	.w6(32'hba101bb4),
	.w7(32'h3aceace5),
	.w8(32'h3b5c6494),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a0bf4),
	.w1(32'h399b36d3),
	.w2(32'hbb9c4a7c),
	.w3(32'h3b8fcfe6),
	.w4(32'h3bd9bf01),
	.w5(32'hbb39e018),
	.w6(32'h3b18f439),
	.w7(32'h3cb65eaa),
	.w8(32'h3a06d449),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71a73a),
	.w1(32'h3b82a990),
	.w2(32'h39502d11),
	.w3(32'hbac84434),
	.w4(32'h3c260502),
	.w5(32'h3b372986),
	.w6(32'h3c31fe80),
	.w7(32'h3c399387),
	.w8(32'hbbf1971f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule