module layer_10_featuremap_484(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c3952),
	.w1(32'h3ac0b1a8),
	.w2(32'h3aeb705d),
	.w3(32'hb944abc2),
	.w4(32'h3afcf483),
	.w5(32'h3b035799),
	.w6(32'h39d622ee),
	.w7(32'h3ae069f9),
	.w8(32'h3b0f291d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d47c0),
	.w1(32'hbb63f4ab),
	.w2(32'hbba6c895),
	.w3(32'hbaa22dcb),
	.w4(32'hbb0ebc09),
	.w5(32'hbb25698d),
	.w6(32'hba6c6b8f),
	.w7(32'hbac36fa0),
	.w8(32'hba8f1089),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7993c9),
	.w1(32'hb9e07474),
	.w2(32'h392b002f),
	.w3(32'hba3f2bf2),
	.w4(32'hbab7af8e),
	.w5(32'hb9f973ca),
	.w6(32'hba68b738),
	.w7(32'hba5c0485),
	.w8(32'h3834faf7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf6a36),
	.w1(32'h3af3c656),
	.w2(32'h3ae6512d),
	.w3(32'h3a1f2bc0),
	.w4(32'h3aad8532),
	.w5(32'hb61b023a),
	.w6(32'hb9e4f16f),
	.w7(32'hba0310cb),
	.w8(32'hba31d886),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379254aa),
	.w1(32'hb6e27e05),
	.w2(32'hb982eac1),
	.w3(32'h379fdeb2),
	.w4(32'h3915dfca),
	.w5(32'hb90c8b39),
	.w6(32'h3a1a197f),
	.w7(32'hb8e23208),
	.w8(32'h39c57463),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1de9fd),
	.w1(32'h3a31fa29),
	.w2(32'h3a29f739),
	.w3(32'h398f72f6),
	.w4(32'h38fe0db2),
	.w5(32'hb892c01d),
	.w6(32'h3a096c91),
	.w7(32'h390941fb),
	.w8(32'h393d9504),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9c594),
	.w1(32'h3919bb0f),
	.w2(32'h3a1cc1d4),
	.w3(32'h3a804138),
	.w4(32'h38306669),
	.w5(32'h3a0edf0e),
	.w6(32'h3a54e262),
	.w7(32'hbaaee6b6),
	.w8(32'hba630685),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a144da7),
	.w1(32'h3a920c7e),
	.w2(32'h3b207366),
	.w3(32'h3b513dad),
	.w4(32'h3a40bf7c),
	.w5(32'hba1134ec),
	.w6(32'hbb0d93b2),
	.w7(32'hbb28bc08),
	.w8(32'hb914ebf9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39073680),
	.w1(32'h3ad5f274),
	.w2(32'h3a884e1f),
	.w3(32'hb9ee5c78),
	.w4(32'h3a551fc3),
	.w5(32'h3a6c7e77),
	.w6(32'h39c5c076),
	.w7(32'h3a976470),
	.w8(32'h3a3b985f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b102f),
	.w1(32'h3b2bde77),
	.w2(32'h390355d5),
	.w3(32'h3c3d0873),
	.w4(32'h3b48c3b7),
	.w5(32'hbacddc97),
	.w6(32'h3c2260ad),
	.w7(32'h3aede867),
	.w8(32'hbaabccab),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47ae3f),
	.w1(32'hba5da9b7),
	.w2(32'hba0a8c1f),
	.w3(32'hba98aabd),
	.w4(32'hba392d4b),
	.w5(32'hb9f744fa),
	.w6(32'hba3d5212),
	.w7(32'hba467001),
	.w8(32'hba8d5a5f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8388fe),
	.w1(32'h3b854135),
	.w2(32'h3aa8a43a),
	.w3(32'h3b4655a6),
	.w4(32'h3b021ae2),
	.w5(32'hb98d710c),
	.w6(32'h3a68e687),
	.w7(32'hba8a396d),
	.w8(32'hbb4cd068),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6567ee),
	.w1(32'h3b4edfba),
	.w2(32'hb7dc6dc3),
	.w3(32'h3c5e422f),
	.w4(32'h3b81a3a9),
	.w5(32'hba4d2f6f),
	.w6(32'h3c28a6e2),
	.w7(32'h3af54cc0),
	.w8(32'hbb02ddb9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc6636),
	.w1(32'h39110005),
	.w2(32'hbb903d3c),
	.w3(32'h3b2a3f6d),
	.w4(32'h3aff1f54),
	.w5(32'hbb789ad4),
	.w6(32'h3ad48dab),
	.w7(32'h3afea8e4),
	.w8(32'hba1d6cba),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a978d82),
	.w1(32'hba467f46),
	.w2(32'hba17b35a),
	.w3(32'hbaa29d56),
	.w4(32'hbb0b39b7),
	.w5(32'hb95918a8),
	.w6(32'hba1fffad),
	.w7(32'hb9a56f90),
	.w8(32'hba593e9d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc00363),
	.w1(32'h3a83b510),
	.w2(32'h39aaa8a6),
	.w3(32'h3b9fa0f0),
	.w4(32'h3b05ba3b),
	.w5(32'hb96be302),
	.w6(32'h3ba9e2d9),
	.w7(32'h3b004453),
	.w8(32'h3a469861),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba930fb7),
	.w1(32'h3981d46a),
	.w2(32'hb5df9da4),
	.w3(32'hbafd367f),
	.w4(32'h3a4a8f70),
	.w5(32'h3a862629),
	.w6(32'hbac01d13),
	.w7(32'h3ab20522),
	.w8(32'h3acb3eb3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1874a8),
	.w1(32'h3bdf47b9),
	.w2(32'h3bd7806d),
	.w3(32'h3c1ed37e),
	.w4(32'h3aae2fea),
	.w5(32'h3bc33528),
	.w6(32'h3baea863),
	.w7(32'h38e0763e),
	.w8(32'h3bb21112),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9aa45),
	.w1(32'h3b733369),
	.w2(32'h3b8ed74d),
	.w3(32'h3bdb4a56),
	.w4(32'h3b7dc7aa),
	.w5(32'h3b9e4687),
	.w6(32'h3b9044c2),
	.w7(32'h3ada58e9),
	.w8(32'h3b1576ac),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d01cd),
	.w1(32'h3adc2307),
	.w2(32'h3aff0876),
	.w3(32'h3a5ad62c),
	.w4(32'h3a9c5cb6),
	.w5(32'h3b0aeab8),
	.w6(32'h3a9df234),
	.w7(32'h3a60f132),
	.w8(32'h3ad08f21),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4bf50),
	.w1(32'hb96ab592),
	.w2(32'hba207dba),
	.w3(32'h3ade682f),
	.w4(32'h39019caf),
	.w5(32'hba5e5d7c),
	.w6(32'h3adfb345),
	.w7(32'h39b4c8ea),
	.w8(32'hb9436b7a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81e860),
	.w1(32'hba8a9867),
	.w2(32'hbb383391),
	.w3(32'hba6e49ef),
	.w4(32'hba5a89d5),
	.w5(32'hbb03ec81),
	.w6(32'hba554945),
	.w7(32'hba87dcbd),
	.w8(32'hbb050e6c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c389d7f),
	.w1(32'h3c3c5d06),
	.w2(32'h3c624d34),
	.w3(32'h3c0337c5),
	.w4(32'h3c585108),
	.w5(32'h3c1a7ad3),
	.w6(32'h3bd485d9),
	.w7(32'h3aa12735),
	.w8(32'h3bd044ad),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac6653),
	.w1(32'h38b65393),
	.w2(32'hbac485a9),
	.w3(32'h3b892697),
	.w4(32'hbb12fd37),
	.w5(32'hbba66d1d),
	.w6(32'h3ab0f016),
	.w7(32'hbb43587c),
	.w8(32'hbb8181a8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae477b9),
	.w1(32'hbb8485f3),
	.w2(32'hbb849401),
	.w3(32'hb9ba9ef2),
	.w4(32'hbba9a7e5),
	.w5(32'hbbc5a2cd),
	.w6(32'hba87263a),
	.w7(32'hbbae884c),
	.w8(32'hbbaa6f9f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb851e1ba),
	.w1(32'hba614475),
	.w2(32'hb994f0f9),
	.w3(32'hba68885c),
	.w4(32'hb9f9f497),
	.w5(32'hba5373f9),
	.w6(32'hba17fb03),
	.w7(32'hb9f12adf),
	.w8(32'h38332c86),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9020c20),
	.w1(32'h39fd6501),
	.w2(32'h3929bd04),
	.w3(32'hba00a186),
	.w4(32'h3a3cddea),
	.w5(32'h39454db2),
	.w6(32'hba04b0b9),
	.w7(32'h3a314ce5),
	.w8(32'h38d749e2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d2d7f),
	.w1(32'hbae07e39),
	.w2(32'hbb82ccbc),
	.w3(32'hb96d8ddd),
	.w4(32'hbb4d1047),
	.w5(32'hbb5e6808),
	.w6(32'hb91a07b4),
	.w7(32'hbb2e0350),
	.w8(32'hbb6e74dd),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72ca33),
	.w1(32'hb9375d1e),
	.w2(32'hbb2147a9),
	.w3(32'hbaee7cca),
	.w4(32'hba33399d),
	.w5(32'hbb04cecb),
	.w6(32'hbb127c94),
	.w7(32'hba496889),
	.w8(32'hbb22a402),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51c7ac),
	.w1(32'hb8430c16),
	.w2(32'hbadf8113),
	.w3(32'h3b284cfd),
	.w4(32'h3a23be82),
	.w5(32'hbacfd198),
	.w6(32'h3b25162e),
	.w7(32'h3aba4d50),
	.w8(32'h3ac6c176),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a681aa0),
	.w1(32'h39c1066b),
	.w2(32'hb9437fcb),
	.w3(32'h3a646edb),
	.w4(32'hb9b3f7d3),
	.w5(32'h3900182d),
	.w6(32'h3a28293b),
	.w7(32'hb98c2921),
	.w8(32'hb6674078),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5aeba2),
	.w1(32'h3a03ea7e),
	.w2(32'h3a4bd75f),
	.w3(32'hb9b3efd2),
	.w4(32'h39d368d2),
	.w5(32'h3a8cde86),
	.w6(32'hba6bb4da),
	.w7(32'h387f7166),
	.w8(32'h3a77c4e2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63bb0f),
	.w1(32'hba5b4665),
	.w2(32'hba32e66f),
	.w3(32'h3b4585d0),
	.w4(32'hba85a0db),
	.w5(32'hbac89768),
	.w6(32'h3b39b169),
	.w7(32'hbab9baf1),
	.w8(32'hbafe549a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eac200),
	.w1(32'hba3b5156),
	.w2(32'hbab00cd7),
	.w3(32'hba75548d),
	.w4(32'hb9ff600a),
	.w5(32'hba9870f5),
	.w6(32'hba526bb0),
	.w7(32'hba53ae23),
	.w8(32'hbaf178de),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3755f169),
	.w1(32'hb9ecd499),
	.w2(32'h3a151f1d),
	.w3(32'h38a5cbed),
	.w4(32'hb9eb1156),
	.w5(32'hb9ba03ae),
	.w6(32'hb88511bb),
	.w7(32'hba42c28a),
	.w8(32'hb910fa20),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b556a34),
	.w1(32'h3ab47b2c),
	.w2(32'h3ac8dc5d),
	.w3(32'h3a8911b6),
	.w4(32'hba386950),
	.w5(32'h38c50b10),
	.w6(32'h39ac041b),
	.w7(32'hbaa4431e),
	.w8(32'hb8c81d3b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092a62),
	.w1(32'h3b09f33a),
	.w2(32'h399d627a),
	.w3(32'h3bd4a8b6),
	.w4(32'h3b1603b4),
	.w5(32'h3b32ea67),
	.w6(32'h3b801115),
	.w7(32'h3a0e3240),
	.w8(32'hbab3375a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5c902),
	.w1(32'hbb473977),
	.w2(32'hbc4d5b0e),
	.w3(32'hbbd1da0e),
	.w4(32'hbb1d1a98),
	.w5(32'hbbf10d15),
	.w6(32'hbbec741c),
	.w7(32'hbaf6f539),
	.w8(32'hbba8d5a5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf54c01),
	.w1(32'hbba54b44),
	.w2(32'hbc5cf93a),
	.w3(32'hbc13cb85),
	.w4(32'hbbbb5e9c),
	.w5(32'hbc3e1bcc),
	.w6(32'hbc0f931c),
	.w7(32'hbb180f15),
	.w8(32'hbc026045),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d3408),
	.w1(32'hba31148f),
	.w2(32'h39c78a69),
	.w3(32'hba293018),
	.w4(32'hb8d4d1b6),
	.w5(32'h39835bf0),
	.w6(32'hba34a071),
	.w7(32'h3a6f034d),
	.w8(32'h3a4aba81),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2889ec),
	.w1(32'hb94966eb),
	.w2(32'hb932ea4c),
	.w3(32'hb9d47795),
	.w4(32'hba9f5807),
	.w5(32'hba4fef8f),
	.w6(32'hb9e28844),
	.w7(32'hba1e27d8),
	.w8(32'hb866b370),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64ed1e),
	.w1(32'h3a4fa107),
	.w2(32'h389e6d87),
	.w3(32'hba91dc5f),
	.w4(32'h39ebf3a8),
	.w5(32'h394d83f2),
	.w6(32'hba6d006a),
	.w7(32'h3a25ffa5),
	.w8(32'h39cda771),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c5fac),
	.w1(32'h3ab89725),
	.w2(32'hbaff0eab),
	.w3(32'h3908e266),
	.w4(32'hb9c08f26),
	.w5(32'hbb65b24f),
	.w6(32'h3b0ca5ca),
	.w7(32'h3aa08edd),
	.w8(32'hbb1caf46),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a54ed),
	.w1(32'h3b4c2ff7),
	.w2(32'h3b8cc086),
	.w3(32'h3c1a222b),
	.w4(32'h3bb8d9fc),
	.w5(32'h3aa00c56),
	.w6(32'h3c0e7995),
	.w7(32'h3bb60867),
	.w8(32'h3a303e52),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb7b49),
	.w1(32'h3b154761),
	.w2(32'h381b537d),
	.w3(32'h3b941645),
	.w4(32'h3a2709db),
	.w5(32'hba528aad),
	.w6(32'h3b8ba73a),
	.w7(32'h396f4177),
	.w8(32'hba1ae1fd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c055029),
	.w1(32'h3b24472d),
	.w2(32'hba15eb95),
	.w3(32'h3bde52c4),
	.w4(32'h3b18718c),
	.w5(32'hbb46bcdb),
	.w6(32'h3bb88c83),
	.w7(32'h3abdaefe),
	.w8(32'hbb14da0e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b485d6b),
	.w1(32'h3b01b419),
	.w2(32'h3a749cfb),
	.w3(32'h3aae3a13),
	.w4(32'h3a649331),
	.w5(32'hb9053c04),
	.w6(32'h3a6b7165),
	.w7(32'hba865480),
	.w8(32'hbac56c26),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c468a7a),
	.w1(32'hbaa82f33),
	.w2(32'h39ff858b),
	.w3(32'h3c8764a9),
	.w4(32'h3b318b21),
	.w5(32'h3b0936fd),
	.w6(32'h3c347c0a),
	.w7(32'h3a79d33a),
	.w8(32'hba1965ed),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade6341),
	.w1(32'h3aae7273),
	.w2(32'h3aa20900),
	.w3(32'hbb0c78a3),
	.w4(32'h3acc8a99),
	.w5(32'h3ac6768d),
	.w6(32'hbb0a25c3),
	.w7(32'h3ab77d06),
	.w8(32'h3aff3b15),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed238),
	.w1(32'h3ad7045c),
	.w2(32'h3b007ca6),
	.w3(32'h3ac78c7b),
	.w4(32'h3acb63bf),
	.w5(32'h3ab61ccf),
	.w6(32'h3acccafc),
	.w7(32'h3a54bbbb),
	.w8(32'h3a858a35),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a0ec3),
	.w1(32'hb864b909),
	.w2(32'h38cbe316),
	.w3(32'h3a265908),
	.w4(32'hba193911),
	.w5(32'h3984d969),
	.w6(32'h3993cb48),
	.w7(32'hba5eadd6),
	.w8(32'h39bab5b7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd77b),
	.w1(32'h3a285174),
	.w2(32'hbb5d7078),
	.w3(32'h3bd414c5),
	.w4(32'h3acc9278),
	.w5(32'hbb47e17e),
	.w6(32'h3bd85ebc),
	.w7(32'h3b4b5bdf),
	.w8(32'h399996e7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf8ab8),
	.w1(32'h3a81a9ff),
	.w2(32'h3ad1b22e),
	.w3(32'hb8e7fb10),
	.w4(32'h39b61b5d),
	.w5(32'h3a855c5a),
	.w6(32'hb89d7fed),
	.w7(32'hb7d590e0),
	.w8(32'h3a1454b2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1daf2c),
	.w1(32'h3bd0f74c),
	.w2(32'h3c2e96d5),
	.w3(32'h3c346a9d),
	.w4(32'h3bd0e16d),
	.w5(32'h3beaf871),
	.w6(32'h3b9c2a6a),
	.w7(32'hb9cbfcea),
	.w8(32'h3ab87e55),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1258f),
	.w1(32'hba51c52e),
	.w2(32'hbab584d7),
	.w3(32'h3a37ea27),
	.w4(32'hbaba6847),
	.w5(32'hbacccb11),
	.w6(32'hb8e8cb02),
	.w7(32'hbab2021d),
	.w8(32'hbacfc8ee),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab72b7a),
	.w1(32'h39af1e6e),
	.w2(32'hba082628),
	.w3(32'hbac7a01d),
	.w4(32'hb8eabc26),
	.w5(32'hba5ce348),
	.w6(32'hbab7d0e3),
	.w7(32'hb8708a42),
	.w8(32'hba4835fc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c862c3),
	.w1(32'h3ab56cbd),
	.w2(32'h3ac726bd),
	.w3(32'hb9d502a6),
	.w4(32'h3ad5839a),
	.w5(32'h3b03e73e),
	.w6(32'hba05cb39),
	.w7(32'h3a7a13ec),
	.w8(32'h3ac6c15b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1fbab),
	.w1(32'hbacf1e98),
	.w2(32'hbb04f9d1),
	.w3(32'h3ab6a698),
	.w4(32'hbaff7842),
	.w5(32'hbb1bc414),
	.w6(32'h3a8fe28c),
	.w7(32'hbb11789a),
	.w8(32'hbad73560),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6e032),
	.w1(32'hba87394f),
	.w2(32'hbb4d7258),
	.w3(32'hba3c5d3e),
	.w4(32'hbac6672f),
	.w5(32'hbb59e639),
	.w6(32'hba5420f5),
	.w7(32'hba9732bc),
	.w8(32'hbb29acc0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba011919),
	.w1(32'hba7769b9),
	.w2(32'hba8f5084),
	.w3(32'hb99359d6),
	.w4(32'hb9c678dc),
	.w5(32'hba141434),
	.w6(32'hb8d7a581),
	.w7(32'h389c97d6),
	.w8(32'hba4cbc5e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3137df),
	.w1(32'h3a9c5f4c),
	.w2(32'h3b44fca8),
	.w3(32'h3ba73383),
	.w4(32'h3ac1c330),
	.w5(32'h3a9c703b),
	.w6(32'h3b3d185b),
	.w7(32'hb899126f),
	.w8(32'hba0005cf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4f964),
	.w1(32'h3ad2e24b),
	.w2(32'h3a4657e3),
	.w3(32'hb882c560),
	.w4(32'h398cdf65),
	.w5(32'hb8c1a227),
	.w6(32'h394fa7b7),
	.w7(32'hb7ee4f78),
	.w8(32'h3a9ddf74),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c16b0),
	.w1(32'hba578894),
	.w2(32'hba946ea9),
	.w3(32'hb9fe269f),
	.w4(32'hbaac909c),
	.w5(32'hbaf0f53c),
	.w6(32'hba86377f),
	.w7(32'hba47d36b),
	.w8(32'hbaa033f4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa59e7c),
	.w1(32'h3aadab67),
	.w2(32'h3ae40853),
	.w3(32'hbab370ba),
	.w4(32'h3ab6b457),
	.w5(32'h3af076b7),
	.w6(32'hbaa18fa5),
	.w7(32'h3a52171a),
	.w8(32'h3adfcf4b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e98d4),
	.w1(32'h3af9fbbf),
	.w2(32'h3b18a4ff),
	.w3(32'h3a50f071),
	.w4(32'h3b032346),
	.w5(32'h3b18e6fe),
	.w6(32'h3a8866e5),
	.w7(32'h3aee5f7d),
	.w8(32'h3b238b46),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1c333),
	.w1(32'h3a818578),
	.w2(32'h39cec3c1),
	.w3(32'h3ac233bc),
	.w4(32'h3a690dab),
	.w5(32'h3933d425),
	.w6(32'h3ada45ea),
	.w7(32'h3a4935aa),
	.w8(32'h397a07a3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eead7f),
	.w1(32'hb9b38c37),
	.w2(32'h3b54d076),
	.w3(32'h3a2495d4),
	.w4(32'h3ac3616b),
	.w5(32'h3b9fd378),
	.w6(32'hbad8aab1),
	.w7(32'hbb1596b2),
	.w8(32'h3aa122d9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74d15d),
	.w1(32'h3a6f2e06),
	.w2(32'h3a7be94c),
	.w3(32'h3a9a783f),
	.w4(32'hbb4b4934),
	.w5(32'hbae1cfbe),
	.w6(32'hba049c64),
	.w7(32'hbbaabe5b),
	.w8(32'hbb6f615c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a403611),
	.w1(32'hb982bbc1),
	.w2(32'hbb38862a),
	.w3(32'h3a8ab949),
	.w4(32'hbb67d76c),
	.w5(32'hbb9674ab),
	.w6(32'hbb0166ad),
	.w7(32'hbba32746),
	.w8(32'hbba1fa70),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51f7bf),
	.w1(32'hbc2356fc),
	.w2(32'hbc23fc84),
	.w3(32'hbb72aa57),
	.w4(32'hbc232ccc),
	.w5(32'hbc0696e4),
	.w6(32'hbbd1c333),
	.w7(32'hbc190367),
	.w8(32'hbbbdc05b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fbc49),
	.w1(32'hbb28d8bb),
	.w2(32'hbb1fcbcd),
	.w3(32'hba3eea2b),
	.w4(32'hbb3c99db),
	.w5(32'hbb5deca1),
	.w6(32'hba8fabf5),
	.w7(32'hbb0371e4),
	.w8(32'hbb07fe81),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c92d1),
	.w1(32'h3bb31589),
	.w2(32'h3b7ac60d),
	.w3(32'hbb027f2a),
	.w4(32'h3af82cd5),
	.w5(32'h3b5581f7),
	.w6(32'hbaa79cd2),
	.w7(32'hbb04834a),
	.w8(32'h39c7be5a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6a34c),
	.w1(32'hbb5dba3b),
	.w2(32'hbbaf0e28),
	.w3(32'h3b4dc6de),
	.w4(32'hbabc893c),
	.w5(32'hbb0b9547),
	.w6(32'hba854239),
	.w7(32'hbb163315),
	.w8(32'hbb091e54),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9000d14),
	.w1(32'hbaa6f48a),
	.w2(32'hba7fd168),
	.w3(32'h3af599fc),
	.w4(32'h39806a00),
	.w5(32'hba453767),
	.w6(32'h3ad47a26),
	.w7(32'h3ab5c731),
	.w8(32'h397ee5ab),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1c7a4),
	.w1(32'h3b30e86e),
	.w2(32'h397f7e81),
	.w3(32'hbae1619c),
	.w4(32'h3aab6364),
	.w5(32'h3a470dc2),
	.w6(32'hb8374a1c),
	.w7(32'hbaf0ddb1),
	.w8(32'h3b354510),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55f65b),
	.w1(32'h3b8c8506),
	.w2(32'h3b9a98b1),
	.w3(32'h3b776b6d),
	.w4(32'h3bb745a4),
	.w5(32'h3bdef4d9),
	.w6(32'h3b28f8ac),
	.w7(32'h3a2338ab),
	.w8(32'h3b147d1b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c007b5b),
	.w1(32'hba07b41d),
	.w2(32'h3b05c66b),
	.w3(32'h3c63d1ca),
	.w4(32'hba0afb1b),
	.w5(32'h3b182299),
	.w6(32'h3c21c914),
	.w7(32'hb9c6de7e),
	.w8(32'hbb44717e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb667d7),
	.w1(32'hbb83ddaf),
	.w2(32'hbb9a1fb7),
	.w3(32'h3bc8c802),
	.w4(32'hba71c922),
	.w5(32'hbad79062),
	.w6(32'h3b97b67b),
	.w7(32'h3a480ec0),
	.w8(32'hbb8efcde),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924a370),
	.w1(32'h3928d875),
	.w2(32'h3a6a748a),
	.w3(32'hb8ebde43),
	.w4(32'h39997ca0),
	.w5(32'hba82b866),
	.w6(32'hbb657153),
	.w7(32'h3a81d4ce),
	.w8(32'h3a6fd710),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45af09),
	.w1(32'hbb08fff6),
	.w2(32'hba825b22),
	.w3(32'h3b08aa75),
	.w4(32'hbb243552),
	.w5(32'hbaded33b),
	.w6(32'h3b2d1a3f),
	.w7(32'hbacc4514),
	.w8(32'hba3c2654),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2803f),
	.w1(32'h3b9cec2a),
	.w2(32'h3bb17c9c),
	.w3(32'h399a8fda),
	.w4(32'h3a342dd1),
	.w5(32'hb84614cb),
	.w6(32'hbacf909a),
	.w7(32'h3ba80a4d),
	.w8(32'h3b6f25ff),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c02f5),
	.w1(32'hb9f3a842),
	.w2(32'h39c84575),
	.w3(32'h3bf9ab11),
	.w4(32'h38adbd3a),
	.w5(32'hba1f8655),
	.w6(32'h3c089738),
	.w7(32'h391d2680),
	.w8(32'hbb278c36),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace918b),
	.w1(32'hbaf83f6f),
	.w2(32'hbaec24ab),
	.w3(32'hbb0a4653),
	.w4(32'hba5c05bc),
	.w5(32'hbae94df7),
	.w6(32'hbb0a9d8b),
	.w7(32'h3a04255e),
	.w8(32'h38e1f6b6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66ef54),
	.w1(32'hbabc0814),
	.w2(32'hbb4577d4),
	.w3(32'hbae3319b),
	.w4(32'h3aac7881),
	.w5(32'hba2a2d7f),
	.w6(32'hb9c0441d),
	.w7(32'h38858f5e),
	.w8(32'hbb3472a9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b3f43),
	.w1(32'hba8a9e1a),
	.w2(32'hba8e4796),
	.w3(32'h3a08b6ff),
	.w4(32'hba5da91a),
	.w5(32'hb91a5575),
	.w6(32'hbb0cd7f2),
	.w7(32'hbb370f4f),
	.w8(32'hbb4066a2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb161841),
	.w1(32'hbb678fcd),
	.w2(32'hbaffbc2d),
	.w3(32'h393071e8),
	.w4(32'hbb6a1097),
	.w5(32'h3aeb1fc6),
	.w6(32'hba7d1a68),
	.w7(32'hbac49c7f),
	.w8(32'h3a3d6da7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1c01),
	.w1(32'hbafeae41),
	.w2(32'hbad7fdba),
	.w3(32'hbbb10039),
	.w4(32'hbae6dd91),
	.w5(32'hba8887b4),
	.w6(32'hbb865922),
	.w7(32'hba4b72fd),
	.w8(32'hbb0d35ba),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca92a0),
	.w1(32'h3a1210fb),
	.w2(32'h386d8ad2),
	.w3(32'hbb1f82d4),
	.w4(32'h3ae5092d),
	.w5(32'h3abb8529),
	.w6(32'hbb122311),
	.w7(32'h3989cf80),
	.w8(32'hba040aea),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ec514),
	.w1(32'hb983e27b),
	.w2(32'h3afee751),
	.w3(32'hbae1d055),
	.w4(32'h3830dec9),
	.w5(32'h3a364690),
	.w6(32'hbad365b4),
	.w7(32'hb992c310),
	.w8(32'h3adabe86),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3002cc),
	.w1(32'hbb311c9c),
	.w2(32'h3b77684a),
	.w3(32'h3b8577b7),
	.w4(32'hb8129c0d),
	.w5(32'h3b2aed27),
	.w6(32'h3b6047ad),
	.w7(32'hbac78ce4),
	.w8(32'hba45cd53),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a804db8),
	.w1(32'hbb05a810),
	.w2(32'hbb97ba73),
	.w3(32'hbab1ce02),
	.w4(32'hbac2e73a),
	.w5(32'hbabee8f7),
	.w6(32'hbb63e412),
	.w7(32'hbb280807),
	.w8(32'hbb9fa711),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36653f),
	.w1(32'h3b63e1e3),
	.w2(32'h3ac87dc0),
	.w3(32'h3b2f0e3a),
	.w4(32'h3c187611),
	.w5(32'h3b9648f0),
	.w6(32'h3a821312),
	.w7(32'h3abea2fc),
	.w8(32'h3b366267),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45a215),
	.w1(32'h3abdd83f),
	.w2(32'hbaa00716),
	.w3(32'h3ac327bb),
	.w4(32'hbafb6365),
	.w5(32'hb7a0f9e0),
	.w6(32'hb940ee11),
	.w7(32'hba9cfe5b),
	.w8(32'h3b52cd2e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77ad0c),
	.w1(32'h3b7e6339),
	.w2(32'h3bd21429),
	.w3(32'h3b18591e),
	.w4(32'h3acdf738),
	.w5(32'h3b0b6ee5),
	.w6(32'h3ab692c2),
	.w7(32'hbacce2be),
	.w8(32'h3a228b33),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1f856),
	.w1(32'hbae89160),
	.w2(32'hbb32cc52),
	.w3(32'hba545634),
	.w4(32'hba94f2a7),
	.w5(32'hbadfe254),
	.w6(32'hba840063),
	.w7(32'hbaea6828),
	.w8(32'hba6555b6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f9216),
	.w1(32'hbb125618),
	.w2(32'hbb8bbde9),
	.w3(32'h3a899f23),
	.w4(32'hbb85f7f4),
	.w5(32'hbb5fcb8b),
	.w6(32'h398834ba),
	.w7(32'hbb6910c5),
	.w8(32'hbb3b4281),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98cf8e),
	.w1(32'hba41abdc),
	.w2(32'hbaf972c1),
	.w3(32'hbb901c2e),
	.w4(32'h3ab4764c),
	.w5(32'hbb05b154),
	.w6(32'hbb609d53),
	.w7(32'h38f613e8),
	.w8(32'hbb323167),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd40ab8),
	.w1(32'h384aeccb),
	.w2(32'h3a974e7d),
	.w3(32'h3bba0c74),
	.w4(32'h3a159ec6),
	.w5(32'h3b40de5f),
	.w6(32'h3b90e0fc),
	.w7(32'hbab66b6b),
	.w8(32'h3869d564),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db9f66),
	.w1(32'h3aa5ade6),
	.w2(32'hbab4f9a8),
	.w3(32'h3b22174a),
	.w4(32'h39beab81),
	.w5(32'hbb0a7967),
	.w6(32'hbbdb287c),
	.w7(32'hbb7f7c18),
	.w8(32'hbb8c4030),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae67f15),
	.w1(32'h38373e3e),
	.w2(32'h3b85fa5d),
	.w3(32'h3b3a233f),
	.w4(32'h3b05d770),
	.w5(32'hb9a88c89),
	.w6(32'h3a5e66af),
	.w7(32'hba24661e),
	.w8(32'hbadc29b9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc051286),
	.w1(32'hbbe02ac3),
	.w2(32'hbc6268f4),
	.w3(32'hbc014c8f),
	.w4(32'hbafcb7d8),
	.w5(32'hbc300070),
	.w6(32'hbc3945a5),
	.w7(32'hbb1a7ddd),
	.w8(32'hbc0be68c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92605d),
	.w1(32'h3afbfdb3),
	.w2(32'h3ae95d1b),
	.w3(32'h3ab570d2),
	.w4(32'h3b269434),
	.w5(32'h3b9269e9),
	.w6(32'h39d0b989),
	.w7(32'h3b6bb39e),
	.w8(32'h3ad15152),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba31486),
	.w1(32'h3a05ef76),
	.w2(32'hb8771fdd),
	.w3(32'h3c190542),
	.w4(32'h3a662952),
	.w5(32'hba5cfd12),
	.w6(32'h3b8279af),
	.w7(32'hbaac44c7),
	.w8(32'hbb68e9a8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64005c),
	.w1(32'hbb350e18),
	.w2(32'hba295d40),
	.w3(32'hbaefa146),
	.w4(32'hbb7749c3),
	.w5(32'hbb023b8a),
	.w6(32'hbb31f499),
	.w7(32'hbb1440dd),
	.w8(32'hbb093a97),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35061f),
	.w1(32'h3b8c24ef),
	.w2(32'h3bcd4c64),
	.w3(32'h398167e9),
	.w4(32'hbaee9ee5),
	.w5(32'h3abeb0a5),
	.w6(32'hbbdfb859),
	.w7(32'hbb9244de),
	.w8(32'hbb71c074),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fca2a),
	.w1(32'h3b0a96e1),
	.w2(32'hbb25725f),
	.w3(32'h3be8d7dd),
	.w4(32'h3af489e3),
	.w5(32'hbb3973cc),
	.w6(32'h3bb6a781),
	.w7(32'hb89b08be),
	.w8(32'hbb8d9cf8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e41f3),
	.w1(32'hbb269fa2),
	.w2(32'hbb76a48d),
	.w3(32'hba780880),
	.w4(32'hba8f6f5d),
	.w5(32'hbb17db9d),
	.w6(32'h37e31e83),
	.w7(32'hb9f303be),
	.w8(32'hb9ca5057),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafe2cb),
	.w1(32'h3963fe1f),
	.w2(32'hba5d4cc9),
	.w3(32'hba3d868a),
	.w4(32'hba49aeb6),
	.w5(32'h38dd56d6),
	.w6(32'h39c42706),
	.w7(32'hbb339b60),
	.w8(32'hbad073d4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be038f5),
	.w1(32'h3b4535fa),
	.w2(32'hba42353a),
	.w3(32'h3c0b3060),
	.w4(32'h3b4b041f),
	.w5(32'h3b06adc6),
	.w6(32'h3be383ce),
	.w7(32'h3b158d9e),
	.w8(32'hbb26d25c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87f700),
	.w1(32'h3c096c78),
	.w2(32'h3b5ccaf1),
	.w3(32'h3ba5e9c2),
	.w4(32'h3bbffc7c),
	.w5(32'h3c157d5f),
	.w6(32'h3b12a62b),
	.w7(32'hba906ac7),
	.w8(32'h3ae8bfdc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94b79c),
	.w1(32'hba358b39),
	.w2(32'h39b8c0a2),
	.w3(32'h3b995671),
	.w4(32'h3b07c6aa),
	.w5(32'h3bc907fa),
	.w6(32'hbaa3a296),
	.w7(32'h3b1ce75c),
	.w8(32'h3b2642d2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cd14d),
	.w1(32'hbaed3424),
	.w2(32'h3aded83b),
	.w3(32'h3b84c53d),
	.w4(32'hbad3fd6c),
	.w5(32'h3a020002),
	.w6(32'hba5de87c),
	.w7(32'h3aa99ebd),
	.w8(32'h3aab1797),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56da33),
	.w1(32'h3a400bee),
	.w2(32'hbb4b43af),
	.w3(32'h3ad24daa),
	.w4(32'h39eb4514),
	.w5(32'hbb43d41e),
	.w6(32'hbae7d235),
	.w7(32'h3ac203e3),
	.w8(32'h3a4191ec),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80a924),
	.w1(32'hba5bc373),
	.w2(32'h38a5488f),
	.w3(32'h3ae9752d),
	.w4(32'h3b3e2e7e),
	.w5(32'hba8434df),
	.w6(32'h3b7d8bf3),
	.w7(32'h3a0de93b),
	.w8(32'hba32104c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e1bf3),
	.w1(32'hba808f0a),
	.w2(32'hbb75bbe8),
	.w3(32'h3aac65b9),
	.w4(32'hb942809b),
	.w5(32'hbb54bbef),
	.w6(32'h3b712e34),
	.w7(32'hba93cee6),
	.w8(32'h38927983),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44c067),
	.w1(32'hba22e28f),
	.w2(32'hbb085a86),
	.w3(32'hbb5714b9),
	.w4(32'hb89e3715),
	.w5(32'hbb64e2a6),
	.w6(32'h37983e65),
	.w7(32'hb9a7dc67),
	.w8(32'hbb13c6bd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc4493),
	.w1(32'h3abe94cf),
	.w2(32'hba4cdf08),
	.w3(32'hba6cbe03),
	.w4(32'h3b16e1c7),
	.w5(32'h3a55a12c),
	.w6(32'hba4d8b9f),
	.w7(32'hbb1fb9b3),
	.w8(32'hbadb80c0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa47c93),
	.w1(32'h3b540e84),
	.w2(32'h3baef840),
	.w3(32'h3adca29d),
	.w4(32'h3b9d87c4),
	.w5(32'h3bb5cae1),
	.w6(32'h3a369721),
	.w7(32'h3b23c58b),
	.w8(32'h3bb22681),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eda17),
	.w1(32'h392633fd),
	.w2(32'hba230e81),
	.w3(32'h3b2a321e),
	.w4(32'hba7241ef),
	.w5(32'hba50d45f),
	.w6(32'h3afb5da3),
	.w7(32'h39c2af43),
	.w8(32'hba62dcb5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97ba9b),
	.w1(32'h3ba8b7fc),
	.w2(32'h3aa81327),
	.w3(32'h3b053012),
	.w4(32'h3982a641),
	.w5(32'h394a5971),
	.w6(32'hb7fbd50a),
	.w7(32'hb933646b),
	.w8(32'hb9f16504),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad7e83),
	.w1(32'hb7224c97),
	.w2(32'h37d93d8e),
	.w3(32'h3a419780),
	.w4(32'h3ac89286),
	.w5(32'h3a7002a6),
	.w6(32'h3a8740ab),
	.w7(32'h3a886d43),
	.w8(32'h3ad63ef2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9259b),
	.w1(32'hba4bd862),
	.w2(32'hb9fcd10b),
	.w3(32'h3bb8987c),
	.w4(32'hba7826a9),
	.w5(32'hbb8f27c4),
	.w6(32'h3b93b155),
	.w7(32'hbaea00a4),
	.w8(32'hbaae3f72),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95aa5a),
	.w1(32'hbb96c5cc),
	.w2(32'hbbd91567),
	.w3(32'hbb97808f),
	.w4(32'hbb64fc94),
	.w5(32'hbbf7481b),
	.w6(32'hba18450e),
	.w7(32'hbaaf450a),
	.w8(32'hbb2951e2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04f37c),
	.w1(32'h3b5a10b3),
	.w2(32'h3bc997d7),
	.w3(32'hbb3a5481),
	.w4(32'h3af26982),
	.w5(32'h3b859c11),
	.w6(32'hbaf2edea),
	.w7(32'h3b90a63e),
	.w8(32'h3b16a15c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26ba4f),
	.w1(32'h3bfab804),
	.w2(32'h3ba7b587),
	.w3(32'h3b20bfaa),
	.w4(32'h3ba4dd26),
	.w5(32'h3bcdd3b5),
	.w6(32'h3b164534),
	.w7(32'h3b09bc9c),
	.w8(32'h3b356738),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b443252),
	.w1(32'h3b45e250),
	.w2(32'h3aacbbf5),
	.w3(32'h3bb63f05),
	.w4(32'h3b037c55),
	.w5(32'h3b47d6fc),
	.w6(32'h3b0eab38),
	.w7(32'hba00bdfd),
	.w8(32'h3b014460),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8aa66),
	.w1(32'hbba33dbb),
	.w2(32'hbb8dbcc2),
	.w3(32'h3b955bb7),
	.w4(32'hba836b62),
	.w5(32'hba1193ad),
	.w6(32'h3a9a889a),
	.w7(32'h39ea4a22),
	.w8(32'h3a9ea24d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b797d3e),
	.w1(32'h3ba15bb9),
	.w2(32'h3b9a0561),
	.w3(32'h3baccc4a),
	.w4(32'h3ad99504),
	.w5(32'hb9b48fd1),
	.w6(32'h3b4eb924),
	.w7(32'h3785a1e5),
	.w8(32'h3b027f05),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e9866),
	.w1(32'h3b8bfa04),
	.w2(32'h3bc46ee4),
	.w3(32'h3b3e2955),
	.w4(32'h3b3bbb16),
	.w5(32'h3ba9637e),
	.w6(32'h3bb0429e),
	.w7(32'h3a5b5ad3),
	.w8(32'h3b05c2c0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389dfa5c),
	.w1(32'hbb4ba1c5),
	.w2(32'hbaa02194),
	.w3(32'h3ab265ff),
	.w4(32'hbad5dc89),
	.w5(32'hb9b02146),
	.w6(32'hba5b5b34),
	.w7(32'hbb537800),
	.w8(32'hbacb1957),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d163c),
	.w1(32'h3b815b0f),
	.w2(32'hbaa2a617),
	.w3(32'hba726819),
	.w4(32'h3b9f65cd),
	.w5(32'h3b451a2e),
	.w6(32'hbb150bb9),
	.w7(32'hbb338811),
	.w8(32'hbb8c876b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f3ded),
	.w1(32'hb9eb1ad2),
	.w2(32'hba8e9457),
	.w3(32'hb90488a1),
	.w4(32'hbb101658),
	.w5(32'hbb800b1d),
	.w6(32'h3a05bb1f),
	.w7(32'hbb584770),
	.w8(32'hba8d328e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b9656),
	.w1(32'h3ad37437),
	.w2(32'h3b328dd2),
	.w3(32'hb98ac96f),
	.w4(32'h3a906f9c),
	.w5(32'h3b84ce95),
	.w6(32'h3abb04fa),
	.w7(32'h3af92e72),
	.w8(32'h3a941acf),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb780a3e),
	.w1(32'hbb79ee46),
	.w2(32'hbb036018),
	.w3(32'h3a07a614),
	.w4(32'h39a40edc),
	.w5(32'hbae80f98),
	.w6(32'hba418bda),
	.w7(32'h39629aad),
	.w8(32'hb8f05853),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ab335),
	.w1(32'h3c14d155),
	.w2(32'h3bda305a),
	.w3(32'h3bf859cc),
	.w4(32'h3b4090cb),
	.w5(32'h3bbc3510),
	.w6(32'h3bb05f97),
	.w7(32'hbaebb19c),
	.w8(32'h3ac97892),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf5c99),
	.w1(32'hbb85ac29),
	.w2(32'hbbc29692),
	.w3(32'hb9940472),
	.w4(32'hbb1f0fb4),
	.w5(32'hbbc0956d),
	.w6(32'h38e33d83),
	.w7(32'hbb4c103f),
	.w8(32'hbb62066c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384d005a),
	.w1(32'h3ae1282e),
	.w2(32'h3b38f2ba),
	.w3(32'hbb12128d),
	.w4(32'hba352d85),
	.w5(32'hbb6c1f3c),
	.w6(32'hbb40835b),
	.w7(32'hb9dc90b2),
	.w8(32'hba6502b4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c000057),
	.w1(32'h3b958e41),
	.w2(32'h3bb5ec36),
	.w3(32'h3bae21aa),
	.w4(32'h3b3924a0),
	.w5(32'h3b160d45),
	.w6(32'h3b292d15),
	.w7(32'hbba70cdc),
	.w8(32'h3b406fbd),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc5594),
	.w1(32'h3bc4423c),
	.w2(32'h3b8d7fd9),
	.w3(32'h3b589b8b),
	.w4(32'h3ab639bd),
	.w5(32'h3a81885f),
	.w6(32'h399f86cb),
	.w7(32'hbb80f15c),
	.w8(32'hbb8ac210),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd837ba),
	.w1(32'h3a36706f),
	.w2(32'h3b347d11),
	.w3(32'h3bd334d7),
	.w4(32'h3ac2aa5e),
	.w5(32'h3a3acabe),
	.w6(32'h3b1cc3cc),
	.w7(32'hb6814853),
	.w8(32'hb90c1143),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab03321),
	.w1(32'hba2a0feb),
	.w2(32'hba22ec56),
	.w3(32'h3a98e520),
	.w4(32'h398b71f7),
	.w5(32'hbb0d0496),
	.w6(32'h3a17ec5a),
	.w7(32'h3b0324d5),
	.w8(32'h3a3bb9d3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84e215),
	.w1(32'hbb69bfa4),
	.w2(32'hbb99c21e),
	.w3(32'hbb8ca5b7),
	.w4(32'hbbc8618d),
	.w5(32'hbb8e3083),
	.w6(32'hba734750),
	.w7(32'hbb139ff5),
	.w8(32'hbb150ea5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55b724),
	.w1(32'hbacbb7ab),
	.w2(32'hba8485d0),
	.w3(32'hbbc36925),
	.w4(32'h39545184),
	.w5(32'h3af23eeb),
	.w6(32'hbbc6d565),
	.w7(32'hb98e5516),
	.w8(32'hbb171b76),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad96de8),
	.w1(32'hbaa902e8),
	.w2(32'hbab28bda),
	.w3(32'hb994c3a6),
	.w4(32'hb9299e5f),
	.w5(32'h38d0c070),
	.w6(32'hbaefe83a),
	.w7(32'h36371edb),
	.w8(32'hba5d79b3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dad163),
	.w1(32'h3aecf172),
	.w2(32'h3a93c892),
	.w3(32'h3a16cf3c),
	.w4(32'h3b4e8fb2),
	.w5(32'h3b565713),
	.w6(32'h3930589e),
	.w7(32'h3a7158d8),
	.w8(32'h3b0750ab),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c4993),
	.w1(32'hbaaa2e31),
	.w2(32'hbacfb381),
	.w3(32'h3b36b773),
	.w4(32'hbaa12dc0),
	.w5(32'hba3ce229),
	.w6(32'h3a5fad70),
	.w7(32'hbb19f9a1),
	.w8(32'hba1f0189),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb49c8),
	.w1(32'hbb392c04),
	.w2(32'h3a9b2de9),
	.w3(32'hbba3a597),
	.w4(32'hbb7e4306),
	.w5(32'hbb1eb44b),
	.w6(32'hbbb3afa7),
	.w7(32'hbb0ce432),
	.w8(32'hbb911c6c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b6b2e),
	.w1(32'hbb0d83e2),
	.w2(32'hbb21af55),
	.w3(32'h3c3e5e18),
	.w4(32'h3c02defc),
	.w5(32'h3a657547),
	.w6(32'h3c2185ea),
	.w7(32'h3ba0763a),
	.w8(32'hbb577fa4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a3fd5),
	.w1(32'hbaa692f2),
	.w2(32'hbabf0e9e),
	.w3(32'hba998c1e),
	.w4(32'h3ac5f3e6),
	.w5(32'h39000c01),
	.w6(32'hbb12a299),
	.w7(32'h3afa43d3),
	.w8(32'h394e337a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40b405),
	.w1(32'hbb3559f1),
	.w2(32'hbaf12599),
	.w3(32'h3b602f9c),
	.w4(32'hbad87a78),
	.w5(32'hbab759bc),
	.w6(32'h3b65bc41),
	.w7(32'hbadb247f),
	.w8(32'hbb26e9c4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39813bd9),
	.w1(32'hbaf438c7),
	.w2(32'hbacf7646),
	.w3(32'h3af44bc9),
	.w4(32'hba26116b),
	.w5(32'h38d70d68),
	.w6(32'hb9175926),
	.w7(32'hb808a1fd),
	.w8(32'h3b19caac),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb4b0a),
	.w1(32'h39db66de),
	.w2(32'h3ab01917),
	.w3(32'h3c2fe8e9),
	.w4(32'h3ad002ae),
	.w5(32'h3b31aa88),
	.w6(32'h3bafcf56),
	.w7(32'hbb5281ca),
	.w8(32'hb8ce0774),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5839d0),
	.w1(32'hbb41a0aa),
	.w2(32'hbb1f230f),
	.w3(32'hbacdc347),
	.w4(32'hbac140fb),
	.w5(32'h3ae6993d),
	.w6(32'hbae195fb),
	.w7(32'hbb821e5d),
	.w8(32'hbabd966d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe529a4),
	.w1(32'hbb835676),
	.w2(32'hbb9ef959),
	.w3(32'hbb76bcaf),
	.w4(32'hbba5bffa),
	.w5(32'hbb933b9d),
	.w6(32'hbb54d793),
	.w7(32'hba9e5cfc),
	.w8(32'hb9e7c1c2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17eba8),
	.w1(32'hbaa5030a),
	.w2(32'hbaf51085),
	.w3(32'hba482d9b),
	.w4(32'hba8f2815),
	.w5(32'hbb34f7f1),
	.w6(32'h3a8528b4),
	.w7(32'hba50aa0b),
	.w8(32'h3a12f586),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8780a0),
	.w1(32'h3b61db8a),
	.w2(32'hbaa1c500),
	.w3(32'h3b02c9ab),
	.w4(32'h3a5f8c8b),
	.w5(32'hbb8fd124),
	.w6(32'h3b045333),
	.w7(32'hbb1b2d75),
	.w8(32'hbbab1a93),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf66314),
	.w1(32'hbad846a8),
	.w2(32'hbb8a1223),
	.w3(32'hbc1fccda),
	.w4(32'hbb95ac8c),
	.w5(32'hbba4cc33),
	.w6(32'hbc200f69),
	.w7(32'hbbb0cd44),
	.w8(32'hbb8caf69),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ecdc1),
	.w1(32'hbb4b69df),
	.w2(32'hbb80cc39),
	.w3(32'hbb8aaea2),
	.w4(32'hbb321c1f),
	.w5(32'hbb3a62ed),
	.w6(32'hbb828ecf),
	.w7(32'hb9a253bd),
	.w8(32'hba6ca5eb),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b1950),
	.w1(32'h3b1a1496),
	.w2(32'h3b7219f8),
	.w3(32'hba13a95c),
	.w4(32'h3a98b8e8),
	.w5(32'h3b28d9fe),
	.w6(32'hba7f22af),
	.w7(32'hba8524f5),
	.w8(32'h3b25a9b0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab11401),
	.w1(32'h3aef97bb),
	.w2(32'hba438c53),
	.w3(32'h3aef6c80),
	.w4(32'h3aaed18e),
	.w5(32'h35673565),
	.w6(32'h3a916d82),
	.w7(32'hb8c3ccf8),
	.w8(32'h37f0ffe4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eedd0),
	.w1(32'hbb02a8d5),
	.w2(32'h3aa3d314),
	.w3(32'h3b17916b),
	.w4(32'hba5343c4),
	.w5(32'h3a2bd45e),
	.w6(32'h3aafe454),
	.w7(32'hb8a002f5),
	.w8(32'hbad6069d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad628d0),
	.w1(32'hbaa634f0),
	.w2(32'hba648376),
	.w3(32'hbb80a1ff),
	.w4(32'hbaeff2a3),
	.w5(32'hbadc54ff),
	.w6(32'hbb185df8),
	.w7(32'h39b6329f),
	.w8(32'hba2352ea),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ea10e),
	.w1(32'hbb40fecb),
	.w2(32'hbb3205cb),
	.w3(32'h399e2452),
	.w4(32'hbb7ff0f0),
	.w5(32'hbba60911),
	.w6(32'hbaa89cf4),
	.w7(32'hb8dae61d),
	.w8(32'hb98206ae),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d4689),
	.w1(32'h3b1dad20),
	.w2(32'h3aee7ae3),
	.w3(32'hbb44763f),
	.w4(32'h3aec513c),
	.w5(32'h3acbb596),
	.w6(32'hbac171a3),
	.w7(32'hba0b6654),
	.w8(32'h3acd1412),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab3ccb),
	.w1(32'hb9f6e9b7),
	.w2(32'h3a87ee38),
	.w3(32'h3a5b7053),
	.w4(32'hba3d7a9f),
	.w5(32'h3b03ef23),
	.w6(32'hbb56d499),
	.w7(32'hbbc820d9),
	.w8(32'hbb3831f4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbaef8),
	.w1(32'h3ae06ef4),
	.w2(32'h3a54febf),
	.w3(32'h3ba34f26),
	.w4(32'h3b13d19e),
	.w5(32'h3ab71b72),
	.w6(32'h3abdf49a),
	.w7(32'h3a32cea8),
	.w8(32'h3ac270b7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9357f9),
	.w1(32'h3b8e3ea2),
	.w2(32'h3a1af32b),
	.w3(32'hb9aa8e4a),
	.w4(32'h3a7a6ef3),
	.w5(32'h3a3d52a4),
	.w6(32'hb94f7b46),
	.w7(32'hbaf259f9),
	.w8(32'hbae58008),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf83274),
	.w1(32'h3a5eb58f),
	.w2(32'hb84bbbea),
	.w3(32'hbad249aa),
	.w4(32'h3aba8fec),
	.w5(32'hb9ecdf01),
	.w6(32'hbb1270d3),
	.w7(32'hbaa30a18),
	.w8(32'hba34cd96),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2441be),
	.w1(32'h3c126235),
	.w2(32'h3be8381a),
	.w3(32'h3beee9ab),
	.w4(32'h3b6e8fde),
	.w5(32'h3b045575),
	.w6(32'h3ba4d510),
	.w7(32'h3b61505b),
	.w8(32'h3b043b77),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8322e1c),
	.w1(32'h3a4b1774),
	.w2(32'hba1c0624),
	.w3(32'hbaf5338d),
	.w4(32'h39d411e6),
	.w5(32'hbb22874b),
	.w6(32'h3ad4e725),
	.w7(32'hb9e4ed53),
	.w8(32'hbb167421),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a32c5),
	.w1(32'hbb06c04f),
	.w2(32'hbb4ef59c),
	.w3(32'h3b8fdbba),
	.w4(32'hbb2d7f15),
	.w5(32'hbba7ff6b),
	.w6(32'h3b91b7c1),
	.w7(32'hb8e08d70),
	.w8(32'h3a9151a6),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fd125),
	.w1(32'hba29eb3c),
	.w2(32'hba2ad2c2),
	.w3(32'hba0e3e66),
	.w4(32'hb9929029),
	.w5(32'hba116508),
	.w6(32'h3a74b50e),
	.w7(32'hb9c5de9c),
	.w8(32'hbb2061e7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcec96),
	.w1(32'hb9c4f086),
	.w2(32'hba8a5aa9),
	.w3(32'h3baf134a),
	.w4(32'hbab4d835),
	.w5(32'hbb9af1b8),
	.w6(32'h3a57d633),
	.w7(32'hbb158908),
	.w8(32'hbba09a5b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb251cf7),
	.w1(32'hbb23103d),
	.w2(32'hbbad5386),
	.w3(32'hb94a3c35),
	.w4(32'hbb843a51),
	.w5(32'hbb5d9e08),
	.w6(32'hb7cb1a7b),
	.w7(32'hbb904057),
	.w8(32'hbba911b1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba75aef),
	.w1(32'h3be62682),
	.w2(32'h3bd7c501),
	.w3(32'h3ba3312d),
	.w4(32'h3abdc727),
	.w5(32'h3b5e5890),
	.w6(32'h3b1c2e56),
	.w7(32'hba454b40),
	.w8(32'h3b171ed6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6417d2),
	.w1(32'h3af4b465),
	.w2(32'hb980c55b),
	.w3(32'h3abd4cb8),
	.w4(32'hb88d46df),
	.w5(32'hba146dfe),
	.w6(32'h3b1bc900),
	.w7(32'h3a835015),
	.w8(32'hba0d547c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01975b),
	.w1(32'h3a718ecf),
	.w2(32'h3ba87625),
	.w3(32'h3a0fd3ec),
	.w4(32'hba943055),
	.w5(32'h3af1ad5b),
	.w6(32'h390d8ff9),
	.w7(32'hbb2ebd47),
	.w8(32'hba3db71a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c80de),
	.w1(32'h3b0cdd18),
	.w2(32'h3aac7bd9),
	.w3(32'h3a9935f9),
	.w4(32'h3b0c7c56),
	.w5(32'h3b813619),
	.w6(32'hb9d5114f),
	.w7(32'hb9742515),
	.w8(32'h3af9972c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad74a6e),
	.w1(32'hba231eb6),
	.w2(32'h3a816d41),
	.w3(32'h3b3d95f5),
	.w4(32'hb94f40d3),
	.w5(32'h3aa0e550),
	.w6(32'h39f9dc9c),
	.w7(32'h39a5d7c1),
	.w8(32'h3b2bb16e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5a607),
	.w1(32'hbac50313),
	.w2(32'hb9a2d82a),
	.w3(32'hbb381460),
	.w4(32'hbb061555),
	.w5(32'hb9bb28bc),
	.w6(32'hbab54b43),
	.w7(32'hbab616da),
	.w8(32'hb9be1a4a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a317930),
	.w1(32'h38b671b9),
	.w2(32'hba96a4d1),
	.w3(32'h3b822acc),
	.w4(32'hba8c8865),
	.w5(32'hbb0033e8),
	.w6(32'h3a8e4fb5),
	.w7(32'h3a9f0e3a),
	.w8(32'hba92df81),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a82c6),
	.w1(32'hbb8e35f9),
	.w2(32'hbb1ba01d),
	.w3(32'hba5f3d0d),
	.w4(32'hbb24b570),
	.w5(32'hbb54323f),
	.w6(32'hbac5c698),
	.w7(32'hba42f49c),
	.w8(32'hbb5ccf09),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2524f8),
	.w1(32'h3a1b8ec0),
	.w2(32'hbaa58667),
	.w3(32'hbba4b835),
	.w4(32'h3a3aeca5),
	.w5(32'h39afde06),
	.w6(32'hbb769a4e),
	.w7(32'h399120d4),
	.w8(32'hb8917d29),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec1e3f),
	.w1(32'hbb66a673),
	.w2(32'hbac85ce8),
	.w3(32'h3b4d4a0a),
	.w4(32'hbb84a250),
	.w5(32'hbb2588e6),
	.w6(32'h38c843f2),
	.w7(32'hbbb141b9),
	.w8(32'hbb5add9f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64634c),
	.w1(32'h3b181ed2),
	.w2(32'h3af01652),
	.w3(32'h3b14454e),
	.w4(32'h3ac99857),
	.w5(32'hbb2de1ae),
	.w6(32'hbad201d3),
	.w7(32'h3a471fa1),
	.w8(32'h3a01554a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94cda0),
	.w1(32'hbb141366),
	.w2(32'hbb2ce663),
	.w3(32'hba40ffd4),
	.w4(32'hba0a4df4),
	.w5(32'h35fd55f4),
	.w6(32'hba41f9b9),
	.w7(32'h3a562441),
	.w8(32'h3a433f75),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacba942),
	.w1(32'h3aebca64),
	.w2(32'hbab2a068),
	.w3(32'hbae6d341),
	.w4(32'h3b04457d),
	.w5(32'hb94868a9),
	.w6(32'hb97965a0),
	.w7(32'h3a9f61b7),
	.w8(32'hb87e6d0a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2bcfc),
	.w1(32'h3c1dba8f),
	.w2(32'h3bd22dd5),
	.w3(32'h3cdb4335),
	.w4(32'h3c2d2715),
	.w5(32'h3b7b76d4),
	.w6(32'h3c5a6036),
	.w7(32'hbb0373cb),
	.w8(32'hbbb561f8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90557d),
	.w1(32'hbbbbb805),
	.w2(32'hbbe32809),
	.w3(32'hbbc374e2),
	.w4(32'hbb847897),
	.w5(32'hbb0ee544),
	.w6(32'hbc04feb3),
	.w7(32'h39e3ec31),
	.w8(32'h3a8a428f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79c880),
	.w1(32'h3a049dfb),
	.w2(32'hbaab35d2),
	.w3(32'hb977ebb1),
	.w4(32'hbac14195),
	.w5(32'hba56de3c),
	.w6(32'hba9336d5),
	.w7(32'hbb4c7fcb),
	.w8(32'hbb9412eb),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d6f9d),
	.w1(32'hba398cbd),
	.w2(32'hbb224b34),
	.w3(32'hbae5b554),
	.w4(32'h3953f22c),
	.w5(32'hb9b1d40e),
	.w6(32'hbb5efbd2),
	.w7(32'hb8dda12b),
	.w8(32'h3a641af8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8109f6),
	.w1(32'h371988e0),
	.w2(32'h380a95f3),
	.w3(32'hba82249b),
	.w4(32'hbaa54ca3),
	.w5(32'hbb0ca431),
	.w6(32'h38f32ccc),
	.w7(32'h3a8be50b),
	.w8(32'h398c18da),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabcf97),
	.w1(32'h3b1f5594),
	.w2(32'h3b70821d),
	.w3(32'hba8f4897),
	.w4(32'h3a99dae9),
	.w5(32'h3aceadee),
	.w6(32'h39fc938a),
	.w7(32'h3b53db11),
	.w8(32'h3b7c803d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b593e63),
	.w1(32'h3b574d21),
	.w2(32'h3b343920),
	.w3(32'h3b4ec489),
	.w4(32'h3b8d3bc5),
	.w5(32'h3b50c877),
	.w6(32'h3b30907a),
	.w7(32'h3a7af15c),
	.w8(32'h3a30c176),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2583f5),
	.w1(32'h3ba68b23),
	.w2(32'h3bbdd24d),
	.w3(32'h3b5a083e),
	.w4(32'h3b5f967c),
	.w5(32'h3b1478d5),
	.w6(32'hba6036df),
	.w7(32'hba3d21f9),
	.w8(32'hba415681),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9efcb8),
	.w1(32'hbb3f9095),
	.w2(32'hba325549),
	.w3(32'h3b813ce0),
	.w4(32'hb9cd66ec),
	.w5(32'hba4a79db),
	.w6(32'h3ba593e8),
	.w7(32'h3a0e1288),
	.w8(32'hbb312376),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08d5e9),
	.w1(32'hba9e97a9),
	.w2(32'hbadb095a),
	.w3(32'hbb676c2b),
	.w4(32'hb9bf63f2),
	.w5(32'h3933b716),
	.w6(32'hbbb1f6fa),
	.w7(32'hbacbd271),
	.w8(32'hba679d83),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd905cb),
	.w1(32'h3b34b17f),
	.w2(32'hbc03d8bf),
	.w3(32'h3c03fe0d),
	.w4(32'h3b5ae537),
	.w5(32'h39f3db48),
	.w6(32'h3bcdd1eb),
	.w7(32'h39774bbe),
	.w8(32'h3b2f98ef),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3015c),
	.w1(32'h3b249814),
	.w2(32'h3b06cfa9),
	.w3(32'hbaabc0bb),
	.w4(32'h3c065995),
	.w5(32'hbb6e53bf),
	.w6(32'h3b262bc3),
	.w7(32'h3b8e4296),
	.w8(32'h3b9975e8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26c101),
	.w1(32'hbb0bc511),
	.w2(32'hbaa64744),
	.w3(32'h3b27879e),
	.w4(32'hbbdc621c),
	.w5(32'hbc8b29fb),
	.w6(32'h3b37a7de),
	.w7(32'h3b802924),
	.w8(32'h3b5d5ec3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbe226),
	.w1(32'hbbdbbbd5),
	.w2(32'hbc43f388),
	.w3(32'hbbccb1eb),
	.w4(32'hbc173d7b),
	.w5(32'hbc4a3a87),
	.w6(32'h391468aa),
	.w7(32'hbc0d7375),
	.w8(32'hbbb430ab),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf94f88),
	.w1(32'h3a925d5a),
	.w2(32'h3aeaa64a),
	.w3(32'hba34913e),
	.w4(32'hbb2beb8e),
	.w5(32'hbbc48ac5),
	.w6(32'h3b1de9ae),
	.w7(32'h3a1f2255),
	.w8(32'hbbd8c5e7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f800d),
	.w1(32'hbab69fdb),
	.w2(32'h3af85be5),
	.w3(32'h3b1f6a23),
	.w4(32'hbbc34af2),
	.w5(32'hbc5b5283),
	.w6(32'h3ad6a7f8),
	.w7(32'hbbf3c09d),
	.w8(32'hbbe52339),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e2549),
	.w1(32'hbbef0ee0),
	.w2(32'hbc3dac32),
	.w3(32'hbb93df95),
	.w4(32'hbb9a0a03),
	.w5(32'hbbdafc48),
	.w6(32'hbc7c5a5d),
	.w7(32'hbb4702d3),
	.w8(32'hbb52d353),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c6062),
	.w1(32'hbb16edba),
	.w2(32'hba75c76b),
	.w3(32'h3b85590c),
	.w4(32'hbb8e5866),
	.w5(32'h3b4703c0),
	.w6(32'h3aa2c99b),
	.w7(32'hbb975124),
	.w8(32'hba7806ef),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e4dcd),
	.w1(32'h3b00dcaa),
	.w2(32'h3bc92ff0),
	.w3(32'h3bbf0f6c),
	.w4(32'hbb8dc791),
	.w5(32'hbc4cd8ef),
	.w6(32'h3af8ec95),
	.w7(32'h3b54dcab),
	.w8(32'h3b417168),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ebad2),
	.w1(32'h3abf266c),
	.w2(32'hbc17b0b2),
	.w3(32'h3b6b2fe4),
	.w4(32'h3a611b65),
	.w5(32'hbb83fb01),
	.w6(32'hba9f204d),
	.w7(32'hba4823ee),
	.w8(32'hbb486bd7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97f2d7),
	.w1(32'hba7d8c13),
	.w2(32'h3c20707b),
	.w3(32'h3b1b75ef),
	.w4(32'h3ac47564),
	.w5(32'hbb9aa230),
	.w6(32'h3b88b266),
	.w7(32'hbbe5ba0f),
	.w8(32'h3add7ee6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28a975),
	.w1(32'h3c3f4e3e),
	.w2(32'hbbff82b6),
	.w3(32'h3cccab55),
	.w4(32'h3c46cd69),
	.w5(32'h3cafd9d5),
	.w6(32'h3c83bc12),
	.w7(32'h3c35ecef),
	.w8(32'hbb31ca8e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9340d6),
	.w1(32'h3ae0c3c7),
	.w2(32'h3b214e35),
	.w3(32'hbc237524),
	.w4(32'h3ae49161),
	.w5(32'h3b10e24e),
	.w6(32'hbbd1ae27),
	.w7(32'hbad227eb),
	.w8(32'hba91bb80),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae32448),
	.w1(32'h3a211ef8),
	.w2(32'h3b3736b3),
	.w3(32'h3b8fc5ba),
	.w4(32'h3affdfee),
	.w5(32'hbb7a35ea),
	.w6(32'h3b824a1c),
	.w7(32'h3ade92fb),
	.w8(32'hbbbd40e8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a98f),
	.w1(32'hbb4a53b4),
	.w2(32'hbb6458ca),
	.w3(32'h3aa325ba),
	.w4(32'hbaaead88),
	.w5(32'hbc818578),
	.w6(32'h3a8cb5b4),
	.w7(32'h3baa44ce),
	.w8(32'hbaba6fd5),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b387b48),
	.w1(32'h3c0e1af5),
	.w2(32'h3c1e78f4),
	.w3(32'hbb64f18f),
	.w4(32'h3a0edfad),
	.w5(32'hbbcebf30),
	.w6(32'h3bdd3c9b),
	.w7(32'hbaa40078),
	.w8(32'hbb1d6e67),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c209815),
	.w1(32'hbb807cab),
	.w2(32'hbc1f81c3),
	.w3(32'h3bea2e93),
	.w4(32'hbbb51361),
	.w5(32'hbbfe1ddf),
	.w6(32'h3b91ead4),
	.w7(32'h3b2b5656),
	.w8(32'h3bbaefed),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93944c),
	.w1(32'h3bdbc90d),
	.w2(32'h3c65b38c),
	.w3(32'h3c9ab74b),
	.w4(32'h3bfe6959),
	.w5(32'h3c2486b8),
	.w6(32'h3b88a00f),
	.w7(32'hbb56f52c),
	.w8(32'h3c27dc97),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8c706),
	.w1(32'h3beca114),
	.w2(32'h3b834c72),
	.w3(32'h3c12a3f3),
	.w4(32'hba7c63be),
	.w5(32'hbbec2a4a),
	.w6(32'h3b8e330d),
	.w7(32'hbbab570b),
	.w8(32'hbc06208a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40a8c2),
	.w1(32'hbb19886b),
	.w2(32'hbb7550bb),
	.w3(32'hbb984154),
	.w4(32'h3a4e3f17),
	.w5(32'h3b58e789),
	.w6(32'hbb923b24),
	.w7(32'h3b8f24be),
	.w8(32'h39e1b3d7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c5618),
	.w1(32'hbc0c4a57),
	.w2(32'h3b83df46),
	.w3(32'hbbd55842),
	.w4(32'hbc75bb42),
	.w5(32'hbc18f971),
	.w6(32'hbb064626),
	.w7(32'hbb6595e0),
	.w8(32'hbc74d23e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8733c3),
	.w1(32'h389d5183),
	.w2(32'hba3fe4d3),
	.w3(32'h3cbe35dc),
	.w4(32'hbb6394af),
	.w5(32'hbb80f721),
	.w6(32'h3bc90193),
	.w7(32'hbc3d28eb),
	.w8(32'hbbba9314),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f5f0d),
	.w1(32'hbabf094f),
	.w2(32'h3b9859a4),
	.w3(32'hbb335c50),
	.w4(32'h3ba5f799),
	.w5(32'h3befecad),
	.w6(32'h3b0d5478),
	.w7(32'h3b7a784a),
	.w8(32'h3c02d6b5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83c0ca),
	.w1(32'h39585c1a),
	.w2(32'hbafab87a),
	.w3(32'hbbdba3fa),
	.w4(32'hbbc6603b),
	.w5(32'hbbf66af2),
	.w6(32'hbb630193),
	.w7(32'hbbe19415),
	.w8(32'hbc30152c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0eac),
	.w1(32'h3b986953),
	.w2(32'hbb65592b),
	.w3(32'hbc14b17e),
	.w4(32'h3a01ff09),
	.w5(32'h3a9a8617),
	.w6(32'hbb853dfb),
	.w7(32'h3ab71185),
	.w8(32'hbb220acb),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bebe3),
	.w1(32'hba822265),
	.w2(32'h3c09fa22),
	.w3(32'hbbda3acf),
	.w4(32'h3b6c075b),
	.w5(32'hbc332066),
	.w6(32'h3b43d1d5),
	.w7(32'hba0278ee),
	.w8(32'h3c5e1f79),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91530dd),
	.w1(32'hbaa334a3),
	.w2(32'h3b9da833),
	.w3(32'h3bd1c533),
	.w4(32'h3baa3751),
	.w5(32'hbc2d7121),
	.w6(32'h3b3ad4d4),
	.w7(32'h3bc1123a),
	.w8(32'h3bb23c1c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b13e58),
	.w1(32'hbaa0c0ac),
	.w2(32'hba9550b4),
	.w3(32'h3b596167),
	.w4(32'h3bbba4bb),
	.w5(32'hbc9186b9),
	.w6(32'h3ba2d7f8),
	.w7(32'h3b27370d),
	.w8(32'hba3e0d71),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e8dea),
	.w1(32'hb9273c78),
	.w2(32'hba9a392f),
	.w3(32'h3af1c963),
	.w4(32'hbb15a8b3),
	.w5(32'hbcad640f),
	.w6(32'h3bce46b5),
	.w7(32'hba04d0db),
	.w8(32'hbbef27e6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c539653),
	.w1(32'hbba90acb),
	.w2(32'h3a0ec78d),
	.w3(32'h3ca7492e),
	.w4(32'hbbba85cd),
	.w5(32'hbb68fddb),
	.w6(32'h3b4f06de),
	.w7(32'hbc26fa81),
	.w8(32'hbbab6af1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e1e26),
	.w1(32'h3be27d7f),
	.w2(32'h3c83dc11),
	.w3(32'h3c4a2757),
	.w4(32'hba0291fb),
	.w5(32'hbbfc8b5d),
	.w6(32'h3acf897d),
	.w7(32'h3a42bc7f),
	.w8(32'hbb5669b2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eae7a),
	.w1(32'h3b0399ce),
	.w2(32'h3b88020f),
	.w3(32'hb80742cd),
	.w4(32'h3ba2f5df),
	.w5(32'hbc2bcead),
	.w6(32'hbad62c82),
	.w7(32'h3b027226),
	.w8(32'hbb88f65a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89869e7),
	.w1(32'hbb3b0150),
	.w2(32'h3b4a9c87),
	.w3(32'hbbe39582),
	.w4(32'hbb8a64ad),
	.w5(32'hbc4ed165),
	.w6(32'h3a8ca17e),
	.w7(32'hb8f489c6),
	.w8(32'hbb9de791),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8186b6),
	.w1(32'hbb902516),
	.w2(32'hb96f1b1c),
	.w3(32'h3cc68f31),
	.w4(32'hbb939668),
	.w5(32'hbc5eee83),
	.w6(32'h3b3ed732),
	.w7(32'hbbd971ac),
	.w8(32'hbc5be743),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd27330),
	.w1(32'h3b105e08),
	.w2(32'h3bde1217),
	.w3(32'hba1cf0df),
	.w4(32'hbbeabba2),
	.w5(32'hbc13f785),
	.w6(32'h3b2ae387),
	.w7(32'hbbfe96a6),
	.w8(32'hbba92afc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47be07),
	.w1(32'hbb5dda81),
	.w2(32'h3b725d36),
	.w3(32'h3c0a6954),
	.w4(32'hb983f76b),
	.w5(32'hbc5f268f),
	.w6(32'hba239203),
	.w7(32'hbb6609bf),
	.w8(32'h3a8f8116),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be088b3),
	.w1(32'hba2f065c),
	.w2(32'hbb54d076),
	.w3(32'hbb653baf),
	.w4(32'hbaf58b91),
	.w5(32'hbb16f70e),
	.w6(32'h3baeec26),
	.w7(32'hbbaf13a8),
	.w8(32'hbb7ac469),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af08e52),
	.w1(32'hbb4e4e01),
	.w2(32'hbad63a66),
	.w3(32'hbbdc4381),
	.w4(32'h3be8010e),
	.w5(32'h3b9118b2),
	.w6(32'hba9b4753),
	.w7(32'h3bdc0688),
	.w8(32'h3adcaccc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2159f4),
	.w1(32'hbc021369),
	.w2(32'hbc1b522b),
	.w3(32'h3b3119f8),
	.w4(32'hbb15d7bf),
	.w5(32'h3b640216),
	.w6(32'hb9ce519c),
	.w7(32'hbab40ab0),
	.w8(32'h3a0f482c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02874a),
	.w1(32'hbbcb4bd0),
	.w2(32'hb955bb21),
	.w3(32'hbb2fb5a2),
	.w4(32'hbb9149ce),
	.w5(32'hbc09a231),
	.w6(32'h3b363753),
	.w7(32'hbc0d3c8b),
	.w8(32'hbb02a069),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba381a2),
	.w1(32'hbacd71be),
	.w2(32'hb9a37be8),
	.w3(32'h3c05e43f),
	.w4(32'h3b122f04),
	.w5(32'hbc61a1ea),
	.w6(32'h3aa07648),
	.w7(32'hbba234aa),
	.w8(32'hbb7c1dc4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8464f1),
	.w1(32'hbbf0143e),
	.w2(32'hbc24c00e),
	.w3(32'hba2f4f93),
	.w4(32'hbba746a1),
	.w5(32'h3c00ccc5),
	.w6(32'hbbef7c40),
	.w7(32'hbb9ebd4d),
	.w8(32'hbb93ae95),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82d897),
	.w1(32'h3a174653),
	.w2(32'h3c088677),
	.w3(32'h3c1c84df),
	.w4(32'h3b233227),
	.w5(32'hbc750990),
	.w6(32'hbbe6947d),
	.w7(32'h3ab4fc1d),
	.w8(32'hbab37839),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42191a),
	.w1(32'hbb040645),
	.w2(32'hbb47f182),
	.w3(32'h3bbc888d),
	.w4(32'hbb83bfef),
	.w5(32'hbc014f31),
	.w6(32'h3c107ba8),
	.w7(32'hbba15f8f),
	.w8(32'hbc118de5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1815e2),
	.w1(32'hbb51e650),
	.w2(32'hbbe36b4e),
	.w3(32'h3b12ac76),
	.w4(32'hbb78746e),
	.w5(32'hbbbf64f3),
	.w6(32'hbba23fbe),
	.w7(32'hbb4852eb),
	.w8(32'hbc3d2991),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a458574),
	.w1(32'h38f26f16),
	.w2(32'hbbf6b8b0),
	.w3(32'hbc495eb4),
	.w4(32'h3aa0ca9a),
	.w5(32'hb9b04b2b),
	.w6(32'hbb797d9a),
	.w7(32'hba9363ed),
	.w8(32'hbb13cff3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf03e7d),
	.w1(32'hbb5e95af),
	.w2(32'hbb387404),
	.w3(32'hbc04e933),
	.w4(32'hbc2935dc),
	.w5(32'hbbd3336c),
	.w6(32'hbafc572d),
	.w7(32'hbbf4b16a),
	.w8(32'hbb85dff2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f2f57),
	.w1(32'hbc0d71e1),
	.w2(32'hbbabcab5),
	.w3(32'hba38c190),
	.w4(32'hbb18be0d),
	.w5(32'hbb40fed5),
	.w6(32'hbab4f1ef),
	.w7(32'hbb7196ca),
	.w8(32'hbb77f3c2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d1813),
	.w1(32'hbb2a1be5),
	.w2(32'h3b2f1676),
	.w3(32'hbb4ac2a3),
	.w4(32'hba9795e0),
	.w5(32'h3b79ee19),
	.w6(32'hbaa48ca6),
	.w7(32'hbbdddd0f),
	.w8(32'hbb1e884f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79c0a),
	.w1(32'h3b3a79b5),
	.w2(32'h3beb8c22),
	.w3(32'h3942ec7c),
	.w4(32'hbb48b4e9),
	.w5(32'hbbf190bd),
	.w6(32'hbb55392e),
	.w7(32'hbb1195c9),
	.w8(32'hb9441a1d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6fc43),
	.w1(32'hbb368dc9),
	.w2(32'h397a0ba5),
	.w3(32'h3a0a5364),
	.w4(32'hbbcd09df),
	.w5(32'hbb8f111b),
	.w6(32'hb914c26e),
	.w7(32'hbbc8edf1),
	.w8(32'h3b733e91),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c257013),
	.w1(32'h3ace7262),
	.w2(32'hbba974ef),
	.w3(32'h3bf3cf91),
	.w4(32'h3af6f1c0),
	.w5(32'h3ad226f5),
	.w6(32'h3b9c6fb8),
	.w7(32'h3bdc44ac),
	.w8(32'hbb7aa929),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb201768),
	.w1(32'hbbe2be67),
	.w2(32'h3ac8edc0),
	.w3(32'hbb68ca04),
	.w4(32'hba8d288a),
	.w5(32'h3c8c5483),
	.w6(32'hbab0561a),
	.w7(32'hbaa095f7),
	.w8(32'hbb9311fc),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cab78),
	.w1(32'h3affdd8a),
	.w2(32'h3a8d3d16),
	.w3(32'hbbc19377),
	.w4(32'h3be10a5d),
	.w5(32'hbb97eab8),
	.w6(32'hbac19b13),
	.w7(32'h3b74478d),
	.w8(32'h3b85aceb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b84fe),
	.w1(32'hbbb4937c),
	.w2(32'hbb2950a0),
	.w3(32'h3bd31980),
	.w4(32'hbb2f2237),
	.w5(32'hbb036245),
	.w6(32'h3a57c7b0),
	.w7(32'hbb9fde53),
	.w8(32'hbb5226be),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38942a),
	.w1(32'hbb3c4332),
	.w2(32'h3bb0a1c2),
	.w3(32'h3b8c5d32),
	.w4(32'hbb0985c9),
	.w5(32'hbbe1b743),
	.w6(32'hbb48a105),
	.w7(32'h39924fe8),
	.w8(32'h3a85afe4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941b2e),
	.w1(32'hbbd4cec2),
	.w2(32'h3b018051),
	.w3(32'h3b3ac3ce),
	.w4(32'h3ad78554),
	.w5(32'hbc13eda8),
	.w6(32'hbba0f1ee),
	.w7(32'hbb7a6699),
	.w8(32'h3a343da1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d5661),
	.w1(32'hbc6d0c49),
	.w2(32'hbbcc2c56),
	.w3(32'h3afc9638),
	.w4(32'hbbd6c9bb),
	.w5(32'hbc3ec81d),
	.w6(32'hbae810ea),
	.w7(32'hbc48b7dc),
	.w8(32'h394e172a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e85fb),
	.w1(32'h3b00227e),
	.w2(32'hb7857f38),
	.w3(32'hbc3ef7ca),
	.w4(32'h39f16b5d),
	.w5(32'hbba34af0),
	.w6(32'hbc3a686d),
	.w7(32'h3a9917b1),
	.w8(32'h39748900),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule