module layer_8_featuremap_7(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4c7a2),
	.w1(32'hbc9304d4),
	.w2(32'h3c25a35a),
	.w3(32'h3c3a0ff3),
	.w4(32'hbc30743b),
	.w5(32'h3c7740c6),
	.w6(32'h3b7bfd45),
	.w7(32'hbb8b9df6),
	.w8(32'h3c83592f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99e559),
	.w1(32'h3b054282),
	.w2(32'h39e7964c),
	.w3(32'hbbb2ad9c),
	.w4(32'h3bb662a4),
	.w5(32'h3b518880),
	.w6(32'hbc1013b7),
	.w7(32'hbb840500),
	.w8(32'hbad87f20),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25a56e),
	.w1(32'h3ba73956),
	.w2(32'hbbc43baf),
	.w3(32'hbbbfe510),
	.w4(32'h3b85c7a5),
	.w5(32'hbbcb8b04),
	.w6(32'hbc01e55c),
	.w7(32'h3aa9e19e),
	.w8(32'hbc05a089),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14ae39),
	.w1(32'hbcf1524e),
	.w2(32'h3c98c920),
	.w3(32'h3cc5ae74),
	.w4(32'hbca29934),
	.w5(32'h3bf2292b),
	.w6(32'h3c7e19ee),
	.w7(32'h3cf08eb3),
	.w8(32'h3c640d65),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31f80e),
	.w1(32'hbb757a4f),
	.w2(32'h3c88fef1),
	.w3(32'h3ca2aedb),
	.w4(32'h3b4f50c6),
	.w5(32'h3cb40a5c),
	.w6(32'h3ce3cbad),
	.w7(32'hbbc970dd),
	.w8(32'h3c602cbc),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0e2c6),
	.w1(32'hbd1ee65f),
	.w2(32'hbc760da5),
	.w3(32'h3ca1334d),
	.w4(32'hbc72e996),
	.w5(32'hbcc95ebf),
	.w6(32'hbc9af89e),
	.w7(32'h3cba4e58),
	.w8(32'h3c1c322b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7142e),
	.w1(32'h3ae0f2cb),
	.w2(32'h3b1eb381),
	.w3(32'h3c110a84),
	.w4(32'hbb59f53f),
	.w5(32'hbb68fdc2),
	.w6(32'h3aefa556),
	.w7(32'hbb976c89),
	.w8(32'hbba4ee77),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6239f),
	.w1(32'h3ad64641),
	.w2(32'hbbe6cdfe),
	.w3(32'hbc1650cc),
	.w4(32'h3c1a9f38),
	.w5(32'h3bc4eafe),
	.w6(32'hbb8ce982),
	.w7(32'h387f46e2),
	.w8(32'hbc890d51),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25e466),
	.w1(32'h3ae3eb60),
	.w2(32'h3a72d449),
	.w3(32'h3cb68964),
	.w4(32'h3b251938),
	.w5(32'h3b4b844a),
	.w6(32'hbc9e6cd7),
	.w7(32'hbb79100d),
	.w8(32'hbb84d2e3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c571e),
	.w1(32'hbcb10f86),
	.w2(32'hbd121092),
	.w3(32'hbca4496e),
	.w4(32'h3ceef604),
	.w5(32'h3d189a90),
	.w6(32'hbaf38e56),
	.w7(32'hbbd76c7b),
	.w8(32'hbbc78837),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2012ad),
	.w1(32'hbc7b4981),
	.w2(32'hbb7b51f1),
	.w3(32'h3cd9f148),
	.w4(32'hbc185442),
	.w5(32'hbc3872ff),
	.w6(32'hbc39c1c3),
	.w7(32'h3c703f9c),
	.w8(32'hbb3534b2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf8ba2),
	.w1(32'h3b4a78a7),
	.w2(32'h3c3beab6),
	.w3(32'h3b7dba30),
	.w4(32'h3cb4de1c),
	.w5(32'h3c0a78ae),
	.w6(32'hbbce9a91),
	.w7(32'h3c01a34d),
	.w8(32'h3c26c59b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f1d8),
	.w1(32'h3cbb6c61),
	.w2(32'h3c992cb1),
	.w3(32'h3a10a68e),
	.w4(32'hbd163e2a),
	.w5(32'hbd114c04),
	.w6(32'hbc0192b4),
	.w7(32'h3c9f18b2),
	.w8(32'h3ca209d0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c8b6b),
	.w1(32'h3b3be69e),
	.w2(32'hbacdb73e),
	.w3(32'hbcc616e8),
	.w4(32'hba63d319),
	.w5(32'hbb7892a4),
	.w6(32'h3d2243a9),
	.w7(32'h3bb0bd5c),
	.w8(32'h3bd9aef2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43795),
	.w1(32'hba7c4552),
	.w2(32'h3b538ab4),
	.w3(32'hbbb53bbe),
	.w4(32'hbb9b9dc9),
	.w5(32'hbb9a7507),
	.w6(32'h3b82af63),
	.w7(32'hb8e2421c),
	.w8(32'h3a95454e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc90c70),
	.w1(32'h3a3bd892),
	.w2(32'h385e6e53),
	.w3(32'hbb61254d),
	.w4(32'hbc23cd21),
	.w5(32'hbb9ddfc4),
	.w6(32'h3ac07dcb),
	.w7(32'h3c0b3842),
	.w8(32'h3c360859),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec62c6),
	.w1(32'h3afb8972),
	.w2(32'h3bdd18c9),
	.w3(32'hbbbc91ce),
	.w4(32'hbccb89d3),
	.w5(32'hbc70ea1a),
	.w6(32'h3a07f785),
	.w7(32'h3b7c9b43),
	.w8(32'h3d16deb0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb571682),
	.w1(32'h3bea2ae3),
	.w2(32'hbb6fbb74),
	.w3(32'hbc8b17ab),
	.w4(32'h3bdcafc9),
	.w5(32'h3b3426d4),
	.w6(32'h3ca26e1f),
	.w7(32'hbbc9595d),
	.w8(32'h3c39ccfb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d140e30),
	.w1(32'hbd6daff1),
	.w2(32'hbc8a41f8),
	.w3(32'h3b5a4cf9),
	.w4(32'hbb140ff7),
	.w5(32'hbc270d2f),
	.w6(32'hbd68ebe7),
	.w7(32'h3d3c49f8),
	.w8(32'h3c3bd6b8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10b9ef),
	.w1(32'h3ca49985),
	.w2(32'h3c07af7f),
	.w3(32'h3c49c79c),
	.w4(32'h3c37ed37),
	.w5(32'h3c8053e6),
	.w6(32'h3bf1fb31),
	.w7(32'hbcfc3e5f),
	.w8(32'hbba79b82),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82978a),
	.w1(32'hbac9e377),
	.w2(32'hbb951c20),
	.w3(32'h3c23af57),
	.w4(32'hbbbc3183),
	.w5(32'hbb27d1f4),
	.w6(32'hbce9ea77),
	.w7(32'hbc7006a2),
	.w8(32'h3b8f0866),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18858c),
	.w1(32'hbb8b2b87),
	.w2(32'h3aba9d23),
	.w3(32'hba79a07c),
	.w4(32'h3bf8bc36),
	.w5(32'h3c7bd21c),
	.w6(32'hba07ae2b),
	.w7(32'hbc50f013),
	.w8(32'hbc9fbec4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b158be7),
	.w1(32'hbca8ae75),
	.w2(32'hbc90d49e),
	.w3(32'hbcec1f85),
	.w4(32'h3b22829d),
	.w5(32'h3aa27473),
	.w6(32'hbd5d0c5b),
	.w7(32'h3cf85626),
	.w8(32'h3d33a57b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e642c),
	.w1(32'h3c4e235f),
	.w2(32'h3c5b2bc9),
	.w3(32'h3b813c84),
	.w4(32'h3a3dc074),
	.w5(32'h3afabd4d),
	.w6(32'h3c74700a),
	.w7(32'hbc79ac15),
	.w8(32'hbc884aec),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2883d3),
	.w1(32'h3b8907d7),
	.w2(32'h3bf3a385),
	.w3(32'h3ab17652),
	.w4(32'h3b3bfdf1),
	.w5(32'h3b67848b),
	.w6(32'hbbe37c32),
	.w7(32'h3c0e052d),
	.w8(32'h3bf3777a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8b04),
	.w1(32'hbc325e39),
	.w2(32'hbbd8851a),
	.w3(32'hb868e38a),
	.w4(32'hbb321b9f),
	.w5(32'hbc25f60f),
	.w6(32'hbcba1b06),
	.w7(32'h3adfd98d),
	.w8(32'h3bf71807),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb975d55e),
	.w1(32'hbacf4e6f),
	.w2(32'h399d01e5),
	.w3(32'hbbad92ac),
	.w4(32'hbbed5ff4),
	.w5(32'hbb88bb11),
	.w6(32'hbbcbb665),
	.w7(32'hbbc55fad),
	.w8(32'hbb662568),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e429cfe),
	.w1(32'h3beee692),
	.w2(32'hbe194312),
	.w3(32'h3d87c33f),
	.w4(32'h3dd37e11),
	.w5(32'hbda13d14),
	.w6(32'hbe27f346),
	.w7(32'hbd15140e),
	.w8(32'h3e4c991c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb6312),
	.w1(32'hbc4cdd41),
	.w2(32'hbc53d15a),
	.w3(32'hbc2289e3),
	.w4(32'hbbf13866),
	.w5(32'hbc878398),
	.w6(32'h3cfc6556),
	.w7(32'h3b0c21fa),
	.w8(32'h3ba55118),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc062990),
	.w1(32'h3ac99010),
	.w2(32'h39cad07a),
	.w3(32'hbc1cb0da),
	.w4(32'hbb6ce06f),
	.w5(32'hbba73416),
	.w6(32'h3ba66921),
	.w7(32'h3baf9382),
	.w8(32'h3bb0c805),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5770ce),
	.w1(32'h3c08fa1b),
	.w2(32'h3c0c5a3f),
	.w3(32'hbbb5aba2),
	.w4(32'h3b11c6b0),
	.w5(32'h3bb7db4e),
	.w6(32'h3b152e5c),
	.w7(32'hbbdeb51b),
	.w8(32'hbc3dc27d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c058388),
	.w1(32'h3b053260),
	.w2(32'h3c323204),
	.w3(32'h3ab3d5bd),
	.w4(32'h3b5e94b4),
	.w5(32'h3b4beec8),
	.w6(32'hbbacd8e5),
	.w7(32'hbc2dd4e3),
	.w8(32'hb9abebfe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ed5fb),
	.w1(32'h3a1c3062),
	.w2(32'h3a95176b),
	.w3(32'h3a012a0c),
	.w4(32'hbae16ec0),
	.w5(32'hbb40a05f),
	.w6(32'hbc0f6792),
	.w7(32'hbb57a2ce),
	.w8(32'hbb23fbfb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49ce72),
	.w1(32'h3bfdf66b),
	.w2(32'h3c26b85c),
	.w3(32'hbb76a08a),
	.w4(32'hbb9086d4),
	.w5(32'hbbe3ebb8),
	.w6(32'hbb0db190),
	.w7(32'hbbcf3d28),
	.w8(32'hbc5f88a3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca539f8),
	.w1(32'h3c7a112e),
	.w2(32'h3c2f6e2e),
	.w3(32'hbb2cdc2b),
	.w4(32'h3c4599bd),
	.w5(32'h3c67e69a),
	.w6(32'hbc16985f),
	.w7(32'hbb3050f1),
	.w8(32'h3b9884b3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c801497),
	.w1(32'hba24ef30),
	.w2(32'hbc8b2143),
	.w3(32'hbbce6be0),
	.w4(32'h3bf44349),
	.w5(32'h3b66bb42),
	.w6(32'hbc8b3f65),
	.w7(32'h396f9a7f),
	.w8(32'h3ca6ebaa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba55811),
	.w1(32'h3bf72003),
	.w2(32'h3c9edaa2),
	.w3(32'hb9ee02ef),
	.w4(32'hbab9ad5f),
	.w5(32'hbb967750),
	.w6(32'h3b80e9bf),
	.w7(32'hbcbee0c9),
	.w8(32'hbcba70cf),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ae844),
	.w1(32'h3b7702da),
	.w2(32'h3b3a5e21),
	.w3(32'h3bc85708),
	.w4(32'h3cb1cb5c),
	.w5(32'h3c307e85),
	.w6(32'hbc599ea2),
	.w7(32'hbab11edd),
	.w8(32'hbbe64f96),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a943d4b),
	.w1(32'hbd0055d6),
	.w2(32'hbcd45b10),
	.w3(32'h3c0b1423),
	.w4(32'hbcad6f13),
	.w5(32'hbc95ee47),
	.w6(32'h3c0710d9),
	.w7(32'h3cc67a2b),
	.w8(32'h3d07c8b8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd03338),
	.w1(32'h3a4f3bd3),
	.w2(32'h39c8df80),
	.w3(32'hbc1d4222),
	.w4(32'h3b4d42db),
	.w5(32'hbbd35951),
	.w6(32'h3d047de9),
	.w7(32'hbc3c3fbb),
	.w8(32'hbbd41983),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca4bc5),
	.w1(32'hbc8299e3),
	.w2(32'h3a01deda),
	.w3(32'hbb0c6ed0),
	.w4(32'hbc43f289),
	.w5(32'hbc17d92b),
	.w6(32'hbbfd3ac7),
	.w7(32'h3cfe37fa),
	.w8(32'h3d166a00),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39859c6a),
	.w1(32'hbbadc296),
	.w2(32'h3b0ae853),
	.w3(32'hbb6593d3),
	.w4(32'hbbe7ca61),
	.w5(32'h3aa6ce8a),
	.w6(32'h3c14b139),
	.w7(32'h3b4f96f7),
	.w8(32'hbaef7f43),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b224ee9),
	.w1(32'hbb536166),
	.w2(32'hbba31cdb),
	.w3(32'h3aa8ae1d),
	.w4(32'h3b050591),
	.w5(32'hb9ac083f),
	.w6(32'h39e7fa40),
	.w7(32'h3b8bbba9),
	.w8(32'h3b9d068b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad693b),
	.w1(32'hbcd421fc),
	.w2(32'hbc8b4e28),
	.w3(32'h3bcd27d9),
	.w4(32'hbcb4ebfe),
	.w5(32'hbd07f49c),
	.w6(32'hbad3ec06),
	.w7(32'h3c169548),
	.w8(32'h3b86b6d5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcebf6d),
	.w1(32'hbcb6d2db),
	.w2(32'hbbf5038d),
	.w3(32'hbb5a6eb4),
	.w4(32'hbd1a59d5),
	.w5(32'hbd39f5f8),
	.w6(32'hbc95475c),
	.w7(32'h3d368180),
	.w8(32'h3d97873f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38038f),
	.w1(32'hbb28bc58),
	.w2(32'h3c17fef5),
	.w3(32'hbcc93542),
	.w4(32'h3c80d5ef),
	.w5(32'h3d0cd8d9),
	.w6(32'h3d3450d1),
	.w7(32'hbcb74b32),
	.w8(32'hbd07e8f5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d3f58),
	.w1(32'h3cbea728),
	.w2(32'h3c9d50b1),
	.w3(32'h3cb389aa),
	.w4(32'h3c0613ca),
	.w5(32'hbb54aefd),
	.w6(32'hbcd6b5f1),
	.w7(32'hbc76ceac),
	.w8(32'hbc4b05bd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07eebc),
	.w1(32'hbb7aac4f),
	.w2(32'h3ba9a14e),
	.w3(32'hbbdd31e5),
	.w4(32'hbb5da5e9),
	.w5(32'hbc6daa32),
	.w6(32'hbd6144c1),
	.w7(32'h3ad4c30c),
	.w8(32'h3c8a5062),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6bf1c),
	.w1(32'hbafa0164),
	.w2(32'hbad4f748),
	.w3(32'hbba1aeaf),
	.w4(32'h3962c3aa),
	.w5(32'hbb0d0553),
	.w6(32'hbbf4fb11),
	.w7(32'hbba2dbad),
	.w8(32'hbb7249b4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dc696),
	.w1(32'hbc2661de),
	.w2(32'h3cc774ff),
	.w3(32'h3cefd7d4),
	.w4(32'h3a1712cc),
	.w5(32'h37d568a8),
	.w6(32'h3c214ead),
	.w7(32'h3d0d271d),
	.w8(32'h3bce4fe0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3b55f),
	.w1(32'h3a68b83f),
	.w2(32'h3c8077a9),
	.w3(32'hbc8112e5),
	.w4(32'h3bfd7f34),
	.w5(32'h3caf140b),
	.w6(32'hbce7831e),
	.w7(32'hbc958d62),
	.w8(32'h3b866195),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dfa30),
	.w1(32'hbcf5432e),
	.w2(32'hbb95f2fa),
	.w3(32'h3c01ff4c),
	.w4(32'hbd1b09ad),
	.w5(32'hbca5a917),
	.w6(32'hbcaf4942),
	.w7(32'h3ce0d39d),
	.w8(32'hbc0dd5b1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e78973),
	.w1(32'hbb5f4229),
	.w2(32'hbc812a5b),
	.w3(32'h3b5c0fad),
	.w4(32'hbcbab22d),
	.w5(32'hbc69c0f7),
	.w6(32'h3b7df38b),
	.w7(32'h3cb97a37),
	.w8(32'h3d55dc0e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36f23e),
	.w1(32'h3be5e1b8),
	.w2(32'h3c0122d8),
	.w3(32'hbc54ed16),
	.w4(32'hbc012bfc),
	.w5(32'h3b5d1b82),
	.w6(32'h3d2cc8a5),
	.w7(32'hbc13973a),
	.w8(32'h3c55cf88),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3118a4),
	.w1(32'h3b2d4afe),
	.w2(32'h3c19fde6),
	.w3(32'hbc54172e),
	.w4(32'h3b4c2ae9),
	.w5(32'hb8ab5537),
	.w6(32'h3bc4e993),
	.w7(32'hbbc925b0),
	.w8(32'hbc2e630f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5e647b),
	.w1(32'h3c6468dd),
	.w2(32'hbb0d4743),
	.w3(32'hbcaf07b1),
	.w4(32'h3d08cdb0),
	.w5(32'h3b245996),
	.w6(32'hbd09e0b1),
	.w7(32'h3c471872),
	.w8(32'h3d7c7377),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ad620),
	.w1(32'h3a9c2dae),
	.w2(32'hba985584),
	.w3(32'hbaed2f4e),
	.w4(32'h3b09fa14),
	.w5(32'h3bd79570),
	.w6(32'h3ab6df9c),
	.w7(32'hbbe589f5),
	.w8(32'hbad5bc06),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7499),
	.w1(32'hbce2c0a3),
	.w2(32'hbc7eb35a),
	.w3(32'h3c4c397c),
	.w4(32'hbc279eb9),
	.w5(32'hbb1f83db),
	.w6(32'hbc2935af),
	.w7(32'h3bfbc122),
	.w8(32'hbc4cbaf1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56767),
	.w1(32'hbbd8e0cd),
	.w2(32'hbbb54a8a),
	.w3(32'h3b978207),
	.w4(32'hbbef1b34),
	.w5(32'hbbdb0944),
	.w6(32'hbc67e83c),
	.w7(32'h3afd41d2),
	.w8(32'h3c000717),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d9f27),
	.w1(32'hbcd49f84),
	.w2(32'hbd192943),
	.w3(32'hb8a25914),
	.w4(32'hbcf5a6f3),
	.w5(32'hbb2e35ec),
	.w6(32'h3c9ddab5),
	.w7(32'h3d1bad8f),
	.w8(32'h3ccf1f65),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd786fb),
	.w1(32'h3b823d98),
	.w2(32'h3b84d7e9),
	.w3(32'h3c203fe4),
	.w4(32'hbbfbf721),
	.w5(32'hbc2f1953),
	.w6(32'hba17df4e),
	.w7(32'hbb400c70),
	.w8(32'hbc0d1a06),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25c071),
	.w1(32'h3c7753b1),
	.w2(32'h3c89a813),
	.w3(32'hbc8e3b26),
	.w4(32'h3c16fe4f),
	.w5(32'h3b5d5765),
	.w6(32'hba303821),
	.w7(32'hbc275bab),
	.w8(32'hbc46e3a2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89a81f),
	.w1(32'hbc13ca3b),
	.w2(32'h3b08595e),
	.w3(32'hbc128ddc),
	.w4(32'h3bfcf502),
	.w5(32'h3b2e1921),
	.w6(32'hbc7e5734),
	.w7(32'hbbbc0a44),
	.w8(32'h3a0cef4a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d7be9),
	.w1(32'h3b059cdc),
	.w2(32'hbb9f6a5b),
	.w3(32'hbc14e5ca),
	.w4(32'hbca05771),
	.w5(32'hbc66d127),
	.w6(32'hbc45054e),
	.w7(32'h3c14b64d),
	.w8(32'h3c8cb109),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc195419),
	.w1(32'hbb0ffa10),
	.w2(32'hbb943d02),
	.w3(32'hbb30541c),
	.w4(32'hbacf835f),
	.w5(32'hbba89309),
	.w6(32'h3c89db84),
	.w7(32'h3b8f0f33),
	.w8(32'h3c01b203),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73bd31),
	.w1(32'hbb1eecb6),
	.w2(32'hbbaec46f),
	.w3(32'hbb4ab63d),
	.w4(32'hbbffa6c2),
	.w5(32'hbbfbc3db),
	.w6(32'hbbcd6cbe),
	.w7(32'h3b5cbdba),
	.w8(32'h3bc4c12a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affcae9),
	.w1(32'hba837613),
	.w2(32'h3a968619),
	.w3(32'h3b99b033),
	.w4(32'hbbbc4a6d),
	.w5(32'hbc07e955),
	.w6(32'hbb801d2b),
	.w7(32'h3a0265df),
	.w8(32'hba57789a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9977230),
	.w1(32'hbb99debc),
	.w2(32'hbb765e22),
	.w3(32'hbca5e3b6),
	.w4(32'h39433193),
	.w5(32'hbaf8ea53),
	.w6(32'hbc59c8c4),
	.w7(32'h3c0284e6),
	.w8(32'h3cec9de9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb738272),
	.w1(32'h39d8af0b),
	.w2(32'h39b11340),
	.w3(32'hbbd17275),
	.w4(32'hbc26776a),
	.w5(32'hbc5a8751),
	.w6(32'h3cb35c08),
	.w7(32'hbba4741b),
	.w8(32'hbbd19d8c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5651ed),
	.w1(32'hbc3185e8),
	.w2(32'hbcf8f7fa),
	.w3(32'h3c50d5e9),
	.w4(32'hbcb5c05b),
	.w5(32'hbd464a03),
	.w6(32'hbd35accc),
	.w7(32'h3aa8a401),
	.w8(32'h3d011b72),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7d3d5),
	.w1(32'h3a952aa9),
	.w2(32'h3b887d82),
	.w3(32'h393be1fc),
	.w4(32'h3b3bd42c),
	.w5(32'h3bc92ece),
	.w6(32'h3bdff618),
	.w7(32'h3b9d6351),
	.w8(32'h3c280f7b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad8f79),
	.w1(32'hba51f089),
	.w2(32'h3b254905),
	.w3(32'h3bd4518d),
	.w4(32'h398a139c),
	.w5(32'hbc0891a4),
	.w6(32'h3c135eb0),
	.w7(32'h3ba76d1a),
	.w8(32'h398e6db5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2df737),
	.w1(32'hbb26e220),
	.w2(32'hbac05922),
	.w3(32'hb7997daa),
	.w4(32'hbb6db838),
	.w5(32'hbb4f35de),
	.w6(32'h3a0e0ef1),
	.w7(32'hbba76dcd),
	.w8(32'hbba47061),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98e1cb),
	.w1(32'h3c6a1308),
	.w2(32'hbb40a216),
	.w3(32'hbb413f6e),
	.w4(32'h3d0e1d31),
	.w5(32'h3c903980),
	.w6(32'h3c2843fd),
	.w7(32'hba82bf80),
	.w8(32'h3d021705),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb028ac5),
	.w1(32'hbb140538),
	.w2(32'h3956881a),
	.w3(32'hbb2fd960),
	.w4(32'hbb041faf),
	.w5(32'hba5bc24c),
	.w6(32'h3ae6de8a),
	.w7(32'hbb9abfee),
	.w8(32'hbbb8ac73),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62ad9e),
	.w1(32'hbb23d305),
	.w2(32'h3a211e5c),
	.w3(32'h3b818de7),
	.w4(32'hbc242bf9),
	.w5(32'hbb6ced00),
	.w6(32'h3afbc0cf),
	.w7(32'hbbdce1b8),
	.w8(32'hbb81c615),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a874826),
	.w1(32'h3c0c288c),
	.w2(32'h3c2aa976),
	.w3(32'h3a898694),
	.w4(32'hba64fcbd),
	.w5(32'h3b89927a),
	.w6(32'h3af0a8a9),
	.w7(32'hbcc7d7e8),
	.w8(32'hbc6e819b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3af4e),
	.w1(32'hbcb2faea),
	.w2(32'hbc900653),
	.w3(32'h3c5d0440),
	.w4(32'hbcaa73e4),
	.w5(32'hbcec10d2),
	.w6(32'hbc970a54),
	.w7(32'hbc357d65),
	.w8(32'hbbb4c5af),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8f56b),
	.w1(32'h3c8cfc34),
	.w2(32'h3c47b034),
	.w3(32'hbca8ff6f),
	.w4(32'h3c96469a),
	.w5(32'h3cb2cbf2),
	.w6(32'hbcd7ebed),
	.w7(32'h3c807f8f),
	.w8(32'h3cf2c9a0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1815fb),
	.w1(32'hb945a832),
	.w2(32'hba4c7e00),
	.w3(32'h3b734a13),
	.w4(32'hbace4c0b),
	.w5(32'hbaf4d471),
	.w6(32'h3c418de1),
	.w7(32'h3b184e35),
	.w8(32'h3b74d542),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b8218),
	.w1(32'h3a58c697),
	.w2(32'h3c0a026b),
	.w3(32'hbaa42332),
	.w4(32'h3b82fd6f),
	.w5(32'h3c13dc26),
	.w6(32'h3b9c5cd7),
	.w7(32'hba87f44f),
	.w8(32'h3ba687c4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f1b8),
	.w1(32'hbb28ae51),
	.w2(32'h3c1a28aa),
	.w3(32'h3cc64c41),
	.w4(32'hbba719f2),
	.w5(32'hbc9e5b2a),
	.w6(32'hbb83e23d),
	.w7(32'h3c0eedd5),
	.w8(32'hbc144134),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab52afa),
	.w1(32'hbc80d421),
	.w2(32'h3baefb43),
	.w3(32'hbaca5613),
	.w4(32'hbbe6679a),
	.w5(32'hbc0fc4cd),
	.w6(32'hbca2a712),
	.w7(32'hbc20b3e7),
	.w8(32'hbb85afeb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9600ce),
	.w1(32'h3c61e03d),
	.w2(32'h3d6a8ca7),
	.w3(32'h3cbc5624),
	.w4(32'hbc206e47),
	.w5(32'h3d496954),
	.w6(32'h3d783bc1),
	.w7(32'h3c9513fc),
	.w8(32'hbbcc1513),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d65a3),
	.w1(32'hbcacd498),
	.w2(32'hbbade453),
	.w3(32'h3c928357),
	.w4(32'hbc6f537f),
	.w5(32'hbc9b364d),
	.w6(32'hbc48c697),
	.w7(32'h3c17e919),
	.w8(32'h3b075695),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba620b0),
	.w1(32'hb9c9c998),
	.w2(32'h3c4416ef),
	.w3(32'h3cf75074),
	.w4(32'hbb298ad3),
	.w5(32'hbc8588d6),
	.w6(32'h3c8e466e),
	.w7(32'h3d0dd66e),
	.w8(32'h3a62e252),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ba04),
	.w1(32'hbc1009bf),
	.w2(32'h3c16c5c6),
	.w3(32'hbb3cb98a),
	.w4(32'hba6bb088),
	.w5(32'h3bb409e3),
	.w6(32'h3b3e2072),
	.w7(32'hbab2e4c8),
	.w8(32'h3bfbd645),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbb757),
	.w1(32'h3b31d874),
	.w2(32'h3bc9ad25),
	.w3(32'h3baeee44),
	.w4(32'h3b540234),
	.w5(32'h3be0d946),
	.w6(32'hbb2ced05),
	.w7(32'h3bc3c30e),
	.w8(32'h3c2dd0bf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45066c),
	.w1(32'h3adeac6c),
	.w2(32'h3b9ccb03),
	.w3(32'h3b5105a4),
	.w4(32'hba64b673),
	.w5(32'hb8f84815),
	.w6(32'h3bf8fd62),
	.w7(32'hbb4bbaaa),
	.w8(32'h3b96d432),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d4a99),
	.w1(32'hbb5fa4d1),
	.w2(32'hbbda66c5),
	.w3(32'hba9d0549),
	.w4(32'h3a79f36f),
	.w5(32'h3ab7f243),
	.w6(32'h3a576f7b),
	.w7(32'h3c8e6787),
	.w8(32'h3ca2eb32),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6866d),
	.w1(32'h3a78bf9b),
	.w2(32'h3c2d4ee2),
	.w3(32'hbbbdd791),
	.w4(32'hbbc01ab3),
	.w5(32'hbbb1fbbc),
	.w6(32'h3c2f29bf),
	.w7(32'hbc79b1f2),
	.w8(32'hbb5fdbd8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819ed6),
	.w1(32'h3bd989dd),
	.w2(32'h3aa49985),
	.w3(32'hbbe9d925),
	.w4(32'hbb8464cb),
	.w5(32'hbb88a0ca),
	.w6(32'hbba2e959),
	.w7(32'h3bd2fee8),
	.w8(32'h3b9e7bed),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec08c2),
	.w1(32'h3b7e66b4),
	.w2(32'hbb002b5e),
	.w3(32'h3c5dc825),
	.w4(32'hbc5a11c4),
	.w5(32'hbbba0bee),
	.w6(32'h3c210299),
	.w7(32'hbba91eec),
	.w8(32'hbc7958c9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35ae21),
	.w1(32'hbc00935f),
	.w2(32'hbb69f2e6),
	.w3(32'hbc579447),
	.w4(32'hbb83ed0d),
	.w5(32'hbabcd48e),
	.w6(32'hbc4afd99),
	.w7(32'h3a27e1a8),
	.w8(32'h3b74376a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ecccf),
	.w1(32'h3c07fa71),
	.w2(32'h3ab9dcc8),
	.w3(32'hbbf08c85),
	.w4(32'h3c32f85e),
	.w5(32'h3b8cbbb5),
	.w6(32'hbadce3db),
	.w7(32'h3b2fe486),
	.w8(32'h3b5f4f50),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392207f4),
	.w1(32'h3bcdb96e),
	.w2(32'h3c1dda81),
	.w3(32'hbc82a293),
	.w4(32'hbb281166),
	.w5(32'h3c7d3f6f),
	.w6(32'hbc53d932),
	.w7(32'hb932f51e),
	.w8(32'h3c3104e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66e898),
	.w1(32'hbc1d86bc),
	.w2(32'hba2934f4),
	.w3(32'h3b16c92f),
	.w4(32'hbb8f8fed),
	.w5(32'hbb3c7fff),
	.w6(32'h3beb5adb),
	.w7(32'hbb8fed50),
	.w8(32'hbc00b756),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab96b59),
	.w1(32'h39341d2e),
	.w2(32'hbb9c859b),
	.w3(32'hbb0f065c),
	.w4(32'hb98bc5ac),
	.w5(32'hbab472b4),
	.w6(32'hbafc47ee),
	.w7(32'h3b913f0d),
	.w8(32'h3b3d54cb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1b1ad),
	.w1(32'h395c549c),
	.w2(32'hb983268e),
	.w3(32'hbbde1625),
	.w4(32'hb881f47e),
	.w5(32'hb9a9849e),
	.w6(32'h3aaa3162),
	.w7(32'h39112957),
	.w8(32'hb9fa4fa5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39468cb5),
	.w1(32'hbac71e8a),
	.w2(32'hbb57e209),
	.w3(32'hb9486903),
	.w4(32'h3a759eb2),
	.w5(32'hbaf2d3a1),
	.w6(32'hb9f0f4d9),
	.w7(32'h3b0dc9b2),
	.w8(32'h39d9f935),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a030),
	.w1(32'hbc022d2e),
	.w2(32'hbb688826),
	.w3(32'hbb01bde9),
	.w4(32'hbc0b3d83),
	.w5(32'hbc045c44),
	.w6(32'hba7c6098),
	.w7(32'hbc05737c),
	.w8(32'hbae75a81),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e2458),
	.w1(32'h3a6a0d94),
	.w2(32'h3a35b22b),
	.w3(32'hbc775a6f),
	.w4(32'h3b819390),
	.w5(32'hbad5882b),
	.w6(32'hbc00ea43),
	.w7(32'h3c40c029),
	.w8(32'h3c03aaee),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7d105),
	.w1(32'hba8a73cf),
	.w2(32'hbae35274),
	.w3(32'hbb343d4c),
	.w4(32'hbad63c2f),
	.w5(32'hb8b67e74),
	.w6(32'h3be931c4),
	.w7(32'hbbd0bc67),
	.w8(32'hbbbd41d9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba2902),
	.w1(32'h3c7f8f65),
	.w2(32'h3bb9426f),
	.w3(32'h3c3a8df4),
	.w4(32'hbbeda0a6),
	.w5(32'hbc0275a6),
	.w6(32'hbb7cb4c5),
	.w7(32'hbc2c783a),
	.w8(32'hbc89b1c9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa918a8),
	.w1(32'h3c129aac),
	.w2(32'h3bb2445e),
	.w3(32'h3a168161),
	.w4(32'hbb2797d4),
	.w5(32'hbbb8b02c),
	.w6(32'h3b88ed74),
	.w7(32'h3bd8c279),
	.w8(32'h3b674ced),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b217a),
	.w1(32'hbc3c670a),
	.w2(32'hbc51fe62),
	.w3(32'h3c07ef7a),
	.w4(32'hbc286da3),
	.w5(32'hbce7875f),
	.w6(32'hbc157847),
	.w7(32'hbbbb19cf),
	.w8(32'h39b10563),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02e971),
	.w1(32'hbaca88c1),
	.w2(32'hbae5b525),
	.w3(32'hbba94892),
	.w4(32'h3b1ced88),
	.w5(32'h3ad24d4d),
	.w6(32'hbc11923a),
	.w7(32'h3abf5b1d),
	.w8(32'h3a09ace2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c0cf8),
	.w1(32'h3bbc62e3),
	.w2(32'h3c52e333),
	.w3(32'h3b531757),
	.w4(32'h3ab01f3e),
	.w5(32'h3c1b29d8),
	.w6(32'h3b13e8bf),
	.w7(32'h3ab1df5f),
	.w8(32'h3b32ff23),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37f318),
	.w1(32'hbb95e2f4),
	.w2(32'hbc14a5bf),
	.w3(32'h3bae4bdc),
	.w4(32'hbbf8df71),
	.w5(32'hbc6ce628),
	.w6(32'hb9a4abed),
	.w7(32'hbca2a87d),
	.w8(32'hbc9fc7e5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0cc72),
	.w1(32'h3baa68f2),
	.w2(32'h3bfdb3c3),
	.w3(32'hbcca67aa),
	.w4(32'h3aefa2a7),
	.w5(32'h3aff111b),
	.w6(32'hbcd0480c),
	.w7(32'h3bd3719f),
	.w8(32'h3c1028fa),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b671b78),
	.w1(32'hbb521c55),
	.w2(32'hb9dbd4f0),
	.w3(32'hbc3601ea),
	.w4(32'h3b6e8f57),
	.w5(32'h3c0cb0ea),
	.w6(32'hbbb61e4d),
	.w7(32'hbc086022),
	.w8(32'h3ac045a7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ac94b),
	.w1(32'h3aa0f0d7),
	.w2(32'h3c5725ac),
	.w3(32'h3b170f41),
	.w4(32'h3b98ac28),
	.w5(32'h3bd44435),
	.w6(32'hbb6bb156),
	.w7(32'h3c3943a8),
	.w8(32'h3c2a401a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88c30e),
	.w1(32'h3c42cec9),
	.w2(32'h3c06a2d8),
	.w3(32'h3c3df5e0),
	.w4(32'h3c6121b2),
	.w5(32'h3c14af0b),
	.w6(32'h3b62c3e0),
	.w7(32'h3c8b0e49),
	.w8(32'h3c38a74c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35241f),
	.w1(32'h3bfaced6),
	.w2(32'h3b21cc2c),
	.w3(32'h3bf96303),
	.w4(32'hb9f4fc6f),
	.w5(32'h3aefd78f),
	.w6(32'h3c215863),
	.w7(32'hb9a547c4),
	.w8(32'h3bf44e8e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5368d4),
	.w1(32'h3b0b9d4e),
	.w2(32'h3c2709a0),
	.w3(32'h3b8a26dc),
	.w4(32'h3adb0b72),
	.w5(32'h3bf767b3),
	.w6(32'h3c24b375),
	.w7(32'h3c33b24f),
	.w8(32'h3c2d3554),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7028d5),
	.w1(32'hb9a95233),
	.w2(32'hba36d333),
	.w3(32'hbaacadad),
	.w4(32'h39cc04a3),
	.w5(32'h3a84cc28),
	.w6(32'h3a8975ff),
	.w7(32'h3a6adbe9),
	.w8(32'h39c94afb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a182b79),
	.w1(32'h3bca2602),
	.w2(32'h3c3b895a),
	.w3(32'h39156105),
	.w4(32'h3b923b08),
	.w5(32'h3c0a92b0),
	.w6(32'hbb5ed779),
	.w7(32'hbc169fec),
	.w8(32'hbbcb83be),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69628a),
	.w1(32'hbb61e355),
	.w2(32'hbb951fe6),
	.w3(32'h3c112380),
	.w4(32'h3b14f1dd),
	.w5(32'hbae26036),
	.w6(32'hbbb1fd10),
	.w7(32'h3bf4add5),
	.w8(32'h3ca3f6e2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be82c28),
	.w1(32'hbbf0d280),
	.w2(32'h3b1d64f6),
	.w3(32'h3a12117f),
	.w4(32'hbbfa69ee),
	.w5(32'hbac9a805),
	.w6(32'hba683ebb),
	.w7(32'hb9cf53ac),
	.w8(32'hbb321c47),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf026c3),
	.w1(32'hba3b8931),
	.w2(32'h3a4a9bad),
	.w3(32'h394a7e11),
	.w4(32'hba6c73b8),
	.w5(32'hba872ce0),
	.w6(32'hbb54cf0b),
	.w7(32'hbac8126d),
	.w8(32'hbaa8ac2b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3302f),
	.w1(32'h3c75d8f0),
	.w2(32'h3bf4070a),
	.w3(32'hbbbad5db),
	.w4(32'h3c26fea7),
	.w5(32'h3cb11a2f),
	.w6(32'h3c0cd4c9),
	.w7(32'h39b83736),
	.w8(32'h3c101bd4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf19b7d),
	.w1(32'h3b1a9aeb),
	.w2(32'hbaa2ec17),
	.w3(32'hb9df2b25),
	.w4(32'h3bb3fd68),
	.w5(32'h3916592a),
	.w6(32'h3bda2318),
	.w7(32'h3a8ff8eb),
	.w8(32'hbb349ebe),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aac52),
	.w1(32'hbb0d0f16),
	.w2(32'hbb024a13),
	.w3(32'h3a9035e2),
	.w4(32'hbaeb9151),
	.w5(32'hbab7d2da),
	.w6(32'h36eeb028),
	.w7(32'hbaa792c1),
	.w8(32'hba7f9b73),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb167b39),
	.w1(32'hba46757d),
	.w2(32'h38d59eee),
	.w3(32'hbb1366c6),
	.w4(32'hbbce9906),
	.w5(32'hbb784b54),
	.w6(32'hbaf619c3),
	.w7(32'hbc02f7c2),
	.w8(32'hbc055e04),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e2901),
	.w1(32'h392e8dad),
	.w2(32'hbab607b7),
	.w3(32'hbb2da0c4),
	.w4(32'hba67848d),
	.w5(32'hbbe9de6b),
	.w6(32'hbbe9a0ff),
	.w7(32'h3c20570b),
	.w8(32'h3b5e1833),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce9d995),
	.w1(32'hb9f837b5),
	.w2(32'h3c171852),
	.w3(32'h3c431b48),
	.w4(32'hba220194),
	.w5(32'h3c17f0fc),
	.w6(32'h3cb1e686),
	.w7(32'hbb8cf898),
	.w8(32'h3c2e71c5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28101b),
	.w1(32'h3bb45d48),
	.w2(32'h3ad69ed9),
	.w3(32'hbb225319),
	.w4(32'h3c3c33e2),
	.w5(32'h3bd38dc2),
	.w6(32'hbc11357c),
	.w7(32'h3aa05871),
	.w8(32'h3c18e912),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9404c56),
	.w1(32'hbbcc112b),
	.w2(32'hbad5382a),
	.w3(32'hbbb733c5),
	.w4(32'hbc71a716),
	.w5(32'hbbcdcd3f),
	.w6(32'hbc7704d6),
	.w7(32'hbbd21cb4),
	.w8(32'h3b463dd5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule