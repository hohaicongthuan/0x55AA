module layer_6_featuremap_6(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebe592),
	.w1(32'h3bfd627d),
	.w2(32'h3d3ec8a4),
	.w3(32'hb7e2d794),
	.w4(32'hbc72f4e8),
	.w5(32'hbcaacacd),
	.w6(32'hbbf8fc87),
	.w7(32'h3ca7e376),
	.w8(32'hbcc7dcc0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514290),
	.w1(32'h39180cad),
	.w2(32'hbbee1b7f),
	.w3(32'hbd107307),
	.w4(32'hbc05cdda),
	.w5(32'hbbd3c56f),
	.w6(32'h3affde2f),
	.w7(32'h3b1af901),
	.w8(32'hbb718cdb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801815),
	.w1(32'h3b8ecb7c),
	.w2(32'hbae59a4d),
	.w3(32'hbb12a33e),
	.w4(32'h3b13b668),
	.w5(32'hbba5aec4),
	.w6(32'hbaeae6c5),
	.w7(32'hbb2f9f56),
	.w8(32'hbc022257),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84818e),
	.w1(32'h3c4b7543),
	.w2(32'h3cf97a4b),
	.w3(32'hb506e735),
	.w4(32'h3b955949),
	.w5(32'h3cd1315e),
	.w6(32'hbc7261bb),
	.w7(32'h3bdb7b2e),
	.w8(32'hbc96091f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1de2a3),
	.w1(32'hbbe0f0da),
	.w2(32'hbc0f440c),
	.w3(32'hbc0b3e93),
	.w4(32'hbb11e51e),
	.w5(32'hbb906f04),
	.w6(32'hbb6bc6b6),
	.w7(32'hbb861212),
	.w8(32'hb99dde80),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadebcff),
	.w1(32'hbc11d808),
	.w2(32'hbbfc6a27),
	.w3(32'h3a945ea4),
	.w4(32'hbc31099a),
	.w5(32'hbc517fa7),
	.w6(32'h3ba341b1),
	.w7(32'h3c902666),
	.w8(32'hbb70aa2d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cba8f),
	.w1(32'h3caac47b),
	.w2(32'h3d079d6d),
	.w3(32'hbcc240c6),
	.w4(32'h3c4ab35e),
	.w5(32'h3ccd8131),
	.w6(32'h3c7f5013),
	.w7(32'h3ccf01ab),
	.w8(32'h3c33ebad),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78b4bf),
	.w1(32'hbc83d73c),
	.w2(32'hbb8c902e),
	.w3(32'h3c075be2),
	.w4(32'hbb85099c),
	.w5(32'h3bf1363a),
	.w6(32'hbbb03879),
	.w7(32'h3bb558f7),
	.w8(32'h3ac7d36f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4890b2),
	.w1(32'hbbefa28a),
	.w2(32'hbc2f1e3d),
	.w3(32'h3bb03024),
	.w4(32'hbaca6449),
	.w5(32'h3a799bfd),
	.w6(32'hbbc7d5ff),
	.w7(32'h39cb58eb),
	.w8(32'h3a08a7c2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba858de4),
	.w1(32'h3c9b3dd1),
	.w2(32'h3cc52c35),
	.w3(32'hba0eeea3),
	.w4(32'h3c62d06f),
	.w5(32'h3ca23ff0),
	.w6(32'h3c79d526),
	.w7(32'h3c9a6db4),
	.w8(32'h3c5602b3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77acc2),
	.w1(32'hb88e7d14),
	.w2(32'hbba0aaa4),
	.w3(32'h3c2e662d),
	.w4(32'h3a0124f2),
	.w5(32'h3b1697ac),
	.w6(32'hbb4e5052),
	.w7(32'hbc06368c),
	.w8(32'h3ac6dce3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2994c9),
	.w1(32'h39a60aba),
	.w2(32'h3c4647ff),
	.w3(32'h3b1195d5),
	.w4(32'hbbc6b9ec),
	.w5(32'h3bec61d0),
	.w6(32'hbba39434),
	.w7(32'hbad550be),
	.w8(32'hbba7000e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9513cd),
	.w1(32'h3c0e2db8),
	.w2(32'h3ca467c9),
	.w3(32'hbc01b6bf),
	.w4(32'hbb8e48ca),
	.w5(32'hbc3d68ca),
	.w6(32'h3a19ce98),
	.w7(32'h3c41c454),
	.w8(32'hbc4db667),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb053),
	.w1(32'h3ce9da3c),
	.w2(32'h3d58eec3),
	.w3(32'hbc605871),
	.w4(32'hbbe7d98e),
	.w5(32'hbc137225),
	.w6(32'hbbd2363c),
	.w7(32'h3c13dbec),
	.w8(32'hbc378c47),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88a5ea),
	.w1(32'hbabf1485),
	.w2(32'h3c80b6ec),
	.w3(32'hbcc38720),
	.w4(32'hbaaf4adc),
	.w5(32'hba9c3796),
	.w6(32'h3cb05c95),
	.w7(32'h3bedaea1),
	.w8(32'hbc072b73),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8292c8),
	.w1(32'h3b133964),
	.w2(32'h3c1f95df),
	.w3(32'h3ba65a57),
	.w4(32'h39211090),
	.w5(32'hbc2f4e3b),
	.w6(32'hb9fac4a6),
	.w7(32'hbb2d765e),
	.w8(32'hbc33dc9c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b192a03),
	.w1(32'hbb14ff63),
	.w2(32'h3b8cd3c6),
	.w3(32'hbc460954),
	.w4(32'hbbbf63bb),
	.w5(32'hb84e8f3d),
	.w6(32'hbbe1abf8),
	.w7(32'hbc5ae547),
	.w8(32'hbc29e0d4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7bede),
	.w1(32'hbc61a051),
	.w2(32'hbd0629dc),
	.w3(32'hbb469ad7),
	.w4(32'h39f151fc),
	.w5(32'hbce22ff5),
	.w6(32'hb9afe9de),
	.w7(32'hbc4ee116),
	.w8(32'h3bc6c5ee),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00be9a),
	.w1(32'hbba08d22),
	.w2(32'hbbc5583c),
	.w3(32'h3c9b1780),
	.w4(32'hb962c078),
	.w5(32'hb9a82a6c),
	.w6(32'hbb5f5dce),
	.w7(32'hbb07b873),
	.w8(32'hbab26901),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf8c95),
	.w1(32'h3ba5cab1),
	.w2(32'h3a927846),
	.w3(32'h39e58f89),
	.w4(32'hbc6ba648),
	.w5(32'hbd10439c),
	.w6(32'h3b89ba49),
	.w7(32'hbba63375),
	.w8(32'hbc893763),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb61ba7),
	.w1(32'hbc07f3e0),
	.w2(32'hbc3767e8),
	.w3(32'hbd324a84),
	.w4(32'hbb55f9f5),
	.w5(32'hbc11a819),
	.w6(32'h3a643a78),
	.w7(32'hbba14e3e),
	.w8(32'h3b164e0d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b298000),
	.w1(32'hbbf976ac),
	.w2(32'hbb8fd7a1),
	.w3(32'h3c2f1f87),
	.w4(32'hba117dc6),
	.w5(32'h3a66ede9),
	.w6(32'hbba7a240),
	.w7(32'hbb76be89),
	.w8(32'hbb66b88b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba257447),
	.w1(32'h3aa9cf6e),
	.w2(32'h3b0f8e0b),
	.w3(32'h3abec6cb),
	.w4(32'h3adc0875),
	.w5(32'hb944e6b4),
	.w6(32'h3c23b439),
	.w7(32'h3acc6b5a),
	.w8(32'h3bf2283f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6c8f5),
	.w1(32'hbbe0a884),
	.w2(32'hbbe18b37),
	.w3(32'h39f362b3),
	.w4(32'hbc2c301c),
	.w5(32'hbc901707),
	.w6(32'hbad0da29),
	.w7(32'hbbc707da),
	.w8(32'hbc8d8d1c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc582dbd),
	.w1(32'hbaffb3ab),
	.w2(32'h3c1d81f0),
	.w3(32'hbca38b0e),
	.w4(32'hbc03c043),
	.w5(32'hbc4bb27e),
	.w6(32'h3b674144),
	.w7(32'h3c6df580),
	.w8(32'hbca6b31e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca51010),
	.w1(32'h39977ec8),
	.w2(32'hbc5435f8),
	.w3(32'hbced2e53),
	.w4(32'hbb868941),
	.w5(32'hbc7d05ef),
	.w6(32'h3ba6d729),
	.w7(32'hb99a759c),
	.w8(32'h3c1d8eca),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20347f),
	.w1(32'h3bbe7f1b),
	.w2(32'h3c658aea),
	.w3(32'hba8f8ff3),
	.w4(32'h3ae8cc0f),
	.w5(32'h3c669b7f),
	.w6(32'hbba33896),
	.w7(32'h3a717b26),
	.w8(32'hbb513421),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f9a2),
	.w1(32'h39725656),
	.w2(32'h3c72f00f),
	.w3(32'h3c1b4dd3),
	.w4(32'hbb51b748),
	.w5(32'hbbf85000),
	.w6(32'h3bef6064),
	.w7(32'h3c9bb4af),
	.w8(32'hbb425967),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7944de),
	.w1(32'hbb8dcfd4),
	.w2(32'hba16b574),
	.w3(32'hbc8255c8),
	.w4(32'hbbbed14a),
	.w5(32'hbba50973),
	.w6(32'hbb82bbba),
	.w7(32'hb93abf97),
	.w8(32'hbc68e456),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d0406),
	.w1(32'h3c264ae2),
	.w2(32'h3c70bdf4),
	.w3(32'hbbfa4f97),
	.w4(32'h3b898881),
	.w5(32'h3ca5e1b8),
	.w6(32'hbbfe7c22),
	.w7(32'h3c3be018),
	.w8(32'hbb7f9676),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f1cdf),
	.w1(32'hb672c4be),
	.w2(32'hb664f25c),
	.w3(32'hbb0f0be9),
	.w4(32'hb6010b02),
	.w5(32'h36a8a753),
	.w6(32'h365979e3),
	.w7(32'h376a1fbb),
	.w8(32'h35f714f6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71d3ac8),
	.w1(32'h359c39a0),
	.w2(32'hb6d080cf),
	.w3(32'hb7256b04),
	.w4(32'hb5a401e8),
	.w5(32'h3647dbd7),
	.w6(32'h36c945b2),
	.w7(32'h36b4387f),
	.w8(32'hb6a312f1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809c902),
	.w1(32'h37bcaffc),
	.w2(32'h3718ec7b),
	.w3(32'h383680a2),
	.w4(32'h3809ad30),
	.w5(32'h378d960d),
	.w6(32'h386d5689),
	.w7(32'h381bcec7),
	.w8(32'h37cecaa7),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a55247),
	.w1(32'h37fc0dcd),
	.w2(32'h37fc015f),
	.w3(32'h377d4da6),
	.w4(32'h379d6ea7),
	.w5(32'h370e58ba),
	.w6(32'h35961f80),
	.w7(32'h371cc702),
	.w8(32'h372e83cb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3705c1bf),
	.w1(32'h3759dc0d),
	.w2(32'h36c82fd0),
	.w3(32'h36cd6814),
	.w4(32'h36afe86f),
	.w5(32'h36f030e3),
	.w6(32'h359fbfef),
	.w7(32'h369901cc),
	.w8(32'h36a382cc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c288e),
	.w1(32'h36410d89),
	.w2(32'hb851b696),
	.w3(32'hb856b8dd),
	.w4(32'h37d69c37),
	.w5(32'hb657c19b),
	.w6(32'h38c0af4c),
	.w7(32'h389c9a8e),
	.w8(32'h37c1227f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ec71e),
	.w1(32'hb800ee37),
	.w2(32'hb7ebe3d0),
	.w3(32'hb7a6a14c),
	.w4(32'hb7838418),
	.w5(32'hb7db30dd),
	.w6(32'hb4e2443e),
	.w7(32'h37a3d66e),
	.w8(32'hb78590de),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bfa7c4),
	.w1(32'h388cc990),
	.w2(32'h3846c1b7),
	.w3(32'h38b83f1f),
	.w4(32'h38c05890),
	.w5(32'h38e214f5),
	.w6(32'h392f1a68),
	.w7(32'h391b4f24),
	.w8(32'h3905193b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e6427f),
	.w1(32'hb7ec8648),
	.w2(32'hb789e2ea),
	.w3(32'hb7beda4b),
	.w4(32'hb7c4fcf7),
	.w5(32'hb7810eab),
	.w6(32'hb7a47d13),
	.w7(32'hb7843252),
	.w8(32'hb6ca155c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36511b18),
	.w1(32'h38a32b37),
	.w2(32'h37f8ec5c),
	.w3(32'h395387c9),
	.w4(32'h399b4f33),
	.w5(32'h390b90fb),
	.w6(32'h39a13642),
	.w7(32'h391892a2),
	.w8(32'h38648c5f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8286abc),
	.w1(32'hb74842d1),
	.w2(32'h375c3c1c),
	.w3(32'hb7eecbd9),
	.w4(32'hb584fd46),
	.w5(32'h35045962),
	.w6(32'hb7a02994),
	.w7(32'hb7f7804c),
	.w8(32'hb82b51c4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b936f6),
	.w1(32'hb7f98534),
	.w2(32'hb7eb2566),
	.w3(32'hb7a8deda),
	.w4(32'hb76d5a7e),
	.w5(32'hb7e3790a),
	.w6(32'h381a32df),
	.w7(32'h382893fa),
	.w8(32'h35f3a9be),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63adc21),
	.w1(32'hb626bbd6),
	.w2(32'hb6076b12),
	.w3(32'h34c49d14),
	.w4(32'h34de9200),
	.w5(32'h3483b749),
	.w6(32'h350757d3),
	.w7(32'h356610ff),
	.w8(32'h356370b7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bc715),
	.w1(32'hb7f6147f),
	.w2(32'hb8b98b7f),
	.w3(32'hb97fa155),
	.w4(32'hb896ced1),
	.w5(32'hb7d0259d),
	.w6(32'h39d53e38),
	.w7(32'h39ce3856),
	.w8(32'h39aff41e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7981bc6),
	.w1(32'h37349ba5),
	.w2(32'hb80fd2de),
	.w3(32'h3755bcd2),
	.w4(32'h38f12bb3),
	.w5(32'h386a069e),
	.w6(32'h39432b20),
	.w7(32'h38c9df1c),
	.w8(32'hb75c1e2b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a6e23f),
	.w1(32'hb603ac99),
	.w2(32'hb70e7ac4),
	.w3(32'h34834ad7),
	.w4(32'hb59343e5),
	.w5(32'hb62fc634),
	.w6(32'h35c9f38e),
	.w7(32'hb60cacc5),
	.w8(32'hb695d840),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37301183),
	.w1(32'h372f6c79),
	.w2(32'h37095e7d),
	.w3(32'h3707d9b0),
	.w4(32'h374b1b65),
	.w5(32'h367212af),
	.w6(32'h372011db),
	.w7(32'h36f53b3d),
	.w8(32'h36e7472f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39037d3a),
	.w1(32'h3875a99c),
	.w2(32'h37e536c8),
	.w3(32'h376dad7e),
	.w4(32'hb89e5f1d),
	.w5(32'hb8ce55df),
	.w6(32'h38a8e958),
	.w7(32'hb881ed0e),
	.w8(32'hb91427ff),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bd6170),
	.w1(32'hb8658c44),
	.w2(32'hb7c9e44c),
	.w3(32'hb81e782e),
	.w4(32'hb8672709),
	.w5(32'hb80dd172),
	.w6(32'hb81c5a6a),
	.w7(32'hb894511a),
	.w8(32'hb81f1d2a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b5962c),
	.w1(32'hb7bb9b3a),
	.w2(32'hb5d48f48),
	.w3(32'hb8e8e076),
	.w4(32'hb93c744e),
	.w5(32'hb90f8aae),
	.w6(32'hb82402b4),
	.w7(32'hb90d47bb),
	.w8(32'hb922d3c0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a875c0),
	.w1(32'h38fd0de6),
	.w2(32'h38f1d42a),
	.w3(32'h386b5447),
	.w4(32'h388c66d9),
	.w5(32'h388ca783),
	.w6(32'h388f01bd),
	.w7(32'h388d5cbe),
	.w8(32'h384b9ece),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3796d737),
	.w1(32'h37d4c08d),
	.w2(32'h382a7bc4),
	.w3(32'hb61b696b),
	.w4(32'h380ca845),
	.w5(32'h3707832d),
	.w6(32'h37978aac),
	.w7(32'h37b0afc4),
	.w8(32'hb6c82c1f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378b21ec),
	.w1(32'h369ba288),
	.w2(32'hb7f7d42c),
	.w3(32'h37ef1e98),
	.w4(32'h3730b995),
	.w5(32'hb8c035cd),
	.w6(32'h394e0ea3),
	.w7(32'hb788806e),
	.w8(32'hb97c58d7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a54aa6),
	.w1(32'hb8c5d306),
	.w2(32'hb86d5667),
	.w3(32'hb89688fe),
	.w4(32'hb93ddbc6),
	.w5(32'hb9594040),
	.w6(32'hb8e036ba),
	.w7(32'hb96642be),
	.w8(32'hb934ad87),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b1171),
	.w1(32'hb80f96e4),
	.w2(32'hb84836fd),
	.w3(32'hb8269f97),
	.w4(32'hb81c32c1),
	.w5(32'hb83b77c8),
	.w6(32'hb770d3cd),
	.w7(32'hb82f0885),
	.w8(32'hb8472fe3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384daf36),
	.w1(32'h38d8554b),
	.w2(32'h392769ea),
	.w3(32'h390faa01),
	.w4(32'h3918c0ab),
	.w5(32'h38f07aa4),
	.w6(32'h396e2b9a),
	.w7(32'h3968ecd7),
	.w8(32'h39272c06),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931b3ee),
	.w1(32'hb94a570c),
	.w2(32'hb8989a79),
	.w3(32'hb9bc9839),
	.w4(32'hb96e82ae),
	.w5(32'hb92720b3),
	.w6(32'hb9bb84dc),
	.w7(32'hb9a956e6),
	.w8(32'hb94a7ad6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ed316),
	.w1(32'h39845593),
	.w2(32'h398adfd5),
	.w3(32'h39a59b24),
	.w4(32'h39b2da41),
	.w5(32'h39a0f260),
	.w6(32'h39ba9057),
	.w7(32'h39d896c7),
	.w8(32'h39bb9d83),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3854b205),
	.w1(32'h38b8f209),
	.w2(32'h38a503ce),
	.w3(32'hb79b7a1c),
	.w4(32'hb8d1d6d8),
	.w5(32'hb7a97063),
	.w6(32'hb8c85d35),
	.w7(32'hb8e4be46),
	.w8(32'hb83066ec),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b92d88),
	.w1(32'h39be4e4b),
	.w2(32'h39692b1a),
	.w3(32'h3988d56f),
	.w4(32'h39ed0802),
	.w5(32'h39abb7f4),
	.w6(32'h3906a369),
	.w7(32'h390a0d14),
	.w8(32'h3913f596),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3797e443),
	.w1(32'hb5d64c61),
	.w2(32'hb9113024),
	.w3(32'hb8b3fa0a),
	.w4(32'hb6d47100),
	.w5(32'hb972f332),
	.w6(32'hb987f672),
	.w7(32'hb8e31658),
	.w8(32'h38e10f72),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996c60c),
	.w1(32'hb750202f),
	.w2(32'h39864735),
	.w3(32'h38a80e3b),
	.w4(32'hb7bdd3b4),
	.w5(32'hb93eb816),
	.w6(32'h3a1698c5),
	.w7(32'h3931fb3a),
	.w8(32'h330469b8),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394cfdfd),
	.w1(32'h3c34cf40),
	.w2(32'hbb0ad9ae),
	.w3(32'h399385ec),
	.w4(32'h3bfeec25),
	.w5(32'hbc8e3b7a),
	.w6(32'hbc3eea47),
	.w7(32'hbbb92e39),
	.w8(32'hbc94bf0b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986e62c),
	.w1(32'h3c0f815e),
	.w2(32'hbd5e76c5),
	.w3(32'hbca4db9c),
	.w4(32'hbd1169bd),
	.w5(32'hbcc82cbd),
	.w6(32'hbbd60c0d),
	.w7(32'h3cb21c94),
	.w8(32'hbb3fe497),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule