module layer_10_featuremap_316(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391faa9c),
	.w1(32'hbb2f683c),
	.w2(32'h384a7f32),
	.w3(32'h3b1f58c6),
	.w4(32'h3b1d60ad),
	.w5(32'hbb762e83),
	.w6(32'hbb847d8f),
	.w7(32'hbad49f4b),
	.w8(32'hbb2e1510),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a803da),
	.w1(32'hba608aef),
	.w2(32'hbb36e433),
	.w3(32'hb9915e66),
	.w4(32'h3a9a808e),
	.w5(32'h3bafe450),
	.w6(32'hbb019bec),
	.w7(32'hbb8156d4),
	.w8(32'h3affa00d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63406b),
	.w1(32'hbb7902d8),
	.w2(32'hbb4ad348),
	.w3(32'hb80995ba),
	.w4(32'hbae78935),
	.w5(32'hbb8876b8),
	.w6(32'hbb3b5d09),
	.w7(32'hbb6d2601),
	.w8(32'hbb7f5325),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dc31a),
	.w1(32'hbb177782),
	.w2(32'hbac8763e),
	.w3(32'hbb4b5218),
	.w4(32'hbb01d18d),
	.w5(32'hbb96f721),
	.w6(32'hbb28299f),
	.w7(32'hba4986b3),
	.w8(32'hbbe96412),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb71caf),
	.w1(32'hbb89396a),
	.w2(32'hbb95f03e),
	.w3(32'hbb48f6f7),
	.w4(32'hbb9a1ed9),
	.w5(32'h3a73ad9c),
	.w6(32'hbbfa8186),
	.w7(32'hbbf8253a),
	.w8(32'h3ac7491a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1db590),
	.w1(32'h3b57363f),
	.w2(32'h3b5d1789),
	.w3(32'h380adc49),
	.w4(32'h3b86e92a),
	.w5(32'hbb84ef12),
	.w6(32'h3ad0e5d5),
	.w7(32'h3b789b0f),
	.w8(32'hbb8ce43a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298d0a),
	.w1(32'hbb431efc),
	.w2(32'hbb812930),
	.w3(32'hbb287bbc),
	.w4(32'hbb7049c1),
	.w5(32'hbaf82088),
	.w6(32'hbaa1b772),
	.w7(32'hbb9b2d19),
	.w8(32'hbb785c37),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2868f2),
	.w1(32'hbba0d569),
	.w2(32'h38f24c8e),
	.w3(32'hbbb1ea44),
	.w4(32'hbbbb019a),
	.w5(32'h3b8bc7da),
	.w6(32'hbb95ec14),
	.w7(32'hbb992a53),
	.w8(32'hbb0720aa),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5405c6),
	.w1(32'h3af35520),
	.w2(32'h3a7ed87f),
	.w3(32'h3af9541f),
	.w4(32'h3b96a162),
	.w5(32'hbaa60ebe),
	.w6(32'h3b5dc299),
	.w7(32'h3b51183d),
	.w8(32'hba6725e5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53ee21),
	.w1(32'h3acd1dc9),
	.w2(32'h3a444a61),
	.w3(32'hb9bf1e95),
	.w4(32'h3a9d3c83),
	.w5(32'hbb4c3574),
	.w6(32'h3a438443),
	.w7(32'h3ad131e4),
	.w8(32'hbb0fff1e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89594f),
	.w1(32'hbafcf6a7),
	.w2(32'hbabad2cb),
	.w3(32'hbb26efbb),
	.w4(32'hbb17e72a),
	.w5(32'h3989f820),
	.w6(32'hbb25df1c),
	.w7(32'hbaa8a700),
	.w8(32'hb9c25c03),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a345a77),
	.w1(32'hbab5c726),
	.w2(32'h3ac11f97),
	.w3(32'h3a0fb1da),
	.w4(32'hba8ce381),
	.w5(32'hbb04868f),
	.w6(32'h392900d8),
	.w7(32'hbae650aa),
	.w8(32'hbacfbc32),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f48ee),
	.w1(32'h3a042aed),
	.w2(32'hbb368d9a),
	.w3(32'h3ae72cf9),
	.w4(32'hba609465),
	.w5(32'hbbd2a953),
	.w6(32'hbab75419),
	.w7(32'hbb061d97),
	.w8(32'hbba8f7d6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbfd92),
	.w1(32'h3bc98141),
	.w2(32'h3b1e70c2),
	.w3(32'h3ba9f87c),
	.w4(32'h397da862),
	.w5(32'hbb000598),
	.w6(32'h3c10e9e0),
	.w7(32'h3a34f276),
	.w8(32'hbae3f43c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9c1fd),
	.w1(32'hbb1b4436),
	.w2(32'hbad790b1),
	.w3(32'hb9481023),
	.w4(32'h3a922410),
	.w5(32'hbbd217b1),
	.w6(32'h3a726f79),
	.w7(32'h3b023b04),
	.w8(32'hbbd4284d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc093ef8),
	.w1(32'hba0d528d),
	.w2(32'hbb69f810),
	.w3(32'hba96e28e),
	.w4(32'hbbce5fca),
	.w5(32'h3c08a073),
	.w6(32'hba33c12f),
	.w7(32'hbbdd6324),
	.w8(32'h3b91e408),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9dd52),
	.w1(32'h3b67f19b),
	.w2(32'h3be289a3),
	.w3(32'h3ba62ac3),
	.w4(32'h3c036582),
	.w5(32'h3a72932a),
	.w6(32'hba81efda),
	.w7(32'h3b8b14c5),
	.w8(32'h39a73b21),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9fb58),
	.w1(32'hbadc1a94),
	.w2(32'hbb0aa7ce),
	.w3(32'hbb25dee0),
	.w4(32'hb90ced06),
	.w5(32'h39876f1b),
	.w6(32'hbb123bbe),
	.w7(32'hbb48f017),
	.w8(32'hbb0ee89b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3e47c),
	.w1(32'hba56711e),
	.w2(32'h39cc56a1),
	.w3(32'hba64b556),
	.w4(32'h3a184ec1),
	.w5(32'hbaeeff2e),
	.w6(32'hbaf486bc),
	.w7(32'hba456d1a),
	.w8(32'h39cb3263),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b571ccb),
	.w1(32'h3c06038d),
	.w2(32'h3ad63de8),
	.w3(32'h3b7b0ec8),
	.w4(32'h3b1ec2ee),
	.w5(32'hbbf55222),
	.w6(32'h3bdb4373),
	.w7(32'hb93c893a),
	.w8(32'hbc1b74fc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb1b65),
	.w1(32'hbb1a8da1),
	.w2(32'hbb50702f),
	.w3(32'h3a842496),
	.w4(32'hbbb3c5b8),
	.w5(32'hba886eaf),
	.w6(32'hbb094ef3),
	.w7(32'hbbb57b20),
	.w8(32'hba714ace),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03bf0e),
	.w1(32'h39bb571f),
	.w2(32'h3b1abb9f),
	.w3(32'h3aacf46d),
	.w4(32'h3b4a1d31),
	.w5(32'h3ac9c168),
	.w6(32'hba471072),
	.w7(32'h3ad79481),
	.w8(32'h3af06ce9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f1ffe),
	.w1(32'hbb8dd8b0),
	.w2(32'hbac3c2be),
	.w3(32'hbb9fed30),
	.w4(32'h3908a7eb),
	.w5(32'hbc280cf1),
	.w6(32'hbb8ff8e9),
	.w7(32'h3ae8e68e),
	.w8(32'hbc6601c8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51db16),
	.w1(32'hbb353bb2),
	.w2(32'hbbf7d20f),
	.w3(32'hbb86cd61),
	.w4(32'hbc1acfda),
	.w5(32'hba8d0b62),
	.w6(32'hbaf2fce3),
	.w7(32'hbbe0cef2),
	.w8(32'hbb62853e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb154d07),
	.w1(32'hbb04a32a),
	.w2(32'hbb897fe2),
	.w3(32'hbaee6c28),
	.w4(32'hbb657b98),
	.w5(32'hbb2fe904),
	.w6(32'hbbc6f5c6),
	.w7(32'hbba6d058),
	.w8(32'hbb88470c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0edb94),
	.w1(32'hbb40960f),
	.w2(32'h3888b739),
	.w3(32'hba197733),
	.w4(32'h3ac25dd6),
	.w5(32'hba8b443f),
	.w6(32'hbac200d3),
	.w7(32'hba20450a),
	.w8(32'hbaa9de0d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f77135),
	.w1(32'hbb32d25a),
	.w2(32'hb9d8c848),
	.w3(32'hbb638aca),
	.w4(32'hbaa72e33),
	.w5(32'h3be868d7),
	.w6(32'hbb479503),
	.w7(32'hba91f8f0),
	.w8(32'h3baae0dc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14df6b),
	.w1(32'h3ba3ff58),
	.w2(32'h3b4f7a25),
	.w3(32'h3bea76fe),
	.w4(32'h3c22e16e),
	.w5(32'hbac21d2f),
	.w6(32'h3be0b848),
	.w7(32'h3b761b02),
	.w8(32'hba84946c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d9aba),
	.w1(32'h3b0dd691),
	.w2(32'hb8ff9dec),
	.w3(32'h3b0c1e30),
	.w4(32'hbb17337a),
	.w5(32'hbb3d6b12),
	.w6(32'h3b4c5255),
	.w7(32'hbb24705d),
	.w8(32'hbb5fdc98),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3adc79),
	.w1(32'hbb92df4d),
	.w2(32'hbb860cca),
	.w3(32'h3aa5922d),
	.w4(32'hb9c08564),
	.w5(32'hbbb7fb6c),
	.w6(32'hbb00a1d2),
	.w7(32'hb9d09678),
	.w8(32'h3ba82a13),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45a04c),
	.w1(32'h3a81bb53),
	.w2(32'hbb452daa),
	.w3(32'hbc13f59b),
	.w4(32'hbb8b3d5e),
	.w5(32'h3b85b52a),
	.w6(32'h3bb7b1e0),
	.w7(32'h3ab2035d),
	.w8(32'h3a23dcd8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050f57),
	.w1(32'hbbb8b8ea),
	.w2(32'hbb6fdc86),
	.w3(32'h3a95bd96),
	.w4(32'hbb05257a),
	.w5(32'h3a9413a3),
	.w6(32'hbb2a28a4),
	.w7(32'hbb16d156),
	.w8(32'h3aa435bd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bc957),
	.w1(32'hbb4a0216),
	.w2(32'hbabe43c6),
	.w3(32'hbb371111),
	.w4(32'hb9ceed2b),
	.w5(32'hbafeb5cd),
	.w6(32'hbaa1d2a5),
	.w7(32'hba4dc507),
	.w8(32'hba6514e9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25af92),
	.w1(32'hbb048eb0),
	.w2(32'hbabb20c8),
	.w3(32'hbb2330ad),
	.w4(32'hb81c6a1d),
	.w5(32'h3b02cece),
	.w6(32'hbb1df20d),
	.w7(32'hbac2e15c),
	.w8(32'hb9f91867),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4e139),
	.w1(32'hba274d9c),
	.w2(32'h39f2470c),
	.w3(32'h3a9d45e3),
	.w4(32'h37cf08bf),
	.w5(32'hba4453cd),
	.w6(32'hba2a10fa),
	.w7(32'h39cd9eeb),
	.w8(32'hbb57a89e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5586a0),
	.w1(32'hbae29343),
	.w2(32'hba194f0c),
	.w3(32'hbba0a144),
	.w4(32'hbb9f50e5),
	.w5(32'h3b0df961),
	.w6(32'hbba4333b),
	.w7(32'hbb587f71),
	.w8(32'h3a8173fb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895620),
	.w1(32'hbab1b109),
	.w2(32'h3b2d4c75),
	.w3(32'hbb78c14a),
	.w4(32'hba8bf3b5),
	.w5(32'h3b76cf50),
	.w6(32'hbae6f7f2),
	.w7(32'hba1a1c8a),
	.w8(32'hbb66991f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe7f08),
	.w1(32'hbb05bf4f),
	.w2(32'h3a81be61),
	.w3(32'h3958d814),
	.w4(32'h3b326901),
	.w5(32'h3abe9ca9),
	.w6(32'hbacb299f),
	.w7(32'h3b45a420),
	.w8(32'h3c0dee22),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bfa48),
	.w1(32'h3bcca180),
	.w2(32'hb8fd119a),
	.w3(32'h3ba63db2),
	.w4(32'h3bbc579e),
	.w5(32'hbb9ee28a),
	.w6(32'h3b96c934),
	.w7(32'h3b558c40),
	.w8(32'hbb03ac97),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf76aa9),
	.w1(32'h3a8eb289),
	.w2(32'h3bb7edf9),
	.w3(32'h3a53a158),
	.w4(32'h399ccab5),
	.w5(32'h3af60df2),
	.w6(32'hba1c8f44),
	.w7(32'h390e78e7),
	.w8(32'h3b8b574a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2667cf),
	.w1(32'h3bdf5edb),
	.w2(32'h3b8952fe),
	.w3(32'h3b3b4c7d),
	.w4(32'h3b27052b),
	.w5(32'hbb7de27a),
	.w6(32'h3bca93ad),
	.w7(32'h3b9e8017),
	.w8(32'hbbb83035),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93284a),
	.w1(32'hbba88de0),
	.w2(32'hbaf4f47a),
	.w3(32'hbb6045b0),
	.w4(32'hba9ee9a1),
	.w5(32'hba6574e9),
	.w6(32'hbbc7b8e0),
	.w7(32'hbb895e10),
	.w8(32'hba70d22e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c631d),
	.w1(32'h3b3aaa5c),
	.w2(32'h3a58ca80),
	.w3(32'hb69f53a5),
	.w4(32'h3b3bff4c),
	.w5(32'hb9affcaf),
	.w6(32'h3952d94e),
	.w7(32'h3b01a3ef),
	.w8(32'h3a611d53),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af59b0b),
	.w1(32'hb9dfd2ca),
	.w2(32'hbacf3a74),
	.w3(32'hbc078183),
	.w4(32'hb9d1a374),
	.w5(32'hbb046500),
	.w6(32'hbb8d4893),
	.w7(32'hb99f94ad),
	.w8(32'hba1f312c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf8f12),
	.w1(32'hbb5ad7d1),
	.w2(32'hbb6ff911),
	.w3(32'hbb58d365),
	.w4(32'hbb967263),
	.w5(32'h3ad1c2ad),
	.w6(32'hbb5b1cba),
	.w7(32'hbb095ffa),
	.w8(32'h3a9912f5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164062),
	.w1(32'hbb21baec),
	.w2(32'hb9982791),
	.w3(32'hbb1e7c83),
	.w4(32'hbaddb1e3),
	.w5(32'hbaf827eb),
	.w6(32'hbb85d6c7),
	.w7(32'hbb4885af),
	.w8(32'hbb61fd7c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb574442),
	.w1(32'hbb66a03c),
	.w2(32'hbb2d5171),
	.w3(32'hbb896da6),
	.w4(32'hbad54a0d),
	.w5(32'h3b66e91c),
	.w6(32'hbb725067),
	.w7(32'hbb1c1354),
	.w8(32'h3b0baab2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b970bb7),
	.w1(32'h3b3f9792),
	.w2(32'h3a12dee3),
	.w3(32'h3b419a2c),
	.w4(32'h3bb5a93f),
	.w5(32'hbb595d65),
	.w6(32'h3b203ecd),
	.w7(32'h3b08f618),
	.w8(32'hbb829317),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9227c2a),
	.w1(32'hba288ca4),
	.w2(32'hbb8421b8),
	.w3(32'hbb7509b6),
	.w4(32'hbb682e19),
	.w5(32'hbb1bc0e1),
	.w6(32'hbb18ccc9),
	.w7(32'hbb63c38b),
	.w8(32'hbb86a3a7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a3910),
	.w1(32'hbb6d0e51),
	.w2(32'h3a2f6ae1),
	.w3(32'h3894144d),
	.w4(32'h3ab397e3),
	.w5(32'hbaf4054a),
	.w6(32'hba797ae6),
	.w7(32'hb945db89),
	.w8(32'hbb958169),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90e4a4),
	.w1(32'hbb7c1b27),
	.w2(32'hbaf363b0),
	.w3(32'hbb91e198),
	.w4(32'h3a246107),
	.w5(32'h3aca2d1b),
	.w6(32'hbba669ff),
	.w7(32'hbb07fdc7),
	.w8(32'h3b36d941),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabc872),
	.w1(32'h3a3a952d),
	.w2(32'hb9b85db4),
	.w3(32'hbb3b6d17),
	.w4(32'hbaa02386),
	.w5(32'hbbd2a44d),
	.w6(32'hba2cb378),
	.w7(32'hb9a0f179),
	.w8(32'hbbaf1392),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba466cc),
	.w1(32'hbabc85c9),
	.w2(32'hbb16c5e3),
	.w3(32'hbb427176),
	.w4(32'hbbbf056b),
	.w5(32'hba4416ee),
	.w6(32'hbb44679a),
	.w7(32'hbb476b7a),
	.w8(32'hb90f9e12),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8614d4),
	.w1(32'hbb74199a),
	.w2(32'h3b2330cc),
	.w3(32'hbb134c4c),
	.w4(32'hbb7a4022),
	.w5(32'hba64c755),
	.w6(32'hb9e9f791),
	.w7(32'hba6cf253),
	.w8(32'h39ff388f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84138e9),
	.w1(32'h3b1c36de),
	.w2(32'hbaa0216a),
	.w3(32'h3a293e66),
	.w4(32'h3aae8456),
	.w5(32'hbaa0174b),
	.w6(32'h3ad5fab2),
	.w7(32'hba844d7a),
	.w8(32'hbb9bfc89),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28d587),
	.w1(32'hbb3aa4b4),
	.w2(32'hbb3aad68),
	.w3(32'h39e2552b),
	.w4(32'hba4c7c5e),
	.w5(32'h3b96ba46),
	.w6(32'hbb285dfe),
	.w7(32'hbaf89b64),
	.w8(32'h3ba0f912),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc64675),
	.w1(32'h3bf12c6b),
	.w2(32'h3b840777),
	.w3(32'h3ba33fe3),
	.w4(32'h3b4771d7),
	.w5(32'hbab72bc2),
	.w6(32'h3bbde0cd),
	.w7(32'h3b99f678),
	.w8(32'hbaef9cb3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e1ae7),
	.w1(32'h3a1f4688),
	.w2(32'h3aa6f480),
	.w3(32'h3b98ba68),
	.w4(32'hbabbed4b),
	.w5(32'hbaf8175e),
	.w6(32'h3b35955a),
	.w7(32'hba7b9a3d),
	.w8(32'hbb7725a6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae69a07),
	.w1(32'hbb7dc9ef),
	.w2(32'h3ab088c0),
	.w3(32'h39f1bf7d),
	.w4(32'h3a94199f),
	.w5(32'h3be04460),
	.w6(32'h3a68a156),
	.w7(32'h3a0ed2fd),
	.w8(32'h3bad56c9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9af78a),
	.w1(32'hb80ae6a3),
	.w2(32'h37f121d8),
	.w3(32'hba568f02),
	.w4(32'h39abf6cf),
	.w5(32'hbb5e462c),
	.w6(32'hbba24b8f),
	.w7(32'hbb139298),
	.w8(32'h3acbe9e1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01741a),
	.w1(32'h3ae3d3a4),
	.w2(32'hba1018ea),
	.w3(32'hbae8568c),
	.w4(32'h3b3989bf),
	.w5(32'hbb815e00),
	.w6(32'hba2cbb3f),
	.w7(32'hb989f4c6),
	.w8(32'hbb2ca612),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919dc1),
	.w1(32'hba60472e),
	.w2(32'hba4ad8fc),
	.w3(32'hbb47271d),
	.w4(32'hba988c46),
	.w5(32'hbb1dbf40),
	.w6(32'hb9a63b75),
	.w7(32'hbaeeb7a4),
	.w8(32'hba96f562),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f9f66),
	.w1(32'hb99cc2a5),
	.w2(32'hbacd55ee),
	.w3(32'hbb4fd776),
	.w4(32'hbb838963),
	.w5(32'h39743a63),
	.w6(32'hbb6728fe),
	.w7(32'hbb6817c7),
	.w8(32'h37ea37d0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ca542),
	.w1(32'h3a14face),
	.w2(32'h3a9b93b4),
	.w3(32'h38a957e8),
	.w4(32'h38d431e6),
	.w5(32'h3b2ed54f),
	.w6(32'h3aa3b9fe),
	.w7(32'h3ab9e4ec),
	.w8(32'h3acc304b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a829ffd),
	.w1(32'h3a1689b9),
	.w2(32'hbb49d0a2),
	.w3(32'h3b0ee084),
	.w4(32'hba356bab),
	.w5(32'hbb84b3e5),
	.w6(32'h3a64921e),
	.w7(32'hba9d82c4),
	.w8(32'hbbb71675),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2842a1),
	.w1(32'hbb721b59),
	.w2(32'hbb86dd9f),
	.w3(32'hbba131a9),
	.w4(32'hbb622877),
	.w5(32'hba4bad3b),
	.w6(32'hbbea46fe),
	.w7(32'hbb8c1796),
	.w8(32'hba3cd241),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961d26),
	.w1(32'h3ae56165),
	.w2(32'h3bc923c4),
	.w3(32'h3a93723f),
	.w4(32'h39f901cc),
	.w5(32'h3b36d3c2),
	.w6(32'h3b6faa1d),
	.w7(32'h3b52a903),
	.w8(32'h3b7a41e4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e322a),
	.w1(32'h3b1cd180),
	.w2(32'h3b9698b0),
	.w3(32'hba977183),
	.w4(32'h3acb1037),
	.w5(32'h3b62b11a),
	.w6(32'h3bc83def),
	.w7(32'h3ba9e88b),
	.w8(32'hba08d501),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38198d2f),
	.w1(32'hbab63f08),
	.w2(32'hba66b545),
	.w3(32'h3b2a32fd),
	.w4(32'h3aa4be47),
	.w5(32'h3b0aaf7d),
	.w6(32'h3a9a3539),
	.w7(32'hbb04f722),
	.w8(32'h3af8ae8a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdf075),
	.w1(32'h3a4c13ff),
	.w2(32'h3b08c736),
	.w3(32'hbb3cc1ca),
	.w4(32'h3b3e8208),
	.w5(32'hba81c574),
	.w6(32'hbb719c21),
	.w7(32'h3a854ac1),
	.w8(32'hb7a9b078),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82cf76e),
	.w1(32'hbac0cf6e),
	.w2(32'hb8e5f95a),
	.w3(32'hba8c76e4),
	.w4(32'hb7c79251),
	.w5(32'h3a00b52a),
	.w6(32'hbadd43d4),
	.w7(32'h39d224b6),
	.w8(32'hba678ef1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3be02),
	.w1(32'h3be3e616),
	.w2(32'h3b9cf42d),
	.w3(32'h3bed83a3),
	.w4(32'hbb3927a7),
	.w5(32'h3b73bb71),
	.w6(32'h3beeedd6),
	.w7(32'hb8ceeee1),
	.w8(32'h3bf051a4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b0a6e),
	.w1(32'h3bfd9378),
	.w2(32'h3bb98cc4),
	.w3(32'h3a696c36),
	.w4(32'h3b120d10),
	.w5(32'h3afb09e1),
	.w6(32'h3bf0c9c4),
	.w7(32'h3c07a3ce),
	.w8(32'h3b9d97a4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d2942),
	.w1(32'h3b12b730),
	.w2(32'hbb388349),
	.w3(32'hb98f9a97),
	.w4(32'hba3adb9c),
	.w5(32'hba164ef3),
	.w6(32'h39705c05),
	.w7(32'hbba8abde),
	.w8(32'h3a9e4635),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a775cf7),
	.w1(32'h3aed05e2),
	.w2(32'h3b6b373b),
	.w3(32'hb843df5d),
	.w4(32'h3b0504c2),
	.w5(32'h3b6673db),
	.w6(32'h3a5153ea),
	.w7(32'h3b6215b4),
	.w8(32'h3b49884b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb124c3),
	.w1(32'h3b1fd900),
	.w2(32'hbb819f8b),
	.w3(32'h39e85d8a),
	.w4(32'hba6efc5d),
	.w5(32'hbad95f24),
	.w6(32'hba1d944e),
	.w7(32'hbb412151),
	.w8(32'hbafb3aee),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62354b),
	.w1(32'hbb144cc2),
	.w2(32'hbb2c63aa),
	.w3(32'hbb9db296),
	.w4(32'hbb0cdbaf),
	.w5(32'h3a036aac),
	.w6(32'hbb84bdca),
	.w7(32'hbac90fa2),
	.w8(32'hbb0605b7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa0c8e),
	.w1(32'h39bf61bc),
	.w2(32'h3aec3c54),
	.w3(32'hb98f3f72),
	.w4(32'h3aabb9db),
	.w5(32'h3ab36f00),
	.w6(32'hba46f9af),
	.w7(32'h3b0a3a81),
	.w8(32'h3b008827),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb075213),
	.w1(32'hba7335c7),
	.w2(32'h3a040cfb),
	.w3(32'hbae23319),
	.w4(32'hbb4d5a28),
	.w5(32'h3b413d78),
	.w6(32'h3aabd906),
	.w7(32'hba819299),
	.w8(32'h3b7b9f60),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eeb330),
	.w1(32'h3b03597d),
	.w2(32'h3b30d847),
	.w3(32'h3a464a9c),
	.w4(32'h3b545a18),
	.w5(32'hbb1e96e1),
	.w6(32'h3b38d589),
	.w7(32'h3ac0c2f9),
	.w8(32'hbbf125b2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f1943),
	.w1(32'hbab43306),
	.w2(32'hb98b3e99),
	.w3(32'hb9a451f9),
	.w4(32'hba999629),
	.w5(32'h3b126a8e),
	.w6(32'hbb01800e),
	.w7(32'h3aa70150),
	.w8(32'h3b6ec40a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2c4ef),
	.w1(32'h3b8a50a0),
	.w2(32'hb91d0061),
	.w3(32'h3a68aa6b),
	.w4(32'h3a335b8e),
	.w5(32'h3aecec50),
	.w6(32'h3b013d1b),
	.w7(32'hba9db5d1),
	.w8(32'h3af86194),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8b22d),
	.w1(32'hba98756e),
	.w2(32'h39c84640),
	.w3(32'hba32c8fd),
	.w4(32'hba246200),
	.w5(32'hbbcc0880),
	.w6(32'hb8a71e5f),
	.w7(32'hba2fdd3d),
	.w8(32'hbbb7119a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96bf75),
	.w1(32'hbb645b13),
	.w2(32'hbaf3abdf),
	.w3(32'hbbb46a64),
	.w4(32'hbb5b12a1),
	.w5(32'h3b57721c),
	.w6(32'hbb72bffa),
	.w7(32'hba65c42d),
	.w8(32'h3b26014c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a692f3b),
	.w1(32'hbb0ebf59),
	.w2(32'hbb0bd181),
	.w3(32'h39c06a57),
	.w4(32'h398a4732),
	.w5(32'h3a3d3a97),
	.w6(32'hbab7c83a),
	.w7(32'hba4d9c08),
	.w8(32'h3b435e90),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a8388),
	.w1(32'hba7cb809),
	.w2(32'hbb9170dd),
	.w3(32'hbabe105a),
	.w4(32'hbb7b0069),
	.w5(32'h3aba1b2d),
	.w6(32'h3a524799),
	.w7(32'hbb54b18e),
	.w8(32'h3aa8defb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f6957),
	.w1(32'hba2cbb39),
	.w2(32'h3b1f2137),
	.w3(32'h3b13ab09),
	.w4(32'h36bb3344),
	.w5(32'hbb735b3c),
	.w6(32'h3a3cede0),
	.w7(32'hbad917be),
	.w8(32'hba8c7901),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2565a),
	.w1(32'hb8d63d1d),
	.w2(32'hba82848c),
	.w3(32'hbb451309),
	.w4(32'h38438825),
	.w5(32'hb88985ec),
	.w6(32'hbb0d1334),
	.w7(32'hba948949),
	.w8(32'hb88eb770),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fc6ad),
	.w1(32'hba086dfe),
	.w2(32'h38a3e8c1),
	.w3(32'hb8fc658a),
	.w4(32'h3b2ce93d),
	.w5(32'hbbc9633b),
	.w6(32'h3a91fc7c),
	.w7(32'h3b2034c4),
	.w8(32'hbbfa462a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf9f61),
	.w1(32'hbbb96838),
	.w2(32'hbb5ccb94),
	.w3(32'hbae16f7c),
	.w4(32'hba190613),
	.w5(32'hbb26108e),
	.w6(32'hbbb3228c),
	.w7(32'hbb159e19),
	.w8(32'hbae947f6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac542f6),
	.w1(32'hbb933ebd),
	.w2(32'hba80fffd),
	.w3(32'hbb9740e2),
	.w4(32'h3b733ca1),
	.w5(32'hbbb8945f),
	.w6(32'hbb25ef25),
	.w7(32'hb8ac3232),
	.w8(32'hbb9d5ab0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedd197),
	.w1(32'hbbad04eb),
	.w2(32'hba9fd5e8),
	.w3(32'hbba2bd0f),
	.w4(32'h397b8130),
	.w5(32'h397f0f89),
	.w6(32'hbb2606b8),
	.w7(32'h3a5b0b40),
	.w8(32'hbb6ddc7a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7464b8),
	.w1(32'hbc0aa6a9),
	.w2(32'hbba0b4a6),
	.w3(32'hbabeaca5),
	.w4(32'hbb65c65c),
	.w5(32'hbb1c6260),
	.w6(32'hbbd10c0f),
	.w7(32'hbbddc645),
	.w8(32'hbb751628),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7e713),
	.w1(32'hbc1244f5),
	.w2(32'hbb5d81ad),
	.w3(32'hbc025548),
	.w4(32'hbb3a2b8e),
	.w5(32'h3b388a04),
	.w6(32'hbbc4875a),
	.w7(32'hbb6cab31),
	.w8(32'h38bd248b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae43d42),
	.w1(32'h3a4ecb34),
	.w2(32'h3b1b2c7f),
	.w3(32'h3b8c9296),
	.w4(32'h3ac171a7),
	.w5(32'h3b4b5a38),
	.w6(32'h3ba24513),
	.w7(32'h3b1d4aa6),
	.w8(32'h3a8dd2e2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b777b0c),
	.w1(32'h39c18cce),
	.w2(32'h3b035cdb),
	.w3(32'hba624e70),
	.w4(32'h3b7cc878),
	.w5(32'hbadb27d4),
	.w6(32'h3b164d3e),
	.w7(32'h3bd24c6f),
	.w8(32'h3af0c0da),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a2644),
	.w1(32'h3aef745a),
	.w2(32'hba881c1d),
	.w3(32'h3a0d695a),
	.w4(32'hbaa3f9c2),
	.w5(32'h3acc5d61),
	.w6(32'hb6917836),
	.w7(32'hbb284f3d),
	.w8(32'h3a5fdacd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c75f9),
	.w1(32'h39c6114e),
	.w2(32'hbafd5b83),
	.w3(32'hbadde9da),
	.w4(32'h3aaadd30),
	.w5(32'hbc21d9ee),
	.w6(32'h3b07224e),
	.w7(32'h3b0dd998),
	.w8(32'hbc211e45),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941754),
	.w1(32'h38d3939f),
	.w2(32'hbb151a1d),
	.w3(32'hbb0ddb5b),
	.w4(32'hbaa3bcf8),
	.w5(32'hbc6a7ddc),
	.w6(32'hb9a1981c),
	.w7(32'hbb83adb0),
	.w8(32'hbc401c3e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d071b),
	.w1(32'h3c18478c),
	.w2(32'h3c551451),
	.w3(32'hbc95afb7),
	.w4(32'h3b9e6257),
	.w5(32'hbbbac84f),
	.w6(32'hbc9d6ae1),
	.w7(32'h3c9e89d2),
	.w8(32'hbcb2cc92),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b457029),
	.w1(32'h3c1dd286),
	.w2(32'h3c4a1f59),
	.w3(32'hbbef77b5),
	.w4(32'h3b8330c6),
	.w5(32'hbb586fe4),
	.w6(32'hbbc3bc55),
	.w7(32'h3be0c4c0),
	.w8(32'h3baee0c5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bf0b2),
	.w1(32'h3ad949e1),
	.w2(32'h3bc27348),
	.w3(32'h3b3852d1),
	.w4(32'hbc04ebc2),
	.w5(32'hbbbfe901),
	.w6(32'hbc1006c0),
	.w7(32'h3bdf3fa3),
	.w8(32'hbbade0c3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadba49),
	.w1(32'h3b65c6d7),
	.w2(32'h3ba88b9b),
	.w3(32'hbb8e63a1),
	.w4(32'h3bacfc92),
	.w5(32'hbbfd8451),
	.w6(32'h3ba173a7),
	.w7(32'h3c17f899),
	.w8(32'hbc86b4ca),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ae11d),
	.w1(32'h3b8727ac),
	.w2(32'h3cfc7fc8),
	.w3(32'hbc3d1102),
	.w4(32'h3ba85c8e),
	.w5(32'hbb89b6ba),
	.w6(32'hbc8e2927),
	.w7(32'h3ca9ed91),
	.w8(32'h3a6e4526),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a1bd1),
	.w1(32'h3b9fbff2),
	.w2(32'h3b7f61dd),
	.w3(32'h3aafc1da),
	.w4(32'hbbec7652),
	.w5(32'hbc3cde57),
	.w6(32'h3c044526),
	.w7(32'h3caa974d),
	.w8(32'hbc86b5d2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0574e6),
	.w1(32'hbb1d1a55),
	.w2(32'h3be7dfae),
	.w3(32'hbc15e9fb),
	.w4(32'h3b18539b),
	.w5(32'hbcb4b463),
	.w6(32'hbc66e5e7),
	.w7(32'h39b25b1e),
	.w8(32'hbc83acd0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc833bd7),
	.w1(32'hbc454066),
	.w2(32'h3c4d95fd),
	.w3(32'hbc1310b7),
	.w4(32'hba280f50),
	.w5(32'hb9560f6a),
	.w6(32'hbc159f6c),
	.w7(32'h3b99fcae),
	.w8(32'hba52cc6d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e63c4),
	.w1(32'h398d839f),
	.w2(32'h3ab986f0),
	.w3(32'h39734348),
	.w4(32'hbac8423b),
	.w5(32'hbce7251c),
	.w6(32'h3a7a638e),
	.w7(32'h3adf1468),
	.w8(32'hbccf6aa3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91363b),
	.w1(32'hbba6128b),
	.w2(32'hb90c671a),
	.w3(32'hbc7594e2),
	.w4(32'hbbda8429),
	.w5(32'h3ab7c290),
	.w6(32'hbc5ca5ab),
	.w7(32'hbb99f0bd),
	.w8(32'h3b04601f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e3a3e),
	.w1(32'hbb9bd4cc),
	.w2(32'hbbf1bc1f),
	.w3(32'h3bb6bfd5),
	.w4(32'hbb7a3a3e),
	.w5(32'hb9fb151a),
	.w6(32'h3b7935e1),
	.w7(32'hbb0a3207),
	.w8(32'hbae63f2d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b268e3),
	.w1(32'hbac12c81),
	.w2(32'h3ac5c16b),
	.w3(32'hbb08c7a8),
	.w4(32'hbbfe4877),
	.w5(32'hbb19b57f),
	.w6(32'h36c0f799),
	.w7(32'h3b7b856e),
	.w8(32'h3ac09693),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea9989),
	.w1(32'hbb32cd42),
	.w2(32'hbb6889ac),
	.w3(32'hbb0a295c),
	.w4(32'hbb7ceb08),
	.w5(32'h3c8b743a),
	.w6(32'hbb0957f9),
	.w7(32'hbb83f7ed),
	.w8(32'h3cbee555),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be555c2),
	.w1(32'hbc0cd69f),
	.w2(32'hbcdbd6d9),
	.w3(32'h3c254779),
	.w4(32'hbbd572cc),
	.w5(32'h3b3b7831),
	.w6(32'h3c4c2a0f),
	.w7(32'hbcbbbfc8),
	.w8(32'hbbe1b456),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f47a3),
	.w1(32'h3bf90d8e),
	.w2(32'h3af2bd2d),
	.w3(32'hbb7e010c),
	.w4(32'hbaca90c1),
	.w5(32'h39608b3b),
	.w6(32'hbbff2253),
	.w7(32'hba12615c),
	.w8(32'hba964ba3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44864c),
	.w1(32'h3b5ea8fd),
	.w2(32'h3c7cfd9d),
	.w3(32'hbbb91c18),
	.w4(32'hba795571),
	.w5(32'hb8e3a9f8),
	.w6(32'hbc71c01e),
	.w7(32'h3c14163a),
	.w8(32'h39f1c21d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d831c),
	.w1(32'hbb09345b),
	.w2(32'hbb10d485),
	.w3(32'h3a19a94c),
	.w4(32'h3a5ca6bb),
	.w5(32'h3a1fc9f5),
	.w6(32'hbc15ebb6),
	.w7(32'h3a59a8b9),
	.w8(32'hbb703d6f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5fee2),
	.w1(32'hbaa4849a),
	.w2(32'hbbdc6a47),
	.w3(32'hbb4a30f2),
	.w4(32'h3a77217b),
	.w5(32'hbc28bb30),
	.w6(32'hbb8236e0),
	.w7(32'hbb799b2f),
	.w8(32'hbb624311),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84554c),
	.w1(32'h3b7eb8d5),
	.w2(32'h3c2c4437),
	.w3(32'hb923e5e6),
	.w4(32'hbb13f435),
	.w5(32'h39fea1d0),
	.w6(32'hbb213020),
	.w7(32'h3c10d67d),
	.w8(32'hbb891991),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda2382),
	.w1(32'h3adb1298),
	.w2(32'hbc291d88),
	.w3(32'h3b5db49c),
	.w4(32'hbbcd0d02),
	.w5(32'hbca84184),
	.w6(32'h3bc25862),
	.w7(32'hbb58c10b),
	.w8(32'hbcd41d4d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1530b9),
	.w1(32'hbbb21deb),
	.w2(32'h3ae8f360),
	.w3(32'hbc3e3e28),
	.w4(32'hbb22ffce),
	.w5(32'h3b2da406),
	.w6(32'hbcb8a850),
	.w7(32'hbb20ffff),
	.w8(32'h3bbeb8de),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d8edf),
	.w1(32'h3afafc0c),
	.w2(32'h3bac0b51),
	.w3(32'hb9ec9071),
	.w4(32'h3bc77dfe),
	.w5(32'hbaf9f775),
	.w6(32'hbc01adb5),
	.w7(32'h3c302008),
	.w8(32'hbbadae70),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc013e9e),
	.w1(32'hbbc8a9bf),
	.w2(32'hbbb7d8a0),
	.w3(32'h3bdb4d3e),
	.w4(32'h39e20605),
	.w5(32'h3b5d3670),
	.w6(32'h3bd4e738),
	.w7(32'h390cc356),
	.w8(32'h3c4c2c35),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94cffd),
	.w1(32'h39be9d58),
	.w2(32'hbc5fdcae),
	.w3(32'h3c42a19b),
	.w4(32'hbb8cbd3e),
	.w5(32'h3a2f9d49),
	.w6(32'h3bafc64c),
	.w7(32'hbc1f7364),
	.w8(32'h3bff30f8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5f34f),
	.w1(32'hbc1e937f),
	.w2(32'hbc6732c7),
	.w3(32'hba0d968b),
	.w4(32'hbc4a8a6a),
	.w5(32'hbbb75d41),
	.w6(32'h3ba0daee),
	.w7(32'hbc3545f6),
	.w8(32'h3c473246),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98ecab),
	.w1(32'h3bb78e73),
	.w2(32'hbc747cdd),
	.w3(32'h39e10d78),
	.w4(32'hbb486f69),
	.w5(32'h3c2b50a1),
	.w6(32'h3c2fbff3),
	.w7(32'hbae8f590),
	.w8(32'h3c0f3255),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0d888),
	.w1(32'h3a8d74d0),
	.w2(32'hbb218dd7),
	.w3(32'h3abee898),
	.w4(32'hbb89e3e9),
	.w5(32'hbb7bb40a),
	.w6(32'hbb34a8d7),
	.w7(32'h387163d6),
	.w8(32'hbb5122c7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb57e15),
	.w1(32'hbbe24d54),
	.w2(32'hbc58c2c7),
	.w3(32'h39f75201),
	.w4(32'hbbcca8bf),
	.w5(32'h3bfb8fe5),
	.w6(32'h3b9f4ed1),
	.w7(32'hbac63303),
	.w8(32'hbb0d2b44),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd986e),
	.w1(32'h3c18841e),
	.w2(32'h3c605187),
	.w3(32'h3b2485de),
	.w4(32'h3a347c79),
	.w5(32'hbae0d329),
	.w6(32'hbb94b5a2),
	.w7(32'h3afd4b4b),
	.w8(32'h3b0df264),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecf994),
	.w1(32'hbc466513),
	.w2(32'hbc8494ad),
	.w3(32'hbb8b7dd8),
	.w4(32'hbc7e2c2f),
	.w5(32'h3b96e2c0),
	.w6(32'hbbfc63ce),
	.w7(32'hbc85c466),
	.w8(32'h3bfa479e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae91a8f),
	.w1(32'h3ad678b9),
	.w2(32'hbc717f27),
	.w3(32'h3b004de4),
	.w4(32'h3b74c1ee),
	.w5(32'hbb8dfc1a),
	.w6(32'h3c454cdb),
	.w7(32'h3a00986a),
	.w8(32'hbb15ccc0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c154890),
	.w1(32'h399ee02d),
	.w2(32'h391b33d0),
	.w3(32'hbaba68b7),
	.w4(32'hbb20b129),
	.w5(32'hbba9dbfa),
	.w6(32'hbb914273),
	.w7(32'hbbf072a5),
	.w8(32'hb79722d8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bee78f),
	.w1(32'hbb7f8aae),
	.w2(32'hbc1037da),
	.w3(32'h3a7a0ad6),
	.w4(32'hbb0fca20),
	.w5(32'h3bcf4e48),
	.w6(32'h3b4c1b72),
	.w7(32'hbbd45357),
	.w8(32'hbae04b4b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0c5fb),
	.w1(32'h3bb00b63),
	.w2(32'h3bc82201),
	.w3(32'h3afcda9b),
	.w4(32'h3c3443e5),
	.w5(32'h3b1bd5d2),
	.w6(32'hbc32254c),
	.w7(32'h3bbebf25),
	.w8(32'h3c13b01f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab10134),
	.w1(32'h3b1de81f),
	.w2(32'hbbd436ba),
	.w3(32'h3c30b862),
	.w4(32'hbaa44727),
	.w5(32'h3a94b5e1),
	.w6(32'h3c43fc36),
	.w7(32'h39063f6b),
	.w8(32'h3beb1a82),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c121d),
	.w1(32'hbb998afa),
	.w2(32'hbc8d2dd7),
	.w3(32'h39aa837f),
	.w4(32'hbb9cb6d2),
	.w5(32'hbb6bf14b),
	.w6(32'h3b854a93),
	.w7(32'hbc3a7040),
	.w8(32'hbba667e9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50b635),
	.w1(32'hbb9a0e0b),
	.w2(32'hbbdcc9f3),
	.w3(32'hbb6843d1),
	.w4(32'hbb360cf7),
	.w5(32'h3c0a0a4e),
	.w6(32'hbba2830e),
	.w7(32'hbb7bf687),
	.w8(32'h3c6f4682),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4717ad),
	.w1(32'hbbead4be),
	.w2(32'hbcb2567e),
	.w3(32'h3b48f2da),
	.w4(32'hbb82c894),
	.w5(32'h3b560ca7),
	.w6(32'h390b569d),
	.w7(32'hbc80e2d4),
	.w8(32'h3bf64252),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23db85),
	.w1(32'h3b952085),
	.w2(32'hbb8b7a00),
	.w3(32'h3c1bd520),
	.w4(32'h3a21caba),
	.w5(32'h3adee99c),
	.w6(32'h3c4346cd),
	.w7(32'h3ac1261e),
	.w8(32'h3bf3316e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b272242),
	.w1(32'h3a9495dd),
	.w2(32'hbbac2290),
	.w3(32'h3c2acf74),
	.w4(32'h3a967538),
	.w5(32'h3b9adea2),
	.w6(32'h3bf90d3b),
	.w7(32'hbba01d51),
	.w8(32'hbb2cc78a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b435d76),
	.w1(32'h3b8c8934),
	.w2(32'h3b8172b9),
	.w3(32'hbb30237e),
	.w4(32'h3bebba1e),
	.w5(32'h3b01e33d),
	.w6(32'hb9f1f66a),
	.w7(32'h3b972f6b),
	.w8(32'h3c85c534),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbbc88),
	.w1(32'h3b7dfe13),
	.w2(32'hbc272568),
	.w3(32'h3c1baba0),
	.w4(32'hbc029f97),
	.w5(32'hbbabd42d),
	.w6(32'h3c594b48),
	.w7(32'hba279182),
	.w8(32'hbb81a4f7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd780),
	.w1(32'hbb0bb22e),
	.w2(32'h3b0cc612),
	.w3(32'hbb2591e7),
	.w4(32'hbaa4138a),
	.w5(32'h39e0d126),
	.w6(32'h3c3acbc5),
	.w7(32'h3c099750),
	.w8(32'h3ae6b19f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f881),
	.w1(32'hbbb38602),
	.w2(32'hbbaf4b64),
	.w3(32'h3b4f58ad),
	.w4(32'hbb8e33bf),
	.w5(32'h3b4592bd),
	.w6(32'h3b68ee9d),
	.w7(32'hbbbc0942),
	.w8(32'h3ab0b938),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd1443),
	.w1(32'hbc33f4fa),
	.w2(32'hbba4fe14),
	.w3(32'hbb189dcb),
	.w4(32'hbacf9709),
	.w5(32'hba8e0c72),
	.w6(32'h3c1d4f63),
	.w7(32'hbbbcba96),
	.w8(32'h3b95ee95),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e5a7d),
	.w1(32'hbb445263),
	.w2(32'hbc101db0),
	.w3(32'h3b89c586),
	.w4(32'h3b4c72d2),
	.w5(32'hbc22c4fe),
	.w6(32'h3be22d37),
	.w7(32'h3b6981ec),
	.w8(32'hbc0c0686),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf13a3),
	.w1(32'h3ab957d4),
	.w2(32'h3b972802),
	.w3(32'hbbaf7c69),
	.w4(32'hbb3f9cf0),
	.w5(32'hbc34682e),
	.w6(32'hbc217c11),
	.w7(32'h3b3e538e),
	.w8(32'hbc44e994),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3b51d),
	.w1(32'h3b9bc12a),
	.w2(32'h3b7c6733),
	.w3(32'hbc5f803e),
	.w4(32'hbc050f68),
	.w5(32'h3b7781b8),
	.w6(32'hbc40d85e),
	.w7(32'h3c5ac094),
	.w8(32'h3b819c79),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b542e),
	.w1(32'hbb84d81f),
	.w2(32'hbb1516a7),
	.w3(32'hbb789b8b),
	.w4(32'hbc23eb48),
	.w5(32'h3b802106),
	.w6(32'hbb9d440f),
	.w7(32'hbbc3f0b3),
	.w8(32'h3b2cdedb),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3822a),
	.w1(32'hbbc5318f),
	.w2(32'hbc6e3dd4),
	.w3(32'hbb90f101),
	.w4(32'hbb68b1e4),
	.w5(32'hbbcb1699),
	.w6(32'h3c26b948),
	.w7(32'hbb8547a1),
	.w8(32'hbc10cdc6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac29d11),
	.w1(32'h3a1b5e28),
	.w2(32'h3b1310d9),
	.w3(32'hbb3b1269),
	.w4(32'h3bb5c681),
	.w5(32'hbbc13fd0),
	.w6(32'hbb9b4644),
	.w7(32'h3b8c0392),
	.w8(32'hbb9a3946),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1892a0),
	.w1(32'h3b6977f4),
	.w2(32'h3b9eff2f),
	.w3(32'hbaac1a27),
	.w4(32'h3b110daa),
	.w5(32'h3bef22aa),
	.w6(32'h3ba2efa9),
	.w7(32'h3b80766a),
	.w8(32'h3ca88a64),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1326e),
	.w1(32'hbc82a9cf),
	.w2(32'hbc168149),
	.w3(32'h3bf9c641),
	.w4(32'hbc0ade48),
	.w5(32'hb9b11d00),
	.w6(32'hbb5bc0e6),
	.w7(32'hbc744b67),
	.w8(32'hbb402840),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba291501),
	.w1(32'hba88c775),
	.w2(32'h3bac3694),
	.w3(32'h3997143e),
	.w4(32'hbb38cabf),
	.w5(32'hbb14060a),
	.w6(32'hbc08d9b4),
	.w7(32'hbaa4eff6),
	.w8(32'hbb205ebf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb6e20),
	.w1(32'h3bcd1585),
	.w2(32'h3abb8d62),
	.w3(32'hbb67495c),
	.w4(32'hba3dad9c),
	.w5(32'hbc402551),
	.w6(32'h3c126313),
	.w7(32'h3a5d93a2),
	.w8(32'hbc599377),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf70c63),
	.w1(32'h3bb8a75a),
	.w2(32'h3c692398),
	.w3(32'hbb85336c),
	.w4(32'h3bebcfeb),
	.w5(32'hb85c7b0b),
	.w6(32'h3a83a1b5),
	.w7(32'h3bf65da2),
	.w8(32'h3b1f9f73),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c678),
	.w1(32'hbc4f7e9e),
	.w2(32'hbc8017fd),
	.w3(32'hbbb21d1c),
	.w4(32'hbc143d59),
	.w5(32'h39dcab88),
	.w6(32'hbb96c738),
	.w7(32'hbc23e8dd),
	.w8(32'h3bbe2927),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb96d7c),
	.w1(32'hbbdaa93b),
	.w2(32'hbb5f68a1),
	.w3(32'hbb770e30),
	.w4(32'hbbea2b51),
	.w5(32'hba8e4b98),
	.w6(32'hba19e6bc),
	.w7(32'hbb730bc3),
	.w8(32'hbb9c4e64),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedcda9),
	.w1(32'hbb9ded4f),
	.w2(32'hbb1593ba),
	.w3(32'h3be7c396),
	.w4(32'hbb8bfa70),
	.w5(32'h3b168612),
	.w6(32'h3b65ae8b),
	.w7(32'h3bb2ac49),
	.w8(32'h3b0fb80b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd73937),
	.w1(32'hbc58326d),
	.w2(32'hbbb586ec),
	.w3(32'h3a71bce3),
	.w4(32'hba4c6cdb),
	.w5(32'hbbc247b4),
	.w6(32'hbc8af2b2),
	.w7(32'hbc1e93f8),
	.w8(32'hbb6165b4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b435357),
	.w1(32'hbbad77f1),
	.w2(32'hbc1738c1),
	.w3(32'hbbfe039e),
	.w4(32'hbac2ae23),
	.w5(32'h3c20a212),
	.w6(32'hbbd9be86),
	.w7(32'hbb8079a9),
	.w8(32'h3b84b2d7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b908cbc),
	.w1(32'h3b95600e),
	.w2(32'h3bbe7ba2),
	.w3(32'hbc4bcafb),
	.w4(32'h3bbfa593),
	.w5(32'hbc526a1c),
	.w6(32'hbca02061),
	.w7(32'h3bc84eee),
	.w8(32'hbc0076fd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7be1c),
	.w1(32'hbb99396d),
	.w2(32'h3b99647e),
	.w3(32'hbc380779),
	.w4(32'h3b15232f),
	.w5(32'hb9771f83),
	.w6(32'hbc35fb44),
	.w7(32'h3c09d0e7),
	.w8(32'h3b78364d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b722b95),
	.w1(32'h3a9e9c1e),
	.w2(32'hbaae3e3a),
	.w3(32'h3b45cbbe),
	.w4(32'hbb6fea86),
	.w5(32'hbbf37dd7),
	.w6(32'hbb9f784b),
	.w7(32'hb9f5fdbf),
	.w8(32'hbc0d27b7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68c72f),
	.w1(32'h3c0d3e68),
	.w2(32'h3c269dae),
	.w3(32'hbbbafbb5),
	.w4(32'h3bc2f0d9),
	.w5(32'h3bb141fe),
	.w6(32'hbbbfabfe),
	.w7(32'h3c077c28),
	.w8(32'hbc1f4a68),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26717d),
	.w1(32'h39dc8d0b),
	.w2(32'h3c737dd2),
	.w3(32'h3b3befbf),
	.w4(32'hbac1de4b),
	.w5(32'h3b740abc),
	.w6(32'hbc2d94cf),
	.w7(32'h3c48f2ab),
	.w8(32'h3bd5b3a7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd41127),
	.w1(32'h3c5e2854),
	.w2(32'h3b889b61),
	.w3(32'h3b50b8a0),
	.w4(32'h3bc63d9c),
	.w5(32'h3ba5d983),
	.w6(32'h3cb39550),
	.w7(32'h3bc60856),
	.w8(32'h3bb97148),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a577),
	.w1(32'hb9db34c3),
	.w2(32'hbc47d519),
	.w3(32'h3c00aa63),
	.w4(32'hbbb53b65),
	.w5(32'hbc185acb),
	.w6(32'h3b889c9f),
	.w7(32'hbc36cf36),
	.w8(32'hbc2f9079),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe169ad),
	.w1(32'hbb7e5186),
	.w2(32'h3bf22be5),
	.w3(32'hbbebebb5),
	.w4(32'hba428e0c),
	.w5(32'hba84a6b9),
	.w6(32'hb8cfda8e),
	.w7(32'h3beb03eb),
	.w8(32'h3aef0d33),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf5e6c),
	.w1(32'h3938176f),
	.w2(32'hbbe959ed),
	.w3(32'hbbfd6003),
	.w4(32'hbc16f534),
	.w5(32'hbb0f8af7),
	.w6(32'h3aa470ae),
	.w7(32'hbbc1b1c7),
	.w8(32'hbbcd07a4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf92b4d),
	.w1(32'h3ae2df84),
	.w2(32'h3aaffbb7),
	.w3(32'h3afa6b5c),
	.w4(32'h3b78e3fc),
	.w5(32'hb9f2d4ff),
	.w6(32'h3c0a7589),
	.w7(32'h3b05a982),
	.w8(32'h3a828b94),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfa947),
	.w1(32'h3b54321c),
	.w2(32'hbb88d979),
	.w3(32'hb9e3fefe),
	.w4(32'hbabaf0e6),
	.w5(32'h3b90bac0),
	.w6(32'hb9b25850),
	.w7(32'hbb9fdb7a),
	.w8(32'h3ba0f667),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c650743),
	.w1(32'h3c8a1834),
	.w2(32'hba96eb7e),
	.w3(32'h3c2bb282),
	.w4(32'h3c453123),
	.w5(32'hbbe13111),
	.w6(32'h3c8db6cf),
	.w7(32'h3bec7500),
	.w8(32'hbc3b0b1a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39357763),
	.w1(32'hbbcb4e6a),
	.w2(32'hb9207bfe),
	.w3(32'hbc4c4431),
	.w4(32'hbbd9afb8),
	.w5(32'hba610711),
	.w6(32'hbc80c010),
	.w7(32'hbbb4e0ab),
	.w8(32'hbbc61635),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82789c),
	.w1(32'hbc4539da),
	.w2(32'h3ae78b76),
	.w3(32'hbbb9fd1c),
	.w4(32'hba4e8438),
	.w5(32'hbc2ded9e),
	.w6(32'hbbf77298),
	.w7(32'h3b84b477),
	.w8(32'hbc7dedfc),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194f48),
	.w1(32'h3ac882e7),
	.w2(32'h3c3937da),
	.w3(32'hbc0d9a16),
	.w4(32'h3be21223),
	.w5(32'h3c4b0be1),
	.w6(32'hbc226ffa),
	.w7(32'h3c3c5cbe),
	.w8(32'h3c85dffc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5de61),
	.w1(32'hbb5dc4bd),
	.w2(32'hbcc207f5),
	.w3(32'h3c3fc1d3),
	.w4(32'hbb26793d),
	.w5(32'h3c51b0ab),
	.w6(32'h3c2f2447),
	.w7(32'hbc9c99a3),
	.w8(32'h3ca55a60),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3b7c9),
	.w1(32'hbbbf4e6d),
	.w2(32'hbccc7b04),
	.w3(32'h3c6e3669),
	.w4(32'hbc0eb799),
	.w5(32'hbb632aa5),
	.w6(32'h3c80de25),
	.w7(32'hbc88354c),
	.w8(32'hbc1ff8a6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac23709),
	.w1(32'h3b0429fc),
	.w2(32'h3b0df419),
	.w3(32'hbbb7fbd2),
	.w4(32'h3b8d2f27),
	.w5(32'hbba1cf67),
	.w6(32'hbb0163e4),
	.w7(32'h3b9cd8d2),
	.w8(32'h3ace71e8),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbdd65),
	.w1(32'h3aa1866e),
	.w2(32'h3b9e3b9a),
	.w3(32'hbb3637f6),
	.w4(32'h3c7c19d5),
	.w5(32'hbc3317d6),
	.w6(32'hbc87e39e),
	.w7(32'h3c0f5b00),
	.w8(32'hbbc82c78),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d764),
	.w1(32'hbaa463ca),
	.w2(32'h3afd729a),
	.w3(32'hbba93ae7),
	.w4(32'h3c101c8a),
	.w5(32'hbb994e9c),
	.w6(32'hbbbc37ef),
	.w7(32'h3b929f78),
	.w8(32'h3911a399),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983a37),
	.w1(32'hbb8cf805),
	.w2(32'hbacae75b),
	.w3(32'hbc390735),
	.w4(32'hbbe9a308),
	.w5(32'h3ad504e4),
	.w6(32'hbbb30010),
	.w7(32'hba84393c),
	.w8(32'hbb5c9279),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e73d),
	.w1(32'hbaf2d1f0),
	.w2(32'h3c862bf2),
	.w3(32'hbb324078),
	.w4(32'h395db1da),
	.w5(32'h3a0757b4),
	.w6(32'h3a6dfd6b),
	.w7(32'h3c6871d6),
	.w8(32'h3b128ff9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880a57d),
	.w1(32'h3af2069e),
	.w2(32'h3aeb3f93),
	.w3(32'hbb37db35),
	.w4(32'hbb28bd4e),
	.w5(32'hbb6f075c),
	.w6(32'hbabad008),
	.w7(32'hba11d578),
	.w8(32'hba7aa747),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d96c),
	.w1(32'h3b1f0029),
	.w2(32'hbbe2ee70),
	.w3(32'hbb4f4a19),
	.w4(32'h3aebe5dd),
	.w5(32'h3b584f72),
	.w6(32'hbbbde7f7),
	.w7(32'hbb948870),
	.w8(32'h3b2eb55a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb56d5c),
	.w1(32'h3a8202e7),
	.w2(32'hbba21f4e),
	.w3(32'hba85e4b9),
	.w4(32'hbb395059),
	.w5(32'hbb5950e6),
	.w6(32'h3acf4e44),
	.w7(32'hbc1b37a3),
	.w8(32'hbb8f211e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf85016),
	.w1(32'hbc4d7ab6),
	.w2(32'h3b42196f),
	.w3(32'hbb2d1359),
	.w4(32'hbb8877d0),
	.w5(32'hbad41125),
	.w6(32'h3a838075),
	.w7(32'h3bfad4db),
	.w8(32'hbc17b0d3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1031f3),
	.w1(32'hbb07358c),
	.w2(32'hba97f15f),
	.w3(32'hbc01da79),
	.w4(32'h3aaa9fbc),
	.w5(32'h3bab8630),
	.w6(32'hbb87624c),
	.w7(32'hbb4a76ec),
	.w8(32'hbc10bc17),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b134ff7),
	.w1(32'h3c002ac1),
	.w2(32'h3b2e8c4c),
	.w3(32'h3b8277e5),
	.w4(32'h3c3cbf95),
	.w5(32'h3bbb81ae),
	.w6(32'hbabe29d2),
	.w7(32'h3b673800),
	.w8(32'h3af276b8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8d604),
	.w1(32'hbb459923),
	.w2(32'hbbfc45c9),
	.w3(32'h3c239662),
	.w4(32'hba5fe18d),
	.w5(32'hbbac201a),
	.w6(32'h3c14c7b4),
	.w7(32'hbba260c2),
	.w8(32'hba01f568),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a0aed),
	.w1(32'hbbc63862),
	.w2(32'hbc21103c),
	.w3(32'hbb783147),
	.w4(32'hbbef8087),
	.w5(32'h3b4a9aec),
	.w6(32'h3c027808),
	.w7(32'hbb19fa90),
	.w8(32'hba95d337),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab38571),
	.w1(32'h3b4ea948),
	.w2(32'hbc114abc),
	.w3(32'h3b52c51b),
	.w4(32'hbb599cac),
	.w5(32'hbc1411c7),
	.w6(32'hbbd641b8),
	.w7(32'hbb46923d),
	.w8(32'hbbb35999),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e0b4c),
	.w1(32'h3b57ca17),
	.w2(32'h3a954165),
	.w3(32'hbb952285),
	.w4(32'h3b563453),
	.w5(32'h3b93c7dd),
	.w6(32'hba7eb863),
	.w7(32'h3b80651b),
	.w8(32'h3b1fdebc),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba707957),
	.w1(32'h3a62ebae),
	.w2(32'hbae428ca),
	.w3(32'hba0f1eb8),
	.w4(32'hbc09d105),
	.w5(32'hbaecc06a),
	.w6(32'h3b3e0598),
	.w7(32'h3ac05af3),
	.w8(32'hbb8ffe26),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0201dd),
	.w1(32'hb8f65ded),
	.w2(32'hbb9764c0),
	.w3(32'hbb69b3c2),
	.w4(32'hbb696c3b),
	.w5(32'hb9a1d1ce),
	.w6(32'hbbc13242),
	.w7(32'hbbb68331),
	.w8(32'h3b16b512),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886099e),
	.w1(32'hbc02f6a5),
	.w2(32'hbc67736d),
	.w3(32'h3c131252),
	.w4(32'hbc140546),
	.w5(32'h3c168c9c),
	.w6(32'h3a69aa80),
	.w7(32'hbc82efef),
	.w8(32'h3c3552fa),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01d85a),
	.w1(32'hbba7b705),
	.w2(32'hbccfbbe4),
	.w3(32'h3c7e956e),
	.w4(32'h3ad502c5),
	.w5(32'h3bf7b092),
	.w6(32'h3ca7631e),
	.w7(32'hbca831db),
	.w8(32'h3c60f3c7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bce0c),
	.w1(32'h3bb034d2),
	.w2(32'h3c5ca10d),
	.w3(32'h39ed6116),
	.w4(32'h3b26b1bd),
	.w5(32'hbb7a1e0d),
	.w6(32'hbb992f88),
	.w7(32'h3c356d65),
	.w8(32'hbc4b7587),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b573266),
	.w1(32'h3b64c7e3),
	.w2(32'h3ba0eae5),
	.w3(32'hba18d388),
	.w4(32'h3b457cfa),
	.w5(32'hbb8bec68),
	.w6(32'hbc1c3684),
	.w7(32'h3ba60e4d),
	.w8(32'hbc4da97d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b88c),
	.w1(32'h3b67c068),
	.w2(32'h3beb398d),
	.w3(32'hbb82c8d1),
	.w4(32'hbb25a58d),
	.w5(32'h3c22a8b0),
	.w6(32'hbbe8bd6a),
	.w7(32'h39c630fa),
	.w8(32'h3bbba90d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82b862),
	.w1(32'hbbf4cb8a),
	.w2(32'hbbdbaa8c),
	.w3(32'hb92a0265),
	.w4(32'hbbaa24fe),
	.w5(32'hb90c3e19),
	.w6(32'h3bb96dbf),
	.w7(32'hbc408bc1),
	.w8(32'h3baedb6f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba527cf),
	.w1(32'hba38e303),
	.w2(32'hbc0c1ae1),
	.w3(32'hb8830c18),
	.w4(32'h3a55683e),
	.w5(32'h3becba44),
	.w6(32'h3c3f6c70),
	.w7(32'hbc2da99d),
	.w8(32'h3bf05208),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20b327),
	.w1(32'hbbca8beb),
	.w2(32'hbbffbeab),
	.w3(32'hba823533),
	.w4(32'hb9b82eaa),
	.w5(32'h3b86ec75),
	.w6(32'hbae8fc98),
	.w7(32'h3b52fc40),
	.w8(32'h3c6d4f2d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fd51a),
	.w1(32'hbbdd7565),
	.w2(32'hbc39d970),
	.w3(32'h3c143761),
	.w4(32'hbbb631cb),
	.w5(32'h3bb59302),
	.w6(32'h3bdb3b01),
	.w7(32'hbc5d9b20),
	.w8(32'h3c34dac7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38437cf8),
	.w1(32'h3b8b9541),
	.w2(32'hbbe3f6ef),
	.w3(32'h3bcc6a31),
	.w4(32'h392fae5e),
	.w5(32'hba7a7508),
	.w6(32'h3bbcc083),
	.w7(32'hba50dc76),
	.w8(32'hbb8a86bf),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b2e58),
	.w1(32'h3b8cf7ae),
	.w2(32'hbad2dc6f),
	.w3(32'hbbb11bbb),
	.w4(32'hbba130bd),
	.w5(32'hbc50e8e6),
	.w6(32'hbb1c8835),
	.w7(32'hbb64f413),
	.w8(32'hbca753a3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc054d73),
	.w1(32'hbb476015),
	.w2(32'h3c54874a),
	.w3(32'hbbf3ffcd),
	.w4(32'h3c1d2c5c),
	.w5(32'h3b21e3a7),
	.w6(32'hbca409e0),
	.w7(32'h3c64cea4),
	.w8(32'h3c640a40),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa43263),
	.w1(32'hbbc47b4d),
	.w2(32'hbc5fe1f9),
	.w3(32'h3a25299c),
	.w4(32'hbc0073ac),
	.w5(32'h3bdfe820),
	.w6(32'hbab92190),
	.w7(32'hbbad3010),
	.w8(32'h3c6b0b98),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e2cc4),
	.w1(32'hbc466758),
	.w2(32'hbcc3df77),
	.w3(32'h3c52a95b),
	.w4(32'hbb6615f5),
	.w5(32'h3c5b611d),
	.w6(32'h3c389819),
	.w7(32'hbc32cad8),
	.w8(32'h3c30f9bb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd43d93),
	.w1(32'hbad9f73b),
	.w2(32'hbc8c9a2a),
	.w3(32'h3bfa49c6),
	.w4(32'hbbfbb4e4),
	.w5(32'hba41f4c4),
	.w6(32'h3bb7d8e7),
	.w7(32'hbc2182b6),
	.w8(32'h3a6c042b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91db91),
	.w1(32'h3a34156d),
	.w2(32'hbbe19e14),
	.w3(32'hbb330b0c),
	.w4(32'hbb83c1b8),
	.w5(32'hbbcf07d7),
	.w6(32'hb9337d64),
	.w7(32'h3b445fbb),
	.w8(32'hbb219559),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0ae5c),
	.w1(32'hbb9c60f8),
	.w2(32'hbb30dd08),
	.w3(32'hbb51d003),
	.w4(32'hba516443),
	.w5(32'hbc606826),
	.w6(32'hbbb523e8),
	.w7(32'h3a65989f),
	.w8(32'hbb880d9b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af135),
	.w1(32'h3b1b81cb),
	.w2(32'h3b68558c),
	.w3(32'h3bdc3076),
	.w4(32'hbb834786),
	.w5(32'hba90bdb2),
	.w6(32'h3cc4bf5a),
	.w7(32'h3a2a3f45),
	.w8(32'hba78ce7e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b454e60),
	.w1(32'h3992a6c0),
	.w2(32'h3989ec34),
	.w3(32'h3b7f5625),
	.w4(32'h3b3edba7),
	.w5(32'h3a99ba3a),
	.w6(32'h3b7dd6d1),
	.w7(32'h3ba629ed),
	.w8(32'h3b32bfa4),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cd58b),
	.w1(32'hbb77b409),
	.w2(32'hbad7eb13),
	.w3(32'h3b7ba0a3),
	.w4(32'hbc3d6b39),
	.w5(32'hba67a3e8),
	.w6(32'h3b875b39),
	.w7(32'hba256194),
	.w8(32'hbc1995d4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad57649),
	.w1(32'h3bc114bd),
	.w2(32'h3c5a086b),
	.w3(32'hbb5330ba),
	.w4(32'hba9a4e00),
	.w5(32'h3b3e57b4),
	.w6(32'h3b7534a0),
	.w7(32'h3bcb5eb0),
	.w8(32'h3b576591),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39aa83),
	.w1(32'h3ab27dec),
	.w2(32'hbc13a091),
	.w3(32'hba0a7a79),
	.w4(32'hbafdf12e),
	.w5(32'h3b792466),
	.w6(32'hbb78d2c0),
	.w7(32'hbbdd3fd3),
	.w8(32'h3c1149aa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aace9bd),
	.w1(32'h3aa2c857),
	.w2(32'hbc43b5bc),
	.w3(32'h3b265389),
	.w4(32'h393aac75),
	.w5(32'hbabdf485),
	.w6(32'h3c02adea),
	.w7(32'hbb90d1ba),
	.w8(32'h3b0ff3f7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8e655),
	.w1(32'hbb2dcb55),
	.w2(32'hbb950fe7),
	.w3(32'h3a8af28f),
	.w4(32'hbc78c0df),
	.w5(32'hbb21e0eb),
	.w6(32'hb938b11e),
	.w7(32'hbc1f85fb),
	.w8(32'h3bcd8767),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e16f9),
	.w1(32'hbc7f0a45),
	.w2(32'hbc3d84cd),
	.w3(32'h3a76ead0),
	.w4(32'hbbff0972),
	.w5(32'hbb8cbead),
	.w6(32'hba8c163a),
	.w7(32'hbc286508),
	.w8(32'hbbd2b08c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38651fa6),
	.w1(32'h3c5d24f1),
	.w2(32'h3c37c157),
	.w3(32'hbc074360),
	.w4(32'h3b92c7f3),
	.w5(32'hbbb61a62),
	.w6(32'hbbd225f4),
	.w7(32'h3c3edf67),
	.w8(32'hbc171b48),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb6c38),
	.w1(32'h3c22e634),
	.w2(32'h3c495443),
	.w3(32'hbbfe389b),
	.w4(32'h3b82b9a2),
	.w5(32'h3b949ed2),
	.w6(32'hbc2eb574),
	.w7(32'h3b4eb12b),
	.w8(32'h3b1c9572),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe52b3),
	.w1(32'hbbb9ce4f),
	.w2(32'hbc82540b),
	.w3(32'h3be0fcee),
	.w4(32'hbbdd5496),
	.w5(32'h3b2f7d16),
	.w6(32'h3c2d4d90),
	.w7(32'hb9c3febc),
	.w8(32'h3b7eefe8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17654b),
	.w1(32'hba81780b),
	.w2(32'h3b2fdf45),
	.w3(32'hb8ca645d),
	.w4(32'hbb8d53bc),
	.w5(32'hbbdf1a8c),
	.w6(32'h3bb0c6ca),
	.w7(32'hbbb165ac),
	.w8(32'hbbe4ac13),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc5fc8),
	.w1(32'h3b6697a7),
	.w2(32'hb9e6382e),
	.w3(32'hbb269dfc),
	.w4(32'hbadc9c8c),
	.w5(32'h3b6a4224),
	.w6(32'h39a0365e),
	.w7(32'hba8c7e07),
	.w8(32'h3c43d339),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f49ab1),
	.w1(32'hbc11b807),
	.w2(32'hbc3d869a),
	.w3(32'hbaedc47f),
	.w4(32'hba8c987c),
	.w5(32'h3c0233e3),
	.w6(32'h3b2569ea),
	.w7(32'hbc00de1d),
	.w8(32'h3bff02f8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954e22a),
	.w1(32'h39110d14),
	.w2(32'h3c328b58),
	.w3(32'hbb1bfa8d),
	.w4(32'hbb6add8e),
	.w5(32'hb8848e14),
	.w6(32'hbc8987bf),
	.w7(32'h3b02db72),
	.w8(32'hb7371646),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b4a3d),
	.w1(32'hba17630b),
	.w2(32'hba27eade),
	.w3(32'hb9d0d167),
	.w4(32'h39153c1a),
	.w5(32'hbabc114f),
	.w6(32'hb953910e),
	.w7(32'h39b18739),
	.w8(32'hba4c7b63),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388cdc04),
	.w1(32'hba54131c),
	.w2(32'hbac135fa),
	.w3(32'h3abda453),
	.w4(32'hb9524550),
	.w5(32'hba06a20b),
	.w6(32'h3a17c2e1),
	.w7(32'hb9dd1b70),
	.w8(32'hba251b1f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28ac21),
	.w1(32'h3828fcd7),
	.w2(32'hba8262aa),
	.w3(32'hbab236ff),
	.w4(32'hba11b34c),
	.w5(32'h39b944ff),
	.w6(32'hba3858fe),
	.w7(32'hb9c350c3),
	.w8(32'hba5e3cb7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba190397),
	.w1(32'hba47a609),
	.w2(32'hbaa83187),
	.w3(32'hb794aa85),
	.w4(32'hb98435b9),
	.w5(32'hb8ad9094),
	.w6(32'hba94bf85),
	.w7(32'hba52c418),
	.w8(32'hb8ca8d36),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d3733),
	.w1(32'hbab4ef45),
	.w2(32'hba274ce1),
	.w3(32'hbb0531e1),
	.w4(32'hb7cedb1e),
	.w5(32'h39ad18cf),
	.w6(32'hbadf3c4b),
	.w7(32'h3815f797),
	.w8(32'hbad81275),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902068b),
	.w1(32'h38af48a5),
	.w2(32'h394eadb8),
	.w3(32'hba4fdf3e),
	.w4(32'hbab5405f),
	.w5(32'hba7bb15f),
	.w6(32'hba92ebff),
	.w7(32'hbab8ba04),
	.w8(32'hbaa48a53),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d8923),
	.w1(32'hbad2c853),
	.w2(32'hba706b05),
	.w3(32'hbaa76f74),
	.w4(32'hba6da684),
	.w5(32'h3881e932),
	.w6(32'hbad6ac9f),
	.w7(32'h39f964ec),
	.w8(32'h39af8ca2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b82989),
	.w1(32'h3867497a),
	.w2(32'hb97d6a50),
	.w3(32'h392f2dd5),
	.w4(32'h3a6275d3),
	.w5(32'hba99ab13),
	.w6(32'h3994dcde),
	.w7(32'hb80195f8),
	.w8(32'hba83e76d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87981e),
	.w1(32'hba3aca88),
	.w2(32'hba824f48),
	.w3(32'hba206ae7),
	.w4(32'h3a4394b1),
	.w5(32'hb998219f),
	.w6(32'hba402085),
	.w7(32'hb9865ed3),
	.w8(32'hb9f35231),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959da6e),
	.w1(32'h3aa59b30),
	.w2(32'hb937f127),
	.w3(32'h39989554),
	.w4(32'hba187df8),
	.w5(32'h3a3b6ea2),
	.w6(32'h3a46cf6d),
	.w7(32'hb9428f6c),
	.w8(32'h3a8b42e7),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73cad0),
	.w1(32'h3901c4e6),
	.w2(32'h39f77000),
	.w3(32'hb94f0ee8),
	.w4(32'h3a8d80c5),
	.w5(32'hba576350),
	.w6(32'h3898bb84),
	.w7(32'h3a3adf5e),
	.w8(32'hba628d9b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19aab0),
	.w1(32'hb9fe5239),
	.w2(32'hba6dc607),
	.w3(32'hbabd0f30),
	.w4(32'hba9db0fe),
	.w5(32'hb9783a59),
	.w6(32'hba2d7e4d),
	.w7(32'hba91e225),
	.w8(32'h371093d6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82269f),
	.w1(32'h39d55cdd),
	.w2(32'h3a8bfe9b),
	.w3(32'h39f0cacf),
	.w4(32'h3aceede0),
	.w5(32'hb90531fd),
	.w6(32'h39bf3a88),
	.w7(32'h3a90d91d),
	.w8(32'h3a42fc76),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4d304),
	.w1(32'h39e35fa5),
	.w2(32'hb95a95a9),
	.w3(32'hba9a27d2),
	.w4(32'hba167ba3),
	.w5(32'h39d48428),
	.w6(32'h39ace5c5),
	.w7(32'h399ae09b),
	.w8(32'h3a9344ba),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7eae6c),
	.w1(32'hba8e5d38),
	.w2(32'h3a721a6e),
	.w3(32'h397bcec2),
	.w4(32'h3b0a3139),
	.w5(32'h39d277cf),
	.w6(32'h3a098ee1),
	.w7(32'h3adb2ee5),
	.w8(32'h3ada736a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac01ce),
	.w1(32'h3a5dbda4),
	.w2(32'hba5db45a),
	.w3(32'h392a7bad),
	.w4(32'h3a142d51),
	.w5(32'hba733410),
	.w6(32'h39202e8f),
	.w7(32'hb9eb9e7d),
	.w8(32'hba9fa730),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd9a9e),
	.w1(32'h39b4a9be),
	.w2(32'h3732da1b),
	.w3(32'hba391a73),
	.w4(32'hba6bb89c),
	.w5(32'h3926431a),
	.w6(32'h3b06821c),
	.w7(32'hba8f2b70),
	.w8(32'h3873eb6a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea64aa),
	.w1(32'hb9218167),
	.w2(32'hb9c012b9),
	.w3(32'hb9af43cb),
	.w4(32'hb9c75025),
	.w5(32'h3a85bdcd),
	.w6(32'hba406468),
	.w7(32'h38ed8b9c),
	.w8(32'h3a810eb1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab553a6),
	.w1(32'h3a07c22f),
	.w2(32'h3a007491),
	.w3(32'h39c16797),
	.w4(32'h3a8ed18a),
	.w5(32'hb735e5a2),
	.w6(32'hb97efe4a),
	.w7(32'h39f23d2f),
	.w8(32'hb98a60eb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b4b8),
	.w1(32'hbb369947),
	.w2(32'hbb46599e),
	.w3(32'hbaaa9d91),
	.w4(32'hbb0af9a5),
	.w5(32'hb9092d6c),
	.w6(32'hbb1e5b09),
	.w7(32'hba0eb321),
	.w8(32'hb9e1c982),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d696c),
	.w1(32'hbab95d6b),
	.w2(32'hbaa3f529),
	.w3(32'hbb373f05),
	.w4(32'hbabb3f99),
	.w5(32'h3a6bf3dd),
	.w6(32'hbb17b7e0),
	.w7(32'hbab00919),
	.w8(32'h3a5012d8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34a1e7),
	.w1(32'h3ab234ec),
	.w2(32'h3a78aef1),
	.w3(32'hba56a593),
	.w4(32'hba76a983),
	.w5(32'hb9ccee18),
	.w6(32'h3a6e2b32),
	.w7(32'hb9578593),
	.w8(32'h3805fc29),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e7910c),
	.w1(32'hb91b1606),
	.w2(32'h39c267ad),
	.w3(32'h3a259f1b),
	.w4(32'hb9e81dfe),
	.w5(32'h3a3cfb4d),
	.w6(32'hb9876a39),
	.w7(32'h3a135bc8),
	.w8(32'h38f9c398),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8397b6),
	.w1(32'hba3596be),
	.w2(32'h39e66c13),
	.w3(32'hba55ee35),
	.w4(32'hba251f49),
	.w5(32'h3aaa6d12),
	.w6(32'h36aefdd0),
	.w7(32'hba01219e),
	.w8(32'hb8eb70b5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff0dae),
	.w1(32'h3a781d05),
	.w2(32'h3a320d1e),
	.w3(32'h3aba180a),
	.w4(32'h3ace387d),
	.w5(32'h3a3d22fa),
	.w6(32'h3a31297d),
	.w7(32'h3a201fea),
	.w8(32'hb892aa8e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39016a27),
	.w1(32'h3ab317e4),
	.w2(32'hb5c0563e),
	.w3(32'h3a0e3203),
	.w4(32'h3a9830af),
	.w5(32'h3a80b3bd),
	.w6(32'h3a8126a7),
	.w7(32'hba0a8162),
	.w8(32'hb95efd74),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d54ca2),
	.w1(32'h38d22a6e),
	.w2(32'h39b437b2),
	.w3(32'h3a628cc8),
	.w4(32'h3a2c7ed5),
	.w5(32'hba293a5a),
	.w6(32'h3a35aa85),
	.w7(32'h39a3db63),
	.w8(32'hba0911ba),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfe520),
	.w1(32'hba6f3962),
	.w2(32'hbb1a0bab),
	.w3(32'hbad1798a),
	.w4(32'h3962e383),
	.w5(32'h395eaf39),
	.w6(32'hbaaed031),
	.w7(32'hbb208aed),
	.w8(32'h3ad6abba),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c6e63),
	.w1(32'h393cce2a),
	.w2(32'h3802419f),
	.w3(32'hb9e1759e),
	.w4(32'hb9b40abe),
	.w5(32'h3a3b4adf),
	.w6(32'hb9888dbb),
	.w7(32'hb9e3ecbb),
	.w8(32'h3a562b06),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38502237),
	.w1(32'hb908ed24),
	.w2(32'hba175cf3),
	.w3(32'hbaf0ef96),
	.w4(32'h3967b39c),
	.w5(32'hb9ef6237),
	.w6(32'h38a63a6d),
	.w7(32'hba894d4d),
	.w8(32'hbb0a6c44),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule