module layer_10_featuremap_297(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a273353),
	.w1(32'h3ac4a93a),
	.w2(32'h3a80c6b7),
	.w3(32'h3a3f2dd5),
	.w4(32'h3a09febb),
	.w5(32'hba0ca63b),
	.w6(32'h3aebe0c1),
	.w7(32'h3ab9f097),
	.w8(32'hba9e33a5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31de96),
	.w1(32'hba93e660),
	.w2(32'h39b54cf3),
	.w3(32'hba34c1c1),
	.w4(32'h3a3af431),
	.w5(32'h3a84da26),
	.w6(32'hbaee4034),
	.w7(32'hb9956018),
	.w8(32'h3abdb5fc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba570e55),
	.w1(32'hba9cfc78),
	.w2(32'hbab3ad7a),
	.w3(32'hb93d3455),
	.w4(32'hb9011f6c),
	.w5(32'h38304048),
	.w6(32'h3a3b7387),
	.w7(32'hb92e5fcb),
	.w8(32'h3a2b4165),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1a71d),
	.w1(32'h3989c072),
	.w2(32'h39122ce1),
	.w3(32'hb9cdbe89),
	.w4(32'h39be16e8),
	.w5(32'hba849ce9),
	.w6(32'h39cba43d),
	.w7(32'h3a20cb78),
	.w8(32'hb92a04b2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90c59b),
	.w1(32'hbb0f8804),
	.w2(32'hbb170d69),
	.w3(32'hba896f07),
	.w4(32'hbaa1cd36),
	.w5(32'hb9b5e4cf),
	.w6(32'hb9b43c6c),
	.w7(32'hba22c9a6),
	.w8(32'hb93ab348),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba035155),
	.w1(32'hb8dd46ee),
	.w2(32'hb9a20c99),
	.w3(32'hb87a28a5),
	.w4(32'hb95b0be6),
	.w5(32'h39ee3675),
	.w6(32'hb816c1bc),
	.w7(32'hb7d4b1d1),
	.w8(32'h379be83f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2f3e6),
	.w1(32'hbaf1a67d),
	.w2(32'hbb786616),
	.w3(32'h391b484d),
	.w4(32'hbb26a45a),
	.w5(32'hbbc61cd8),
	.w6(32'h3a6899d6),
	.w7(32'hba1a488f),
	.w8(32'hbb67c061),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a5efd),
	.w1(32'hbbd625d4),
	.w2(32'hbbc55e30),
	.w3(32'hbba321c8),
	.w4(32'hbbf548c0),
	.w5(32'hba3176a5),
	.w6(32'hbab026a8),
	.w7(32'hbbb0fee2),
	.w8(32'hb829273e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba86a4),
	.w1(32'h3848ae1b),
	.w2(32'hba395435),
	.w3(32'hb9983333),
	.w4(32'hba0a1967),
	.w5(32'hba60b184),
	.w6(32'h3893ce27),
	.w7(32'hb82add75),
	.w8(32'hba11730b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42f1c2),
	.w1(32'hbb19781f),
	.w2(32'hbb9464b7),
	.w3(32'hbb2e5c41),
	.w4(32'hbae69f2e),
	.w5(32'hbb59be4c),
	.w6(32'hba568718),
	.w7(32'hba471511),
	.w8(32'hbaa64b5a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46437b),
	.w1(32'hba6649a6),
	.w2(32'hba430241),
	.w3(32'hba895cad),
	.w4(32'hba8940b7),
	.w5(32'h3a965e6c),
	.w6(32'hba9f6b1b),
	.w7(32'hba37ad58),
	.w8(32'h3a6100df),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b50c7),
	.w1(32'hba921308),
	.w2(32'hbb54e29a),
	.w3(32'h38c2c661),
	.w4(32'hb9c71a33),
	.w5(32'hbb31d084),
	.w6(32'h3b1291f2),
	.w7(32'h3b0150a1),
	.w8(32'hbb2a2f46),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb459668),
	.w1(32'hbb786b27),
	.w2(32'hbbb06c28),
	.w3(32'hba3ab3ac),
	.w4(32'hbaa61ef8),
	.w5(32'hbb8c793b),
	.w6(32'hb98d344b),
	.w7(32'hba86e904),
	.w8(32'hbb96f3a5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb485fa9),
	.w1(32'hbb4c85b5),
	.w2(32'hbb089531),
	.w3(32'hbb2c7d80),
	.w4(32'hbaddb105),
	.w5(32'h39eba774),
	.w6(32'hbad46645),
	.w7(32'hbb141e5e),
	.w8(32'h393209e1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9953e4d),
	.w1(32'hb90e1a6e),
	.w2(32'h39b802a6),
	.w3(32'h394e1bd6),
	.w4(32'h3acbe00c),
	.w5(32'h39a0017f),
	.w6(32'hb9927ec9),
	.w7(32'h3a7b6cf2),
	.w8(32'hb819d542),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e88d8),
	.w1(32'hbac1bdad),
	.w2(32'hbb68d8e3),
	.w3(32'hbaff7adb),
	.w4(32'h3a05a796),
	.w5(32'hba339470),
	.w6(32'hbb255877),
	.w7(32'hba826757),
	.w8(32'h398a295a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803461),
	.w1(32'hba119ccb),
	.w2(32'hb9d2e8a7),
	.w3(32'hba2431c6),
	.w4(32'h38da49b2),
	.w5(32'h3a066978),
	.w6(32'hba998b4d),
	.w7(32'h380c047d),
	.w8(32'h3a0c8261),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3b00a),
	.w1(32'hbbd6d5b0),
	.w2(32'hbbecac44),
	.w3(32'hbb221f0c),
	.w4(32'hbb428ef2),
	.w5(32'hba34592c),
	.w6(32'hbab598ce),
	.w7(32'hbb8917be),
	.w8(32'hba75a3a3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b9b17),
	.w1(32'hbb58c71a),
	.w2(32'hbb3acffe),
	.w3(32'hbab7e848),
	.w4(32'hbabc34e1),
	.w5(32'hba9937f1),
	.w6(32'h3998bd21),
	.w7(32'hbac8761e),
	.w8(32'hbb15d80d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a219e3f),
	.w1(32'hba4d99c9),
	.w2(32'h396cd821),
	.w3(32'h3950cc54),
	.w4(32'h390fcc85),
	.w5(32'hba8c6099),
	.w6(32'hb94dbae1),
	.w7(32'h3a6e0173),
	.w8(32'hba8eb576),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47da35),
	.w1(32'hbae52108),
	.w2(32'hba4067fc),
	.w3(32'hb9e098a2),
	.w4(32'hba6d2770),
	.w5(32'h3a236f9c),
	.w6(32'hbaa6cb8b),
	.w7(32'hba328ac6),
	.w8(32'h3aa78cbb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31ca91),
	.w1(32'h3ad840de),
	.w2(32'h3ae80284),
	.w3(32'h3af373b2),
	.w4(32'h3a8695da),
	.w5(32'hbaad338d),
	.w6(32'h3aea02a4),
	.w7(32'h3abc09f1),
	.w8(32'hbaa273c8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5da86b),
	.w1(32'hbbf6d702),
	.w2(32'hbc015d42),
	.w3(32'hbba3a51c),
	.w4(32'hbb18c800),
	.w5(32'hbb694a65),
	.w6(32'hbbc0ded5),
	.w7(32'hbb92c3a3),
	.w8(32'hbbaaa723),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4408fa),
	.w1(32'hbaee1833),
	.w2(32'hbb4b0f6e),
	.w3(32'hba2efff4),
	.w4(32'hba982ccf),
	.w5(32'hba60aba7),
	.w6(32'hba8e0e86),
	.w7(32'hba885794),
	.w8(32'hba1fd61f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8db66),
	.w1(32'hba3e75f8),
	.w2(32'hba3295df),
	.w3(32'h3b565186),
	.w4(32'h396ad7e3),
	.w5(32'h3a4561bb),
	.w6(32'h3a720baa),
	.w7(32'hbaf92158),
	.w8(32'hba4ef548),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397eefa6),
	.w1(32'h3ac93fbf),
	.w2(32'h3a5c29f7),
	.w3(32'h3a8bf4db),
	.w4(32'h3ac3bfae),
	.w5(32'h3a82f1b5),
	.w6(32'h3a8f6f1a),
	.w7(32'h3aaf6ee9),
	.w8(32'h3a9070de),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d9326),
	.w1(32'h3ac17c33),
	.w2(32'h3ad5f105),
	.w3(32'h3ab86a9c),
	.w4(32'h3addbe62),
	.w5(32'hb8cb8082),
	.w6(32'h3ac6ae89),
	.w7(32'h3af75c11),
	.w8(32'h39b48df7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8efe85),
	.w1(32'hbbc328a1),
	.w2(32'hbc042aed),
	.w3(32'h3c5a62ad),
	.w4(32'hbbf8dcfc),
	.w5(32'hbbf4e3e4),
	.w6(32'h3c79958c),
	.w7(32'hbbc21bea),
	.w8(32'hba1e2dc5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10a934),
	.w1(32'hb93f3eb7),
	.w2(32'h399a68c5),
	.w3(32'h3ad300d3),
	.w4(32'h3a941497),
	.w5(32'hba198b4d),
	.w6(32'h3a579c38),
	.w7(32'h3adfe795),
	.w8(32'h3a6b75ff),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2becf6),
	.w1(32'hba6c78b3),
	.w2(32'hbada51bc),
	.w3(32'h3c038845),
	.w4(32'hba41e323),
	.w5(32'hbb1a9f90),
	.w6(32'h3c0c99d1),
	.w7(32'hba7403eb),
	.w8(32'hba7499b7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812ced8),
	.w1(32'h39fae534),
	.w2(32'h3a850f6e),
	.w3(32'h3a0f2783),
	.w4(32'hb9171436),
	.w5(32'h3a0e758a),
	.w6(32'hba3c7ca2),
	.w7(32'hba0914b4),
	.w8(32'h39c0b927),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0a258),
	.w1(32'hbad2f0e1),
	.w2(32'hb6a50d1a),
	.w3(32'hb993da15),
	.w4(32'h39a48304),
	.w5(32'h3a6c76d4),
	.w6(32'h39d400ef),
	.w7(32'hb9f15d8e),
	.w8(32'h3a703e03),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399151d0),
	.w1(32'h39ddbc55),
	.w2(32'hb9cd7268),
	.w3(32'h399ae83c),
	.w4(32'h3a3405e5),
	.w5(32'hb99fe4a9),
	.w6(32'h3a661a76),
	.w7(32'h3894f822),
	.w8(32'hba2c7a8f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c6ee1),
	.w1(32'hb9a25aa2),
	.w2(32'h3955826f),
	.w3(32'hb95243e5),
	.w4(32'hb9f71f0f),
	.w5(32'hba09b44b),
	.w6(32'hbaa594f4),
	.w7(32'hba84db64),
	.w8(32'hba551f44),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf9319),
	.w1(32'hba6c789e),
	.w2(32'hba9ae1f7),
	.w3(32'hba457e9a),
	.w4(32'hba9afc39),
	.w5(32'hba7be44e),
	.w6(32'h3946c95c),
	.w7(32'hba0a44e8),
	.w8(32'hb9700cea),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf12361),
	.w1(32'hbb452a01),
	.w2(32'hbb32ecfd),
	.w3(32'hba903298),
	.w4(32'hbab84c0f),
	.w5(32'hbb0f39df),
	.w6(32'hbaf8a6f5),
	.w7(32'hbb258e2f),
	.w8(32'hbb05d3cb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f90c7),
	.w1(32'hba6a7f19),
	.w2(32'h38f4c242),
	.w3(32'hbc1c2bbf),
	.w4(32'h3b06c7f3),
	.w5(32'h3b43deff),
	.w6(32'hbc21593c),
	.w7(32'h3b78fd41),
	.w8(32'hb9998bae),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4fd5d),
	.w1(32'hbae08d7f),
	.w2(32'h39b23daa),
	.w3(32'h3be3a370),
	.w4(32'h3a872125),
	.w5(32'hbb266968),
	.w6(32'h3ba60601),
	.w7(32'h3a03209b),
	.w8(32'hbbbdd4fb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e81f3),
	.w1(32'hbb3c6298),
	.w2(32'hbb4de1d4),
	.w3(32'h3c741411),
	.w4(32'hba96ee1c),
	.w5(32'hbc036be5),
	.w6(32'h3c463381),
	.w7(32'hbb6d5504),
	.w8(32'hbc0902e3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a69eb),
	.w1(32'h3b4cbf71),
	.w2(32'h3b10f333),
	.w3(32'h3a02b08f),
	.w4(32'hba6f979f),
	.w5(32'hba8e04d4),
	.w6(32'h3b119600),
	.w7(32'h3a969dce),
	.w8(32'hbaf70975),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1544b),
	.w1(32'hbad26cec),
	.w2(32'hb9e701c2),
	.w3(32'hbb0cdca6),
	.w4(32'hbb0545f7),
	.w5(32'h3a6d6ef8),
	.w6(32'hbaa15500),
	.w7(32'hbacbf354),
	.w8(32'h3ae79003),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0fc55),
	.w1(32'h3b0f7835),
	.w2(32'h3ad5b9e7),
	.w3(32'h3b1fa02d),
	.w4(32'h3ae873dd),
	.w5(32'h3a888356),
	.w6(32'h3b4bc7a7),
	.w7(32'h3afe7a6f),
	.w8(32'h3abd110d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c87df),
	.w1(32'h39fca255),
	.w2(32'h3ae82e40),
	.w3(32'h3a2b0ffe),
	.w4(32'h3a8e968a),
	.w5(32'hb9338a77),
	.w6(32'h3a875e47),
	.w7(32'h3ac34344),
	.w8(32'hba270d2a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3887f2),
	.w1(32'hbbf26967),
	.w2(32'hbc193d0d),
	.w3(32'hbaa89362),
	.w4(32'hbb302958),
	.w5(32'hbb7a5800),
	.w6(32'h39b171bc),
	.w7(32'hbabaa591),
	.w8(32'hbb1b7c7b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51b75a),
	.w1(32'h3abf9292),
	.w2(32'h3b02cf8b),
	.w3(32'h3a22d982),
	.w4(32'h3a0d7c86),
	.w5(32'h3b3cb41e),
	.w6(32'h3ad495a4),
	.w7(32'h39a2f629),
	.w8(32'h3a772780),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1739a),
	.w1(32'h3a147617),
	.w2(32'h3a1b6fc5),
	.w3(32'h3aa67ece),
	.w4(32'h3afd153d),
	.w5(32'h3b0d97b8),
	.w6(32'hbaceceff),
	.w7(32'h3a2cf13b),
	.w8(32'h3a953ad5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39739a7b),
	.w1(32'h3aa18093),
	.w2(32'h39ee8e9d),
	.w3(32'h3abf817d),
	.w4(32'h3b3d4e68),
	.w5(32'h3a353061),
	.w6(32'h3aa15141),
	.w7(32'h3a999612),
	.w8(32'h390120f7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfbc54),
	.w1(32'hbba5751f),
	.w2(32'hbc0ba135),
	.w3(32'hbac48293),
	.w4(32'hba66c791),
	.w5(32'hbb611ac5),
	.w6(32'hba08ee28),
	.w7(32'hbae9779d),
	.w8(32'hbb84f343),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba924e28),
	.w1(32'h374cf1dc),
	.w2(32'h39bd3748),
	.w3(32'hb980bc23),
	.w4(32'h39d9537b),
	.w5(32'h3a8d04e0),
	.w6(32'h398d0955),
	.w7(32'h3a566776),
	.w8(32'h3ac01d5c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b028fcd),
	.w1(32'h3b0c3fee),
	.w2(32'h3a8a65e4),
	.w3(32'h3ab9c558),
	.w4(32'h3a5c8951),
	.w5(32'hbb40d215),
	.w6(32'h3b209901),
	.w7(32'h3a81e735),
	.w8(32'hbb5c48a6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb643b),
	.w1(32'hb98ba775),
	.w2(32'h396e6093),
	.w3(32'hb99fb5eb),
	.w4(32'hb9119efc),
	.w5(32'h3aa50d97),
	.w6(32'hb9e38d9a),
	.w7(32'h3a695524),
	.w8(32'h3a51a901),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901d1b0),
	.w1(32'hbb03924e),
	.w2(32'h3900ca96),
	.w3(32'h3a3951d3),
	.w4(32'h36924237),
	.w5(32'hbaae0988),
	.w6(32'hb812e888),
	.w7(32'hba6b333f),
	.w8(32'hbb15b721),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf387b5),
	.w1(32'hbad8df91),
	.w2(32'hbb05a523),
	.w3(32'hbaa70f4f),
	.w4(32'hbb0cce76),
	.w5(32'h3a57af5b),
	.w6(32'hbae2da16),
	.w7(32'hbb129c39),
	.w8(32'h3a3bc362),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a3776),
	.w1(32'hbba932dd),
	.w2(32'hbbd02fda),
	.w3(32'hba8f4222),
	.w4(32'hbaeeaea3),
	.w5(32'hbb3cfa07),
	.w6(32'h3b83b3ce),
	.w7(32'hb9999e22),
	.w8(32'hbae6d39e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0580f),
	.w1(32'hbad235c6),
	.w2(32'hbac7e507),
	.w3(32'h3abb82ac),
	.w4(32'hba7c4e5f),
	.w5(32'hbae39108),
	.w6(32'h3a7e3724),
	.w7(32'hb98e1be9),
	.w8(32'hbadbe11a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc070e),
	.w1(32'hb91597b1),
	.w2(32'hb9255687),
	.w3(32'hb9eb2666),
	.w4(32'hb8c2818c),
	.w5(32'hb9ed6597),
	.w6(32'h39853bc2),
	.w7(32'h396c9d36),
	.w8(32'hba02b5f0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64b278),
	.w1(32'hba23ef2b),
	.w2(32'hb9e6f3b8),
	.w3(32'hb9e934cd),
	.w4(32'hb8089fcd),
	.w5(32'h3950b404),
	.w6(32'hba2ee772),
	.w7(32'hb9c17666),
	.w8(32'h39c74d30),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad70fae),
	.w1(32'h38c02535),
	.w2(32'hb94eeebe),
	.w3(32'h39ec9ef7),
	.w4(32'hba7ea03f),
	.w5(32'h381c3107),
	.w6(32'h3a4a30df),
	.w7(32'hba677cde),
	.w8(32'h3a19c6de),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfcdf5),
	.w1(32'h3b043ee8),
	.w2(32'h3ae06eaa),
	.w3(32'h3ab51bd1),
	.w4(32'h3a77f51a),
	.w5(32'h3adc977c),
	.w6(32'h3aff3e08),
	.w7(32'h3aa94de6),
	.w8(32'h3b194896),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b442c9c),
	.w1(32'h3ae49403),
	.w2(32'h3aad73d1),
	.w3(32'h3a8b08d3),
	.w4(32'h3ad4be39),
	.w5(32'hba151c6b),
	.w6(32'h3ac0d830),
	.w7(32'h3b2990bc),
	.w8(32'hba01bdb2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbad0b),
	.w1(32'hbb2791cf),
	.w2(32'hbb74288b),
	.w3(32'hba922907),
	.w4(32'hba456743),
	.w5(32'hbadd6638),
	.w6(32'hba5fec7d),
	.w7(32'hba84f00c),
	.w8(32'hbaaa8242),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961f404),
	.w1(32'hbb783cf4),
	.w2(32'hbb5a2a36),
	.w3(32'h3ab961d3),
	.w4(32'hbb358aca),
	.w5(32'hba95ca21),
	.w6(32'h3adeafed),
	.w7(32'hbb481139),
	.w8(32'h3a524195),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba175fe1),
	.w1(32'hbaae774d),
	.w2(32'hbab81d85),
	.w3(32'hba903440),
	.w4(32'hba8038f5),
	.w5(32'hba9ee9d3),
	.w6(32'hb8fa8839),
	.w7(32'hba13e784),
	.w8(32'hba64d73c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5499e6),
	.w1(32'hba19bb71),
	.w2(32'hba3f6103),
	.w3(32'hba889802),
	.w4(32'hba4270f0),
	.w5(32'hba482570),
	.w6(32'hba207153),
	.w7(32'hba8b6052),
	.w8(32'hb901afcc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72a2aa),
	.w1(32'h3a6a56d6),
	.w2(32'h3a3a6e5f),
	.w3(32'h399f86b4),
	.w4(32'h396e9f80),
	.w5(32'hb8e79dc0),
	.w6(32'h39f38c50),
	.w7(32'h39701e3b),
	.w8(32'hba42e041),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c1935),
	.w1(32'hb9ea2a7c),
	.w2(32'hb8ca8654),
	.w3(32'hb9433a1a),
	.w4(32'hb99b12aa),
	.w5(32'hba92fdbb),
	.w6(32'h37bcb013),
	.w7(32'h354ffc93),
	.w8(32'hba6a1a7d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae77596),
	.w1(32'hbb8b2414),
	.w2(32'hbc07b4f4),
	.w3(32'hbaf8155a),
	.w4(32'hbaf0d8e9),
	.w5(32'hbb86b545),
	.w6(32'h3b561186),
	.w7(32'h3b1ce694),
	.w8(32'h3b61860d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910ff2),
	.w1(32'hbb38514c),
	.w2(32'hbb83dafe),
	.w3(32'h3a8f4fa8),
	.w4(32'h3a572226),
	.w5(32'h39df5a84),
	.w6(32'hbbeb2e17),
	.w7(32'hbb2fcb70),
	.w8(32'hbb22b281),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8ca07),
	.w1(32'hba8d7262),
	.w2(32'hbb8b9542),
	.w3(32'h3a90064d),
	.w4(32'h3ab770c1),
	.w5(32'hb9e24513),
	.w6(32'hba8f20d1),
	.w7(32'hbaae142f),
	.w8(32'hbb394842),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc16a52),
	.w1(32'hbaf45d74),
	.w2(32'h3a25fbe0),
	.w3(32'h3be5d1bf),
	.w4(32'h3b02af47),
	.w5(32'h3a9372e2),
	.w6(32'h3aada468),
	.w7(32'hba7170b1),
	.w8(32'hbb4e66df),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4591ae),
	.w1(32'h3a7a3481),
	.w2(32'h3a8b5a89),
	.w3(32'h397dc9a7),
	.w4(32'h3a58599a),
	.w5(32'hbab51933),
	.w6(32'h3a05d357),
	.w7(32'h3a82d1e6),
	.w8(32'hba8379cb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71ec05),
	.w1(32'hbab5aadb),
	.w2(32'hb9ff5115),
	.w3(32'hb9ac2283),
	.w4(32'hbacc8f6e),
	.w5(32'hbaa0298d),
	.w6(32'hba9fb627),
	.w7(32'hbaef9930),
	.w8(32'hba4d5a4f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7f794),
	.w1(32'hbaabadd8),
	.w2(32'hba5bdfd2),
	.w3(32'hb9fe7093),
	.w4(32'hba161e9c),
	.w5(32'h3997c0f2),
	.w6(32'hbac1527b),
	.w7(32'hba8c3be7),
	.w8(32'h3a348e42),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b07c49),
	.w1(32'hba7cbe76),
	.w2(32'hba2eaab0),
	.w3(32'h39f96e34),
	.w4(32'h39ae2abe),
	.w5(32'hbac0c6f8),
	.w6(32'h39999a74),
	.w7(32'h399da19a),
	.w8(32'hbab9c821),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60f782),
	.w1(32'hb99f04b4),
	.w2(32'hba7f229a),
	.w3(32'hba9018d0),
	.w4(32'hba230cf1),
	.w5(32'hba289105),
	.w6(32'hba00d762),
	.w7(32'hb79d4eb0),
	.w8(32'hba24aa23),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e7fef),
	.w1(32'hbb8a6250),
	.w2(32'hbb5356bc),
	.w3(32'hbaea9dcb),
	.w4(32'hba97b842),
	.w5(32'hbb56ce10),
	.w6(32'h39ed4f2d),
	.w7(32'hba46b809),
	.w8(32'hbb151e5e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5de9b),
	.w1(32'hbb8c1861),
	.w2(32'hbbbecfb4),
	.w3(32'hbb893066),
	.w4(32'hbb35f27e),
	.w5(32'hb996c63b),
	.w6(32'hbb02d6d9),
	.w7(32'hbae2d8d7),
	.w8(32'hbb02b473),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84cbb9),
	.w1(32'h3917478b),
	.w2(32'h3b1606e4),
	.w3(32'h3a108aa5),
	.w4(32'h3a189c52),
	.w5(32'h3b096bc0),
	.w6(32'h3afcbe6f),
	.w7(32'h39a67e01),
	.w8(32'h3b46d84c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d28dac),
	.w1(32'h3879c90d),
	.w2(32'hbad7bc7f),
	.w3(32'h3a8b417b),
	.w4(32'h3a8ba13d),
	.w5(32'hb9f2f573),
	.w6(32'h3b11999b),
	.w7(32'h3a9b25c8),
	.w8(32'hbada6f53),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed5671),
	.w1(32'hbafdd260),
	.w2(32'hbb27e204),
	.w3(32'hba134ddd),
	.w4(32'hb93aff0f),
	.w5(32'hbad58372),
	.w6(32'h3a91d31e),
	.w7(32'hb6ff3cf7),
	.w8(32'h3ae24c9d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e5ad6),
	.w1(32'hba92a4b7),
	.w2(32'hbac177a7),
	.w3(32'hba67be91),
	.w4(32'hba8dab88),
	.w5(32'hb7944706),
	.w6(32'hb810e304),
	.w7(32'hb9e9b961),
	.w8(32'hb8cc9539),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a8ed0),
	.w1(32'hbb1502f9),
	.w2(32'hbb1785a2),
	.w3(32'hba82f354),
	.w4(32'hba8634b0),
	.w5(32'hbb3e7a1f),
	.w6(32'hb9f54523),
	.w7(32'hba38b3fb),
	.w8(32'hbb487192),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de4ae),
	.w1(32'h38af427e),
	.w2(32'hbaaa120c),
	.w3(32'hba1e5ca3),
	.w4(32'h374547b8),
	.w5(32'hb90b29c9),
	.w6(32'h3a4e0b9e),
	.w7(32'hb9826a81),
	.w8(32'h3a0e10ec),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a722d),
	.w1(32'h388855e8),
	.w2(32'hba77fe24),
	.w3(32'hba5fa20e),
	.w4(32'hba91f334),
	.w5(32'hba73bf5d),
	.w6(32'hb93133ea),
	.w7(32'hb8d3ee4b),
	.w8(32'hba8ac3e6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba125088),
	.w1(32'h38b9bac9),
	.w2(32'hba58dc2e),
	.w3(32'hba2868ba),
	.w4(32'hb9857cbf),
	.w5(32'hb9e0b636),
	.w6(32'h39fbbdef),
	.w7(32'h3903828b),
	.w8(32'hba3be793),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5cecf),
	.w1(32'hb8f03336),
	.w2(32'h383d8d91),
	.w3(32'h3a83ef32),
	.w4(32'h3a74bd2c),
	.w5(32'hb970ba21),
	.w6(32'h3a5eeab5),
	.w7(32'h3a11297c),
	.w8(32'h39864360),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3770aa4a),
	.w1(32'hb8ee2904),
	.w2(32'h3ad80dee),
	.w3(32'h3882e8c0),
	.w4(32'h3a17afd1),
	.w5(32'h3ab35331),
	.w6(32'hba8049f7),
	.w7(32'h390db5ed),
	.w8(32'hba2bf036),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd5d2e),
	.w1(32'hba586c85),
	.w2(32'hb92353c8),
	.w3(32'h37853f65),
	.w4(32'hb9b01a7d),
	.w5(32'h3a3c9c17),
	.w6(32'h3999789f),
	.w7(32'h3a2e9eb0),
	.w8(32'h39dd6eac),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83fd6a),
	.w1(32'h3913dce0),
	.w2(32'h3ad68f6c),
	.w3(32'h397fc6e6),
	.w4(32'h3a2c130a),
	.w5(32'hb86a9ec2),
	.w6(32'hbaa1d822),
	.w7(32'hb8763d3c),
	.w8(32'hbaad724f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc80004),
	.w1(32'hbb94b5e5),
	.w2(32'hbb81a784),
	.w3(32'hbb74e6a9),
	.w4(32'hbad5e120),
	.w5(32'hba394778),
	.w6(32'hbb89ba1b),
	.w7(32'hbb9470b5),
	.w8(32'hbaf0f7a0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9301),
	.w1(32'hbae70b08),
	.w2(32'hbb182dde),
	.w3(32'h3b945596),
	.w4(32'hbb4dd27d),
	.w5(32'hbb4a5e8b),
	.w6(32'h3b7c9319),
	.w7(32'hbb1dc625),
	.w8(32'hbb2c186c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8967d4),
	.w1(32'h3827e5a0),
	.w2(32'hbb70a7ef),
	.w3(32'hbb2b69d1),
	.w4(32'hb6b08fbf),
	.w5(32'hbb219b3d),
	.w6(32'h3999165f),
	.w7(32'h3b5994ea),
	.w8(32'h3a843387),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ebb6e),
	.w1(32'hba7ae868),
	.w2(32'hbabf01cf),
	.w3(32'h3ac5103b),
	.w4(32'hb8937cd8),
	.w5(32'hbb29c9bb),
	.w6(32'h39d8b52b),
	.w7(32'hbab7cd65),
	.w8(32'hbb7d47b5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60f37b),
	.w1(32'hbb0657eb),
	.w2(32'hbbab9fb4),
	.w3(32'h3a2de572),
	.w4(32'h3ad4544e),
	.w5(32'h3aa68e1e),
	.w6(32'h3a9f783f),
	.w7(32'h372f53cc),
	.w8(32'h3a5b89dc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a802bc3),
	.w1(32'h3a7ad471),
	.w2(32'h3a700756),
	.w3(32'h3b0538fd),
	.w4(32'h3abcca2d),
	.w5(32'h3aeb1efd),
	.w6(32'h3b25306d),
	.w7(32'h3b0ae91b),
	.w8(32'h3b6ffc19),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b969d4b),
	.w1(32'hba94b598),
	.w2(32'hba884a25),
	.w3(32'h3bb0619e),
	.w4(32'h39e469c7),
	.w5(32'hba4ec65b),
	.w6(32'h3bce72f8),
	.w7(32'h3aedf1b6),
	.w8(32'h3b140399),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba050a),
	.w1(32'h3b0ea014),
	.w2(32'h3a361cd8),
	.w3(32'h3a36a943),
	.w4(32'h39e10128),
	.w5(32'hbb08a91d),
	.w6(32'h3af2f6a5),
	.w7(32'h3a967418),
	.w8(32'hbb6a022c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d8296),
	.w1(32'hbb16d6d0),
	.w2(32'hbb99af5a),
	.w3(32'hbb2065db),
	.w4(32'hbb2065b8),
	.w5(32'hbb13fc31),
	.w6(32'hb9af4f20),
	.w7(32'hbb728d76),
	.w8(32'hbb211c06),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9df705),
	.w1(32'hbbebf9fe),
	.w2(32'hbc22aa9a),
	.w3(32'h38fbe523),
	.w4(32'hbbbf4ab9),
	.w5(32'hbb1b635d),
	.w6(32'h3c1526c1),
	.w7(32'hbc002212),
	.w8(32'h3b167cad),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ee123),
	.w1(32'h3c13249d),
	.w2(32'h3b8619bb),
	.w3(32'h3b632e62),
	.w4(32'h3b6dc4c6),
	.w5(32'h3c9cf066),
	.w6(32'hbc1696fd),
	.w7(32'hbbafd77c),
	.w8(32'h3ba8d9c9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f05a2),
	.w1(32'h3b84ec4f),
	.w2(32'h3c9e9632),
	.w3(32'h3b457c90),
	.w4(32'h3c8aa2f1),
	.w5(32'h3b11a605),
	.w6(32'h399706eb),
	.w7(32'hbb074fb4),
	.w8(32'hbb986dd5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8649b6),
	.w1(32'hbb9da004),
	.w2(32'hbb444f93),
	.w3(32'h3c0f6af1),
	.w4(32'hbc0635f6),
	.w5(32'h39a2dc4e),
	.w6(32'h3bcc21c8),
	.w7(32'hbbfe7a70),
	.w8(32'hbaf24330),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad8a4a),
	.w1(32'hb97fc67c),
	.w2(32'hbbc039e9),
	.w3(32'hbbf1776e),
	.w4(32'h3aafb00f),
	.w5(32'hb9e3777e),
	.w6(32'hbb7a4628),
	.w7(32'hbad437dc),
	.w8(32'h3b84e788),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e1ac2),
	.w1(32'h3c35b1e7),
	.w2(32'h374ecc80),
	.w3(32'h3be017fb),
	.w4(32'hba45b864),
	.w5(32'h3b851e44),
	.w6(32'h3b8d385f),
	.w7(32'h3c18a4b6),
	.w8(32'hbbc87352),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf634e5),
	.w1(32'h3ad62192),
	.w2(32'h3c185e80),
	.w3(32'h3c10669d),
	.w4(32'hbb53fef1),
	.w5(32'h3b840f25),
	.w6(32'h3c18d32f),
	.w7(32'hbbae0b76),
	.w8(32'hbaca16d0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcce46),
	.w1(32'hba0f8bf6),
	.w2(32'h3b9bf29d),
	.w3(32'hbb49cf6c),
	.w4(32'hbb220bec),
	.w5(32'hbb79bb6e),
	.w6(32'hbcde9283),
	.w7(32'h3c4586a7),
	.w8(32'hbba14567),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae90bb6),
	.w1(32'h3cd6ddaf),
	.w2(32'hbbe0be97),
	.w3(32'hbaec605f),
	.w4(32'h3bf69ace),
	.w5(32'h3aef3d78),
	.w6(32'h3bbf7ea4),
	.w7(32'h3c93631e),
	.w8(32'hba843589),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d7680),
	.w1(32'h3aebe63a),
	.w2(32'hba39c53d),
	.w3(32'hbade4efe),
	.w4(32'hba1f1ed3),
	.w5(32'hbbc29499),
	.w6(32'h3c37d502),
	.w7(32'hbb62f58f),
	.w8(32'hbbb6437a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed1080),
	.w1(32'hbc0d630c),
	.w2(32'hbc055e8b),
	.w3(32'hbbe91f9d),
	.w4(32'hbbe5816f),
	.w5(32'hbb9f36d1),
	.w6(32'hbc090c06),
	.w7(32'hbbeb3137),
	.w8(32'hbc0d792f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3185eb),
	.w1(32'hbb6ac0c4),
	.w2(32'hba844f55),
	.w3(32'hbac654a5),
	.w4(32'hb9c521f1),
	.w5(32'h3b75add0),
	.w6(32'h38ac4577),
	.w7(32'hbbbd293e),
	.w8(32'hbbe1ad51),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88792),
	.w1(32'hbbadd9b2),
	.w2(32'hbb4b7721),
	.w3(32'h3b3e7232),
	.w4(32'hbc2a8824),
	.w5(32'hbc31f9f8),
	.w6(32'h3c82acc7),
	.w7(32'hbc556156),
	.w8(32'hbb9ef723),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68a92a8),
	.w1(32'h3a8eee2e),
	.w2(32'hbbb3de7c),
	.w3(32'h3b4a90c9),
	.w4(32'h3b0c95db),
	.w5(32'hbc082688),
	.w6(32'h3a89f53e),
	.w7(32'h39b25c77),
	.w8(32'hbc1f9aa6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1eeb),
	.w1(32'hbc36e69d),
	.w2(32'hbc670403),
	.w3(32'hbb81d42e),
	.w4(32'hbc7d1a7d),
	.w5(32'h39df66b4),
	.w6(32'h3b9a88a0),
	.w7(32'hbc93192b),
	.w8(32'h3b03630d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99f904),
	.w1(32'h3bb0048f),
	.w2(32'hbb448c94),
	.w3(32'h3a7ffe3e),
	.w4(32'hbafe8c33),
	.w5(32'h3c1bc02c),
	.w6(32'hbb6da56e),
	.w7(32'h3b9dd475),
	.w8(32'h3c484a1a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695653),
	.w1(32'h3cad538a),
	.w2(32'h3b55a97c),
	.w3(32'hbb1a258f),
	.w4(32'h3bb7eeb2),
	.w5(32'hbb5560ea),
	.w6(32'h3a167d8a),
	.w7(32'hbc14107c),
	.w8(32'h3b4b8c01),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cd3bc),
	.w1(32'h3bd73cc2),
	.w2(32'hbbeb490a),
	.w3(32'hba589214),
	.w4(32'hbb02150f),
	.w5(32'hbb4153fd),
	.w6(32'h3a83add7),
	.w7(32'hbb08dfe0),
	.w8(32'h39a78cbe),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae28108),
	.w1(32'hb96fd434),
	.w2(32'h3b2cf3fa),
	.w3(32'hbac7df1d),
	.w4(32'h3ac7f074),
	.w5(32'h3c0f7adc),
	.w6(32'h3a6f4803),
	.w7(32'h3b101566),
	.w8(32'h3b6a2452),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28495d),
	.w1(32'hbb6ad825),
	.w2(32'h3bb184d3),
	.w3(32'h3ca9fc84),
	.w4(32'h3c0f1e1e),
	.w5(32'hba2f771a),
	.w6(32'h3c5e5ff6),
	.w7(32'h3cb28d0f),
	.w8(32'h3b53b192),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c0fd),
	.w1(32'hb9a571a5),
	.w2(32'hba3e7536),
	.w3(32'h3794b6c1),
	.w4(32'hbad21ed2),
	.w5(32'hbb212cc6),
	.w6(32'h3ab0f139),
	.w7(32'hbc341e45),
	.w8(32'h3b9647dd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcff6a0),
	.w1(32'h3b3b0bfd),
	.w2(32'h37eb4a97),
	.w3(32'hbac08b84),
	.w4(32'h3b07ceeb),
	.w5(32'hbc094c1f),
	.w6(32'hbc99b52b),
	.w7(32'h3c31c4c2),
	.w8(32'hbba01ffc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7086a6),
	.w1(32'h3bfa5d4c),
	.w2(32'h3b3097b6),
	.w3(32'hba1c1efd),
	.w4(32'h3b7d419b),
	.w5(32'hbb2a9b28),
	.w6(32'hbb91055d),
	.w7(32'h3c1adc54),
	.w8(32'hbb9b7a5d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca2e69),
	.w1(32'h3b8aa434),
	.w2(32'hbc01c5a2),
	.w3(32'h3be098a5),
	.w4(32'hbb840c0a),
	.w5(32'hbbaba7a0),
	.w6(32'h3c4137a0),
	.w7(32'hbb9cf630),
	.w8(32'hb9be268e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38ef4c),
	.w1(32'hbbe29c4c),
	.w2(32'hbbb1454f),
	.w3(32'hba9e57b7),
	.w4(32'hbc31e77b),
	.w5(32'hb86854b8),
	.w6(32'h3c5f00db),
	.w7(32'hbbf0d635),
	.w8(32'h3b4d122c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb520ae8),
	.w1(32'hbbbf4971),
	.w2(32'hbbef7387),
	.w3(32'hbb7a0793),
	.w4(32'hbb81c1e4),
	.w5(32'h3bf11952),
	.w6(32'h3bdafaea),
	.w7(32'hbc26d1d0),
	.w8(32'h3b3507ae),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90176f),
	.w1(32'hbb8c7d0d),
	.w2(32'hbbcaf216),
	.w3(32'h3b76d497),
	.w4(32'h3b734f26),
	.w5(32'h3b565fc5),
	.w6(32'h3b17890d),
	.w7(32'hba4e3000),
	.w8(32'h3b9b59c3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad42513),
	.w1(32'h3b359138),
	.w2(32'h3a2a9f33),
	.w3(32'h3bc7d98d),
	.w4(32'hba8b2c65),
	.w5(32'hbb88bcdd),
	.w6(32'h39c51cf0),
	.w7(32'h3b0fe881),
	.w8(32'hbb8452c3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ab1cbe),
	.w1(32'hbb804bbd),
	.w2(32'hbbbaaf19),
	.w3(32'hbacbd16f),
	.w4(32'h3b84f9da),
	.w5(32'h3a7c0298),
	.w6(32'h3c4fd316),
	.w7(32'hbb2b6842),
	.w8(32'h3c4c830a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9bfd9),
	.w1(32'hbabf1b72),
	.w2(32'h3bb1bd1b),
	.w3(32'hba13c28c),
	.w4(32'hbb64875c),
	.w5(32'hbc375fa6),
	.w6(32'hbc7ac588),
	.w7(32'h3b0fea50),
	.w8(32'hbbd27eb1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b9f67),
	.w1(32'hbc519da8),
	.w2(32'hbc419c95),
	.w3(32'hbb95e978),
	.w4(32'hbc42c936),
	.w5(32'hba127fe7),
	.w6(32'h3b1b4b2f),
	.w7(32'hbc7c3d6e),
	.w8(32'h3b43ae45),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba79832),
	.w1(32'h3aea90cd),
	.w2(32'h39dc3ec1),
	.w3(32'h3c695524),
	.w4(32'h3b01854d),
	.w5(32'h3c0ea0d4),
	.w6(32'h3c9bbd57),
	.w7(32'hbb80a056),
	.w8(32'h3bcace0f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf3859),
	.w1(32'h3ca5ce64),
	.w2(32'h3acf234f),
	.w3(32'h3acb3679),
	.w4(32'h3a8ac5bb),
	.w5(32'h3b0d608d),
	.w6(32'h3ac32e00),
	.w7(32'h3bb3919b),
	.w8(32'hbaf3664e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845e26),
	.w1(32'hba572e06),
	.w2(32'hbb314fa8),
	.w3(32'h3af543ca),
	.w4(32'hb93920a1),
	.w5(32'h3b241c96),
	.w6(32'h3c3d4c23),
	.w7(32'hbb99ca90),
	.w8(32'h3c1baf88),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ff8d),
	.w1(32'hbb1714dd),
	.w2(32'hbb882947),
	.w3(32'hbb8f6c40),
	.w4(32'hbb962cd4),
	.w5(32'hb8abba67),
	.w6(32'h3c8bdbed),
	.w7(32'hbbbe38d3),
	.w8(32'hb8584cea),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7654e76),
	.w1(32'hba20c168),
	.w2(32'h3a24b438),
	.w3(32'hba8ada56),
	.w4(32'hba7fca24),
	.w5(32'hbb38a00b),
	.w6(32'h3c20fd42),
	.w7(32'hbb57844f),
	.w8(32'h3b3079e1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe2058),
	.w1(32'h39082d37),
	.w2(32'hbc071c46),
	.w3(32'h3a871b89),
	.w4(32'hb871ca5e),
	.w5(32'hbbe84d54),
	.w6(32'h3c920c5f),
	.w7(32'hbb5a9bbf),
	.w8(32'hbbedb69f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe50791),
	.w1(32'hbb8ba7a1),
	.w2(32'hbae0837b),
	.w3(32'hbb901535),
	.w4(32'hbc130953),
	.w5(32'hbbfd7a64),
	.w6(32'hba6a5a92),
	.w7(32'hbc011d9b),
	.w8(32'hbc0f2c49),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aeafd),
	.w1(32'hbbc4b844),
	.w2(32'hbbeffb69),
	.w3(32'hbc1c253d),
	.w4(32'hbc084cfd),
	.w5(32'hb99447b4),
	.w6(32'hba56738c),
	.w7(32'hbbd4d106),
	.w8(32'h39f0c8d0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a6fe1),
	.w1(32'hbb8ad237),
	.w2(32'hbb58b0a8),
	.w3(32'h39d0d5c2),
	.w4(32'hba636d82),
	.w5(32'h3b787776),
	.w6(32'h3c575b0d),
	.w7(32'hbb7b2f5f),
	.w8(32'h3b511e2b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39076642),
	.w1(32'h3a9d6ef3),
	.w2(32'h3b65ef1b),
	.w3(32'h3a416ffe),
	.w4(32'hbb77c401),
	.w5(32'h3ad36845),
	.w6(32'h3c858b42),
	.w7(32'hbbacaf06),
	.w8(32'h3b9c4059),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ca475),
	.w1(32'h3cad92fd),
	.w2(32'hb6894c16),
	.w3(32'hbc17c3b5),
	.w4(32'h3a02fd8a),
	.w5(32'hbb9fa01a),
	.w6(32'hbb02f40f),
	.w7(32'h3c698873),
	.w8(32'hb8cbf8e7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b219b52),
	.w1(32'h3c2c6247),
	.w2(32'h3b42abdd),
	.w3(32'h3a3b979b),
	.w4(32'hbbaf1cb8),
	.w5(32'hba03e7ed),
	.w6(32'h3c5d5501),
	.w7(32'h3bbfc767),
	.w8(32'hbb832648),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2947c1),
	.w1(32'hbc202189),
	.w2(32'hbb4b2f57),
	.w3(32'h3bde240c),
	.w4(32'hbc187576),
	.w5(32'hbb0f56dd),
	.w6(32'h3badf0ba),
	.w7(32'hbbd0d349),
	.w8(32'hbc00a48f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf90b20),
	.w1(32'h3b51449a),
	.w2(32'h3b9685f1),
	.w3(32'h3a3b8577),
	.w4(32'hbc000f5a),
	.w5(32'hbbbd2353),
	.w6(32'h3c3c8e82),
	.w7(32'hba91aa74),
	.w8(32'hbbea9ff2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d21c2),
	.w1(32'hbbf0eadd),
	.w2(32'hbadf1f43),
	.w3(32'hba4a0c86),
	.w4(32'hbb9daca9),
	.w5(32'hbbd9251a),
	.w6(32'h3c23688b),
	.w7(32'hb94cab02),
	.w8(32'hbb84eb15),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99c066),
	.w1(32'hba5fb6e8),
	.w2(32'h3b5210e7),
	.w3(32'hb71b0f4f),
	.w4(32'hbabb6763),
	.w5(32'hbac9b660),
	.w6(32'h3a582962),
	.w7(32'hbbc89625),
	.w8(32'hbb971603),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a9de7),
	.w1(32'h3a7c3937),
	.w2(32'hbb9d64e1),
	.w3(32'hba47a7cb),
	.w4(32'hbc0c4eef),
	.w5(32'hbb284d0c),
	.w6(32'hbc23aaca),
	.w7(32'h3b3bc12b),
	.w8(32'hbb7ad149),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e0048),
	.w1(32'h3aa53c44),
	.w2(32'hbc100389),
	.w3(32'h3bd4d36d),
	.w4(32'hbb754261),
	.w5(32'hb963d9bf),
	.w6(32'h3c257193),
	.w7(32'h3a8d2878),
	.w8(32'h3a5392fb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb710e94),
	.w1(32'hbb787ded),
	.w2(32'hbb439964),
	.w3(32'h3c18f16f),
	.w4(32'hbb09a5cc),
	.w5(32'h3a96891e),
	.w6(32'h39d39b4b),
	.w7(32'hbb5d7a49),
	.w8(32'hbb746a7f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923b85d),
	.w1(32'hbb2b3349),
	.w2(32'hb910c75f),
	.w3(32'h3b154c61),
	.w4(32'h37eb1227),
	.w5(32'h3b379fbc),
	.w6(32'h3c34eec0),
	.w7(32'h3b0ec9eb),
	.w8(32'h3b046aff),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7be13c),
	.w1(32'hbaf28c8a),
	.w2(32'h3b86e168),
	.w3(32'hbb57f429),
	.w4(32'h3b641332),
	.w5(32'h3b06c3dc),
	.w6(32'hbb4a1a5b),
	.w7(32'h3b3ea424),
	.w8(32'h3b4edbd1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8a1c8),
	.w1(32'h3bf0feb6),
	.w2(32'hbc031e9e),
	.w3(32'h3b3db50b),
	.w4(32'h3b3072e6),
	.w5(32'hbba8e45a),
	.w6(32'h3b81726c),
	.w7(32'h3b593e9c),
	.w8(32'hbb6f3572),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d39e9),
	.w1(32'hbbd47fc9),
	.w2(32'hbac3f1d2),
	.w3(32'hbaf4180d),
	.w4(32'hba347ffb),
	.w5(32'h3bce8918),
	.w6(32'h3c4c7839),
	.w7(32'hbbac1e77),
	.w8(32'h3af897a7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c896333),
	.w1(32'h3b2c5d96),
	.w2(32'hbbe78b5b),
	.w3(32'h3c55b827),
	.w4(32'hbb2caffd),
	.w5(32'hb83ab9d3),
	.w6(32'h3be2c1ea),
	.w7(32'hbc1716e3),
	.w8(32'hbb82c7dc),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2546e9),
	.w1(32'hbaa68fa4),
	.w2(32'h3c20b923),
	.w3(32'hbb4d662c),
	.w4(32'hbb136079),
	.w5(32'h3ba36168),
	.w6(32'h3c5222ef),
	.w7(32'h3b45cfe0),
	.w8(32'hbb4f1967),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad66c10),
	.w1(32'hbb85c5cd),
	.w2(32'h3c0fe9dd),
	.w3(32'hbb058207),
	.w4(32'h3b462f0c),
	.w5(32'hbbb1163d),
	.w6(32'h3a1e2402),
	.w7(32'h3b53bdf8),
	.w8(32'hbc21bf6b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb442f44),
	.w1(32'hbc0311e3),
	.w2(32'hbb88de92),
	.w3(32'hbbf1e1d5),
	.w4(32'hbbb18ad8),
	.w5(32'hba0cef0a),
	.w6(32'hbbcfadaa),
	.w7(32'hbc32e4d7),
	.w8(32'h3b7d65d6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae17404),
	.w1(32'hbb942265),
	.w2(32'hbb8b0e9c),
	.w3(32'h3b6da5f1),
	.w4(32'h3b0e5e65),
	.w5(32'hbbd942b1),
	.w6(32'hbadd1e9b),
	.w7(32'hbbc8c93a),
	.w8(32'hbc614a97),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc606a5),
	.w1(32'hbbfda00c),
	.w2(32'h3b0477ad),
	.w3(32'h3ac12f28),
	.w4(32'h3a11f28d),
	.w5(32'h3c25cc85),
	.w6(32'h3b950642),
	.w7(32'hba36d9b2),
	.w8(32'h3b83937d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23fa72),
	.w1(32'hbbb09b1d),
	.w2(32'hbb351e05),
	.w3(32'h3c578cf5),
	.w4(32'hba469f1f),
	.w5(32'hba489896),
	.w6(32'h3a63d7f7),
	.w7(32'hbaffbcd0),
	.w8(32'h3a8329be),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca6368),
	.w1(32'h3c48aca6),
	.w2(32'h3b503830),
	.w3(32'hb990cad9),
	.w4(32'h3bb7509f),
	.w5(32'h3b0099d7),
	.w6(32'hbc9a3cbf),
	.w7(32'h3b291094),
	.w8(32'h3c843a2d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6d3fb),
	.w1(32'h3bd4b6c5),
	.w2(32'h38837020),
	.w3(32'h3c5fe242),
	.w4(32'h3bc4cdf3),
	.w5(32'h3ac2e78f),
	.w6(32'hbca7da69),
	.w7(32'h3bad1f16),
	.w8(32'h3a019a63),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba732760),
	.w1(32'h3c32389a),
	.w2(32'h3b69f833),
	.w3(32'h3bd0de1f),
	.w4(32'hb88c6fa0),
	.w5(32'hbb4814b3),
	.w6(32'hbc7ae39d),
	.w7(32'h3aac9b56),
	.w8(32'h3b7e5060),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d0fe4),
	.w1(32'h3bc67132),
	.w2(32'h3b8659e1),
	.w3(32'h3bc2f65f),
	.w4(32'hbbef5699),
	.w5(32'h3c96bb8a),
	.w6(32'hbbc421e7),
	.w7(32'hbc12dc2e),
	.w8(32'h3c92e956),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c188439),
	.w1(32'h3c002368),
	.w2(32'hbad9e0b6),
	.w3(32'h39b78776),
	.w4(32'h3b46a439),
	.w5(32'h3c630fd0),
	.w6(32'hbb82dc25),
	.w7(32'h3c2b6c11),
	.w8(32'hbb65728a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50b793),
	.w1(32'hbb74992c),
	.w2(32'hbb89f027),
	.w3(32'h3caa2405),
	.w4(32'h3bb89dba),
	.w5(32'hb9a16929),
	.w6(32'hbc7c07ef),
	.w7(32'h3cbc492a),
	.w8(32'hbbae29d0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6821da),
	.w1(32'hbba8266e),
	.w2(32'hba4cb0fb),
	.w3(32'hbbade32a),
	.w4(32'hbbc436df),
	.w5(32'h3ac22425),
	.w6(32'h3c9633e6),
	.w7(32'hbc0c864d),
	.w8(32'h3bed57f7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b228e68),
	.w1(32'hbbb5a3fb),
	.w2(32'hbb2effed),
	.w3(32'hbc0a31e7),
	.w4(32'hbc25c2f1),
	.w5(32'hbc1ce489),
	.w6(32'h3c1049e4),
	.w7(32'hbbdf498c),
	.w8(32'hbc6c0855),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50ca16),
	.w1(32'hbc28d98b),
	.w2(32'hbbd518a8),
	.w3(32'hbc40b10d),
	.w4(32'hbb9f466d),
	.w5(32'hb99796a2),
	.w6(32'h3a9865c9),
	.w7(32'hbb41b6b7),
	.w8(32'h3c46e85e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba924f0f),
	.w1(32'h39e074fd),
	.w2(32'hbbeea99f),
	.w3(32'hba8031cb),
	.w4(32'hbb849a8f),
	.w5(32'h3b2cd3f7),
	.w6(32'hbc41fdbf),
	.w7(32'h3bcc0f98),
	.w8(32'hbab0f6ee),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e9fa1),
	.w1(32'h3b67c1cb),
	.w2(32'h3c4d6b8e),
	.w3(32'h3999304c),
	.w4(32'h3c273dfb),
	.w5(32'h3a1c0399),
	.w6(32'h3c887ff3),
	.w7(32'h3c12d17d),
	.w8(32'hbc3089cc),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad39d8e),
	.w1(32'hbcb1dca1),
	.w2(32'hbc2bc338),
	.w3(32'hbbf68a80),
	.w4(32'hbc0fd073),
	.w5(32'h3aad0150),
	.w6(32'hbb70193d),
	.w7(32'hbb99cd92),
	.w8(32'h3b9693da),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ef349),
	.w1(32'hbb845d61),
	.w2(32'h3c01bed0),
	.w3(32'h3aa98bf9),
	.w4(32'h3a06fd24),
	.w5(32'hb8e95209),
	.w6(32'h3d097e46),
	.w7(32'hbbbe566c),
	.w8(32'h3ba7eadb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4f55),
	.w1(32'hbb586406),
	.w2(32'hbb03b967),
	.w3(32'h3a08b886),
	.w4(32'h3bb17d1d),
	.w5(32'hbb90c290),
	.w6(32'hbc16f52b),
	.w7(32'hbb337c4e),
	.w8(32'hbbe676db),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42200f),
	.w1(32'h3a94f645),
	.w2(32'h3b06f9eb),
	.w3(32'h3aeb6608),
	.w4(32'h3b77f81e),
	.w5(32'hbc04e9ba),
	.w6(32'h3c055ccb),
	.w7(32'hb9c990ae),
	.w8(32'hbba480d9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc784c9),
	.w1(32'h3b9e09ba),
	.w2(32'h3c01134f),
	.w3(32'hbb442063),
	.w4(32'h3b838cf4),
	.w5(32'hbbb53f1d),
	.w6(32'h38dbc5d3),
	.w7(32'h3c8bd75b),
	.w8(32'h3b8d4a80),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96b7c8),
	.w1(32'hba2a2f76),
	.w2(32'hbab41cd5),
	.w3(32'hbb97ab9c),
	.w4(32'hbb7129cd),
	.w5(32'hbb019224),
	.w6(32'h3c0b8df2),
	.w7(32'hbb823753),
	.w8(32'hbb50a63a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eec60),
	.w1(32'hbb323d2c),
	.w2(32'hbbe27f73),
	.w3(32'hbac92a0d),
	.w4(32'hbbeaf807),
	.w5(32'h3aee29cc),
	.w6(32'h3c17edc3),
	.w7(32'hbb2136f7),
	.w8(32'hb9ad6b4f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fa7d1),
	.w1(32'hbb4b82fd),
	.w2(32'h3bd4ccba),
	.w3(32'hbba1a994),
	.w4(32'h3b265d5c),
	.w5(32'hbc06f905),
	.w6(32'hbbe71f21),
	.w7(32'h385bcd5c),
	.w8(32'h3c1755d3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba266b1),
	.w1(32'h3b6467e8),
	.w2(32'h3ad9e9cc),
	.w3(32'hba2f8c3a),
	.w4(32'hbb1b5e3a),
	.w5(32'hba80e9ca),
	.w6(32'h3bc9dfb0),
	.w7(32'hbc067bf5),
	.w8(32'h3b6de839),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfb5b8),
	.w1(32'h3adc73fb),
	.w2(32'hb98199a8),
	.w3(32'hb9b7a40e),
	.w4(32'h3ba4fa42),
	.w5(32'h3b4e39f6),
	.w6(32'h3bff7250),
	.w7(32'h3b87ef9b),
	.w8(32'hba57a63a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae67430),
	.w1(32'h3ba1ac4e),
	.w2(32'h3b06150b),
	.w3(32'hb9195187),
	.w4(32'h3b27d406),
	.w5(32'hbb35de45),
	.w6(32'h3b80dbec),
	.w7(32'hba4f374e),
	.w8(32'h3b41dce8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b265327),
	.w1(32'h3b80e712),
	.w2(32'h3c95abbb),
	.w3(32'h3c0ca6a6),
	.w4(32'h3ca30976),
	.w5(32'hb9bb65b1),
	.w6(32'hba7fa36f),
	.w7(32'h3d4fd87f),
	.w8(32'h3c032a7b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc45288),
	.w1(32'h39785e85),
	.w2(32'h3a05458f),
	.w3(32'h3b5ba97f),
	.w4(32'hbb556c5c),
	.w5(32'h3b4aa7db),
	.w6(32'hbb04de16),
	.w7(32'hbb194bd5),
	.w8(32'h3bbc4e97),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c59391),
	.w1(32'hbae2fa33),
	.w2(32'h3a16a177),
	.w3(32'h3b5b82d1),
	.w4(32'h3bc4ccba),
	.w5(32'hbb55f8a4),
	.w6(32'hbba7e6ed),
	.w7(32'hbc334416),
	.w8(32'h3aa4dd95),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85b237),
	.w1(32'hbb40b533),
	.w2(32'hbbaa8424),
	.w3(32'hbb28e4af),
	.w4(32'h3ba65149),
	.w5(32'h3a3b348e),
	.w6(32'hbc2ff288),
	.w7(32'h3b8f215f),
	.w8(32'hba357b78),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998e72f),
	.w1(32'hb9819056),
	.w2(32'h3a4e914f),
	.w3(32'h3c8441f0),
	.w4(32'h3a0d376c),
	.w5(32'hbaf33d50),
	.w6(32'h3c98e52f),
	.w7(32'h3c311256),
	.w8(32'hbb35a642),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab36748),
	.w1(32'hbad3a738),
	.w2(32'h3b9e45f3),
	.w3(32'hbafc6f06),
	.w4(32'h396bf153),
	.w5(32'hbb1311c4),
	.w6(32'h3b39fd7f),
	.w7(32'hbaf4f00e),
	.w8(32'hbc72157e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ec943),
	.w1(32'hbc88bdba),
	.w2(32'hbc181aaf),
	.w3(32'hbc847ceb),
	.w4(32'hbbf3194d),
	.w5(32'hbbaba25e),
	.w6(32'hbc2f4495),
	.w7(32'hbc424d07),
	.w8(32'hbbaf04e8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aa7ca),
	.w1(32'hbbe0d390),
	.w2(32'hba84cc52),
	.w3(32'h3aeebb1d),
	.w4(32'hbc1cb50c),
	.w5(32'hbbbf7027),
	.w6(32'h3c775577),
	.w7(32'hbb9b1fa9),
	.w8(32'hbb77406b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47eba1),
	.w1(32'hbc59d044),
	.w2(32'hbc2a07de),
	.w3(32'hbc3b98f2),
	.w4(32'hbc3737e2),
	.w5(32'hb9a23b31),
	.w6(32'h3bfadc92),
	.w7(32'hbb89e354),
	.w8(32'hb9ff615c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab68edd),
	.w1(32'h3aabde93),
	.w2(32'hbb0a2cf0),
	.w3(32'h3a8906aa),
	.w4(32'hbb68032e),
	.w5(32'hbb2dbbb2),
	.w6(32'hbc20353c),
	.w7(32'hbb641846),
	.w8(32'h3c06a10c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6d31e),
	.w1(32'h3b4ec58a),
	.w2(32'hb885c309),
	.w3(32'h3b914401),
	.w4(32'h3b51a723),
	.w5(32'hbb5612e5),
	.w6(32'h3c06854a),
	.w7(32'h3b7945b9),
	.w8(32'hbba78ce5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4c385),
	.w1(32'hbc0f6e97),
	.w2(32'h3b041421),
	.w3(32'h3b09c3ad),
	.w4(32'h398636a2),
	.w5(32'hbb165543),
	.w6(32'hbb729eff),
	.w7(32'hbb858480),
	.w8(32'h3b6efde3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84586e),
	.w1(32'hbbc1e860),
	.w2(32'hbb043496),
	.w3(32'hbb8dd8b4),
	.w4(32'hbb4e464f),
	.w5(32'hba43a13f),
	.w6(32'hbb3dc2a0),
	.w7(32'h3a9d3d8b),
	.w8(32'hbb90bd45),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8334a5),
	.w1(32'h3ab30848),
	.w2(32'hbbc1ea63),
	.w3(32'hbb616ef1),
	.w4(32'hbc2a01bb),
	.w5(32'hba76a7cc),
	.w6(32'h3be8eac1),
	.w7(32'hbbe458a2),
	.w8(32'hbb590122),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c57db),
	.w1(32'hbb44784b),
	.w2(32'h3b266397),
	.w3(32'hbb0ece28),
	.w4(32'hbb61c77f),
	.w5(32'hba0983bc),
	.w6(32'h3c7cdace),
	.w7(32'hbbea29a4),
	.w8(32'h3c4f3feb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d0c27),
	.w1(32'h3b04367d),
	.w2(32'h3c1d8954),
	.w3(32'hbb4edb06),
	.w4(32'h3a825437),
	.w5(32'h3b8e4495),
	.w6(32'hbbecb96e),
	.w7(32'hba8ffbf1),
	.w8(32'hbb32a05c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3798fa45),
	.w1(32'h3b822486),
	.w2(32'h3bd60b13),
	.w3(32'h3b5527b1),
	.w4(32'h3baf5577),
	.w5(32'h3c2ca139),
	.w6(32'h3b247afb),
	.w7(32'h3c4debcb),
	.w8(32'hbb2bbe7f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0445de),
	.w1(32'h3b1ec140),
	.w2(32'h39f6aa15),
	.w3(32'h3c0eeb25),
	.w4(32'h3b8cb96a),
	.w5(32'hbb084775),
	.w6(32'h3a51988d),
	.w7(32'h3b1c532a),
	.w8(32'hbbb067dc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67285e),
	.w1(32'h3c3deba3),
	.w2(32'h3b83cc55),
	.w3(32'h3b2cae7e),
	.w4(32'hbb03204a),
	.w5(32'hbb8b5153),
	.w6(32'h3ca81e27),
	.w7(32'hbb402eb0),
	.w8(32'h3b641e1c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6e165),
	.w1(32'hbb9c3feb),
	.w2(32'hbc2d7bc7),
	.w3(32'hbc4ceeb4),
	.w4(32'hbbc881f9),
	.w5(32'hbb69c3cc),
	.w6(32'h3c11bd60),
	.w7(32'hbbf93efd),
	.w8(32'hbb2f0fc9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191388),
	.w1(32'h3b5d05f7),
	.w2(32'h3bf26e14),
	.w3(32'h3c4bd4b8),
	.w4(32'hbb85b88b),
	.w5(32'hbb0abead),
	.w6(32'hbafbc3fc),
	.w7(32'h3bb28eac),
	.w8(32'hba5ded5d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac930ad),
	.w1(32'h3aa904ae),
	.w2(32'hbb941bcb),
	.w3(32'hb9b1f439),
	.w4(32'hbbf3fe20),
	.w5(32'hbb3abd88),
	.w6(32'h3c45b0b0),
	.w7(32'hbc17c47f),
	.w8(32'h376de9e4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da1f2),
	.w1(32'h3a92bd44),
	.w2(32'hbbe6c471),
	.w3(32'hb9cf6fc3),
	.w4(32'hbbc13411),
	.w5(32'h3b9253d4),
	.w6(32'h3b1f59df),
	.w7(32'h3a6a8c80),
	.w8(32'hba16c2b4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e944c),
	.w1(32'h3a9334ed),
	.w2(32'hbb0e013c),
	.w3(32'hb9d368f4),
	.w4(32'hbab90ca5),
	.w5(32'hbb7a1e3a),
	.w6(32'hb93a6043),
	.w7(32'hbbb27133),
	.w8(32'h3a63aaaa),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e4978),
	.w1(32'h3ba66ab9),
	.w2(32'hbb90a1fe),
	.w3(32'h3be9a9c2),
	.w4(32'hbb58a19e),
	.w5(32'hbb6c3bc2),
	.w6(32'hbb9e39da),
	.w7(32'hb7c5d239),
	.w8(32'h3afa90fd),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca2fdc),
	.w1(32'h3c2eae73),
	.w2(32'hbc641809),
	.w3(32'h3c0bea9d),
	.w4(32'hbc1fa0b4),
	.w5(32'hbbb5a2cc),
	.w6(32'h3cf264b6),
	.w7(32'hbc2dd274),
	.w8(32'hbbf8d205),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8a79f),
	.w1(32'hbbd23120),
	.w2(32'hbba5ef5d),
	.w3(32'hbbf5d699),
	.w4(32'hbc200fd3),
	.w5(32'hbc1cacfd),
	.w6(32'h3b9f20e0),
	.w7(32'hbc1f83f3),
	.w8(32'hbc116ad0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc819331),
	.w1(32'hbc320679),
	.w2(32'hbc1ab17e),
	.w3(32'hbc5b85e5),
	.w4(32'hbc03295f),
	.w5(32'hba89e432),
	.w6(32'h3b800b6f),
	.w7(32'hbc854ed6),
	.w8(32'hbb872bd8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ae964),
	.w1(32'h3b28512c),
	.w2(32'hbb6553e8),
	.w3(32'hbb2fa238),
	.w4(32'hba9801cf),
	.w5(32'hbab8e034),
	.w6(32'hbbfae087),
	.w7(32'h3bb0e6bd),
	.w8(32'hbb3c86fd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3108cc),
	.w1(32'hbb88ea7d),
	.w2(32'h3b9533a1),
	.w3(32'hbc06a86c),
	.w4(32'h389bdb2b),
	.w5(32'h3b1430ce),
	.w6(32'hbbabd3c2),
	.w7(32'hba852cb4),
	.w8(32'hbab6a4c6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95de528),
	.w1(32'h3b528cdb),
	.w2(32'hbae43143),
	.w3(32'h3b4e337e),
	.w4(32'h3ab2ae11),
	.w5(32'h3b2f3eb2),
	.w6(32'h3cbf152c),
	.w7(32'hbb81c445),
	.w8(32'h3b138364),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa3c23),
	.w1(32'hbab831b3),
	.w2(32'hbb4075b6),
	.w3(32'h3b8460d9),
	.w4(32'h3b889abe),
	.w5(32'hbb7d3f06),
	.w6(32'hbc2da4f6),
	.w7(32'hb8d60566),
	.w8(32'hbbc949e1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a70ef3),
	.w1(32'hbc0abb6e),
	.w2(32'hbc11e831),
	.w3(32'hbc1cf057),
	.w4(32'hbbac1cf1),
	.w5(32'h3970688c),
	.w6(32'h3c5ab9f5),
	.w7(32'hbc5aeb1a),
	.w8(32'hba9db929),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade0877),
	.w1(32'h3c6b3c64),
	.w2(32'h3b06fdd2),
	.w3(32'hbae44021),
	.w4(32'h3bc09880),
	.w5(32'hbaf8e5ed),
	.w6(32'h3c32962b),
	.w7(32'h3cf31c81),
	.w8(32'h3b8c7010),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f3039),
	.w1(32'h395fa6f0),
	.w2(32'hba18fb0c),
	.w3(32'h3b72951b),
	.w4(32'hbb29ce03),
	.w5(32'hbbda6c6d),
	.w6(32'hbbf75095),
	.w7(32'hbbaf7ecc),
	.w8(32'hbbe33eaf),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1cc53),
	.w1(32'hbbb4b438),
	.w2(32'hbb2ef3a9),
	.w3(32'hbb940248),
	.w4(32'hbb923400),
	.w5(32'h3beb561c),
	.w6(32'h3b4c06ff),
	.w7(32'hbbb927b3),
	.w8(32'h399fb4a0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4468a5),
	.w1(32'hbbcd2b95),
	.w2(32'hb9a62299),
	.w3(32'hbbb45060),
	.w4(32'hbb3d93e2),
	.w5(32'hbb4d32f1),
	.w6(32'h3b903714),
	.w7(32'h396a399e),
	.w8(32'h3a695f38),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5ab55),
	.w1(32'hbae03a4e),
	.w2(32'hbc1e810c),
	.w3(32'h3bfd5478),
	.w4(32'hbb025d7e),
	.w5(32'hbbcfa272),
	.w6(32'h3c4de6b1),
	.w7(32'hbad7f4f8),
	.w8(32'h3be89afe),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3908a),
	.w1(32'hba93eeda),
	.w2(32'h3b55830f),
	.w3(32'hbb9a91a6),
	.w4(32'hbb904120),
	.w5(32'hbb5443a8),
	.w6(32'hbbeef7d5),
	.w7(32'h3a4b175f),
	.w8(32'h3c48ea79),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38e3f2),
	.w1(32'h3c76c1ec),
	.w2(32'h3ba13584),
	.w3(32'h3c0e65a5),
	.w4(32'h3adbe8fb),
	.w5(32'hba750766),
	.w6(32'hbc55f751),
	.w7(32'hbb4a4136),
	.w8(32'h3b039fba),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd1cba),
	.w1(32'hbc25c3e9),
	.w2(32'hbba1fee2),
	.w3(32'hbb5162dc),
	.w4(32'hba1ff780),
	.w5(32'h3b77b400),
	.w6(32'hbb771423),
	.w7(32'hbc128f67),
	.w8(32'hb98a86aa),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b956122),
	.w1(32'hbabe64ef),
	.w2(32'hbb365724),
	.w3(32'h3a6604de),
	.w4(32'hbb83831c),
	.w5(32'h3a80d17e),
	.w6(32'h3c4d0a23),
	.w7(32'hbbcf436d),
	.w8(32'h3b927819),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11bd4a),
	.w1(32'h3b3b208b),
	.w2(32'h3b8f448b),
	.w3(32'hba6e863a),
	.w4(32'hbc074921),
	.w5(32'hbba75cbf),
	.w6(32'h3c6549cc),
	.w7(32'h3b20423c),
	.w8(32'hb927f13a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e3004),
	.w1(32'h3ae2a2aa),
	.w2(32'hbc58c1c2),
	.w3(32'hbaefd7d9),
	.w4(32'hbbc92af8),
	.w5(32'h3ae3229c),
	.w6(32'h3cab482e),
	.w7(32'hbc0636fc),
	.w8(32'h3ca2de47),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c1471),
	.w1(32'h3bceea0a),
	.w2(32'h3c2d9c81),
	.w3(32'h3be5c0a4),
	.w4(32'h3b2efe28),
	.w5(32'hbbf71ca5),
	.w6(32'hbc83e3c0),
	.w7(32'h3b3a7821),
	.w8(32'h398c8920),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7da20),
	.w1(32'h3c0fe69c),
	.w2(32'h3c565ae6),
	.w3(32'h3ac338bb),
	.w4(32'h3c3dbd54),
	.w5(32'hbabc07cb),
	.w6(32'h3c03fb8b),
	.w7(32'h3c7c7371),
	.w8(32'hbb221e09),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ff760),
	.w1(32'hbcb8c124),
	.w2(32'hbadb496e),
	.w3(32'h3bb5a0e1),
	.w4(32'hbc7e1a56),
	.w5(32'hbcbb4813),
	.w6(32'hbc95f84e),
	.w7(32'hbc399c8f),
	.w8(32'hbc4f8dfc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01dcf1),
	.w1(32'h3b812b63),
	.w2(32'h3b4294e7),
	.w3(32'hbb73496f),
	.w4(32'h3bf47080),
	.w5(32'h3c115875),
	.w6(32'h3beceb4f),
	.w7(32'h3c14c5b4),
	.w8(32'hbb9b775c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedad05),
	.w1(32'hbac6c15d),
	.w2(32'h3b92f954),
	.w3(32'h3b92b941),
	.w4(32'h3b442d88),
	.w5(32'hbaf5192e),
	.w6(32'hbc491fb3),
	.w7(32'hbb64e103),
	.w8(32'hbb18a665),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9862),
	.w1(32'hb9a46eff),
	.w2(32'hba96f245),
	.w3(32'hbc0b2505),
	.w4(32'h3a14a1de),
	.w5(32'h3c1b8ced),
	.w6(32'hbc2cfa64),
	.w7(32'h3b221656),
	.w8(32'h3c35e34d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbedd1),
	.w1(32'hbc838900),
	.w2(32'hbc9250ae),
	.w3(32'h3b8fb05d),
	.w4(32'hbb97b6a8),
	.w5(32'hbc03f41a),
	.w6(32'hbb9a6991),
	.w7(32'hbc8ca7fa),
	.w8(32'hbc8166ad),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62a630),
	.w1(32'h3b0576c7),
	.w2(32'hbc0d3279),
	.w3(32'hbc218dca),
	.w4(32'hbb1a1017),
	.w5(32'h3c3877ae),
	.w6(32'hbc350623),
	.w7(32'hbc620515),
	.w8(32'h3c275bd9),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc494ff8),
	.w1(32'hbcc10a61),
	.w2(32'hbce5917a),
	.w3(32'h3c45dd3a),
	.w4(32'hbc59ed8f),
	.w5(32'hbcab3725),
	.w6(32'hbaf3ef74),
	.w7(32'hbc8bfcd6),
	.w8(32'hbc9047b3),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cd0f3),
	.w1(32'hbcdfbe65),
	.w2(32'hbc0f61e6),
	.w3(32'hbc97ced6),
	.w4(32'hbb56ca7e),
	.w5(32'hbb8b5fe4),
	.w6(32'hbce00b06),
	.w7(32'hbc8c7d18),
	.w8(32'hbbe11414),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f8c89),
	.w1(32'hbc2dcd62),
	.w2(32'h3ae4cced),
	.w3(32'hbb79bb5d),
	.w4(32'hb85afd07),
	.w5(32'hbcb8321a),
	.w6(32'hba63b4a9),
	.w7(32'h3c105a03),
	.w8(32'hbc7854df),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae75e46),
	.w1(32'h3c1748d0),
	.w2(32'h3c5c12db),
	.w3(32'hbc2d0567),
	.w4(32'h3baddc8a),
	.w5(32'hbc4a0aca),
	.w6(32'h3a8cc365),
	.w7(32'h3c52f71e),
	.w8(32'hbc02864e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0dabc),
	.w1(32'h3af1dffa),
	.w2(32'h3baa79e8),
	.w3(32'hbc19bd5b),
	.w4(32'hbb8a1058),
	.w5(32'h3b0e0f3e),
	.w6(32'hbb393586),
	.w7(32'h3bbb1167),
	.w8(32'hbacbdcaa),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92b0e7),
	.w1(32'hba8676a4),
	.w2(32'hbb6879f0),
	.w3(32'hb9e66a22),
	.w4(32'hbc2943d3),
	.w5(32'hb9596cee),
	.w6(32'hbb86ade8),
	.w7(32'hbbc992ce),
	.w8(32'hbba17175),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0da62),
	.w1(32'hbb3984d6),
	.w2(32'h3bc6a4d9),
	.w3(32'hbbb79811),
	.w4(32'h3b1e482c),
	.w5(32'h3c18878a),
	.w6(32'hbbcfee1c),
	.w7(32'h3bde738e),
	.w8(32'h3c3fd1b2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cf4f0),
	.w1(32'h3c2d392a),
	.w2(32'hba9c5ba7),
	.w3(32'h3c06fd2c),
	.w4(32'h3c0dc664),
	.w5(32'hba9c28ce),
	.w6(32'h3c5ea30d),
	.w7(32'h3c11d326),
	.w8(32'h3b159793),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cea80),
	.w1(32'hbbdf685a),
	.w2(32'hbb5cfe32),
	.w3(32'hbb8609fd),
	.w4(32'hbb7e7066),
	.w5(32'h3b703e8e),
	.w6(32'hbab74041),
	.w7(32'hbb72b91f),
	.w8(32'h3c74336f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca2ed1),
	.w1(32'hbc9d1981),
	.w2(32'hbc68c288),
	.w3(32'hbbc4a819),
	.w4(32'hbb587a51),
	.w5(32'h3c0bacc3),
	.w6(32'hbb094e78),
	.w7(32'hbbc28018),
	.w8(32'h387bffdc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba477c02),
	.w1(32'hbaf8cb9d),
	.w2(32'h3bf18394),
	.w3(32'hbb2f5262),
	.w4(32'h3b7d869d),
	.w5(32'hbcac2ce2),
	.w6(32'hbc2838d0),
	.w7(32'h3b1833af),
	.w8(32'hbc606b65),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae554c7),
	.w1(32'h3c5ff79e),
	.w2(32'h3c98d7d2),
	.w3(32'hbc57a777),
	.w4(32'h3bb9a935),
	.w5(32'h3bf8f31a),
	.w6(32'h3b6ac88f),
	.w7(32'h3c984570),
	.w8(32'hbc16ea70),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50217c),
	.w1(32'hb9423fe8),
	.w2(32'hbc09c751),
	.w3(32'h3c9742d0),
	.w4(32'h3bad07f4),
	.w5(32'hbba741b4),
	.w6(32'hbb5ed6a0),
	.w7(32'hbc41d7a9),
	.w8(32'hbb5ebbc1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eca410),
	.w1(32'hbbbcc5bf),
	.w2(32'h3b1bb171),
	.w3(32'hbc144f47),
	.w4(32'h3a1d794f),
	.w5(32'hbaaf100f),
	.w6(32'hbc0923d0),
	.w7(32'h3b65fd34),
	.w8(32'h3b03574b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61be78),
	.w1(32'hbb9dc3c1),
	.w2(32'hbb254f13),
	.w3(32'h3c7421e5),
	.w4(32'h3c2737e2),
	.w5(32'h3b6adc53),
	.w6(32'h3c0efa7d),
	.w7(32'hbb07cf09),
	.w8(32'h3985063b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1a0db),
	.w1(32'hbba2ef41),
	.w2(32'hbbc2b3ad),
	.w3(32'h3bad7b7d),
	.w4(32'h3b11f65b),
	.w5(32'h3c157f81),
	.w6(32'hbb24a714),
	.w7(32'hbbf7deb8),
	.w8(32'h3c18594e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd45799),
	.w1(32'h3b29ec11),
	.w2(32'hba33bb22),
	.w3(32'h3c087962),
	.w4(32'hbb0e6cf0),
	.w5(32'h3cc62396),
	.w6(32'h3c046bad),
	.w7(32'hbb18687a),
	.w8(32'h3c8e85dd),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3862c),
	.w1(32'hbbde9d3e),
	.w2(32'hbbba596b),
	.w3(32'h3c497ff9),
	.w4(32'hba67bba5),
	.w5(32'h3bd71939),
	.w6(32'h3c24341b),
	.w7(32'hbbad6692),
	.w8(32'hba2374af),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5fda4),
	.w1(32'hba9b939c),
	.w2(32'hbc2e4433),
	.w3(32'h3bb31081),
	.w4(32'hbb3820ad),
	.w5(32'h3c7d66b5),
	.w6(32'h3aa6f11b),
	.w7(32'h39407d54),
	.w8(32'h3c848ce6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e41d0),
	.w1(32'h396b9b4d),
	.w2(32'hbb76ebbb),
	.w3(32'h3b6b9a8d),
	.w4(32'hbc2ec686),
	.w5(32'hba04ff94),
	.w6(32'h3b05733b),
	.w7(32'hbc0a76ff),
	.w8(32'h3a4d0631),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c73747),
	.w1(32'hbb03ae4e),
	.w2(32'h3a14fc8c),
	.w3(32'hbbe813ed),
	.w4(32'hba9f2d01),
	.w5(32'hbca135e1),
	.w6(32'h3b8a5c95),
	.w7(32'h3986e756),
	.w8(32'hbb991d98),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba742f2),
	.w1(32'h3b78cf3c),
	.w2(32'h3bb3e8d0),
	.w3(32'hbac14a6b),
	.w4(32'h3c1905c5),
	.w5(32'hba946ade),
	.w6(32'h3c5c3966),
	.w7(32'h3c82111f),
	.w8(32'hb9c398b5),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c89d3),
	.w1(32'hbbd6f69d),
	.w2(32'hbae07456),
	.w3(32'hbc4a60b4),
	.w4(32'hbbb87a2b),
	.w5(32'hb9053afa),
	.w6(32'hbc044ba4),
	.w7(32'hbaf795bf),
	.w8(32'h3c080e43),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule