module layer_10_featuremap_231(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ac251),
	.w1(32'h3ba093a6),
	.w2(32'h3b68a42f),
	.w3(32'hb8455829),
	.w4(32'h3b18303c),
	.w5(32'h3d2795fa),
	.w6(32'hba5cb5a4),
	.w7(32'h3ad3ac63),
	.w8(32'h39b083de),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa77c3f),
	.w1(32'h3c199f04),
	.w2(32'hb9cf14fe),
	.w3(32'hbc08162c),
	.w4(32'h3c89ed96),
	.w5(32'hba8ed4bc),
	.w6(32'hbbdc5fd0),
	.w7(32'h3c20de8c),
	.w8(32'h3c0ad110),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9e0ca),
	.w1(32'hb9e84332),
	.w2(32'hbcbcc168),
	.w3(32'h3b131c7c),
	.w4(32'h3c74e005),
	.w5(32'h3a3756d4),
	.w6(32'hbb56cac3),
	.w7(32'h3b0a5c70),
	.w8(32'h3b50a5f4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae7c46),
	.w1(32'hbbb6b790),
	.w2(32'h3accc0d0),
	.w3(32'hbbacdc2f),
	.w4(32'h3afd89ea),
	.w5(32'hbc27e4fe),
	.w6(32'hbc22bcb3),
	.w7(32'h3a965d01),
	.w8(32'hbc0d5e5b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37b8aa),
	.w1(32'h3a60350d),
	.w2(32'hbb3da571),
	.w3(32'hbb638dbc),
	.w4(32'hbb93e8fb),
	.w5(32'h3b771f5d),
	.w6(32'hbc375ab3),
	.w7(32'hbc514964),
	.w8(32'hbb50349c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10f787),
	.w1(32'h3b6402ef),
	.w2(32'hbb93e91a),
	.w3(32'h397834eb),
	.w4(32'h39e4ac1a),
	.w5(32'h3c80c318),
	.w6(32'h3b90f15c),
	.w7(32'hbc1a540d),
	.w8(32'hbc233644),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76bdf2),
	.w1(32'hbc217d6c),
	.w2(32'hbc6a81cc),
	.w3(32'hbbf62617),
	.w4(32'h3be1586d),
	.w5(32'h3bedafe6),
	.w6(32'hbb025206),
	.w7(32'h3c28ec8f),
	.w8(32'hbacc4e6f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb747810),
	.w1(32'h3c63ef92),
	.w2(32'hbc43a7ea),
	.w3(32'hbbd5a7af),
	.w4(32'h3c0ed58a),
	.w5(32'h3a89d3d6),
	.w6(32'hbbb4dca2),
	.w7(32'h392205e2),
	.w8(32'h3bff9bb2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4888bf),
	.w1(32'hb9baf1c0),
	.w2(32'h3a373ba5),
	.w3(32'h3b24c1ab),
	.w4(32'h3b1c38a2),
	.w5(32'hbb877325),
	.w6(32'hb9207b5e),
	.w7(32'h3bae1f4f),
	.w8(32'hbaad4eb7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92b04a),
	.w1(32'hba28d5b5),
	.w2(32'hbc87cc69),
	.w3(32'hbc1a6325),
	.w4(32'h3b549fe1),
	.w5(32'h3ad25e50),
	.w6(32'h3b6d449a),
	.w7(32'hbac2d092),
	.w8(32'hbafaee0b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3eaead),
	.w1(32'h3b053152),
	.w2(32'hbc179727),
	.w3(32'h3c869d81),
	.w4(32'hbc52a101),
	.w5(32'h3ba7b267),
	.w6(32'hbbc96a97),
	.w7(32'hbba2f901),
	.w8(32'hbbcfab19),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba22e71),
	.w1(32'hbbfc5192),
	.w2(32'hbb53a589),
	.w3(32'h3b690134),
	.w4(32'h3c169331),
	.w5(32'hba67e286),
	.w6(32'h3b2b63e8),
	.w7(32'h3929cb78),
	.w8(32'h3cc1f7af),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97a5e5),
	.w1(32'hbb8c1a04),
	.w2(32'h3a8caf02),
	.w3(32'h3b5c67ad),
	.w4(32'hbb96e1bb),
	.w5(32'h3c079061),
	.w6(32'h3b82f52e),
	.w7(32'h39c24917),
	.w8(32'hbb59ba63),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf02455),
	.w1(32'h3b85038a),
	.w2(32'hbc05615a),
	.w3(32'h3a85db3e),
	.w4(32'h3b892bdc),
	.w5(32'h3b85d0ea),
	.w6(32'hbb609405),
	.w7(32'h3bbb594c),
	.w8(32'h3b88c420),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10372d),
	.w1(32'hbb9348e8),
	.w2(32'hbbcb3211),
	.w3(32'hbbcbe1b7),
	.w4(32'hbc071e26),
	.w5(32'h3c179ab0),
	.w6(32'hbc5174ab),
	.w7(32'h3c194c01),
	.w8(32'h3b113dd8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bbbfd),
	.w1(32'hbbd640ed),
	.w2(32'hbc6dc67e),
	.w3(32'h3b714f01),
	.w4(32'hbaa8368b),
	.w5(32'hba6c994d),
	.w6(32'h3b0260ec),
	.w7(32'hbb2844ba),
	.w8(32'h3b7c9ad5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06ea8c),
	.w1(32'h3a8e3170),
	.w2(32'hbb01fe9a),
	.w3(32'hbb2acbf3),
	.w4(32'hb7e7d2bd),
	.w5(32'hba0b2a1f),
	.w6(32'h3a58df17),
	.w7(32'h3a6690f2),
	.w8(32'hba69dcf6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb928190),
	.w1(32'hb858da7a),
	.w2(32'h3aff67ef),
	.w3(32'hbba56e1c),
	.w4(32'hbae75148),
	.w5(32'h3a4a8f54),
	.w6(32'h3c170977),
	.w7(32'h3b6f4a21),
	.w8(32'hbb97449e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a88bb),
	.w1(32'h3a0a66a1),
	.w2(32'hba74f946),
	.w3(32'hbc18f939),
	.w4(32'hbc294a10),
	.w5(32'hbb6d9ba5),
	.w6(32'hba1b8f2c),
	.w7(32'h3c50218b),
	.w8(32'h3ab1ca72),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82df536),
	.w1(32'hb892468b),
	.w2(32'h3c0d9c54),
	.w3(32'hbc136147),
	.w4(32'hba98f7d4),
	.w5(32'hbbf9a246),
	.w6(32'hbb7c7fd4),
	.w7(32'hbba2de92),
	.w8(32'hbc1fd9ea),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19f0e7),
	.w1(32'hba6d3072),
	.w2(32'hb9c45a57),
	.w3(32'hbb09c0e1),
	.w4(32'hbbdc188b),
	.w5(32'hbc5d9d02),
	.w6(32'hbba576d4),
	.w7(32'h3aeee979),
	.w8(32'h3a9acd5d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd37e7),
	.w1(32'h3a8923ab),
	.w2(32'hbb24fbbc),
	.w3(32'hbaa3edb5),
	.w4(32'h3b3af0b0),
	.w5(32'hbab31b8c),
	.w6(32'hb9a37724),
	.w7(32'h392f77cf),
	.w8(32'hbc22b186),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a1322),
	.w1(32'hba5d3984),
	.w2(32'h3b111e74),
	.w3(32'hbb88b3ed),
	.w4(32'hbb3ae234),
	.w5(32'h3c5af39d),
	.w6(32'h3ace09f9),
	.w7(32'hbc06556b),
	.w8(32'hbaff0659),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba568014),
	.w1(32'h3bb27815),
	.w2(32'h3bd50441),
	.w3(32'hbb9784d7),
	.w4(32'hbbae1c88),
	.w5(32'hbc2eff03),
	.w6(32'hbc0eb8b2),
	.w7(32'h3a5205aa),
	.w8(32'hbaf5b7ec),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf784d7),
	.w1(32'hb96938fe),
	.w2(32'hbb1ae141),
	.w3(32'h3c64fb4a),
	.w4(32'hbc001b12),
	.w5(32'h3b188fc7),
	.w6(32'hbc3b1c52),
	.w7(32'h3c16d196),
	.w8(32'h3c0f44d3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f2d46),
	.w1(32'h3ab69045),
	.w2(32'h3c87eb02),
	.w3(32'hb939ff71),
	.w4(32'h3cd1e03d),
	.w5(32'h3b723dd6),
	.w6(32'h3acc9d95),
	.w7(32'h3b87fee2),
	.w8(32'hbbbabac8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caaf6b3),
	.w1(32'hbbd9e02b),
	.w2(32'hb8542812),
	.w3(32'h3ba4f2bb),
	.w4(32'h39a76672),
	.w5(32'h3b003094),
	.w6(32'h3c1519ac),
	.w7(32'h3c1d0ae6),
	.w8(32'hbadd557d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49b41d),
	.w1(32'hbc7e60bd),
	.w2(32'h3bb21883),
	.w3(32'hbb689f93),
	.w4(32'h3c3b8ff8),
	.w5(32'hbc148ca8),
	.w6(32'hbbb07bfc),
	.w7(32'h3c441060),
	.w8(32'h3ca5b051),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81ba14),
	.w1(32'h3c11a42b),
	.w2(32'hba7db097),
	.w3(32'h3a96cf47),
	.w4(32'h3b0f48f4),
	.w5(32'h3bbf3854),
	.w6(32'hbb0ed117),
	.w7(32'hbc1a0411),
	.w8(32'hbcc738cb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c887413),
	.w1(32'hbb8335a4),
	.w2(32'hbceb89a3),
	.w3(32'hbcf1249d),
	.w4(32'h3bc2800c),
	.w5(32'hbc8dc7b4),
	.w6(32'h3cc8d41f),
	.w7(32'h3b4eca9e),
	.w8(32'hbd4984c6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19d7ff),
	.w1(32'hbc27a52b),
	.w2(32'h3c1829df),
	.w3(32'hb93d2d37),
	.w4(32'hbb5757bb),
	.w5(32'hbac1e061),
	.w6(32'hbb4cb3ca),
	.w7(32'h3c579ce0),
	.w8(32'h3ce4261f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9981c5),
	.w1(32'hbd1e0796),
	.w2(32'hbba0deec),
	.w3(32'hbcb3a43e),
	.w4(32'hbc07c7c9),
	.w5(32'h3c46b417),
	.w6(32'h3abd41fb),
	.w7(32'h3c1d7fe4),
	.w8(32'h3b1c6412),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b7b7),
	.w1(32'h3d31fda5),
	.w2(32'h3ce5b599),
	.w3(32'hbc5ffd2a),
	.w4(32'hba7b24dc),
	.w5(32'hbd3f4f1c),
	.w6(32'hbcdf8b8a),
	.w7(32'hbd04f1e8),
	.w8(32'hbae5549f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86004e),
	.w1(32'h39a85d20),
	.w2(32'hb8eae832),
	.w3(32'h3bc6ad2a),
	.w4(32'h3c10bd4d),
	.w5(32'hba1884b9),
	.w6(32'h3bc55b1e),
	.w7(32'hbc7166fe),
	.w8(32'hbb28e0ce),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdb339),
	.w1(32'hbc38d8c7),
	.w2(32'hbcce2703),
	.w3(32'hbc2843db),
	.w4(32'hbae87f17),
	.w5(32'h3d0b9fcb),
	.w6(32'h3aa8e9f1),
	.w7(32'h3b45fc0b),
	.w8(32'h3bc9be8c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d577b),
	.w1(32'h3bb729a2),
	.w2(32'hbcf8f096),
	.w3(32'hbcc609ad),
	.w4(32'h3c639526),
	.w5(32'hbc2706b4),
	.w6(32'h3ba44056),
	.w7(32'hbc5a2b35),
	.w8(32'hbcf14e07),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89dbe3),
	.w1(32'hbc45f1f1),
	.w2(32'hbcc1914f),
	.w3(32'h3b772380),
	.w4(32'h3a28fa92),
	.w5(32'h3c0019c0),
	.w6(32'h3b78ae82),
	.w7(32'hba8fba03),
	.w8(32'h3bd19bed),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16340e),
	.w1(32'h3b257ea4),
	.w2(32'hbd0e47bf),
	.w3(32'h3bd1048d),
	.w4(32'h3b8762a1),
	.w5(32'hba3d731a),
	.w6(32'h3bbe3918),
	.w7(32'h3ca51981),
	.w8(32'hbd3fadcb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a0744),
	.w1(32'hbcaddbba),
	.w2(32'h3b809145),
	.w3(32'hbbd29094),
	.w4(32'hbc51bfee),
	.w5(32'hbc339356),
	.w6(32'hba8a1963),
	.w7(32'hbc1c1061),
	.w8(32'hbbaf4d7e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd07f13),
	.w1(32'hbba918e2),
	.w2(32'h3b95bbae),
	.w3(32'hbbc9480d),
	.w4(32'hbb374e1f),
	.w5(32'hbc0c6bbe),
	.w6(32'h3c1e175a),
	.w7(32'h3c9fd702),
	.w8(32'h3bd99c59),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3620acde),
	.w1(32'h3b68166b),
	.w2(32'h3c47c64b),
	.w3(32'h3bea3377),
	.w4(32'h3b8e3dab),
	.w5(32'hbc42c5a0),
	.w6(32'h3beaf0d0),
	.w7(32'h3c00f031),
	.w8(32'hbc259d41),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31af18),
	.w1(32'h3ac31c52),
	.w2(32'h3c67375b),
	.w3(32'hbbdf382d),
	.w4(32'h3b23baa4),
	.w5(32'hbbca2bd9),
	.w6(32'h3c262cee),
	.w7(32'h3c51f572),
	.w8(32'h3bc75f45),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978c61),
	.w1(32'h3c9edfdc),
	.w2(32'h3b62642a),
	.w3(32'hbc1abdb3),
	.w4(32'h3c0e5b3e),
	.w5(32'hbc67a667),
	.w6(32'hbcbf9543),
	.w7(32'hbc863902),
	.w8(32'hbbb3325b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d9fdc),
	.w1(32'h3962f8bd),
	.w2(32'hbca60255),
	.w3(32'hbb9b5f4b),
	.w4(32'hbca73082),
	.w5(32'hbc2c0872),
	.w6(32'h3c5e7553),
	.w7(32'h3c1ae308),
	.w8(32'hba18fa91),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc853f62),
	.w1(32'hba934daa),
	.w2(32'hbc2a205e),
	.w3(32'hbb90043b),
	.w4(32'hbc345b6e),
	.w5(32'hbaab6096),
	.w6(32'hbbd76c6a),
	.w7(32'h3cc05370),
	.w8(32'hb903643f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c96a0),
	.w1(32'h3c88ada1),
	.w2(32'hba204eb0),
	.w3(32'hbb9d700d),
	.w4(32'hbc162171),
	.w5(32'h3b9911c2),
	.w6(32'hbadacbd4),
	.w7(32'hbb9cba66),
	.w8(32'hbc4ecfc1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd3a7b),
	.w1(32'hb9e91050),
	.w2(32'hbd322f27),
	.w3(32'h3c73ec72),
	.w4(32'h3c8e2e96),
	.w5(32'hbb329330),
	.w6(32'h3aa618f4),
	.w7(32'hbc7a68fa),
	.w8(32'hbb87a915),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd957ffa),
	.w1(32'hbc5dece8),
	.w2(32'h3ca83919),
	.w3(32'hbcc89397),
	.w4(32'h3ba45005),
	.w5(32'h3c074070),
	.w6(32'h3c89e19d),
	.w7(32'hbc17df4b),
	.w8(32'hbbc06aa0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76bea0),
	.w1(32'hbc944157),
	.w2(32'hbbb1741f),
	.w3(32'h3bd4c9b5),
	.w4(32'hbb4bfbcb),
	.w5(32'hbbf45327),
	.w6(32'hbb1560f5),
	.w7(32'hbcc4ad7e),
	.w8(32'hb821744c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ce6b2),
	.w1(32'h3b799ec1),
	.w2(32'hbbcda75a),
	.w3(32'h3c5c9b52),
	.w4(32'hba46358b),
	.w5(32'h3b3645c9),
	.w6(32'hbbb1014b),
	.w7(32'h3a1306fc),
	.w8(32'h3bf0e9bf),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fff7ee),
	.w1(32'hb91200f7),
	.w2(32'h3c10ef22),
	.w3(32'hbba8455b),
	.w4(32'hbc114558),
	.w5(32'h3a078d4a),
	.w6(32'hbc22bd85),
	.w7(32'h3bb2c645),
	.w8(32'hbb2848e6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36d151),
	.w1(32'h3ba46393),
	.w2(32'hbc97e32d),
	.w3(32'hba758e23),
	.w4(32'hbc8bb69c),
	.w5(32'hbbe807c6),
	.w6(32'h3cade760),
	.w7(32'hbc2a7fad),
	.w8(32'hbc09f0f3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba2eb2),
	.w1(32'hbbddaf6f),
	.w2(32'hbc890a21),
	.w3(32'hbd229355),
	.w4(32'hbc26fd97),
	.w5(32'hbbcc6721),
	.w6(32'hbb85bcce),
	.w7(32'hbc092357),
	.w8(32'h398e5f02),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad423b),
	.w1(32'hbcbd9c16),
	.w2(32'h3bd49127),
	.w3(32'h3c96658c),
	.w4(32'h3b5a36c2),
	.w5(32'h3b37eedc),
	.w6(32'hbcecbb4f),
	.w7(32'hbaa8c041),
	.w8(32'h3c72d059),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696e6a),
	.w1(32'hbc68dbf3),
	.w2(32'hbc85597c),
	.w3(32'h3c77a8b4),
	.w4(32'hbb61ace2),
	.w5(32'h3b53a1c9),
	.w6(32'hbbd9322b),
	.w7(32'hb7f1420a),
	.w8(32'hbb077bdf),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76348b),
	.w1(32'h3a7e3452),
	.w2(32'h3af7a972),
	.w3(32'hbb74a73c),
	.w4(32'hbb8ed098),
	.w5(32'h3b3e6f98),
	.w6(32'hbaba4b5e),
	.w7(32'h3a816f8c),
	.w8(32'hbc1503e0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a245f0f),
	.w1(32'h3bcdc051),
	.w2(32'hbab5aeba),
	.w3(32'h3c1b6dda),
	.w4(32'h3a5535b4),
	.w5(32'h3c584d39),
	.w6(32'h3ba6af39),
	.w7(32'h3ac09c9e),
	.w8(32'h3b155063),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab79d08),
	.w1(32'hbae26c27),
	.w2(32'h3c13de6e),
	.w3(32'hbb14256a),
	.w4(32'h3ca435ba),
	.w5(32'hbb895b63),
	.w6(32'h3ab8929f),
	.w7(32'hbb16eccd),
	.w8(32'h3b0d342b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd33a5),
	.w1(32'h3b3781f4),
	.w2(32'h3abb2512),
	.w3(32'hbbaf4573),
	.w4(32'h3aa85bc6),
	.w5(32'h3aaa7e0c),
	.w6(32'h3bdae5bd),
	.w7(32'hbb7bfc68),
	.w8(32'h3cb6fddf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7733b8),
	.w1(32'hba57bba8),
	.w2(32'hbaa2dfc8),
	.w3(32'hbbff0490),
	.w4(32'h3b967d4a),
	.w5(32'h3b086e86),
	.w6(32'h3954243a),
	.w7(32'h3ba445c7),
	.w8(32'hbba39921),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8bbd3),
	.w1(32'h3c755697),
	.w2(32'hbb87ed99),
	.w3(32'hbb0ce169),
	.w4(32'hba9e4b4b),
	.w5(32'h3c7e6eb5),
	.w6(32'hbc733a71),
	.w7(32'hbb9d98a0),
	.w8(32'hbbc7710e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb472a51),
	.w1(32'hbb8a80e7),
	.w2(32'hb9da3e15),
	.w3(32'h3a7f8161),
	.w4(32'hbab8b9d8),
	.w5(32'hbc1340c7),
	.w6(32'hbb036d60),
	.w7(32'hbaf9a854),
	.w8(32'h3b473812),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f17d7),
	.w1(32'h37dc418d),
	.w2(32'h3c3f6b32),
	.w3(32'h3bb5b8a7),
	.w4(32'h3b132ba1),
	.w5(32'h38b46b94),
	.w6(32'h3bbd4ba2),
	.w7(32'hbb61ca48),
	.w8(32'hbb19dbea),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb894691),
	.w1(32'hbbb71fcd),
	.w2(32'hbb98b76a),
	.w3(32'hbab63582),
	.w4(32'h3bf38f68),
	.w5(32'h3aa3a2cc),
	.w6(32'hbc4c366f),
	.w7(32'h3b084f61),
	.w8(32'h3acc4a28),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb388d4d),
	.w1(32'h3a100331),
	.w2(32'hbb5bfecd),
	.w3(32'hbbd9cf18),
	.w4(32'hbb35f449),
	.w5(32'hbc00fe1b),
	.w6(32'h3c4b0575),
	.w7(32'h3b30ca1f),
	.w8(32'hbaa72e94),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49fcd6),
	.w1(32'hbc3f3cd5),
	.w2(32'hba8c85f9),
	.w3(32'hbb624817),
	.w4(32'hbb7e8d40),
	.w5(32'hba52d497),
	.w6(32'hbb18384c),
	.w7(32'h3c014ade),
	.w8(32'h3c1631dd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc137ab7),
	.w1(32'hbc6147c7),
	.w2(32'hba824f5f),
	.w3(32'hbb52ee42),
	.w4(32'h3b444c30),
	.w5(32'h3bbbf423),
	.w6(32'h3aef9e08),
	.w7(32'hbb964d28),
	.w8(32'hbb6c0942),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd8d67),
	.w1(32'hbb419fe9),
	.w2(32'h3a6e6336),
	.w3(32'h3b52e51b),
	.w4(32'hb9dcafbb),
	.w5(32'hbb88dab4),
	.w6(32'h3988f4a7),
	.w7(32'hbb8d445f),
	.w8(32'hba2787fd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2399),
	.w1(32'hbbec1a2e),
	.w2(32'h3ad6cbc7),
	.w3(32'hbb532312),
	.w4(32'h3991b7f7),
	.w5(32'hbac38a1a),
	.w6(32'hbbdb36c0),
	.w7(32'h3bc66097),
	.w8(32'hbb6ae966),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2745c),
	.w1(32'hba8e8cd4),
	.w2(32'h3b8a8278),
	.w3(32'h38f229d0),
	.w4(32'hba942385),
	.w5(32'hbb405a7d),
	.w6(32'h3aaaacc7),
	.w7(32'hbae378a8),
	.w8(32'h3b80e8a1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad503a1),
	.w1(32'hbb2908f6),
	.w2(32'h3b50f812),
	.w3(32'h3b64bccf),
	.w4(32'h3b7dfc50),
	.w5(32'hbba8bd83),
	.w6(32'h39255c32),
	.w7(32'hbb51cfe1),
	.w8(32'h3b3cbd1d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab22576),
	.w1(32'hbb0c71e6),
	.w2(32'h3baf781c),
	.w3(32'hbbeb6273),
	.w4(32'hba4c3278),
	.w5(32'hbab40f53),
	.w6(32'h39a9495e),
	.w7(32'h39297fa9),
	.w8(32'hba47f358),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceb4e1),
	.w1(32'hba14ec47),
	.w2(32'hba5266d1),
	.w3(32'hbba6fa6c),
	.w4(32'h3c7a5ec8),
	.w5(32'hbba151d1),
	.w6(32'h3a8bd8a0),
	.w7(32'h3b8bd080),
	.w8(32'h3a788f53),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918966f),
	.w1(32'hb84ddf11),
	.w2(32'h3a942e27),
	.w3(32'h3a8438b7),
	.w4(32'h3b73d3b8),
	.w5(32'h3b354c45),
	.w6(32'hbb255dff),
	.w7(32'h3b0d35f5),
	.w8(32'h3b38c04f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b447bf2),
	.w1(32'h3aa0dc8e),
	.w2(32'h38a175ab),
	.w3(32'hbc23089f),
	.w4(32'hbbfac97b),
	.w5(32'h3bb28de8),
	.w6(32'h3bc44d4d),
	.w7(32'hba18159c),
	.w8(32'h3b0a1084),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a4dcf),
	.w1(32'hbb92ce0b),
	.w2(32'hbbe03a92),
	.w3(32'h3baa1d3e),
	.w4(32'h3bc18399),
	.w5(32'h3b88e4ef),
	.w6(32'hbb9207e2),
	.w7(32'h39fa511a),
	.w8(32'hbb0baa7d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbb7f0),
	.w1(32'hba15d637),
	.w2(32'hbb57d3d8),
	.w3(32'hbb98aca1),
	.w4(32'hba1a7e58),
	.w5(32'h3ab93e55),
	.w6(32'h3c48d047),
	.w7(32'h3c28fe70),
	.w8(32'hba08b04b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb4676),
	.w1(32'h3a82d5b3),
	.w2(32'hbafc0168),
	.w3(32'hbb812b16),
	.w4(32'h3bc7622b),
	.w5(32'h3b80c3fd),
	.w6(32'h3b86e7b1),
	.w7(32'h3b4605df),
	.w8(32'hbbdf6ef6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e07d4),
	.w1(32'hba6ee9b9),
	.w2(32'hb8f56f61),
	.w3(32'h3b347761),
	.w4(32'h38bca6af),
	.w5(32'h3b19f6e3),
	.w6(32'h3c965eeb),
	.w7(32'hbb991ab5),
	.w8(32'hbb88f894),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c4fab),
	.w1(32'hbac27ce5),
	.w2(32'h3b06278c),
	.w3(32'h3a0e9b27),
	.w4(32'h3c1b5cbf),
	.w5(32'h3b453957),
	.w6(32'h39fea942),
	.w7(32'h3be6fcbd),
	.w8(32'h3b79f960),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcddccf),
	.w1(32'hbc175aa2),
	.w2(32'hbbda9b7d),
	.w3(32'h3951c6f5),
	.w4(32'h391739ac),
	.w5(32'hbaca792a),
	.w6(32'hbb61c330),
	.w7(32'h3c5b1870),
	.w8(32'h3b0da6e0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44c169),
	.w1(32'hbc5d45d1),
	.w2(32'h3bdb9d17),
	.w3(32'hbb05e1d7),
	.w4(32'hb9c8aadf),
	.w5(32'h3c5011b9),
	.w6(32'h3bf2c13e),
	.w7(32'h3b0907ef),
	.w8(32'hbbce00e2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf28b4d),
	.w1(32'h3c6c9784),
	.w2(32'h3a7b551b),
	.w3(32'h3b39e749),
	.w4(32'h3b88e87e),
	.w5(32'h3af98613),
	.w6(32'hbbd92533),
	.w7(32'hbb60fa17),
	.w8(32'h3c87b379),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb192d9c),
	.w1(32'hbb76f7de),
	.w2(32'hbb4e6354),
	.w3(32'hba875d5d),
	.w4(32'h3ad21f9d),
	.w5(32'hbae7733a),
	.w6(32'hbbc7dd15),
	.w7(32'h3c76bc87),
	.w8(32'h3c912d8b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d05e2),
	.w1(32'h3bbf6033),
	.w2(32'hbb5480f2),
	.w3(32'h391d4193),
	.w4(32'h3b48b17f),
	.w5(32'h3c5f19b0),
	.w6(32'h3a38879f),
	.w7(32'h3b82bab5),
	.w8(32'h3b57003f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4d1ec),
	.w1(32'h3b932660),
	.w2(32'h3c0a6ee0),
	.w3(32'hbb68b63b),
	.w4(32'h3b6a6e4d),
	.w5(32'h3a9d0e6b),
	.w6(32'h3c94f90d),
	.w7(32'hbb8ab50c),
	.w8(32'hba3e8b65),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80cc5a),
	.w1(32'h3ae78ee8),
	.w2(32'h3c9a1aa1),
	.w3(32'h3bfeb893),
	.w4(32'h3b8efa6f),
	.w5(32'h3c136973),
	.w6(32'h3b849ac9),
	.w7(32'hbbb2a01f),
	.w8(32'h3c2167cc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2ce15),
	.w1(32'hba50ba04),
	.w2(32'h3b9d01f4),
	.w3(32'h3bf3ddce),
	.w4(32'h3af6f5ae),
	.w5(32'hbc18e9b2),
	.w6(32'h3c029bbb),
	.w7(32'h3b58c580),
	.w8(32'hbbd28845),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bd8a6),
	.w1(32'hbb8fcf58),
	.w2(32'hbbb938a1),
	.w3(32'h3a98080f),
	.w4(32'h3c00f553),
	.w5(32'hbb0de525),
	.w6(32'h3b602881),
	.w7(32'hbc122d32),
	.w8(32'h3ba0a983),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ebfaa),
	.w1(32'h3c5a97a4),
	.w2(32'hbbfcc0c3),
	.w3(32'h3a092e5b),
	.w4(32'h3a47189d),
	.w5(32'h3b4cf957),
	.w6(32'h3d0e0718),
	.w7(32'hbab977bd),
	.w8(32'h3a531b12),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0f128),
	.w1(32'hbaef922d),
	.w2(32'h3bd379f2),
	.w3(32'h3a2bf0df),
	.w4(32'hbb51c60e),
	.w5(32'h39d768de),
	.w6(32'hbb796a6b),
	.w7(32'h3b07fd7c),
	.w8(32'h3c2bcdf6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82dd02),
	.w1(32'hba4a1e96),
	.w2(32'hbc7b54d5),
	.w3(32'h3b2f3742),
	.w4(32'h3c014299),
	.w5(32'hbc09f3f2),
	.w6(32'h3bbbdffa),
	.w7(32'h3c000c0f),
	.w8(32'h3b9f4eb0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f443),
	.w1(32'h3c0fd690),
	.w2(32'h3c90828a),
	.w3(32'hbc3e640e),
	.w4(32'hbb9721bc),
	.w5(32'h3abf6f1e),
	.w6(32'hbb456a4f),
	.w7(32'h3c1d2147),
	.w8(32'hbaa93029),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b612),
	.w1(32'h3b88fe75),
	.w2(32'hbb95bddd),
	.w3(32'hb8b92fd6),
	.w4(32'h3c353279),
	.w5(32'hbbb09684),
	.w6(32'h3bfaab89),
	.w7(32'hb8ea6586),
	.w8(32'hba59d7ce),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2eed5),
	.w1(32'h3a86185c),
	.w2(32'hb8ea2683),
	.w3(32'h3b461138),
	.w4(32'hbc145e55),
	.w5(32'hbb32aac0),
	.w6(32'hbaa77e8a),
	.w7(32'h3bf2426b),
	.w8(32'hbb5f1d76),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc253007),
	.w1(32'h3c22ae4a),
	.w2(32'h3b3b1a3a),
	.w3(32'h3c4668a8),
	.w4(32'hbb090613),
	.w5(32'h3b1bea41),
	.w6(32'h3cb0b8ef),
	.w7(32'hbc3812c7),
	.w8(32'h3bf72d97),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cba3e9),
	.w1(32'hbb600333),
	.w2(32'h3b5cc48b),
	.w3(32'h3bd8a8c3),
	.w4(32'h393ca1b2),
	.w5(32'hbafe080f),
	.w6(32'h3a100291),
	.w7(32'h3964a3b4),
	.w8(32'h36e3e074),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8df734),
	.w1(32'hbc252b80),
	.w2(32'h3b5ef09a),
	.w3(32'hba6b9667),
	.w4(32'hbb049fae),
	.w5(32'h3b378e47),
	.w6(32'hbb96443e),
	.w7(32'h3c1663e2),
	.w8(32'h3b4e5899),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ac62f),
	.w1(32'h3acf3602),
	.w2(32'h3c19d823),
	.w3(32'h3a77da46),
	.w4(32'h3b280ba9),
	.w5(32'hbc385806),
	.w6(32'h3b4212e2),
	.w7(32'h3b296c5a),
	.w8(32'h3be57376),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb611175),
	.w1(32'h3bc4625c),
	.w2(32'hba7cbb48),
	.w3(32'h3bcadc02),
	.w4(32'h3c839489),
	.w5(32'hbba364a4),
	.w6(32'h3c0445bd),
	.w7(32'hbc530f33),
	.w8(32'h3c01b845),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9831bd5),
	.w1(32'h39e4bf4a),
	.w2(32'h3b514341),
	.w3(32'h3c346d8e),
	.w4(32'hba1067a7),
	.w5(32'h3baeab9d),
	.w6(32'h3b444905),
	.w7(32'h3b087cb9),
	.w8(32'h3c46c800),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9340d4),
	.w1(32'hbaaf74f1),
	.w2(32'hbb4e41ab),
	.w3(32'h3b4be937),
	.w4(32'hbb060b72),
	.w5(32'hb8ea8e2e),
	.w6(32'hbc0c998e),
	.w7(32'hbb386210),
	.w8(32'h3c1005c9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce951ef),
	.w1(32'hbb84e4a3),
	.w2(32'hbc3afb71),
	.w3(32'h3ad1b695),
	.w4(32'h3a279306),
	.w5(32'hbb099cb8),
	.w6(32'h3b9ce098),
	.w7(32'h3b7b0fd6),
	.w8(32'hbc604f12),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92ffb0),
	.w1(32'h3916b3a9),
	.w2(32'h3b10a64a),
	.w3(32'hb9e0ea0a),
	.w4(32'hbaeb2f81),
	.w5(32'hba0d0e5f),
	.w6(32'h3c18d91f),
	.w7(32'h3bd83f1b),
	.w8(32'hbc25b528),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee14d2),
	.w1(32'h3a842fba),
	.w2(32'h3c40efd5),
	.w3(32'h3bbc388f),
	.w4(32'hbbe60287),
	.w5(32'hbc0b2c67),
	.w6(32'h3c118507),
	.w7(32'h3c41f3ff),
	.w8(32'h3bf668a1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a88d2),
	.w1(32'h3c1506a0),
	.w2(32'hb9e86ba4),
	.w3(32'h3a4b6307),
	.w4(32'h3bf2eacc),
	.w5(32'hbb10b88a),
	.w6(32'h3b4cc2bd),
	.w7(32'hbb45edcd),
	.w8(32'h3bcb6e29),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac69eb),
	.w1(32'hbb9d347a),
	.w2(32'hbb41d6bb),
	.w3(32'hbba19c70),
	.w4(32'hb9e7bb04),
	.w5(32'h3865fb3b),
	.w6(32'h3c5f6185),
	.w7(32'h3b851084),
	.w8(32'hb84fdd36),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb773),
	.w1(32'hbb4af7b6),
	.w2(32'h388b3bbc),
	.w3(32'h3abfd293),
	.w4(32'h3b46dfbe),
	.w5(32'h3b1baa72),
	.w6(32'h3b692653),
	.w7(32'hbadb6ea0),
	.w8(32'hbbe80241),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39532421),
	.w1(32'h3bdbf035),
	.w2(32'h3c3d7dc5),
	.w3(32'h3b7b709e),
	.w4(32'h3bd2b588),
	.w5(32'h3b49564a),
	.w6(32'h3b7e071a),
	.w7(32'hb63bad4e),
	.w8(32'h3b83581f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc71c74),
	.w1(32'h3b8ca48d),
	.w2(32'hbba21b92),
	.w3(32'hbb558e94),
	.w4(32'h3cbb71a2),
	.w5(32'hbba59ba0),
	.w6(32'h39143512),
	.w7(32'h3b12d295),
	.w8(32'h3b7511ac),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ae1bbf),
	.w1(32'hbc8feb34),
	.w2(32'hba776dae),
	.w3(32'h3b0421f0),
	.w4(32'h3c448a3d),
	.w5(32'h3c85ffb0),
	.w6(32'h3bd4ccc3),
	.w7(32'h3c12f93e),
	.w8(32'h3c47198d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd48527),
	.w1(32'h3c37b5b1),
	.w2(32'hbc0dd725),
	.w3(32'h3c0c01aa),
	.w4(32'h3a4342e0),
	.w5(32'h3b648c9c),
	.w6(32'h3b9db205),
	.w7(32'h3cacf057),
	.w8(32'h3b903a16),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82cadd),
	.w1(32'hbcea31ba),
	.w2(32'hbc0de1a5),
	.w3(32'hbaa974e7),
	.w4(32'hbbd58109),
	.w5(32'h3bf9e761),
	.w6(32'h3bd12c2e),
	.w7(32'hba45245c),
	.w8(32'hbc064dec),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80879a),
	.w1(32'h3c15d1fc),
	.w2(32'hb90bffd4),
	.w3(32'hbca1ec22),
	.w4(32'hbb0fa465),
	.w5(32'h3b261cf1),
	.w6(32'hbb80a58b),
	.w7(32'hbac94f64),
	.w8(32'hb9124d38),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7be1b4),
	.w1(32'h3c1a65e5),
	.w2(32'hba95363c),
	.w3(32'hbc1c2c99),
	.w4(32'hb9010577),
	.w5(32'h3d5ebdec),
	.w6(32'h3b2fef4d),
	.w7(32'hbad17ff7),
	.w8(32'hbb87734e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d3bf7),
	.w1(32'hb8feed1f),
	.w2(32'hbc1e35d3),
	.w3(32'hbb170c02),
	.w4(32'hba2e13dd),
	.w5(32'hba07d83e),
	.w6(32'hbb9fdde9),
	.w7(32'h3bbca5e3),
	.w8(32'hb7ac648f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3338f3),
	.w1(32'hb8f8ae51),
	.w2(32'h3a1a7bf1),
	.w3(32'hba762acf),
	.w4(32'h3a111999),
	.w5(32'h3bbd0ce8),
	.w6(32'h3cd8b0a7),
	.w7(32'h3c73ae68),
	.w8(32'h3d1d25e7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c7d24),
	.w1(32'hbb208953),
	.w2(32'hbaff56ed),
	.w3(32'hbc9eba58),
	.w4(32'h39d46dc1),
	.w5(32'hba731560),
	.w6(32'h3c6e9fdf),
	.w7(32'h3c143b6d),
	.w8(32'hbc7c31f5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b031d3c),
	.w1(32'h3ae2a530),
	.w2(32'h3a0c966e),
	.w3(32'h3c22b878),
	.w4(32'hba9992a2),
	.w5(32'hbbf11fab),
	.w6(32'hb94eda92),
	.w7(32'hbaa7e1d0),
	.w8(32'hbaba883c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdeeff),
	.w1(32'h3b736a51),
	.w2(32'h3b6ab9cb),
	.w3(32'hbc459bca),
	.w4(32'h3b87f5db),
	.w5(32'hbb7a9f86),
	.w6(32'hbb46a08d),
	.w7(32'hbb5c8db0),
	.w8(32'hbb73587f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d72c1),
	.w1(32'h3ba1340a),
	.w2(32'h3b33d5e5),
	.w3(32'hbc03fd8b),
	.w4(32'h3b337bdd),
	.w5(32'hbac77a37),
	.w6(32'hbbb0d0d3),
	.w7(32'h3cc1329b),
	.w8(32'h3b2841f9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfe251),
	.w1(32'hbc36c600),
	.w2(32'hbc737ae2),
	.w3(32'hbadf6ee9),
	.w4(32'h3b9edf80),
	.w5(32'hbc0225a0),
	.w6(32'h3bc10321),
	.w7(32'hbad8c709),
	.w8(32'hbbb6ffb0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27da34),
	.w1(32'hba13651a),
	.w2(32'hbb02bf84),
	.w3(32'hbc941b7b),
	.w4(32'hbbd23707),
	.w5(32'h3b82d88e),
	.w6(32'hbb1c470f),
	.w7(32'h3b7dbf4d),
	.w8(32'hbbbb2ec7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a275f),
	.w1(32'hbba23ba5),
	.w2(32'hbbbf62cf),
	.w3(32'h388c5eed),
	.w4(32'h38a59360),
	.w5(32'hbb0f4f14),
	.w6(32'h3c3ded7a),
	.w7(32'hbb1af1b1),
	.w8(32'hbc13d8d5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbab056),
	.w1(32'hbad2e753),
	.w2(32'hba96cd0b),
	.w3(32'hbb8cf88b),
	.w4(32'hbb083c8c),
	.w5(32'hbc2f8727),
	.w6(32'hb9fe7df3),
	.w7(32'hbd3a8daa),
	.w8(32'h3b219afd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8296e3),
	.w1(32'hb5aac3d5),
	.w2(32'hba31a0b0),
	.w3(32'hbb901fca),
	.w4(32'h3c7e34e2),
	.w5(32'hbba29a1e),
	.w6(32'h3b5656ce),
	.w7(32'hbab317b6),
	.w8(32'h3b0d69e9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8bff3),
	.w1(32'h3a9af083),
	.w2(32'hbba85a1b),
	.w3(32'h3a3829b6),
	.w4(32'hbbd40c79),
	.w5(32'hbd189ea9),
	.w6(32'h3a778cfd),
	.w7(32'hbbca211a),
	.w8(32'h3bf2f2b4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e4d3b),
	.w1(32'hbb048c87),
	.w2(32'hbbb48713),
	.w3(32'h3c9e1c31),
	.w4(32'h3b71cf73),
	.w5(32'h3d06f385),
	.w6(32'h3c0fc6ee),
	.w7(32'hbc2edaae),
	.w8(32'h3a39d54e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9141ae),
	.w1(32'hbb51c984),
	.w2(32'h3afcbf40),
	.w3(32'h3bab478c),
	.w4(32'h3c34ffcb),
	.w5(32'h3bf57760),
	.w6(32'h3b0e67b9),
	.w7(32'h3b30615b),
	.w8(32'h3b29116a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22b341),
	.w1(32'hbb58ee2e),
	.w2(32'h3b804192),
	.w3(32'h3b9d2651),
	.w4(32'h3b0a66c8),
	.w5(32'h38fd0bb2),
	.w6(32'hbc099550),
	.w7(32'h3a0e9820),
	.w8(32'hbba0217e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3edcaa),
	.w1(32'hbbce13fc),
	.w2(32'h383ad763),
	.w3(32'h3afdfd0f),
	.w4(32'hbb881bd4),
	.w5(32'hbb812a6c),
	.w6(32'hb8d43222),
	.w7(32'hbae2e377),
	.w8(32'h3bc1bd09),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8821f0),
	.w1(32'hbb50e7c2),
	.w2(32'hba6c1aa9),
	.w3(32'hbb20989b),
	.w4(32'hbc712a7c),
	.w5(32'hbc4829c3),
	.w6(32'hbbdb14b5),
	.w7(32'h38815f3e),
	.w8(32'hbbf92350),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b352868),
	.w1(32'hbb0aa48d),
	.w2(32'h3b96bf50),
	.w3(32'hbc93337c),
	.w4(32'h3b6581eb),
	.w5(32'hbd26ddd1),
	.w6(32'h3b6e8579),
	.w7(32'h3d4982ca),
	.w8(32'hbbc9f03a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f3f57),
	.w1(32'h3b3bfebb),
	.w2(32'hbb957258),
	.w3(32'h3996164f),
	.w4(32'h3c07685d),
	.w5(32'h3b2d49a5),
	.w6(32'h3c18a0ac),
	.w7(32'h3bc97fe6),
	.w8(32'h3b1e80b2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c256d),
	.w1(32'hba580a73),
	.w2(32'h3cc57383),
	.w3(32'hbb8923da),
	.w4(32'hbc8a0fc9),
	.w5(32'hbc9cb927),
	.w6(32'h3b7957a2),
	.w7(32'h3bafdc6a),
	.w8(32'hb8e92d08),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f9cde),
	.w1(32'hb8c1a505),
	.w2(32'h3c21621e),
	.w3(32'h3c84517f),
	.w4(32'hbb4695f6),
	.w5(32'hbc57bcc7),
	.w6(32'hbb5fb25f),
	.w7(32'h39141358),
	.w8(32'hbbc322df),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5d82e),
	.w1(32'hbb85681f),
	.w2(32'hbbcb9a15),
	.w3(32'h39234aa1),
	.w4(32'h3c444742),
	.w5(32'hbbe984fc),
	.w6(32'h394e6cc0),
	.w7(32'h3d0a353e),
	.w8(32'hbb76413a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc712e44),
	.w1(32'h3ccb987f),
	.w2(32'hba618cc9),
	.w3(32'hbba665ef),
	.w4(32'h3a8b51ef),
	.w5(32'h3b78b2c5),
	.w6(32'hbb397676),
	.w7(32'h3c0d1412),
	.w8(32'hbb8e279d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ca7d8),
	.w1(32'hbb717af8),
	.w2(32'hbd0946e5),
	.w3(32'hbb592779),
	.w4(32'hbabb75b0),
	.w5(32'h3bbd396f),
	.w6(32'hbae19a1f),
	.w7(32'h3a9acdb9),
	.w8(32'hbc60a90d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb799f93),
	.w1(32'hbbcbfc5d),
	.w2(32'h3a9a9ca8),
	.w3(32'hbbc0b1cb),
	.w4(32'h3baa60f5),
	.w5(32'hbbba2d6b),
	.w6(32'hbbde84ee),
	.w7(32'hbaf4cf9f),
	.w8(32'h3be37064),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b072f35),
	.w1(32'hba09e02d),
	.w2(32'h39f9e713),
	.w3(32'h3c4dca13),
	.w4(32'h3b250a24),
	.w5(32'h3a4b1d82),
	.w6(32'hbaf8db0e),
	.w7(32'hbb04d419),
	.w8(32'hb9ccf83d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c18fa),
	.w1(32'h3c3c87fe),
	.w2(32'hbb84221c),
	.w3(32'hbaa08d5a),
	.w4(32'h3c51bd5d),
	.w5(32'h3a269354),
	.w6(32'h3add69f2),
	.w7(32'hbc2e3f23),
	.w8(32'hb916721b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f83c91),
	.w1(32'hbb585928),
	.w2(32'h39be30e0),
	.w3(32'hbbf9c0ea),
	.w4(32'h3b6c543f),
	.w5(32'h37cac629),
	.w6(32'h3a3af041),
	.w7(32'hbb93c6b1),
	.w8(32'hbb27d4c2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b809a32),
	.w1(32'hbb842f5f),
	.w2(32'hbba0b921),
	.w3(32'hbba01d1d),
	.w4(32'hbb1afc4a),
	.w5(32'h3a34cb43),
	.w6(32'h3b0437a2),
	.w7(32'h3c083e04),
	.w8(32'hbc3e3aa6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c63b4),
	.w1(32'hb97075d1),
	.w2(32'h3c5863c5),
	.w3(32'h3b7f87f5),
	.w4(32'hbb1d55f4),
	.w5(32'hbbd2324b),
	.w6(32'hba8bcf2d),
	.w7(32'hbaff9c09),
	.w8(32'h3c6866b4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30f7ec),
	.w1(32'hbc23f306),
	.w2(32'h3c9ea25d),
	.w3(32'hbb360062),
	.w4(32'hba115326),
	.w5(32'h3813be07),
	.w6(32'h3b567c15),
	.w7(32'h3b3b0156),
	.w8(32'h3b882a11),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8e27e),
	.w1(32'hbb5daf95),
	.w2(32'h3b4c1517),
	.w3(32'hbbb54ef2),
	.w4(32'hbb2ff766),
	.w5(32'hbbb14d65),
	.w6(32'h3a53023c),
	.w7(32'h3bef2c2c),
	.w8(32'h3b2ffccb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13d09d),
	.w1(32'h3b23bd2d),
	.w2(32'h3b503455),
	.w3(32'h3b6ac534),
	.w4(32'hbba926b7),
	.w5(32'h3ac2f284),
	.w6(32'h3a8814a3),
	.w7(32'hbbc48ccb),
	.w8(32'h38358f57),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa16821),
	.w1(32'hbb08f2d6),
	.w2(32'hbd00b12e),
	.w3(32'h3a7892a2),
	.w4(32'hba3ede85),
	.w5(32'hbbd0349b),
	.w6(32'hbb1e1a80),
	.w7(32'h3b583ba5),
	.w8(32'h3ae55761),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6adb0a),
	.w1(32'hbaa0d30b),
	.w2(32'hba333fc6),
	.w3(32'h3ba13cca),
	.w4(32'hbc080622),
	.w5(32'h3b9558ee),
	.w6(32'h3bc4a8ca),
	.w7(32'hbbbff351),
	.w8(32'h3ade24d9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb602aef),
	.w1(32'h3af4ff68),
	.w2(32'h3b970799),
	.w3(32'h3ae5b403),
	.w4(32'hbbd49b42),
	.w5(32'h3bb51bb7),
	.w6(32'hbb2ff182),
	.w7(32'hbc8b32a5),
	.w8(32'h3bc443bd),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1288fb),
	.w1(32'h3c17d3ab),
	.w2(32'hbba2491e),
	.w3(32'h3ad358e5),
	.w4(32'h3bb9c45c),
	.w5(32'h3ac3ab4a),
	.w6(32'hba9349f1),
	.w7(32'h3a7f569e),
	.w8(32'h3b93bef7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba245433),
	.w1(32'h3b23c16b),
	.w2(32'hbb878adc),
	.w3(32'h3bc39359),
	.w4(32'h3b8b8ba0),
	.w5(32'h3b4a4f1b),
	.w6(32'h3aa560f6),
	.w7(32'hbb5f35d5),
	.w8(32'h3bdabef0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f906),
	.w1(32'hbae070fb),
	.w2(32'hbcb1e001),
	.w3(32'hb93bce56),
	.w4(32'h3af7018f),
	.w5(32'h388169a2),
	.w6(32'h3b15fa6a),
	.w7(32'hbb2ef98e),
	.w8(32'hbbc09e2a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bee87f),
	.w1(32'hb9946aac),
	.w2(32'hbb924e70),
	.w3(32'h3ad9db1f),
	.w4(32'hbb7df7ac),
	.w5(32'h3c3b9868),
	.w6(32'hbbc5208f),
	.w7(32'h3b35a9f2),
	.w8(32'h3bef9348),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a583e22),
	.w1(32'hbbc68db9),
	.w2(32'hbb398675),
	.w3(32'hbb974525),
	.w4(32'h3a32b0f4),
	.w5(32'h3c035c1f),
	.w6(32'h3a74a1e0),
	.w7(32'hbb808620),
	.w8(32'h3c094494),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6247cb),
	.w1(32'h3a0ebb43),
	.w2(32'hbb732f72),
	.w3(32'hbafd3e41),
	.w4(32'hbbf66896),
	.w5(32'h3aef9c3b),
	.w6(32'hbc679b90),
	.w7(32'hbad96562),
	.w8(32'h3bc9decf),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6b6e1),
	.w1(32'h39fae2a0),
	.w2(32'hba8ecda2),
	.w3(32'h3a8c9004),
	.w4(32'h38b45a46),
	.w5(32'hbbe5f539),
	.w6(32'h3baf3b95),
	.w7(32'h3b130219),
	.w8(32'h3b45da77),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884b222),
	.w1(32'hbba70d37),
	.w2(32'h37b46203),
	.w3(32'h3c30c5a6),
	.w4(32'hbb650936),
	.w5(32'hbc4fddf3),
	.w6(32'hba8c6370),
	.w7(32'h3c0f4a1e),
	.w8(32'hbba38f41),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695524),
	.w1(32'h3b9d1ffe),
	.w2(32'h3bea5d83),
	.w3(32'h38c18d7c),
	.w4(32'hba4aaffa),
	.w5(32'h3cd592f9),
	.w6(32'hbb999c77),
	.w7(32'hbd048702),
	.w8(32'h3a0e6b01),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39938920),
	.w1(32'hbb6be01a),
	.w2(32'hbb985e39),
	.w3(32'hbb77e98e),
	.w4(32'hbb3601c9),
	.w5(32'h3c31f24d),
	.w6(32'h3ad52a64),
	.w7(32'hb9984390),
	.w8(32'hbae9fd6b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb501a4),
	.w1(32'hbb16c3ce),
	.w2(32'hbce69ef1),
	.w3(32'h3a4afe5e),
	.w4(32'h3b9d8dbd),
	.w5(32'hba9d04dd),
	.w6(32'hbc5ff411),
	.w7(32'h3b8626a1),
	.w8(32'h3bdf2b35),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7580ff),
	.w1(32'hbb30be75),
	.w2(32'h3a09c89e),
	.w3(32'hba9735ba),
	.w4(32'h3b5071af),
	.w5(32'hbb8c7653),
	.w6(32'hbb6304d0),
	.w7(32'hbb339056),
	.w8(32'hbd33f9f8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aefb3),
	.w1(32'hb7bbd1fc),
	.w2(32'hbb750d61),
	.w3(32'hbb614cde),
	.w4(32'h3c53df5e),
	.w5(32'hb799dcc0),
	.w6(32'h3b6fb985),
	.w7(32'h3bed8e73),
	.w8(32'h3a8d8477),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb657ad4),
	.w1(32'h3ab706ae),
	.w2(32'hb90872cb),
	.w3(32'hbaf3ae21),
	.w4(32'hb903d933),
	.w5(32'h3b5cab2e),
	.w6(32'h3b3c0817),
	.w7(32'hb9ee5cfc),
	.w8(32'h3d73da01),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f7d80),
	.w1(32'h3a42427c),
	.w2(32'hba7ed870),
	.w3(32'hbbb69b97),
	.w4(32'hbaf57d16),
	.w5(32'hbc431af7),
	.w6(32'h3c0c4b8f),
	.w7(32'hbb1d07a5),
	.w8(32'hbb1a5373),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a64cf),
	.w1(32'h3c61ff1b),
	.w2(32'hbc010cd5),
	.w3(32'hba945864),
	.w4(32'hb7c2e8af),
	.w5(32'h3b113974),
	.w6(32'hbb5d4988),
	.w7(32'hbb99975e),
	.w8(32'h3adef06f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a9f3d),
	.w1(32'hbbabf0cf),
	.w2(32'hbbac8905),
	.w3(32'h3c47d5ff),
	.w4(32'hba80579f),
	.w5(32'h3a0fcc04),
	.w6(32'hbbdb081a),
	.w7(32'hbb7ebd57),
	.w8(32'h3bc01755),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf62ca2),
	.w1(32'h3b138eb0),
	.w2(32'hbb130174),
	.w3(32'hba64ed28),
	.w4(32'hba319a27),
	.w5(32'hbb55d9ec),
	.w6(32'hbc1e4713),
	.w7(32'hbc913311),
	.w8(32'hbc8068c9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80cc7),
	.w1(32'hbb9a3e7e),
	.w2(32'hba4a977a),
	.w3(32'hbb30a2a1),
	.w4(32'hbb03a11a),
	.w5(32'hbc909d83),
	.w6(32'hb9fc27dc),
	.w7(32'hbc0b7e2f),
	.w8(32'h3caebce9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7f8017),
	.w1(32'hb99b551c),
	.w2(32'hbb4fe7ec),
	.w3(32'hbabc3a2e),
	.w4(32'hbc42a295),
	.w5(32'hbb9cb100),
	.w6(32'h3893a41b),
	.w7(32'hbbdadfe7),
	.w8(32'h3d39ed2d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a43e8),
	.w1(32'hbb33ac82),
	.w2(32'h3cdb8e61),
	.w3(32'h3aa50783),
	.w4(32'h3baff56d),
	.w5(32'h3aaa3ce2),
	.w6(32'hbb93d6ab),
	.w7(32'hbb068978),
	.w8(32'hbc0088d9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ab396),
	.w1(32'h3bc33393),
	.w2(32'h3c05c474),
	.w3(32'hbaa6ebfc),
	.w4(32'h389c2901),
	.w5(32'hbb66fe8b),
	.w6(32'hbb3d7998),
	.w7(32'h3c12bf40),
	.w8(32'h3bdf23c5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e323f),
	.w1(32'hbba5fd07),
	.w2(32'h3b2c399f),
	.w3(32'hbc38d61c),
	.w4(32'hba5c989a),
	.w5(32'hbbd0bfae),
	.w6(32'hb94d0ba2),
	.w7(32'hbb4aa695),
	.w8(32'hb90cb723),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8da6ea),
	.w1(32'h3a770c07),
	.w2(32'hbba84f11),
	.w3(32'h3cfb2342),
	.w4(32'h39ae51f7),
	.w5(32'hbc80c687),
	.w6(32'h3bcfbc03),
	.w7(32'hba512758),
	.w8(32'hbb4f826b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb360c99),
	.w1(32'h39a66b4e),
	.w2(32'h3ad28d46),
	.w3(32'h3bc9ef35),
	.w4(32'h3862a4bc),
	.w5(32'hbc0f8e1d),
	.w6(32'hbc28c3c8),
	.w7(32'h3a906dda),
	.w8(32'hbc446179),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc836e28),
	.w1(32'hbb17490e),
	.w2(32'hbb5f13ef),
	.w3(32'hbb3a93a2),
	.w4(32'h3acf6b9d),
	.w5(32'hbc04a1d5),
	.w6(32'h3a8224b9),
	.w7(32'h3c67cba5),
	.w8(32'h3b8df67d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cbfbb),
	.w1(32'h3bd226d2),
	.w2(32'hbbf60e3d),
	.w3(32'h3c10e006),
	.w4(32'h3c80b4d1),
	.w5(32'hbbb138df),
	.w6(32'hbc2bcb5c),
	.w7(32'h3c8ca7e6),
	.w8(32'hbbedb7f0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e1678),
	.w1(32'hbb22bad6),
	.w2(32'hbc9b25fd),
	.w3(32'hbbe525f8),
	.w4(32'hbb147fa9),
	.w5(32'h3b32423c),
	.w6(32'hbb480333),
	.w7(32'hbb1f4540),
	.w8(32'hbb944871),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1518da),
	.w1(32'hbc9254a8),
	.w2(32'h3c33d3ae),
	.w3(32'hbb52d80d),
	.w4(32'hba69a97c),
	.w5(32'hbab49204),
	.w6(32'h3be34d57),
	.w7(32'hbb31aa54),
	.w8(32'h3d10a9a6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8d0d3),
	.w1(32'h3b59b439),
	.w2(32'hb9374f5b),
	.w3(32'hbbe7c63a),
	.w4(32'h3b8af277),
	.w5(32'hbc465de9),
	.w6(32'h3bab2011),
	.w7(32'h3b2003da),
	.w8(32'h3bdb1113),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85691e),
	.w1(32'h3aa2daee),
	.w2(32'hbbdcf2ac),
	.w3(32'h3bd6a32b),
	.w4(32'hb97d6dd9),
	.w5(32'hbb9d797e),
	.w6(32'hbbbc43e9),
	.w7(32'hbad9123b),
	.w8(32'hbb884624),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a59aa),
	.w1(32'h3bf08845),
	.w2(32'hbc668ad1),
	.w3(32'h3c443bba),
	.w4(32'hbad5fb88),
	.w5(32'hb895496b),
	.w6(32'h35f2285f),
	.w7(32'hbb538b02),
	.w8(32'hbb1d14b3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd13e7f),
	.w1(32'h3b28df77),
	.w2(32'hbcd83103),
	.w3(32'hbb919413),
	.w4(32'h3b80cde6),
	.w5(32'hbc593609),
	.w6(32'hbafbbba1),
	.w7(32'hbc6d527c),
	.w8(32'hbcdf14e5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c586310),
	.w1(32'h3b388955),
	.w2(32'hbc6a5e38),
	.w3(32'hbcb558a3),
	.w4(32'hbc0de1e9),
	.w5(32'hbb0ab4fc),
	.w6(32'hbc6d2205),
	.w7(32'hbc1550d7),
	.w8(32'hbbec269e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf0f67),
	.w1(32'h3b1c39e9),
	.w2(32'hbc2393db),
	.w3(32'hbba008b2),
	.w4(32'h3bfdb93f),
	.w5(32'h3ad66494),
	.w6(32'hbb6435bd),
	.w7(32'hba01ab59),
	.w8(32'hbb5a90d9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b723a),
	.w1(32'h3a1e7568),
	.w2(32'hbb8de634),
	.w3(32'h3b6515a0),
	.w4(32'hbb2b4f70),
	.w5(32'hbb8ef8b7),
	.w6(32'hb9e34d2d),
	.w7(32'h3d03a5c8),
	.w8(32'hbb2d01d0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9291a2),
	.w1(32'hbbed984a),
	.w2(32'hbba99250),
	.w3(32'h396988ed),
	.w4(32'h3b8a462b),
	.w5(32'h38c52ce6),
	.w6(32'hbb992b48),
	.w7(32'hbba8493f),
	.w8(32'hba096688),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee12e7),
	.w1(32'hbcec9a1d),
	.w2(32'hbb3df954),
	.w3(32'h3bb3ac3c),
	.w4(32'h3a022e2b),
	.w5(32'hbb194c8e),
	.w6(32'hbbcfa3e6),
	.w7(32'hbbc62358),
	.w8(32'hbb76a9b5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dcfdb),
	.w1(32'h3b2d4f59),
	.w2(32'hbcfaf492),
	.w3(32'hbb520fc8),
	.w4(32'h3ad6d611),
	.w5(32'hbbb5360d),
	.w6(32'hbc6a3dc4),
	.w7(32'hbb9e6a40),
	.w8(32'h3bc5003c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcde286),
	.w1(32'h3caffd7e),
	.w2(32'hbbe8f7d3),
	.w3(32'h3cf35c5f),
	.w4(32'h3aee2080),
	.w5(32'hb900492c),
	.w6(32'hbbc34619),
	.w7(32'hbc093848),
	.w8(32'hbc1e1b8d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc106d42),
	.w1(32'hbca410e5),
	.w2(32'h3bbec943),
	.w3(32'hba94a195),
	.w4(32'h3b965fd6),
	.w5(32'hbb1114c0),
	.w6(32'h3ba4d384),
	.w7(32'hbb46b45b),
	.w8(32'h3cbd79f0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc0b34),
	.w1(32'hbbffc733),
	.w2(32'hbc0f0669),
	.w3(32'h3a21a76a),
	.w4(32'h3a2c2afe),
	.w5(32'h3927ae29),
	.w6(32'h382bfa28),
	.w7(32'hb9a8ac68),
	.w8(32'hba82d51b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a310db4),
	.w1(32'h3cd29a2b),
	.w2(32'h3cfca61f),
	.w3(32'h3b9cca6f),
	.w4(32'h3ab9b099),
	.w5(32'h3a96fdf9),
	.w6(32'hbbd367c5),
	.w7(32'hbcb76d7c),
	.w8(32'hbbcdf60c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ac2f5),
	.w1(32'h3b7affc3),
	.w2(32'hbbe8bbfb),
	.w3(32'h3a3769c5),
	.w4(32'h39ac22dc),
	.w5(32'h3b99bc04),
	.w6(32'h3d084920),
	.w7(32'h3b97675d),
	.w8(32'h3ba54516),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023cd1),
	.w1(32'h3a75ac74),
	.w2(32'h3b41db29),
	.w3(32'hbd23a241),
	.w4(32'hbb16502a),
	.w5(32'hbb511093),
	.w6(32'hbbe1b458),
	.w7(32'h3d25aa1d),
	.w8(32'hbb8af459),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72cbbd),
	.w1(32'h3bcef79b),
	.w2(32'hbc416eba),
	.w3(32'hbbe41429),
	.w4(32'hbc12508c),
	.w5(32'hbb17c69a),
	.w6(32'hbb870489),
	.w7(32'h3b06875d),
	.w8(32'h3ae3a659),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1212ca),
	.w1(32'h3b450448),
	.w2(32'hbca3f70a),
	.w3(32'h3b620d0d),
	.w4(32'hbaf5cf54),
	.w5(32'hbbc6d90b),
	.w6(32'hbbd62c15),
	.w7(32'h398826a1),
	.w8(32'hbb3702ef),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ac2a9),
	.w1(32'hbc6c8ef8),
	.w2(32'h3c0a0ede),
	.w3(32'h3b9a405b),
	.w4(32'hbc205953),
	.w5(32'hbae72f47),
	.w6(32'h3b4016a8),
	.w7(32'h3b7cf2de),
	.w8(32'hbc0078b7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a6007),
	.w1(32'hbc03b542),
	.w2(32'h3bb20fd8),
	.w3(32'hbb2b8643),
	.w4(32'hbc1dce90),
	.w5(32'hbb689db2),
	.w6(32'h3b4c991e),
	.w7(32'h3978a661),
	.w8(32'h3a3c76b7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59d3b2),
	.w1(32'h3aa906a8),
	.w2(32'hbad33ee1),
	.w3(32'h3d149ffa),
	.w4(32'h3b856834),
	.w5(32'h3b8764f0),
	.w6(32'hb87be2ab),
	.w7(32'hbb1abf51),
	.w8(32'h3bc6ffaa),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef858a),
	.w1(32'hbd123d62),
	.w2(32'h3b3034e7),
	.w3(32'h3bb0d7a1),
	.w4(32'hba67b7c8),
	.w5(32'hbc80d46c),
	.w6(32'h3afaf8f6),
	.w7(32'hbc35e376),
	.w8(32'h3a9bfa12),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba259f45),
	.w1(32'hba574393),
	.w2(32'h3bc3636e),
	.w3(32'hb9d787e4),
	.w4(32'hbc7bb913),
	.w5(32'hbba04d32),
	.w6(32'h3d00cb8d),
	.w7(32'hb964932b),
	.w8(32'h3aaaa1a0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba57d32),
	.w1(32'hbaef7846),
	.w2(32'h392632b6),
	.w3(32'h3bc6ef6b),
	.w4(32'h3b93bcdb),
	.w5(32'h3b9cf921),
	.w6(32'hbb5db560),
	.w7(32'hbac0e5a7),
	.w8(32'hb992ce18),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae50da1),
	.w1(32'hbb021fed),
	.w2(32'h3bab64cb),
	.w3(32'hbba79f0e),
	.w4(32'hbb090312),
	.w5(32'h3a8aa07a),
	.w6(32'hbbca86a4),
	.w7(32'h3a85777f),
	.w8(32'h3b758291),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b7f3),
	.w1(32'hba883128),
	.w2(32'h3be1eccc),
	.w3(32'hbb0ccada),
	.w4(32'h3b132ee9),
	.w5(32'hba02fb23),
	.w6(32'h3a48cdeb),
	.w7(32'hbb2a6f41),
	.w8(32'hbb714414),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b848e),
	.w1(32'h3a519719),
	.w2(32'hbc5e51f1),
	.w3(32'h3b4c8af2),
	.w4(32'hba444b0c),
	.w5(32'h3ad1b034),
	.w6(32'h39e97731),
	.w7(32'hb9f11d41),
	.w8(32'h3afa9b5f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad613b3),
	.w1(32'hbb8fe16d),
	.w2(32'hbc0d3e17),
	.w3(32'h3b7123e7),
	.w4(32'hbcc652d7),
	.w5(32'hbbfc2054),
	.w6(32'h3b3789c8),
	.w7(32'h3bb78f1b),
	.w8(32'h3c3bcb93),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380318ca),
	.w1(32'hbc4bdad8),
	.w2(32'hbbc1f814),
	.w3(32'h3cea7199),
	.w4(32'h379c22bf),
	.w5(32'hba168efb),
	.w6(32'hbade1e55),
	.w7(32'h3c11789f),
	.w8(32'hbc173fda),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba654a0b),
	.w1(32'hbaa59851),
	.w2(32'h3b8a298c),
	.w3(32'hbb00457e),
	.w4(32'h3aebffbe),
	.w5(32'hbb8441d0),
	.w6(32'h3a0ea2fa),
	.w7(32'h3c962371),
	.w8(32'h3a61ddb7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75537e),
	.w1(32'h3be26994),
	.w2(32'hb68e8e5e),
	.w3(32'hbb968271),
	.w4(32'hbbf1e98d),
	.w5(32'h3cace2d2),
	.w6(32'h39f5e880),
	.w7(32'h3cf76d1a),
	.w8(32'hbb11b6ef),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba496817),
	.w1(32'hbbc81c4d),
	.w2(32'h3bcc2154),
	.w3(32'h3b0c9e83),
	.w4(32'hbba7406c),
	.w5(32'hbc2ef18c),
	.w6(32'h3a9b200f),
	.w7(32'h3b8d602a),
	.w8(32'hbba17932),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc806b6),
	.w1(32'hbc1cd98d),
	.w2(32'h3bf32805),
	.w3(32'hbd4073f3),
	.w4(32'h3c1fbebb),
	.w5(32'h3b8d19e1),
	.w6(32'h3c8baa9c),
	.w7(32'hbd6451eb),
	.w8(32'hbb2ae8da),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd665e),
	.w1(32'hbbc75541),
	.w2(32'hbc12bbbe),
	.w3(32'h3c841896),
	.w4(32'h3a8f0087),
	.w5(32'hbc27b307),
	.w6(32'hbb0a8337),
	.w7(32'hbb7bc55a),
	.w8(32'h3b2b3f17),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97bf3a),
	.w1(32'hb9ee0b75),
	.w2(32'h3a809dbd),
	.w3(32'hbbf52802),
	.w4(32'hbb97fa9e),
	.w5(32'h3b9941a7),
	.w6(32'h3aff5159),
	.w7(32'hbb1dd1f2),
	.w8(32'hbb01c52d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb82e),
	.w1(32'h3bd43ef1),
	.w2(32'hbb1f1a79),
	.w3(32'h3ae80ba5),
	.w4(32'hba6054c8),
	.w5(32'h3bea9f37),
	.w6(32'hbb8a3ccd),
	.w7(32'hb7f2667c),
	.w8(32'hbc04f4e5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16a70a),
	.w1(32'h3bea87e0),
	.w2(32'h3cb71b77),
	.w3(32'hbae64c37),
	.w4(32'hbc6b62ec),
	.w5(32'hbc34e686),
	.w6(32'hbbe0da1c),
	.w7(32'hbb321d07),
	.w8(32'hb9e01b60),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ceb17),
	.w1(32'hbbee4434),
	.w2(32'h3be2ce9e),
	.w3(32'h3bdd29f0),
	.w4(32'h3bd28e5a),
	.w5(32'h3a81154c),
	.w6(32'hbbf4b8bf),
	.w7(32'h3af36126),
	.w8(32'h3cf17bb6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17ec2f),
	.w1(32'h3bcfa739),
	.w2(32'hbb273fd9),
	.w3(32'hbcd05332),
	.w4(32'h3a941a3f),
	.w5(32'hb799055c),
	.w6(32'hbb07b0dc),
	.w7(32'hbbb4bfa7),
	.w8(32'h3a661597),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cf095),
	.w1(32'hb9139c46),
	.w2(32'h3c4e6e26),
	.w3(32'hbbe3e3ed),
	.w4(32'h3b404ca8),
	.w5(32'hbbf1db1d),
	.w6(32'hbacba6c8),
	.w7(32'h3ab036c7),
	.w8(32'hbb83236d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8bd9e),
	.w1(32'h3b2f96dc),
	.w2(32'hb9b3557d),
	.w3(32'h3acbaa50),
	.w4(32'h3bb4b28a),
	.w5(32'hbae0bcb3),
	.w6(32'hbaa29d5c),
	.w7(32'hbba40dd4),
	.w8(32'hbaf6d3b5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c120bcf),
	.w1(32'hbade15c4),
	.w2(32'hbc06a018),
	.w3(32'hbc230f75),
	.w4(32'h390b448c),
	.w5(32'hbce8824d),
	.w6(32'h3b2e5942),
	.w7(32'hbaa99a73),
	.w8(32'h3b37c28d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983681),
	.w1(32'hb7e9e24c),
	.w2(32'h3c11dce9),
	.w3(32'hbb8168f8),
	.w4(32'hba135df6),
	.w5(32'hbb812f7c),
	.w6(32'h3be42228),
	.w7(32'hbb78085d),
	.w8(32'h3bc63562),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedc115),
	.w1(32'h3b4d89d0),
	.w2(32'hbc1ca588),
	.w3(32'h3998955f),
	.w4(32'h3a9c3745),
	.w5(32'h3bbbc2c9),
	.w6(32'hb9cf4bbd),
	.w7(32'h3c4a95c0),
	.w8(32'h3a50c2de),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83838d),
	.w1(32'hba9f8fca),
	.w2(32'hbaf75a87),
	.w3(32'hbbbfbeb7),
	.w4(32'hbb7771e8),
	.w5(32'h3c73e932),
	.w6(32'h3b2438d4),
	.w7(32'hbb24d7fd),
	.w8(32'hba5c1b19),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc633d1),
	.w1(32'h3bf38a59),
	.w2(32'h3b253622),
	.w3(32'hbbdbe250),
	.w4(32'h3c11918f),
	.w5(32'h3c16a5f9),
	.w6(32'hbb452529),
	.w7(32'h3ac73259),
	.w8(32'hbb4fe592),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e41c4),
	.w1(32'h3a43577a),
	.w2(32'h3b244b29),
	.w3(32'h3b1f5cef),
	.w4(32'h3cdb186e),
	.w5(32'hbc15f006),
	.w6(32'hbb20b475),
	.w7(32'hbc51ba31),
	.w8(32'h3c4551ff),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd018f6),
	.w1(32'hbb55d472),
	.w2(32'h3c14ed80),
	.w3(32'h3c67b4a5),
	.w4(32'h3c42c8d7),
	.w5(32'h3b798bd3),
	.w6(32'h3b314c81),
	.w7(32'h3aa7ba45),
	.w8(32'hbbb93cde),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9acbd),
	.w1(32'h3c300506),
	.w2(32'hbb89c901),
	.w3(32'hbb1ad785),
	.w4(32'hb8d32421),
	.w5(32'h3c0a4e27),
	.w6(32'h3c3415a3),
	.w7(32'h3b525f32),
	.w8(32'h3b4f54b8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b13ce),
	.w1(32'h3b8c2561),
	.w2(32'h3b9458c4),
	.w3(32'h3c971937),
	.w4(32'hbbe004f3),
	.w5(32'h3bf6f914),
	.w6(32'h3ae41e61),
	.w7(32'h3ac0a47b),
	.w8(32'hbb2a8af5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15dc2e),
	.w1(32'h3b1bf05b),
	.w2(32'h3b73614e),
	.w3(32'h3a34e02e),
	.w4(32'h3c03ce70),
	.w5(32'hbc2ba66f),
	.w6(32'h3ac392bd),
	.w7(32'hbc4c5ab7),
	.w8(32'hbc1890ac),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedc769),
	.w1(32'hba304662),
	.w2(32'h3bcc4baf),
	.w3(32'h3bf5c472),
	.w4(32'h3c670797),
	.w5(32'h398749fc),
	.w6(32'hba2fd8a8),
	.w7(32'hbb561a13),
	.w8(32'hb9dfb6eb),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae0b8e),
	.w1(32'h3b1ac332),
	.w2(32'h3a8c462e),
	.w3(32'hbb399726),
	.w4(32'hbc2c1bc9),
	.w5(32'h399c8431),
	.w6(32'hbbb8cd76),
	.w7(32'h3c1383f2),
	.w8(32'hbc094379),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4efea2),
	.w1(32'h3c9342f5),
	.w2(32'h3c297f79),
	.w3(32'h3c404b8e),
	.w4(32'h3c50c540),
	.w5(32'hbb70da76),
	.w6(32'hbb495141),
	.w7(32'hbb5f4503),
	.w8(32'hbcfe7aa7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc313560),
	.w1(32'h3b9354e9),
	.w2(32'h3b31a169),
	.w3(32'hba91cfdb),
	.w4(32'h3be63b31),
	.w5(32'hbb89d2ec),
	.w6(32'h3b1e674c),
	.w7(32'h3b8725f7),
	.w8(32'h3c3a4e98),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76f5d6),
	.w1(32'hbb3c9bfd),
	.w2(32'hbb4d12ce),
	.w3(32'h3b152d94),
	.w4(32'hbb9345bf),
	.w5(32'h3b81f6af),
	.w6(32'hb99fae2d),
	.w7(32'hbc1bc756),
	.w8(32'hbac6862b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc58847),
	.w1(32'hbb2dcb7e),
	.w2(32'h3ba46071),
	.w3(32'hbb32c4be),
	.w4(32'hba3f4018),
	.w5(32'h3b943685),
	.w6(32'h3c96e34a),
	.w7(32'h3c80d2d9),
	.w8(32'hb81fbdaa),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8660),
	.w1(32'h3baa5233),
	.w2(32'h3b00b3ba),
	.w3(32'h3bd7c74c),
	.w4(32'hbb39d184),
	.w5(32'h3b435e37),
	.w6(32'hbc4b94e7),
	.w7(32'h3b3f9fd3),
	.w8(32'hba8f00bf),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52725),
	.w1(32'hbc020036),
	.w2(32'h3c909b63),
	.w3(32'h3b80ccb7),
	.w4(32'hbc339e26),
	.w5(32'h3bad2d5f),
	.w6(32'hbb2ee01c),
	.w7(32'h3b46b775),
	.w8(32'h3c6d57f0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed30a3),
	.w1(32'hbb6e4a7e),
	.w2(32'hba65b78f),
	.w3(32'hb9977cf8),
	.w4(32'hbba16b0b),
	.w5(32'h3b63f217),
	.w6(32'hbc1045ba),
	.w7(32'hbbb3dea9),
	.w8(32'hbc1f224d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98eafd7),
	.w1(32'hbc18c0b2),
	.w2(32'hba921f4a),
	.w3(32'hbb9225fd),
	.w4(32'h3aa3e0b4),
	.w5(32'h3a9f0497),
	.w6(32'hbc5c06f9),
	.w7(32'hbc3f8f41),
	.w8(32'hbb45f0a0),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fb29),
	.w1(32'h3c0a46b1),
	.w2(32'h3a05e127),
	.w3(32'h3a437117),
	.w4(32'h3b3f1ad0),
	.w5(32'h3af7c090),
	.w6(32'h3ce85673),
	.w7(32'h3c841e5b),
	.w8(32'hbbcd4144),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a03c9),
	.w1(32'hbb058f9e),
	.w2(32'hbb8148ea),
	.w3(32'h3bb5f229),
	.w4(32'hbb13c0a9),
	.w5(32'hbb6e0b3c),
	.w6(32'hbb264355),
	.w7(32'hba97901c),
	.w8(32'h3ab4e33d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16f944),
	.w1(32'h3bb68fdd),
	.w2(32'hbb146ae5),
	.w3(32'hba88f39e),
	.w4(32'hbb617368),
	.w5(32'hbadbbf51),
	.w6(32'hbb9e0966),
	.w7(32'h3bce7912),
	.w8(32'h3a2a4e25),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5141f25),
	.w1(32'hb724e349),
	.w2(32'hbb8b494f),
	.w3(32'hbb5c7a69),
	.w4(32'hbb193c27),
	.w5(32'hbbfa30ba),
	.w6(32'h3c4ebfd8),
	.w7(32'hbae7c4f8),
	.w8(32'hba6e0df5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78505b),
	.w1(32'hb9936d0e),
	.w2(32'hbbcd2106),
	.w3(32'hbc29e910),
	.w4(32'hbbf66412),
	.w5(32'h3c2ceee9),
	.w6(32'hbbca64c9),
	.w7(32'hba5be4c9),
	.w8(32'hba3bd18a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe490b),
	.w1(32'h3ba91029),
	.w2(32'hbbb53e17),
	.w3(32'h3c1e3ff4),
	.w4(32'h383c7cd4),
	.w5(32'hbbc3c7e4),
	.w6(32'hbbba02b1),
	.w7(32'h3a589204),
	.w8(32'hbb0450a4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b956802),
	.w1(32'h3c5a81cb),
	.w2(32'hbbfdd394),
	.w3(32'h3b6a390d),
	.w4(32'h3c113b7a),
	.w5(32'hbbdb9390),
	.w6(32'h3b4fd28a),
	.w7(32'h3c769c7c),
	.w8(32'hbbfc77e7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10cf21),
	.w1(32'hbba5918a),
	.w2(32'hbaf0c6c0),
	.w3(32'hbb64602d),
	.w4(32'h3c03496b),
	.w5(32'h3bb9fe46),
	.w6(32'h39790a43),
	.w7(32'h3bb04edd),
	.w8(32'h3bef5c0e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdca57f),
	.w1(32'hba38b5e1),
	.w2(32'hbc093043),
	.w3(32'hb959c4ab),
	.w4(32'hbbc9cb12),
	.w5(32'h3817f241),
	.w6(32'h3b403933),
	.w7(32'hba0b30e9),
	.w8(32'hb9ced4a9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72cc84),
	.w1(32'hbc5d61ac),
	.w2(32'hbbf2611f),
	.w3(32'hbb04e27f),
	.w4(32'h3c5e4b9a),
	.w5(32'hba523fff),
	.w6(32'h3c32ada0),
	.w7(32'hbb8a2872),
	.w8(32'hbc9d240a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ff06c),
	.w1(32'hbb4928ee),
	.w2(32'hbc0cc639),
	.w3(32'h3c10f79f),
	.w4(32'h3af2d08c),
	.w5(32'h3bcf6578),
	.w6(32'hb906c150),
	.w7(32'hb99bd8b8),
	.w8(32'h3b981f6e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b772dcf),
	.w1(32'hbb562050),
	.w2(32'hbc886b5f),
	.w3(32'h3bc15a59),
	.w4(32'hbbcd20f9),
	.w5(32'h3b8cabcb),
	.w6(32'h3aecdf68),
	.w7(32'hbc3cd51f),
	.w8(32'h3c501601),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5d8be),
	.w1(32'h3c033b42),
	.w2(32'hbb476efd),
	.w3(32'h3b1723e1),
	.w4(32'h3a399199),
	.w5(32'h3c235fa5),
	.w6(32'hbc0ce9fd),
	.w7(32'h3b2dfbac),
	.w8(32'h3c0c7323),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9eba8),
	.w1(32'hbb6b26ba),
	.w2(32'h3c7e8f63),
	.w3(32'h3a8fce9c),
	.w4(32'h3c5f35d0),
	.w5(32'hbb13c8dc),
	.w6(32'hbc8e5889),
	.w7(32'h3be46b71),
	.w8(32'h3baca894),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc165751),
	.w1(32'hbb94ece1),
	.w2(32'hba416b40),
	.w3(32'h3c38aee2),
	.w4(32'h3b9e3db3),
	.w5(32'h3bc6ab8d),
	.w6(32'hbc00ee86),
	.w7(32'hbb4538d6),
	.w8(32'hbc907a96),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule