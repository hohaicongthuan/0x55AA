module layer_10_featuremap_3(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4513c),
	.w1(32'hbb42b021),
	.w2(32'h3a64bb7c),
	.w3(32'h3be0c3b5),
	.w4(32'h3bc77088),
	.w5(32'hbbf48c7c),
	.w6(32'h3ab9a77b),
	.w7(32'h3a538605),
	.w8(32'hbc4bed64),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca9a1a),
	.w1(32'h3b270a68),
	.w2(32'hbc2edc7b),
	.w3(32'h3b82dd40),
	.w4(32'h3c12e307),
	.w5(32'hbc8ee617),
	.w6(32'hbbd4835d),
	.w7(32'h3c2980de),
	.w8(32'hbc22b912),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb160c3d),
	.w1(32'hbb83d965),
	.w2(32'hbc8027ca),
	.w3(32'hbc5eabca),
	.w4(32'hbbb75eea),
	.w5(32'hbc17738d),
	.w6(32'hbb28711c),
	.w7(32'hbbe416c4),
	.w8(32'hbbb28134),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3afef0),
	.w1(32'h3b89a423),
	.w2(32'hbc7ed274),
	.w3(32'hbcd6c930),
	.w4(32'hbc4cbdec),
	.w5(32'hbc1f9dab),
	.w6(32'hbc4f4bae),
	.w7(32'hbc54a0a5),
	.w8(32'hbbcaec85),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc5624),
	.w1(32'hbb72e13f),
	.w2(32'hbc15087b),
	.w3(32'hbc545970),
	.w4(32'hbb75e08c),
	.w5(32'h3b517476),
	.w6(32'hbbb607d9),
	.w7(32'hbb873dde),
	.w8(32'hbb9d0298),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c5e16),
	.w1(32'h3bf5dd3f),
	.w2(32'hbc2257b9),
	.w3(32'hbb2a2cd6),
	.w4(32'h3b3e3806),
	.w5(32'hbc2b197a),
	.w6(32'hbb07d1d6),
	.w7(32'h39b0b884),
	.w8(32'hbc216cfd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a4020),
	.w1(32'hbbd75219),
	.w2(32'hbb2f32a9),
	.w3(32'h3c2c11a8),
	.w4(32'hbb3a3a99),
	.w5(32'h3be8c01d),
	.w6(32'h3c313480),
	.w7(32'hbb252f72),
	.w8(32'h3b0d9ec9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0ff73),
	.w1(32'hbb4b48c1),
	.w2(32'h3b8d95e0),
	.w3(32'h3b48be85),
	.w4(32'h3c2acd48),
	.w5(32'h3bb576b9),
	.w6(32'h3c2507ed),
	.w7(32'hbb887d01),
	.w8(32'hba8c7658),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2b757),
	.w1(32'hbbc2c7c1),
	.w2(32'hbc1f4795),
	.w3(32'h3a1d0da4),
	.w4(32'hbbf9c15c),
	.w5(32'hbc22da71),
	.w6(32'h3a701c1e),
	.w7(32'hbb449bb1),
	.w8(32'hbc690441),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7a59e),
	.w1(32'hbc371916),
	.w2(32'hbbde2e82),
	.w3(32'hbb591f17),
	.w4(32'hbc082aef),
	.w5(32'hbbed3de1),
	.w6(32'hbb2b2f5f),
	.w7(32'hbbf5812b),
	.w8(32'hbb8b3357),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf0daf),
	.w1(32'hbae3c21b),
	.w2(32'hbc232eb4),
	.w3(32'hbb4d98f1),
	.w4(32'hbb4bb3ec),
	.w5(32'hbc54f5fd),
	.w6(32'h3a72fed8),
	.w7(32'hba64c033),
	.w8(32'hbbb0823d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bc791),
	.w1(32'hb98fc574),
	.w2(32'hbbfef46d),
	.w3(32'hbca72a31),
	.w4(32'hbc5f08e4),
	.w5(32'hbbdc4ce4),
	.w6(32'hbc87f764),
	.w7(32'hbc700b8e),
	.w8(32'hbb77b109),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e8c63),
	.w1(32'hbb8144a0),
	.w2(32'hbbf59079),
	.w3(32'h3be765b0),
	.w4(32'h3af61891),
	.w5(32'h39ca86b6),
	.w6(32'h3c2e2e14),
	.w7(32'h3bb910c1),
	.w8(32'hbbbcfa61),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c300651),
	.w1(32'h3b7c0676),
	.w2(32'hbb86af64),
	.w3(32'h3c91e066),
	.w4(32'h3c4eb3fd),
	.w5(32'h3ba46dd8),
	.w6(32'h3c4982be),
	.w7(32'h3b03f308),
	.w8(32'hbac137cf),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca389c1),
	.w1(32'hbae182f3),
	.w2(32'hbb6a2c45),
	.w3(32'hbc0b9691),
	.w4(32'h3c2a3e23),
	.w5(32'hbbdc8256),
	.w6(32'h3c05d46d),
	.w7(32'h3b7541bb),
	.w8(32'h39059fd7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da682),
	.w1(32'hbbc41afe),
	.w2(32'hbc052444),
	.w3(32'hbc01e965),
	.w4(32'hbba3d89d),
	.w5(32'hbb955005),
	.w6(32'hbb308518),
	.w7(32'hbb5ae55b),
	.w8(32'hbbe7a860),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba860940),
	.w1(32'hbb098305),
	.w2(32'h3b76ae07),
	.w3(32'h38995fd4),
	.w4(32'hba81f5fe),
	.w5(32'h3c0178f3),
	.w6(32'h3ad45612),
	.w7(32'hb90efc00),
	.w8(32'h3b14136d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf3088),
	.w1(32'hbb9e2c48),
	.w2(32'hbb726646),
	.w3(32'h3c5978c9),
	.w4(32'h3b95004c),
	.w5(32'hbb3c7e91),
	.w6(32'h3c317264),
	.w7(32'h3bf40da2),
	.w8(32'hbb9438f9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c412164),
	.w1(32'h3b9c24bd),
	.w2(32'hbc9a9b27),
	.w3(32'h3c45e9e2),
	.w4(32'h3c0be844),
	.w5(32'hbc008096),
	.w6(32'h3c645f5a),
	.w7(32'h3beb6363),
	.w8(32'hbbe6e21e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a6ce7),
	.w1(32'hbb339bf6),
	.w2(32'h3b23e454),
	.w3(32'hbcc7eba5),
	.w4(32'hbc84504b),
	.w5(32'h3ac037ac),
	.w6(32'hbc711e63),
	.w7(32'hbc6fd10b),
	.w8(32'hbb6f502e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a986ad5),
	.w1(32'hba64b4a7),
	.w2(32'h3aed2cda),
	.w3(32'h37ec5713),
	.w4(32'h3a037d36),
	.w5(32'hbb239a15),
	.w6(32'hbaeda43f),
	.w7(32'hba4b8191),
	.w8(32'hbbbf64de),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982f41),
	.w1(32'h3c00be89),
	.w2(32'h3b1cb3d5),
	.w3(32'hbc3c8562),
	.w4(32'h3bd58394),
	.w5(32'h3be9de0b),
	.w6(32'hbae08015),
	.w7(32'h3be7e878),
	.w8(32'h3c406f29),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2310cd),
	.w1(32'hbb3dc53c),
	.w2(32'hbbde7700),
	.w3(32'h3a8df6e9),
	.w4(32'h3b668109),
	.w5(32'hba927052),
	.w6(32'h3c082b39),
	.w7(32'hb6afe5d9),
	.w8(32'h3b8d612a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d9959),
	.w1(32'h3b512eff),
	.w2(32'hbbbac85a),
	.w3(32'h3bd43821),
	.w4(32'h3b38d738),
	.w5(32'h3b21b7f2),
	.w6(32'h3c3c6739),
	.w7(32'h3c170394),
	.w8(32'hbacca36b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4e6fe),
	.w1(32'h3b956e42),
	.w2(32'hbc2d5c48),
	.w3(32'h3c5ef0b8),
	.w4(32'h3c33acff),
	.w5(32'hbb5437e0),
	.w6(32'h3c05c7dd),
	.w7(32'h3c23b317),
	.w8(32'hbc26c06d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd28e84),
	.w1(32'hbc62fa71),
	.w2(32'hba8b19c3),
	.w3(32'hbc94819f),
	.w4(32'hbb7195e5),
	.w5(32'hbc2b3a90),
	.w6(32'hbc3e4754),
	.w7(32'hbaf27ed5),
	.w8(32'hbc556897),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72806b),
	.w1(32'hbc86ac1c),
	.w2(32'h38c53453),
	.w3(32'hbd2158a8),
	.w4(32'hbcc04edc),
	.w5(32'h3a28f0bd),
	.w6(32'hbcbae8d9),
	.w7(32'hbb01af92),
	.w8(32'h39a144a8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd63ead),
	.w1(32'h395a0761),
	.w2(32'hb9f91dff),
	.w3(32'hbb98995f),
	.w4(32'hbb041f48),
	.w5(32'h3b98b3f7),
	.w6(32'hbbdf6e93),
	.w7(32'hbbe8c0c5),
	.w8(32'h3b225f74),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33514b),
	.w1(32'hb9f57a7f),
	.w2(32'hbb32fecb),
	.w3(32'h3b8bb5f9),
	.w4(32'h3b9520bb),
	.w5(32'hba60c780),
	.w6(32'h3ba1b35e),
	.w7(32'h3c12e964),
	.w8(32'h3bf2b8b5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc0bfe),
	.w1(32'h3bd2c13b),
	.w2(32'hbb0ba36a),
	.w3(32'hbc6051d6),
	.w4(32'h3b2005c1),
	.w5(32'hbaf1504a),
	.w6(32'hbc61d209),
	.w7(32'hbac8c359),
	.w8(32'hbb3eabe2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba961f78),
	.w1(32'hba609778),
	.w2(32'hbc34a83d),
	.w3(32'hbb76dbc7),
	.w4(32'hbafb2f8c),
	.w5(32'hbc874ca0),
	.w6(32'hbb3afafa),
	.w7(32'hbb880f34),
	.w8(32'hbc749e5d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52570c),
	.w1(32'hbbe63b3d),
	.w2(32'hbc2e1e61),
	.w3(32'hbd072c4d),
	.w4(32'hbcf51de2),
	.w5(32'hbc9d7207),
	.w6(32'hbce77d44),
	.w7(32'hbca218a7),
	.w8(32'hbbdb622a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6c7d5),
	.w1(32'hbae6a465),
	.w2(32'hbbe945a4),
	.w3(32'hbc212669),
	.w4(32'hbbcdd2df),
	.w5(32'hbbc073b9),
	.w6(32'hbbf7fc1e),
	.w7(32'hbb1f79f1),
	.w8(32'h3a8df9f1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0444be),
	.w1(32'h3aabf916),
	.w2(32'hbc2c4f43),
	.w3(32'hbbd827ae),
	.w4(32'h3af87faf),
	.w5(32'hbc30d5de),
	.w6(32'hbaa1a540),
	.w7(32'h3bb77dac),
	.w8(32'hbc1e671e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c6b85),
	.w1(32'hbc2a1f4a),
	.w2(32'hbbe81b08),
	.w3(32'hbce31ef0),
	.w4(32'hbc782679),
	.w5(32'hbbec9105),
	.w6(32'hbcea5470),
	.w7(32'hbc6853b4),
	.w8(32'hbaede3f1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd8c6),
	.w1(32'hbb36f8cb),
	.w2(32'h3c0c913b),
	.w3(32'hba04519e),
	.w4(32'hbb1f49bd),
	.w5(32'h3a953f16),
	.w6(32'h3b850681),
	.w7(32'h3bb31c7d),
	.w8(32'hbb74b9cd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83d08e),
	.w1(32'hbab275ae),
	.w2(32'hbc10aa9b),
	.w3(32'h3c1d7fce),
	.w4(32'hbb96ad66),
	.w5(32'hbc22faed),
	.w6(32'h3b9ecb6b),
	.w7(32'h3bcaa0c5),
	.w8(32'hbb2824a4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cc7c9),
	.w1(32'h3c10fb9a),
	.w2(32'h3b4377d7),
	.w3(32'hbbfb6eec),
	.w4(32'h3c09d19f),
	.w5(32'h39b7328f),
	.w6(32'hbba37be1),
	.w7(32'h3be0fb87),
	.w8(32'h3bd77f1c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb824769),
	.w1(32'h3c4d61d4),
	.w2(32'h3c04d750),
	.w3(32'hbcb5109f),
	.w4(32'h3b4f5e82),
	.w5(32'h3c9ed361),
	.w6(32'hbc6d0daa),
	.w7(32'h3ab1163e),
	.w8(32'h3c8aff2a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9e962),
	.w1(32'hbbb68aeb),
	.w2(32'h3b92d9c3),
	.w3(32'h3c816b11),
	.w4(32'h3b85efaf),
	.w5(32'h3bed9029),
	.w6(32'h3c578dac),
	.w7(32'h3c01b091),
	.w8(32'h3b8ef3cd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed1658),
	.w1(32'h3b15d2fa),
	.w2(32'hbbc8be39),
	.w3(32'h3b9424ce),
	.w4(32'h3acc99ee),
	.w5(32'hbc3e5c67),
	.w6(32'h3bff6baa),
	.w7(32'h3ba45592),
	.w8(32'hba99ef29),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b5912),
	.w1(32'hbb6c470b),
	.w2(32'hbc28c853),
	.w3(32'hbcc0b480),
	.w4(32'hbb96b127),
	.w5(32'hbc3448e1),
	.w6(32'hbc9770fd),
	.w7(32'h3b02e90a),
	.w8(32'hba439e5d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc412eff),
	.w1(32'h3c2119a3),
	.w2(32'hb9e5bf68),
	.w3(32'hbc8417a6),
	.w4(32'h3b5fe3a8),
	.w5(32'hba90de4f),
	.w6(32'hbc2c5160),
	.w7(32'h3b971043),
	.w8(32'h3add86b9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacea3e0),
	.w1(32'hba1c243b),
	.w2(32'hbc8ab9ba),
	.w3(32'h3b03f17f),
	.w4(32'h3b311ce7),
	.w5(32'hbbaf6918),
	.w6(32'h3bdd0683),
	.w7(32'h3b668a28),
	.w8(32'h3b715ae0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0e234),
	.w1(32'h3c3480d0),
	.w2(32'hbcaf55aa),
	.w3(32'hbc017658),
	.w4(32'h3c665132),
	.w5(32'hbc64da61),
	.w6(32'hbc0e2880),
	.w7(32'h3a94a789),
	.w8(32'hbc2ebe70),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc564547),
	.w1(32'hbc014c2f),
	.w2(32'h3cd05be3),
	.w3(32'hbc1993f0),
	.w4(32'hbb0d7c9b),
	.w5(32'h3d1fd19c),
	.w6(32'hbb6df809),
	.w7(32'hbaacb2ba),
	.w8(32'h3c9095b2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1293be),
	.w1(32'h3caad4fe),
	.w2(32'h3b65feb4),
	.w3(32'h3d7fb86e),
	.w4(32'h3d213f58),
	.w5(32'h3c8a0079),
	.w6(32'h3d442d60),
	.w7(32'h3d0c6350),
	.w8(32'h3bcd3f0f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c602fcc),
	.w1(32'h3b834b38),
	.w2(32'hbc02c9a8),
	.w3(32'h3d16597c),
	.w4(32'h3c892ef0),
	.w5(32'hbbb5e5f2),
	.w6(32'h3cd3f2ce),
	.w7(32'h3c2310a7),
	.w8(32'hbbf01b08),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8509b4),
	.w1(32'h3b1653d6),
	.w2(32'hbb92482a),
	.w3(32'h3b317b2a),
	.w4(32'h3b29f8c8),
	.w5(32'hbc76001e),
	.w6(32'h3a93f643),
	.w7(32'h3b444fa1),
	.w8(32'hbc28de4a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4af25e),
	.w1(32'hbc3e01cf),
	.w2(32'h3b65a3b0),
	.w3(32'hbc93f31a),
	.w4(32'hbc97e1ed),
	.w5(32'hbb233caf),
	.w6(32'hbc16a16f),
	.w7(32'hbb0a87ad),
	.w8(32'hbb4509f0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b533cfa),
	.w1(32'h3b66682c),
	.w2(32'hbd00b6c7),
	.w3(32'hbc05061e),
	.w4(32'h3c0b6a04),
	.w5(32'hbca7597a),
	.w6(32'hbbb1fabb),
	.w7(32'h3c6a90f5),
	.w8(32'hbc97e12b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca757ac),
	.w1(32'hbc44f60a),
	.w2(32'h3c282e40),
	.w3(32'hbcc66197),
	.w4(32'hbbd836d8),
	.w5(32'h3c3ff111),
	.w6(32'hbc7331f8),
	.w7(32'hbc51c309),
	.w8(32'h3c01440b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64013a),
	.w1(32'h3ba62704),
	.w2(32'hbb7a020b),
	.w3(32'h3c3f4890),
	.w4(32'h3c6e8eaa),
	.w5(32'hbb6a954b),
	.w6(32'h3c4159a7),
	.w7(32'h3c631b7c),
	.w8(32'h3b40d911),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd20a0),
	.w1(32'hbad916f9),
	.w2(32'hbb32ec50),
	.w3(32'hbb0391c4),
	.w4(32'h3b816f36),
	.w5(32'hbbc80c18),
	.w6(32'h3bee06a9),
	.w7(32'h3c210a04),
	.w8(32'hbc01da76),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf57b6c),
	.w1(32'h3a063bfd),
	.w2(32'h3b0ac482),
	.w3(32'hbc1575c7),
	.w4(32'hbb114feb),
	.w5(32'hbba0b906),
	.w6(32'hbbf1f794),
	.w7(32'hbb1fe738),
	.w8(32'h3b2ec787),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee6514),
	.w1(32'hbb4627a0),
	.w2(32'h3c78ac4d),
	.w3(32'hbc902895),
	.w4(32'hbc40dd01),
	.w5(32'h3cd47efb),
	.w6(32'hbc2c0f71),
	.w7(32'hbae2abf6),
	.w8(32'h3c830753),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad26e3),
	.w1(32'h3b33eb9e),
	.w2(32'h3c0583d1),
	.w3(32'h3cf62c17),
	.w4(32'h3c2f6744),
	.w5(32'h3b9c61a8),
	.w6(32'h3c8358a4),
	.w7(32'h3c32ea9c),
	.w8(32'h3bd13e85),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf751a1),
	.w1(32'hbbd24c02),
	.w2(32'hbad0779b),
	.w3(32'hb928f3df),
	.w4(32'hbba4b48c),
	.w5(32'h3a7a008f),
	.w6(32'h3b86f5da),
	.w7(32'hbb53416c),
	.w8(32'h3bc87c54),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3529dc),
	.w1(32'hb8aa0207),
	.w2(32'h3b120ff8),
	.w3(32'h3b530981),
	.w4(32'h39e6a757),
	.w5(32'hbb4b3d78),
	.w6(32'h3bf68bbf),
	.w7(32'h3b234c98),
	.w8(32'hba47a5c1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba26b1d),
	.w1(32'h3b667021),
	.w2(32'h3b9972ea),
	.w3(32'hb9e4c763),
	.w4(32'hb7b3655a),
	.w5(32'h3b973377),
	.w6(32'h3aa6af52),
	.w7(32'h3af5da49),
	.w8(32'h3be7f2ba),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed0655),
	.w1(32'hba76bf8d),
	.w2(32'h3b167a80),
	.w3(32'h3b41735f),
	.w4(32'hbc30f205),
	.w5(32'h3b9e0639),
	.w6(32'h3be78dbf),
	.w7(32'h3b75aa8c),
	.w8(32'h3ba26121),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b81d3),
	.w1(32'h3c96f5d1),
	.w2(32'hbc9649d0),
	.w3(32'h3cb83988),
	.w4(32'h3cc95f47),
	.w5(32'hbc60fe20),
	.w6(32'h3c8ed468),
	.w7(32'h3c07f17f),
	.w8(32'hbc056711),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7aa7),
	.w1(32'h3c236d08),
	.w2(32'hbc53d2f9),
	.w3(32'hbceff545),
	.w4(32'hbc253cc0),
	.w5(32'hbc545a3c),
	.w6(32'hbc5143ff),
	.w7(32'hbc5fe605),
	.w8(32'hbbd4d131),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf19ef),
	.w1(32'hbb476229),
	.w2(32'h3ae35012),
	.w3(32'hbc0db22a),
	.w4(32'hbc28c198),
	.w5(32'h3c0ce95b),
	.w6(32'hbbca4748),
	.w7(32'hbbaa364d),
	.w8(32'h3c08eac7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa21b4e),
	.w1(32'hbb134641),
	.w2(32'h3be0546a),
	.w3(32'h3c980c12),
	.w4(32'h3be25835),
	.w5(32'h3b910038),
	.w6(32'h3caad9ea),
	.w7(32'h3c00374d),
	.w8(32'h3b5b94c3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae1351),
	.w1(32'h3afc85f0),
	.w2(32'h3b21baf7),
	.w3(32'h3b1ba289),
	.w4(32'h3b53cc7a),
	.w5(32'h3a33db25),
	.w6(32'h3b34da99),
	.w7(32'h3b99bf55),
	.w8(32'h3b93d8a4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab232ad),
	.w1(32'h3a4b6457),
	.w2(32'hbc8ee61d),
	.w3(32'hb95100a7),
	.w4(32'h3b7a19a0),
	.w5(32'hbc8de736),
	.w6(32'h3b2b66fa),
	.w7(32'hbb2fffa5),
	.w8(32'hbc0e6da6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca331),
	.w1(32'h3b05e216),
	.w2(32'h3aa3af72),
	.w3(32'hbc9bf242),
	.w4(32'hbb95065c),
	.w5(32'h3be0a1ea),
	.w6(32'h3a8a3015),
	.w7(32'h3bc69649),
	.w8(32'h3b83e19b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a83f),
	.w1(32'h3b7f0c03),
	.w2(32'hba30e85a),
	.w3(32'h3c88c79a),
	.w4(32'h3c33e120),
	.w5(32'h3b3fc7fd),
	.w6(32'h3c927ea3),
	.w7(32'h3c831ad6),
	.w8(32'h392eaebd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980bd43),
	.w1(32'h3b9139c7),
	.w2(32'hba9f8ab3),
	.w3(32'hb93e86ee),
	.w4(32'h3bd8fac5),
	.w5(32'h3ac0f6e7),
	.w6(32'hbb3350e5),
	.w7(32'h3bb3f620),
	.w8(32'hbbce2550),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b183ceb),
	.w1(32'h3bae3f74),
	.w2(32'h3aebe238),
	.w3(32'h3b33b15d),
	.w4(32'hbaa798f0),
	.w5(32'h3bc70e4b),
	.w6(32'hba8dbd07),
	.w7(32'hbac38c94),
	.w8(32'h3bd319dd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a9b9a),
	.w1(32'hbbfcd4f9),
	.w2(32'h3bf8b7d3),
	.w3(32'hbbc1a2c8),
	.w4(32'hbc085b0e),
	.w5(32'h3c14ac77),
	.w6(32'h3acd9abd),
	.w7(32'hbbeeaa1b),
	.w8(32'h3c4de809),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23b1ac),
	.w1(32'h3c7548a3),
	.w2(32'h3a6f23f1),
	.w3(32'h3ccdfe53),
	.w4(32'h3c84c812),
	.w5(32'h3c57a0e4),
	.w6(32'h3ccbc69e),
	.w7(32'h3c4e82a2),
	.w8(32'h3bcbd03f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c961a71),
	.w1(32'h3c537ef0),
	.w2(32'hbb2da2da),
	.w3(32'h3d00d41d),
	.w4(32'h3ce9ce05),
	.w5(32'hbbbd9d4a),
	.w6(32'h3c995274),
	.w7(32'h3cdcc0e3),
	.w8(32'hbba4633f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39c703),
	.w1(32'hb9baf991),
	.w2(32'hbc91db41),
	.w3(32'hbb389fd7),
	.w4(32'hbba54ca8),
	.w5(32'hbc544af5),
	.w6(32'hbaacd18d),
	.w7(32'h3a7f2e48),
	.w8(32'hbbaaa635),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc874196),
	.w1(32'hbc2e2c88),
	.w2(32'hbc7bc8d5),
	.w3(32'hbc1698af),
	.w4(32'hbb4d95f2),
	.w5(32'hbbcbad8f),
	.w6(32'hbb8ffa8d),
	.w7(32'hb9c490d7),
	.w8(32'hbbed7246),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a8f7),
	.w1(32'hbb648ab0),
	.w2(32'hbc82cff5),
	.w3(32'h3c0970b3),
	.w4(32'hbc00864a),
	.w5(32'hbcb044a6),
	.w6(32'hbaaff8f1),
	.w7(32'hbb0ef91e),
	.w8(32'hbc6bad71),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab5949),
	.w1(32'hbc9001cb),
	.w2(32'h3c8c14a0),
	.w3(32'hbcba42ae),
	.w4(32'hbc8a5222),
	.w5(32'h3ce08e06),
	.w6(32'hbc7fc741),
	.w7(32'hbca4aa8f),
	.w8(32'h3c7221f8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccfcbd0),
	.w1(32'h3be867dd),
	.w2(32'hba16f8a1),
	.w3(32'h3d130d79),
	.w4(32'h3cb03bda),
	.w5(32'h3b8bda75),
	.w6(32'h3ce94b24),
	.w7(32'h3c861501),
	.w8(32'hba3bc779),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eb653),
	.w1(32'hbb4ed53c),
	.w2(32'h3b643a39),
	.w3(32'h3ac8ae76),
	.w4(32'h39b8f9d3),
	.w5(32'hb8dae8bf),
	.w6(32'hbb0ccbd8),
	.w7(32'hbb867def),
	.w8(32'hbb589dd7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d2250),
	.w1(32'hbb599a92),
	.w2(32'hbc15a822),
	.w3(32'h3b9af90b),
	.w4(32'hbb89035e),
	.w5(32'hbbdc0417),
	.w6(32'h3ab3ea88),
	.w7(32'hbafb865c),
	.w8(32'hbb738f03),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b193b),
	.w1(32'hbb871880),
	.w2(32'h3c4dc487),
	.w3(32'hbad2325a),
	.w4(32'hba2949d5),
	.w5(32'h3c7c9ce9),
	.w6(32'h3b21a50b),
	.w7(32'hb98f2927),
	.w8(32'h3bfdf334),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21b7b0),
	.w1(32'h3bfe15f6),
	.w2(32'h3c878ac4),
	.w3(32'h3c3f9f23),
	.w4(32'h3acd3e75),
	.w5(32'h3c94521e),
	.w6(32'h3c4cd7e3),
	.w7(32'hbb3d93c9),
	.w8(32'h3c72a5e3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03a66b),
	.w1(32'h3cbab197),
	.w2(32'h3c64804e),
	.w3(32'h3d48c2bb),
	.w4(32'h3d03e124),
	.w5(32'h3cbed4dc),
	.w6(32'h3d0aa230),
	.w7(32'h3ceade2d),
	.w8(32'h3c173beb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e11db),
	.w1(32'h3c319b65),
	.w2(32'hbbc91dab),
	.w3(32'h3ce380f5),
	.w4(32'h3cd1976e),
	.w5(32'hbbc3ebc8),
	.w6(32'h3ccb2307),
	.w7(32'h3c7ad87e),
	.w8(32'hbb8d6cc9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06910f),
	.w1(32'h3bc9d435),
	.w2(32'hbbc46f4b),
	.w3(32'hbc19f6fe),
	.w4(32'h37d47695),
	.w5(32'hbba2ebc6),
	.w6(32'hbc4660d2),
	.w7(32'h389910bc),
	.w8(32'hbb430120),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbba11d),
	.w1(32'hbb1267f1),
	.w2(32'hb95901e5),
	.w3(32'hbc01ec51),
	.w4(32'hbb747a79),
	.w5(32'hba89c5d1),
	.w6(32'hbbfb6528),
	.w7(32'hbbcaa165),
	.w8(32'hba1b239b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89dea3),
	.w1(32'h3a1e65bd),
	.w2(32'h3c193de4),
	.w3(32'h39b6cb20),
	.w4(32'h3a9ecdd8),
	.w5(32'h3bd93eb4),
	.w6(32'h3ae35a2a),
	.w7(32'h3b6bd6bf),
	.w8(32'h3b076796),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ff774),
	.w1(32'h3b955f89),
	.w2(32'hbbfeed22),
	.w3(32'hbc0c72a1),
	.w4(32'h3b7ad4cb),
	.w5(32'hbcab57ca),
	.w6(32'h3b4a9c08),
	.w7(32'h3c76c7a6),
	.w8(32'hbc8721f4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d3313),
	.w1(32'hbc169fe1),
	.w2(32'h3aeb89d2),
	.w3(32'hbd08a684),
	.w4(32'hbcb10fcf),
	.w5(32'h3b280f0d),
	.w6(32'hbcc4746e),
	.w7(32'hbc1be6ff),
	.w8(32'h3b0adbd7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad491),
	.w1(32'h3b9971a9),
	.w2(32'h3c56387a),
	.w3(32'h3ba53cf7),
	.w4(32'h3c14edc5),
	.w5(32'h3c5a2f54),
	.w6(32'h3bbad116),
	.w7(32'h3c168b05),
	.w8(32'h3c15e306),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3912da),
	.w1(32'h3b46261a),
	.w2(32'hbbb6ac8a),
	.w3(32'h3cb7d43a),
	.w4(32'h3bcaa7de),
	.w5(32'hba58d2d2),
	.w6(32'h3c86ed09),
	.w7(32'h3a701ff6),
	.w8(32'hbad76707),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27aec4),
	.w1(32'h3ad18998),
	.w2(32'h3b455c00),
	.w3(32'hb9ea4660),
	.w4(32'h3b044132),
	.w5(32'h3ba1a460),
	.w6(32'h3a9177a3),
	.w7(32'h3b6208ed),
	.w8(32'h3b6533fd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab77b0),
	.w1(32'hbb0cff5e),
	.w2(32'h3bb13452),
	.w3(32'h3be6c090),
	.w4(32'h3a902a2e),
	.w5(32'h3c534ae6),
	.w6(32'h3bd045d9),
	.w7(32'hba917337),
	.w8(32'h3b2c0912),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14eba5),
	.w1(32'h3c09021b),
	.w2(32'hbb00eab3),
	.w3(32'h3c7e6864),
	.w4(32'h3bc9c64c),
	.w5(32'hbb8cbdb0),
	.w6(32'h3c3f299b),
	.w7(32'h3c044d6f),
	.w8(32'h3b944a30),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b32f3),
	.w1(32'hbc148e92),
	.w2(32'hbb2ce4a1),
	.w3(32'hbc9f7f3f),
	.w4(32'hbc99bd69),
	.w5(32'hbc54a455),
	.w6(32'hb9af7171),
	.w7(32'h3bf446e6),
	.w8(32'h3aa4f8ae),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fa2c8),
	.w1(32'hbc279efb),
	.w2(32'hbc6fbe2b),
	.w3(32'hbcb7692c),
	.w4(32'hbc3927cb),
	.w5(32'hbc1feb77),
	.w6(32'hbbf81058),
	.w7(32'h3b39ee56),
	.w8(32'hbb585514),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31a34f),
	.w1(32'hbb305559),
	.w2(32'hbc9c63d1),
	.w3(32'hbc421f46),
	.w4(32'hbbd15c02),
	.w5(32'hbd334323),
	.w6(32'hbc7d3f11),
	.w7(32'hbc45b9cf),
	.w8(32'hbcfe7bc8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7ce24),
	.w1(32'hbcefc50d),
	.w2(32'hbbe8627e),
	.w3(32'hbd623bac),
	.w4(32'hbd19e0dd),
	.w5(32'hbafd4aeb),
	.w6(32'hbd2ff987),
	.w7(32'hbcd4c164),
	.w8(32'hbb523170),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be5b2),
	.w1(32'h3b0e9bde),
	.w2(32'h3bdcd56f),
	.w3(32'h3c121915),
	.w4(32'h3c015acd),
	.w5(32'h3c85f67c),
	.w6(32'h3c107eeb),
	.w7(32'h3c3f3e01),
	.w8(32'h3ca6de80),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8aed76),
	.w1(32'h3c2dcc0b),
	.w2(32'h3c2c927e),
	.w3(32'h3cabe54e),
	.w4(32'h3cbb567e),
	.w5(32'h3c457451),
	.w6(32'h3c6f5343),
	.w7(32'h3c913784),
	.w8(32'h3be65d89),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c061d25),
	.w1(32'h3be64fce),
	.w2(32'hb78f3a1d),
	.w3(32'h3ca1dc03),
	.w4(32'h3c42f280),
	.w5(32'hbb829ba9),
	.w6(32'h3c01db26),
	.w7(32'h3c8c47a2),
	.w8(32'h39fee931),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb011301),
	.w1(32'hbb65fa0d),
	.w2(32'hbc3a8569),
	.w3(32'h3af153aa),
	.w4(32'h3aaf081f),
	.w5(32'hbc4a39b8),
	.w6(32'h3b111d6e),
	.w7(32'h3b876650),
	.w8(32'hbc070935),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79403d),
	.w1(32'h3b27e46f),
	.w2(32'h3c80cfef),
	.w3(32'hbc095303),
	.w4(32'hbc068138),
	.w5(32'h3c8919b7),
	.w6(32'hbbeac9db),
	.w7(32'hbb7983f2),
	.w8(32'h3bed7fe0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb48bc3),
	.w1(32'hb9b66883),
	.w2(32'hbbb355e5),
	.w3(32'h3cbe6cf2),
	.w4(32'h3c7747ad),
	.w5(32'hbc43c177),
	.w6(32'h3c9ae6c3),
	.w7(32'h3c759e1e),
	.w8(32'hbbbecfce),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4586de),
	.w1(32'hbbcc73c5),
	.w2(32'h3a9c8d1e),
	.w3(32'hb9951ae5),
	.w4(32'hbbc8afa5),
	.w5(32'hbb27cdf1),
	.w6(32'h3bc98c5d),
	.w7(32'h3b9ee0d4),
	.w8(32'hbba9d2e5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881aea),
	.w1(32'hbb8fd9a8),
	.w2(32'h3b5250ee),
	.w3(32'h3bd9e46a),
	.w4(32'hbb9fcd5b),
	.w5(32'h3bdfb90c),
	.w6(32'h3ba0e5e9),
	.w7(32'hb900bb22),
	.w8(32'h3bc44296),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45a5d1),
	.w1(32'hbc278a0d),
	.w2(32'h3c52e4a9),
	.w3(32'h3b589e3c),
	.w4(32'hbbb72459),
	.w5(32'h3cc83753),
	.w6(32'h3b88f88f),
	.w7(32'h3b6c713d),
	.w8(32'h3c8aa876),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f6e77),
	.w1(32'hbb8f6ac2),
	.w2(32'hbc3147f5),
	.w3(32'h3cdfca13),
	.w4(32'h3b924521),
	.w5(32'hbc9ec54a),
	.w6(32'h3ca0897f),
	.w7(32'h3c5335fc),
	.w8(32'hbc0592ee),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93177f),
	.w1(32'hbc01ec79),
	.w2(32'hbc85fd40),
	.w3(32'hbcdf7885),
	.w4(32'hbc530fe0),
	.w5(32'hbc0b6fad),
	.w6(32'hbc80216b),
	.w7(32'hbb95802a),
	.w8(32'h3b9011e5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc075d55),
	.w1(32'h3bcdb0b3),
	.w2(32'h3c0b0fc7),
	.w3(32'hbcafd503),
	.w4(32'h3b2673f5),
	.w5(32'h3bf6c02e),
	.w6(32'hbca03a99),
	.w7(32'hbc084ecd),
	.w8(32'hb9270564),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34126d),
	.w1(32'hbb786775),
	.w2(32'h397054d7),
	.w3(32'h3c69073d),
	.w4(32'hbb6c1a8c),
	.w5(32'hbc87834f),
	.w6(32'h3b9bd339),
	.w7(32'hbadaf4db),
	.w8(32'hbb8ce56d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f7bd),
	.w1(32'h37e4f40c),
	.w2(32'hbc121611),
	.w3(32'hbc7bedc8),
	.w4(32'hbc40b4de),
	.w5(32'hbc23cc24),
	.w6(32'hbc869e0b),
	.w7(32'hbb74bf5a),
	.w8(32'hbbc0487d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57b261),
	.w1(32'hbc84d346),
	.w2(32'h3b06270f),
	.w3(32'hbc81a300),
	.w4(32'hbb99409a),
	.w5(32'hbc476f78),
	.w6(32'hbba182c8),
	.w7(32'hbbe0e0ff),
	.w8(32'hbc050058),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33e834),
	.w1(32'hbc26ea48),
	.w2(32'h3b2d4646),
	.w3(32'hbcb824c0),
	.w4(32'hbc538508),
	.w5(32'h3c07885d),
	.w6(32'hbc3e2895),
	.w7(32'hbc0a0fb2),
	.w8(32'h3bf9c2a5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b445eb6),
	.w1(32'hb9ece171),
	.w2(32'h3c03e99c),
	.w3(32'h3c2063df),
	.w4(32'h3bd343ca),
	.w5(32'h3bc61aca),
	.w6(32'h3c26e3a3),
	.w7(32'h3c0afa0f),
	.w8(32'h3b351dfc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd373e5),
	.w1(32'h3b56643a),
	.w2(32'hbafecf3d),
	.w3(32'h3bd33a45),
	.w4(32'h3b87a6ca),
	.w5(32'hbb7f5df6),
	.w6(32'h3b94df77),
	.w7(32'h3b8efe5c),
	.w8(32'h3b8abec6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374e9018),
	.w1(32'h3b0fd682),
	.w2(32'hbcb63762),
	.w3(32'hbb1373b4),
	.w4(32'hb9a4d233),
	.w5(32'hbcdff3ed),
	.w6(32'h3bc26932),
	.w7(32'h3c3ae8e6),
	.w8(32'hbc90fad0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc06b27),
	.w1(32'hbc50f141),
	.w2(32'h3bfa2fa2),
	.w3(32'hbd03dbf9),
	.w4(32'hbcfb0e2f),
	.w5(32'h3c9d9649),
	.w6(32'hbc910036),
	.w7(32'hbcacb9af),
	.w8(32'h3c329297),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4436c8),
	.w1(32'h3c2af313),
	.w2(32'hbb3f8afe),
	.w3(32'h3d0008f1),
	.w4(32'h3cc841f3),
	.w5(32'hb9d19045),
	.w6(32'h3cbb2d6a),
	.w7(32'h3cc12681),
	.w8(32'h3bd4a742),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcebd20),
	.w1(32'h3ba092f5),
	.w2(32'hb92649eb),
	.w3(32'hbcc8d676),
	.w4(32'hbbdb8419),
	.w5(32'h38a085c6),
	.w6(32'hbc3f7549),
	.w7(32'hbc0bcb36),
	.w8(32'hba44ca26),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a0417),
	.w1(32'hba0460dd),
	.w2(32'hbbb66db6),
	.w3(32'h3a5216c5),
	.w4(32'hbb28460f),
	.w5(32'hbb430d31),
	.w6(32'h3b232bd8),
	.w7(32'hbb0e2317),
	.w8(32'hbaf53e62),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe93db9),
	.w1(32'h3b038fe0),
	.w2(32'h3c008d7a),
	.w3(32'hbbebabd3),
	.w4(32'h3b0f1eb3),
	.w5(32'h3c2d25c3),
	.w6(32'hbbc58135),
	.w7(32'h3b098468),
	.w8(32'h3b3ed74c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23a78f),
	.w1(32'hbb3ba825),
	.w2(32'h3b331937),
	.w3(32'h3c24fce2),
	.w4(32'h3bb9749e),
	.w5(32'h3a9a1e43),
	.w6(32'h3c099670),
	.w7(32'hbac3ebf3),
	.w8(32'h3b535053),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81518b),
	.w1(32'h3bb2725a),
	.w2(32'hbca0fbe2),
	.w3(32'h3b8be04f),
	.w4(32'h3b09bdc6),
	.w5(32'hbc6f3ed3),
	.w6(32'h3b2364c4),
	.w7(32'h376c5421),
	.w8(32'hbc557800),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8772c9),
	.w1(32'hbc152beb),
	.w2(32'hbc14cab7),
	.w3(32'hbcfd4306),
	.w4(32'hbc7ee8c2),
	.w5(32'hbba05e5f),
	.w6(32'hbcb22168),
	.w7(32'hbbea4f52),
	.w8(32'hbb46f01a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35f82e),
	.w1(32'h3bf551b1),
	.w2(32'hbc2b1cb8),
	.w3(32'hbbb41147),
	.w4(32'hb9401cdd),
	.w5(32'hbc2ad065),
	.w6(32'hbbfe871c),
	.w7(32'hba8fb715),
	.w8(32'hbbe61e05),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03576b),
	.w1(32'hbc064b7d),
	.w2(32'hbb6ec113),
	.w3(32'hbc838b8f),
	.w4(32'hbc886b06),
	.w5(32'h3c2c6e35),
	.w6(32'hbafbc525),
	.w7(32'h3b8f4567),
	.w8(32'h3c3517bd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c6fa),
	.w1(32'h3c2283a1),
	.w2(32'h3b1c726d),
	.w3(32'h3c9d8d36),
	.w4(32'h3c4cd89e),
	.w5(32'h3cb00ab2),
	.w6(32'h3c502bf2),
	.w7(32'h3c060b70),
	.w8(32'h3c8e27a1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09ed7b),
	.w1(32'hbbe7eb6d),
	.w2(32'hbc520316),
	.w3(32'h3b29baf9),
	.w4(32'hbc3f5680),
	.w5(32'hbb882cab),
	.w6(32'h3c8056cb),
	.w7(32'hbbad8eff),
	.w8(32'hbb8ad9f3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30be2d),
	.w1(32'hbb22f4ce),
	.w2(32'h3c0f2537),
	.w3(32'hbc20b55e),
	.w4(32'h3b568d4d),
	.w5(32'h3bcbb35b),
	.w6(32'hbc0c386c),
	.w7(32'hbc81a31a),
	.w8(32'h3b89eb82),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b2988),
	.w1(32'h3c887e1c),
	.w2(32'hbc363007),
	.w3(32'h3bf97306),
	.w4(32'h3c67b543),
	.w5(32'hbc823712),
	.w6(32'h3ba9ed8c),
	.w7(32'h3b840075),
	.w8(32'hbbc8bf98),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9908db),
	.w1(32'hbc7aed21),
	.w2(32'hbc157517),
	.w3(32'hbc966843),
	.w4(32'hbc4b4a42),
	.w5(32'hbac130b2),
	.w6(32'hbbd1e894),
	.w7(32'hbc450a60),
	.w8(32'hbb6eb120),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc230077),
	.w1(32'h3ab840c1),
	.w2(32'hbc01608b),
	.w3(32'hbc121b8c),
	.w4(32'h39ae1f10),
	.w5(32'hbc02e954),
	.w6(32'hbc92ab0c),
	.w7(32'hb6b77ff8),
	.w8(32'hbb8f0b24),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a496f76),
	.w1(32'hbc1170fc),
	.w2(32'hbbf7f648),
	.w3(32'h3b056f24),
	.w4(32'hbbf8590d),
	.w5(32'hbc4517c2),
	.w6(32'h3b67ec09),
	.w7(32'hbb901594),
	.w8(32'hbb9d97f4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ac3eb),
	.w1(32'h3c2ec07c),
	.w2(32'h3bc0aa83),
	.w3(32'hbb6a4a85),
	.w4(32'h3be573b3),
	.w5(32'h3aec7865),
	.w6(32'h3b34cbda),
	.w7(32'h3c518843),
	.w8(32'h3b716391),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a9f8b),
	.w1(32'hbba18ad2),
	.w2(32'hbafd81d1),
	.w3(32'h3bb8a464),
	.w4(32'h3ac1855c),
	.w5(32'h3bb6b7c1),
	.w6(32'h3b3fa90e),
	.w7(32'h3b8e8080),
	.w8(32'h3b5d7d7c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb470a73),
	.w1(32'hbc0b856d),
	.w2(32'hbbaa8212),
	.w3(32'h3c1f80ed),
	.w4(32'hbb4d60aa),
	.w5(32'hbafc9389),
	.w6(32'h3bb40275),
	.w7(32'hbb33964f),
	.w8(32'hbae741c5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3aa0c7),
	.w1(32'h3b5b98ca),
	.w2(32'h3c0130d9),
	.w3(32'h3b927ad1),
	.w4(32'h3bab16c7),
	.w5(32'h3bd458f8),
	.w6(32'h3bb8a8b6),
	.w7(32'h3bc3d2a3),
	.w8(32'h3c14085d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae5af4),
	.w1(32'h3c7f8dd5),
	.w2(32'hbc013c14),
	.w3(32'h3c52b797),
	.w4(32'h3c9db302),
	.w5(32'hbbb61c66),
	.w6(32'h3bc1e0d4),
	.w7(32'h3c226561),
	.w8(32'hbc28a304),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2160a6),
	.w1(32'hbbb157ac),
	.w2(32'h3bcc9106),
	.w3(32'hbb833859),
	.w4(32'hbbb3e2cd),
	.w5(32'h3bbfb66d),
	.w6(32'hbbae13b0),
	.w7(32'hbba9f4a0),
	.w8(32'h3ada80bf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaa15a),
	.w1(32'h3b5b78fa),
	.w2(32'h3b2c52e9),
	.w3(32'h3bfeb281),
	.w4(32'h3c4c2bed),
	.w5(32'h3b86e85a),
	.w6(32'h3bdbcc66),
	.w7(32'h3bb35a03),
	.w8(32'h3b80d2ed),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb78b03),
	.w1(32'h3b12cc12),
	.w2(32'hba524a0a),
	.w3(32'hb9223188),
	.w4(32'h3b6df28b),
	.w5(32'hbb1eff50),
	.w6(32'hbb0158f1),
	.w7(32'h3c24bf5a),
	.w8(32'h396a2d84),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb173a9b),
	.w1(32'hbae94f41),
	.w2(32'hbb14e43e),
	.w3(32'hb96b7edd),
	.w4(32'hbbbdf06a),
	.w5(32'hbab8eed7),
	.w6(32'h3bd17183),
	.w7(32'h3bdf690a),
	.w8(32'hbb1be6e5),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fda12),
	.w1(32'hbabc56f9),
	.w2(32'hbc319b48),
	.w3(32'h3ad7442c),
	.w4(32'h39befcf1),
	.w5(32'hbbb63b4c),
	.w6(32'h3a0a3e11),
	.w7(32'hbb02ff74),
	.w8(32'hbbb02739),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd15a1),
	.w1(32'hb923c813),
	.w2(32'hba877822),
	.w3(32'hbc00e9e0),
	.w4(32'hbb7de663),
	.w5(32'h3c024652),
	.w6(32'hbc23eaa3),
	.w7(32'hbc067fa5),
	.w8(32'h3b06ae50),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14b722),
	.w1(32'h3ac488da),
	.w2(32'hba19334a),
	.w3(32'hbb6b4bdb),
	.w4(32'h3b9bf536),
	.w5(32'h3b48ed0c),
	.w6(32'hbab22864),
	.w7(32'hbb8571a8),
	.w8(32'h3bda766e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c4031),
	.w1(32'hbb1f47f6),
	.w2(32'hbb8f39c8),
	.w3(32'hbbd0a8ab),
	.w4(32'h3a9c189b),
	.w5(32'hbba844b2),
	.w6(32'hbc0a5784),
	.w7(32'h3b0fce78),
	.w8(32'hbbbff1e8),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3d3ba),
	.w1(32'hbb14c90c),
	.w2(32'hbc4c2d9f),
	.w3(32'hbb0bef8a),
	.w4(32'hbbd9e25f),
	.w5(32'hbc37b845),
	.w6(32'hbba2523f),
	.w7(32'hbb9ba26c),
	.w8(32'h3aa7af65),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70d45d),
	.w1(32'hbc4954c7),
	.w2(32'hbb55b6d9),
	.w3(32'hbc8b45c4),
	.w4(32'hbb7f7b4b),
	.w5(32'hbb20671b),
	.w6(32'hbc386b4a),
	.w7(32'hbc5182d9),
	.w8(32'hbb12c33e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef3504),
	.w1(32'hbb9e0195),
	.w2(32'hba5ebdda),
	.w3(32'h3c6d8775),
	.w4(32'h3c3ba98e),
	.w5(32'h3af46c5a),
	.w6(32'h3b49415d),
	.w7(32'h3c2a8e11),
	.w8(32'h3a0ddb9b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b132cfd),
	.w1(32'h3aa515d2),
	.w2(32'h3bb692df),
	.w3(32'h3be332b8),
	.w4(32'h3b3ae8fa),
	.w5(32'h3c8f98b6),
	.w6(32'h3b9d180e),
	.w7(32'h3b3d678d),
	.w8(32'h3c01890f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a3f24),
	.w1(32'h3c28ef84),
	.w2(32'hbc203877),
	.w3(32'h3c5bc283),
	.w4(32'h3c529977),
	.w5(32'hba861f21),
	.w6(32'h3c6a8fdf),
	.w7(32'h3b9b2777),
	.w8(32'hbb1b2b91),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6de1f2),
	.w1(32'hbba2b50a),
	.w2(32'hb9ca0e79),
	.w3(32'hbc24ec36),
	.w4(32'hbc3459e1),
	.w5(32'hbb1ba17f),
	.w6(32'hbc4f564b),
	.w7(32'h3913d5df),
	.w8(32'hbb109312),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ef52a),
	.w1(32'hbbaadd35),
	.w2(32'h3b32d691),
	.w3(32'h3b5eba6c),
	.w4(32'hbb4d0032),
	.w5(32'hbb5b0df8),
	.w6(32'h3b70ff0d),
	.w7(32'hbb4e50ef),
	.w8(32'h3b0a7b03),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9266b2),
	.w1(32'h3b3c4a45),
	.w2(32'hbc71280f),
	.w3(32'hba360370),
	.w4(32'hbb2dc3ef),
	.w5(32'hbc7d6eb3),
	.w6(32'h3a3e55bb),
	.w7(32'h3a969250),
	.w8(32'hbc4e87a0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73c1e7),
	.w1(32'hbbf70d4b),
	.w2(32'hbc33bbaf),
	.w3(32'h3b2bdc22),
	.w4(32'hbb65c2bc),
	.w5(32'h3a2a108d),
	.w6(32'h3a620926),
	.w7(32'hbba0b366),
	.w8(32'h3b442c5a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68d259),
	.w1(32'hbc79df4b),
	.w2(32'hbab3287f),
	.w3(32'h393dcbc4),
	.w4(32'hbb19dc90),
	.w5(32'hbadf2261),
	.w6(32'h3be87452),
	.w7(32'h3bb7c65e),
	.w8(32'hba9e373e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fe202),
	.w1(32'hbb443a37),
	.w2(32'h3bbcea74),
	.w3(32'hb9bd5cf7),
	.w4(32'hbaaa3fc0),
	.w5(32'h3c88edca),
	.w6(32'hbaabcd1d),
	.w7(32'hbb453724),
	.w8(32'h3c2bcb7c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bffdd),
	.w1(32'h3c4160b3),
	.w2(32'h3b6c2acf),
	.w3(32'h3cd31f3c),
	.w4(32'h3c8dbd2e),
	.w5(32'h3bb68f16),
	.w6(32'h3caf9926),
	.w7(32'h3c70c40a),
	.w8(32'h3bf20526),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c339d48),
	.w1(32'h3a25af9d),
	.w2(32'hbbabd731),
	.w3(32'h3c6475f6),
	.w4(32'h3c8d78d6),
	.w5(32'hbb2afef9),
	.w6(32'h3c535eda),
	.w7(32'h3b756450),
	.w8(32'hbbbcacac),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b3047),
	.w1(32'hbb8c5cd6),
	.w2(32'h3b306c4a),
	.w3(32'h3a1bd52f),
	.w4(32'h3b283002),
	.w5(32'h3c41d0fa),
	.w6(32'hbb2cd3aa),
	.w7(32'hbb3eb8ce),
	.w8(32'h3b75dfd2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bdc93),
	.w1(32'hbbf9cd35),
	.w2(32'hbb9b5a54),
	.w3(32'hbbfcd250),
	.w4(32'hbc7111ec),
	.w5(32'hbb2a4d61),
	.w6(32'hbb54a11f),
	.w7(32'hbc3954b4),
	.w8(32'hbb9bdca6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1101fe),
	.w1(32'hb9981a3a),
	.w2(32'hbcc52007),
	.w3(32'hba719a00),
	.w4(32'h3b32f0fe),
	.w5(32'hbb55a082),
	.w6(32'hba63939d),
	.w7(32'h3af20216),
	.w8(32'h3bb61a5d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb001de),
	.w1(32'hbca13a88),
	.w2(32'hbc711707),
	.w3(32'hbb242628),
	.w4(32'hbb7809dd),
	.w5(32'hbb863b4d),
	.w6(32'h3c93d5de),
	.w7(32'h3c804da2),
	.w8(32'hbc059045),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb19cb),
	.w1(32'hbb38f32c),
	.w2(32'h3be768ee),
	.w3(32'h3c3af903),
	.w4(32'h3c7538fb),
	.w5(32'h3bdfc6ce),
	.w6(32'h3bc6b10c),
	.w7(32'h3c0113ee),
	.w8(32'h3c371b18),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a562da),
	.w1(32'hba1e4eee),
	.w2(32'hbb903038),
	.w3(32'h3c627afe),
	.w4(32'h3bf1ba61),
	.w5(32'hbc147bda),
	.w6(32'h3c5d8b14),
	.w7(32'h3c65ebf8),
	.w8(32'hbaaf4863),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510047),
	.w1(32'h3b8d22f0),
	.w2(32'h399306b1),
	.w3(32'h3c0d9a31),
	.w4(32'h3c507056),
	.w5(32'hba721c1b),
	.w6(32'h3c107929),
	.w7(32'h3c443db4),
	.w8(32'h3b479732),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a2568),
	.w1(32'h3b4f3990),
	.w2(32'h3bbb1ca1),
	.w3(32'h3baec06c),
	.w4(32'h3b7e7749),
	.w5(32'h3c267dfd),
	.w6(32'h3c55d6a8),
	.w7(32'h3c508044),
	.w8(32'h3b06d389),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7d792),
	.w1(32'h3c3a4af6),
	.w2(32'hba282e78),
	.w3(32'h3c7e3c0d),
	.w4(32'h3c854b08),
	.w5(32'h3c5c4da5),
	.w6(32'h3bd9143c),
	.w7(32'h3b60b47c),
	.w8(32'h3b8523a1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba44eea),
	.w1(32'h3bc7c017),
	.w2(32'hbbc08e0c),
	.w3(32'h3c9065e8),
	.w4(32'h3c51bd0c),
	.w5(32'hb991b8bc),
	.w6(32'h3cc76d54),
	.w7(32'h3c8ed868),
	.w8(32'hba93b715),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68d90b),
	.w1(32'hbb457f41),
	.w2(32'hbc0efb01),
	.w3(32'h3b7abc3c),
	.w4(32'h3b021c52),
	.w5(32'hbba0333b),
	.w6(32'h3b95f14d),
	.w7(32'h3b9b928b),
	.w8(32'h3bc0da65),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f93f),
	.w1(32'h3b5a5d9f),
	.w2(32'hbc41d010),
	.w3(32'h3b277c1a),
	.w4(32'h3a0ba4ff),
	.w5(32'hbbafc935),
	.w6(32'h3c17e658),
	.w7(32'h3b687f70),
	.w8(32'hba87534e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21fb89),
	.w1(32'hbc2807c5),
	.w2(32'hbd17dce2),
	.w3(32'h3b3d453d),
	.w4(32'h3b12f6da),
	.w5(32'hbd3ecca6),
	.w6(32'h3beab6cd),
	.w7(32'h3b4f1350),
	.w8(32'hbce1923e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd30a107),
	.w1(32'hbce33ddf),
	.w2(32'hba944d71),
	.w3(32'hbd80a32a),
	.w4(32'hbd511936),
	.w5(32'h3c067c95),
	.w6(32'hbd3bbde6),
	.w7(32'hbd1d6bb8),
	.w8(32'h3ae29196),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81d3e2a),
	.w1(32'h3a8a074d),
	.w2(32'hbb86f199),
	.w3(32'h3adc95f7),
	.w4(32'hbb063ac4),
	.w5(32'hba1133af),
	.w6(32'h3c863062),
	.w7(32'h3c0ca322),
	.w8(32'hbb25b06b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57e13a),
	.w1(32'h3b18df54),
	.w2(32'hbbb78dd9),
	.w3(32'h3b53f771),
	.w4(32'h3bc2ced0),
	.w5(32'hbbb3becb),
	.w6(32'h3acd7064),
	.w7(32'h3bd046c8),
	.w8(32'hbb978c2b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9678b7),
	.w1(32'h3bbda415),
	.w2(32'hbb0a5f93),
	.w3(32'h3abbf8df),
	.w4(32'h393c6fa5),
	.w5(32'hbcc7bc9f),
	.w6(32'hbc2b3519),
	.w7(32'h390b8b85),
	.w8(32'hbcc6b4f2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb94117),
	.w1(32'hbce094cd),
	.w2(32'hbb87ece0),
	.w3(32'hbd3f47b9),
	.w4(32'hbd1602cf),
	.w5(32'hbc26fb68),
	.w6(32'hbcddbb90),
	.w7(32'hbc706ad0),
	.w8(32'hbb140372),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf45e1b),
	.w1(32'hbc3ec994),
	.w2(32'h3b76e3b6),
	.w3(32'hbbe3687a),
	.w4(32'hba054566),
	.w5(32'hbc21a32d),
	.w6(32'h3bebb0a7),
	.w7(32'h3b855f0b),
	.w8(32'hbc36fd41),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67234c),
	.w1(32'hbc7fbffe),
	.w2(32'hbb6ba2c4),
	.w3(32'hbcf83347),
	.w4(32'hbc9e575a),
	.w5(32'h3b52b730),
	.w6(32'hbc9edb58),
	.w7(32'hbbe3afe3),
	.w8(32'hbc134e30),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3811b),
	.w1(32'hbadad90f),
	.w2(32'hbbbefd80),
	.w3(32'h3c209915),
	.w4(32'h3b222a9b),
	.w5(32'h3b44e970),
	.w6(32'hbb1899ea),
	.w7(32'hbc11a58a),
	.w8(32'h3c01c5c9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41fdd3),
	.w1(32'h3a152dae),
	.w2(32'h393de92a),
	.w3(32'h3b8dc889),
	.w4(32'h3b10570a),
	.w5(32'h3b770dc2),
	.w6(32'h3c862ced),
	.w7(32'h3be69b31),
	.w8(32'h3bdaa7f1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54067),
	.w1(32'hbb65f2ca),
	.w2(32'hbbcf06c4),
	.w3(32'h3b6d045b),
	.w4(32'h3b0ccd32),
	.w5(32'hbca16264),
	.w6(32'h3c3b16c1),
	.w7(32'h3b6bdaea),
	.w8(32'hbb6c2c5c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb162d67),
	.w1(32'h3b3bd235),
	.w2(32'hbcb2a383),
	.w3(32'hbc071dbf),
	.w4(32'hbbd05807),
	.w5(32'hbc2b80f9),
	.w6(32'hbbdf2833),
	.w7(32'hbbb3a21c),
	.w8(32'hbc0e72f6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a453),
	.w1(32'hbc081560),
	.w2(32'hbc097c65),
	.w3(32'h3ac7356d),
	.w4(32'h3be23b21),
	.w5(32'hbbc4061a),
	.w6(32'h3bb7917c),
	.w7(32'h3c244ab3),
	.w8(32'h3b79e681),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07902e),
	.w1(32'h3c856aff),
	.w2(32'hbb491157),
	.w3(32'hbb00e9f6),
	.w4(32'h3cc95b08),
	.w5(32'hbac4e0d2),
	.w6(32'h3b7addae),
	.w7(32'h3d02afb9),
	.w8(32'h3a55b846),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c45741),
	.w1(32'hbbe7b0e8),
	.w2(32'hbcb26d67),
	.w3(32'h3c0d11d7),
	.w4(32'h39eb91cf),
	.w5(32'hbc80b25a),
	.w6(32'h3c7212f3),
	.w7(32'h3c02090b),
	.w8(32'hbc546564),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90b4cd),
	.w1(32'hbb730e3e),
	.w2(32'hbc60ba9d),
	.w3(32'h3b923743),
	.w4(32'h3b95d134),
	.w5(32'hbbd7562a),
	.w6(32'hbaca28f9),
	.w7(32'h3b0bd7cc),
	.w8(32'hbaa2711c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6abf44),
	.w1(32'hbc00dd17),
	.w2(32'h3b701121),
	.w3(32'hbc8db445),
	.w4(32'hbbcb81ef),
	.w5(32'h3c360301),
	.w6(32'hbaa0a932),
	.w7(32'hbaa068b0),
	.w8(32'h3c413221),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c358d),
	.w1(32'h3bc2c2c8),
	.w2(32'hba4e67b1),
	.w3(32'h3bfdf6ef),
	.w4(32'h3c0e4615),
	.w5(32'hbb42f15b),
	.w6(32'h3c6db46a),
	.w7(32'h3c465036),
	.w8(32'hbbfbc5d0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8eac5),
	.w1(32'h3b768d58),
	.w2(32'hbac8902f),
	.w3(32'h3b07e089),
	.w4(32'h3b7c0e5d),
	.w5(32'hba9c1ad7),
	.w6(32'hbaea913c),
	.w7(32'hbb608dc8),
	.w8(32'h3b272875),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e7cbc),
	.w1(32'hbac46c8d),
	.w2(32'hbb4fcd17),
	.w3(32'h3c1b8e6f),
	.w4(32'h3bef0c0a),
	.w5(32'hba391317),
	.w6(32'h3b9d2cf7),
	.w7(32'h3a8a3799),
	.w8(32'hbad7d365),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984933b),
	.w1(32'hbbba2630),
	.w2(32'hbc48ed3d),
	.w3(32'h3b434dcb),
	.w4(32'hbb46c60b),
	.w5(32'hbbf4ba05),
	.w6(32'h3ba6af9f),
	.w7(32'h3ab1c273),
	.w8(32'hbbd60249),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12df81),
	.w1(32'hbc0084bc),
	.w2(32'hbca96115),
	.w3(32'h3962735f),
	.w4(32'h3a66d23f),
	.w5(32'hbd0b72ad),
	.w6(32'h3af62dc7),
	.w7(32'h3ad16509),
	.w8(32'hbcbcd408),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd17f7d2),
	.w1(32'hbcc71e11),
	.w2(32'h3b5dbb78),
	.w3(32'hbd7d91e1),
	.w4(32'hbd200ce4),
	.w5(32'h3c3840f1),
	.w6(32'hbd1895f0),
	.w7(32'hbc9f85cb),
	.w8(32'h3c201734),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a4140),
	.w1(32'hb98bd432),
	.w2(32'hbb1377cb),
	.w3(32'h3bbc0278),
	.w4(32'h3c238f60),
	.w5(32'hbb9aaf70),
	.w6(32'h3bd75a62),
	.w7(32'h3c043143),
	.w8(32'hbb81b7e1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c369142),
	.w1(32'hbb0099e7),
	.w2(32'hbcb0bf6f),
	.w3(32'h3c31ec42),
	.w4(32'hbb3a5143),
	.w5(32'hbc57846a),
	.w6(32'h3c57010b),
	.w7(32'hbad8abed),
	.w8(32'hbc379c47),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8241c),
	.w1(32'hbbbfedca),
	.w2(32'h3b8ef213),
	.w3(32'h3ba96e8d),
	.w4(32'h39891b8c),
	.w5(32'hbb1a4095),
	.w6(32'h3c108555),
	.w7(32'h3ade6909),
	.w8(32'hbb89c199),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2431a2),
	.w1(32'h3b8814c8),
	.w2(32'hbd01f945),
	.w3(32'h3b64883d),
	.w4(32'hb9ff61c8),
	.w5(32'hbd304dcd),
	.w6(32'h3bad7bf4),
	.w7(32'hb98d87dd),
	.w8(32'hbcaa18f5),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd40dc24),
	.w1(32'hbcc62345),
	.w2(32'hbc56d5d1),
	.w3(32'hbd94ea28),
	.w4(32'hbd438aed),
	.w5(32'hbaec0b02),
	.w6(32'hbd4d5d92),
	.w7(32'hbd11d799),
	.w8(32'hbc207e60),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafba8ca),
	.w1(32'hbb90bfec),
	.w2(32'hbbdfdaae),
	.w3(32'h3cc607b8),
	.w4(32'h3c86aa36),
	.w5(32'hbb93d2c4),
	.w6(32'hba9cfc5b),
	.w7(32'h3ba00edb),
	.w8(32'hbb8f8ac5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5473b),
	.w1(32'hbb65547e),
	.w2(32'hbc3f72bc),
	.w3(32'hba03eff1),
	.w4(32'h3afa3625),
	.w5(32'hbc83c5ff),
	.w6(32'hbb2bede3),
	.w7(32'h3aaf3538),
	.w8(32'hbc4f7433),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc804d08),
	.w1(32'hbc36d662),
	.w2(32'h3bc71b11),
	.w3(32'hbc936666),
	.w4(32'hbc44d022),
	.w5(32'h3c8b9830),
	.w6(32'hbc7bfc3f),
	.w7(32'hbc33bf63),
	.w8(32'h3c6e6e15),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d9592),
	.w1(32'h3c23e571),
	.w2(32'h3c06f50c),
	.w3(32'h3c34a50d),
	.w4(32'h3c5d7896),
	.w5(32'h3c37866f),
	.w6(32'h3b3ec64c),
	.w7(32'h3b6d0904),
	.w8(32'h3b762357),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee1025),
	.w1(32'h3bf24274),
	.w2(32'hbb2a7549),
	.w3(32'h3c62e547),
	.w4(32'h3c8aeb91),
	.w5(32'hbae16edf),
	.w6(32'h3b893595),
	.w7(32'hba0f5a26),
	.w8(32'h3b2b095c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012000),
	.w1(32'h3bb836ad),
	.w2(32'h3ab5931b),
	.w3(32'hbc0d6726),
	.w4(32'hbbfb1e1c),
	.w5(32'hb726f364),
	.w6(32'h3b0dfa5e),
	.w7(32'hbb46f860),
	.w8(32'h3b0479ff),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53ae07),
	.w1(32'hba340915),
	.w2(32'h3b3e86e6),
	.w3(32'h3c8e5876),
	.w4(32'hbb04c686),
	.w5(32'h3bda8aac),
	.w6(32'h3c53c07e),
	.w7(32'hbacbd9b9),
	.w8(32'h3be3a503),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77c991),
	.w1(32'h3bb7bf0e),
	.w2(32'h39699e73),
	.w3(32'h3c045763),
	.w4(32'h3c3a1fe9),
	.w5(32'hba69b1e7),
	.w6(32'h3c8b074b),
	.w7(32'h3c5012be),
	.w8(32'h39dfc801),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab39d5d),
	.w1(32'hbb164d7f),
	.w2(32'h3c22be62),
	.w3(32'h3b4c3ef2),
	.w4(32'hbaa80191),
	.w5(32'h3c77f1fc),
	.w6(32'h3b724311),
	.w7(32'hbb58c1b5),
	.w8(32'h3bba1100),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb0ac3),
	.w1(32'h393e6339),
	.w2(32'hbc545ee2),
	.w3(32'h3b4f0c85),
	.w4(32'h3bcf89d8),
	.w5(32'hbc7bf76a),
	.w6(32'h3b6efcba),
	.w7(32'h3bde2d09),
	.w8(32'hbba32ec9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c0d0a),
	.w1(32'hbc9a9731),
	.w2(32'hbcf002a2),
	.w3(32'hbc968320),
	.w4(32'hbcea2ebd),
	.w5(32'hbd0e4923),
	.w6(32'hbafc7fc8),
	.w7(32'hbc3a6fff),
	.w8(32'hbc75b13b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfdb9c),
	.w1(32'hbc83d708),
	.w2(32'hbc51084f),
	.w3(32'hbd408a13),
	.w4(32'hbd1c5a14),
	.w5(32'hbcab53a1),
	.w6(32'hbcc65c83),
	.w7(32'hbcd6f76d),
	.w8(32'hbbaead2c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc808da5),
	.w1(32'hbb74253f),
	.w2(32'h3a2cd91f),
	.w3(32'hbcabf596),
	.w4(32'h39875242),
	.w5(32'h3b5ab9df),
	.w6(32'hbb38545c),
	.w7(32'h3bb2d931),
	.w8(32'h3bb18d56),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba24a90),
	.w1(32'hbb928b16),
	.w2(32'hbb9cffb8),
	.w3(32'hbb103227),
	.w4(32'h3a64aba9),
	.w5(32'hbb86d132),
	.w6(32'hbb9b093b),
	.w7(32'hbb30c204),
	.w8(32'hbb9670fd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9787e6),
	.w1(32'h3aaef5ad),
	.w2(32'h3bd7efc5),
	.w3(32'hb9f66e2c),
	.w4(32'h3add2b8e),
	.w5(32'hbcaed69b),
	.w6(32'hba1f3daf),
	.w7(32'h3aff846b),
	.w8(32'hbc89264d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c2990),
	.w1(32'hbcddc330),
	.w2(32'hbb05382b),
	.w3(32'hbd31a56f),
	.w4(32'hbce93627),
	.w5(32'h3bd5b079),
	.w6(32'hbcbffd06),
	.w7(32'hbc2ef645),
	.w8(32'hbb8f0f77),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa9ab0),
	.w1(32'hbb4e0761),
	.w2(32'hbcd104f4),
	.w3(32'h3c9ad197),
	.w4(32'h3c2cb469),
	.w5(32'hbcb1f1e5),
	.w6(32'h3c5d1e7f),
	.w7(32'h3c7f82ae),
	.w8(32'hba04b386),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba62699),
	.w1(32'hbc5c6169),
	.w2(32'hbcdce106),
	.w3(32'h3ba4b6b3),
	.w4(32'hba793e49),
	.w5(32'hbc8bbdfd),
	.w6(32'h3cac778f),
	.w7(32'h3c4e63d9),
	.w8(32'hbc9bfd33),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d5e5b),
	.w1(32'hbc6f481b),
	.w2(32'h3b715a72),
	.w3(32'hb8d83b60),
	.w4(32'h3a9835d1),
	.w5(32'h3a2902c9),
	.w6(32'h3b1696ee),
	.w7(32'h3b93c0bf),
	.w8(32'hbaba1136),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b9072),
	.w1(32'h3c883825),
	.w2(32'hbb7b1e87),
	.w3(32'h3bb0314d),
	.w4(32'h3c2bc239),
	.w5(32'h3799b720),
	.w6(32'h3b4c6d81),
	.w7(32'h3bbfe2ae),
	.w8(32'h3afd35cb),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb647d2c),
	.w1(32'hb98d296e),
	.w2(32'h3c956846),
	.w3(32'hbb060bc9),
	.w4(32'h3b06ab8e),
	.w5(32'h3c872028),
	.w6(32'hba851da7),
	.w7(32'h3b1a4471),
	.w8(32'h3c2d61c7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b0169),
	.w1(32'h3c26c347),
	.w2(32'h3ba3b27b),
	.w3(32'hbaf8fb40),
	.w4(32'h3bd136e4),
	.w5(32'hb9913411),
	.w6(32'h3b8f3b4b),
	.w7(32'h3b8ab5e9),
	.w8(32'hbbe24a49),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c807a86),
	.w1(32'h3bda76c7),
	.w2(32'h3980732e),
	.w3(32'hbb603cfa),
	.w4(32'hbc0d2f0a),
	.w5(32'h3c0e4783),
	.w6(32'hbc8063a3),
	.w7(32'hbc8c42c8),
	.w8(32'h3a197a0d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9e600),
	.w1(32'hbb69b6d4),
	.w2(32'hbc1b7785),
	.w3(32'hb936c031),
	.w4(32'h3b27f551),
	.w5(32'hbbff7d26),
	.w6(32'hbb10140d),
	.w7(32'hb6f90429),
	.w8(32'h3bc274ae),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a2da),
	.w1(32'h3a06a67a),
	.w2(32'h3c1ecef4),
	.w3(32'hbcc4dd22),
	.w4(32'hbc8d0a46),
	.w5(32'h3ba5a15a),
	.w6(32'hbaaa696c),
	.w7(32'hbc38e30c),
	.w8(32'hbb8e9936),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b806c),
	.w1(32'h3b93e3c4),
	.w2(32'hbb9f3825),
	.w3(32'h3c7e771d),
	.w4(32'h3900e7fe),
	.w5(32'hb9c26f5b),
	.w6(32'h3c054846),
	.w7(32'hbb7c7431),
	.w8(32'h3ba5f65c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4d9ef),
	.w1(32'h3bfac958),
	.w2(32'h3b3a2685),
	.w3(32'h3abd9ab7),
	.w4(32'h3c5abb81),
	.w5(32'h3c6154f4),
	.w6(32'h3bd0b974),
	.w7(32'h3c5fbfb1),
	.w8(32'h3b9a209e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b281c),
	.w1(32'h3c0ab624),
	.w2(32'h3abc42c0),
	.w3(32'h3d15d329),
	.w4(32'h3cc70206),
	.w5(32'h3c583f51),
	.w6(32'h3c903d0f),
	.w7(32'h3cae70e7),
	.w8(32'h3c049867),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90a6f7),
	.w1(32'h3c5c3066),
	.w2(32'hbbdfe896),
	.w3(32'h3d1d86c8),
	.w4(32'h3ceedfdd),
	.w5(32'hb9df34cb),
	.w6(32'h3c907055),
	.w7(32'h3c699b8f),
	.w8(32'hbbc49eeb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaad240),
	.w1(32'hbae485f6),
	.w2(32'hbb82aa72),
	.w3(32'h3c40fd9e),
	.w4(32'h3ba9189b),
	.w5(32'hbb123986),
	.w6(32'h3c06c4b3),
	.w7(32'h3bccaa74),
	.w8(32'h3af053f3),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b400d99),
	.w1(32'h3ab08008),
	.w2(32'hbca39d33),
	.w3(32'h3bc8f367),
	.w4(32'h39d9e6bc),
	.w5(32'hbd10b464),
	.w6(32'h3bcdd672),
	.w7(32'hba958587),
	.w8(32'hbca3d788),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa78aa),
	.w1(32'hbced8d35),
	.w2(32'hbacbaeb8),
	.w3(32'hbd5547b7),
	.w4(32'hbd3524c7),
	.w5(32'hbafe3a15),
	.w6(32'hbd107eee),
	.w7(32'hbd01173a),
	.w8(32'hb9cc148e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba810973),
	.w1(32'hbad2d1f8),
	.w2(32'hbacdba04),
	.w3(32'h3b4a1670),
	.w4(32'h3a679684),
	.w5(32'hbadb55b4),
	.w6(32'h3bb2c1f7),
	.w7(32'hba17b50d),
	.w8(32'h39e653f4),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87193b),
	.w1(32'h3ba49544),
	.w2(32'h3a39f883),
	.w3(32'h3bba5312),
	.w4(32'h3bad878a),
	.w5(32'hbafbd422),
	.w6(32'h3bca774c),
	.w7(32'h3baf23b6),
	.w8(32'h3bc2d00d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147948),
	.w1(32'h3bb2daaa),
	.w2(32'hbcaefd8f),
	.w3(32'hbba02142),
	.w4(32'hbb3f8e3b),
	.w5(32'hbd1197fa),
	.w6(32'h3b801814),
	.w7(32'h3a84cd13),
	.w8(32'hbc5bc67f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95698d),
	.w1(32'hbc172725),
	.w2(32'h3a9fc944),
	.w3(32'hbd1e3ecb),
	.w4(32'hbca15f6a),
	.w5(32'h3c5c0eed),
	.w6(32'hbd07f410),
	.w7(32'hbcbfc9fb),
	.w8(32'h39b22923),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a2ba4),
	.w1(32'h3c75b780),
	.w2(32'hbb6b4b88),
	.w3(32'h3cd4672a),
	.w4(32'h3cb74733),
	.w5(32'hbb314ade),
	.w6(32'h3c80e539),
	.w7(32'h3c9b838c),
	.w8(32'h3b9927a4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa031a7),
	.w1(32'h3ba1cebd),
	.w2(32'hbc2163be),
	.w3(32'hbc2c00eb),
	.w4(32'h3a5187b8),
	.w5(32'hbcb644b1),
	.w6(32'hbb93f660),
	.w7(32'h3b23e2e4),
	.w8(32'hbc71e7d3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5f59a),
	.w1(32'hbcd5cedb),
	.w2(32'hbb72cc6e),
	.w3(32'hbce8c0cf),
	.w4(32'hbca335ea),
	.w5(32'h3c0577b7),
	.w6(32'hbc9c24de),
	.w7(32'hbc6a688d),
	.w8(32'hbc0916dd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c314f4b),
	.w1(32'h3b84d538),
	.w2(32'h3b1d7dfb),
	.w3(32'h3b890507),
	.w4(32'hbb8980f8),
	.w5(32'hba5420a5),
	.w6(32'hbb9c9509),
	.w7(32'hbbeaaa69),
	.w8(32'h3a73299a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4ec7e),
	.w1(32'h3b8558ea),
	.w2(32'hbb19ac28),
	.w3(32'h3c6a1a5b),
	.w4(32'h3c0e2916),
	.w5(32'hbb252e5e),
	.w6(32'h3c8d3156),
	.w7(32'h3c1d18cf),
	.w8(32'hbb241960),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc221a6),
	.w1(32'hba14d418),
	.w2(32'h38e26375),
	.w3(32'hbbb886a8),
	.w4(32'hbc559049),
	.w5(32'h39dfc82a),
	.w6(32'h3b8cf126),
	.w7(32'hbbb8dcf5),
	.w8(32'hbb63fd2d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cc584),
	.w1(32'h3a29fbb3),
	.w2(32'hbc4866d0),
	.w3(32'h3a7bacde),
	.w4(32'h3a2bf5a5),
	.w5(32'hbbb0ba0a),
	.w6(32'hbbaf8a81),
	.w7(32'hbbc27100),
	.w8(32'hbc10752c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4d9e0),
	.w1(32'h3a42c427),
	.w2(32'hbb88bf55),
	.w3(32'h3c1fb78b),
	.w4(32'h3c384db9),
	.w5(32'h3b1599a7),
	.w6(32'h3b598875),
	.w7(32'h3b3b6396),
	.w8(32'h3b657caa),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c6823),
	.w1(32'hbb49c470),
	.w2(32'h3b0ffd6a),
	.w3(32'h3c0ff52d),
	.w4(32'h3bf33f17),
	.w5(32'h3c0749ff),
	.w6(32'h3b8858a7),
	.w7(32'hba7a02ee),
	.w8(32'h3c15da71),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2067b2),
	.w1(32'h3beb37a8),
	.w2(32'hb8ce370d),
	.w3(32'h3cf6546f),
	.w4(32'h3cbfd217),
	.w5(32'h3c5da548),
	.w6(32'h3cb89478),
	.w7(32'h3c8e6a50),
	.w8(32'hba09dcb9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e9b20),
	.w1(32'h3c72e2c5),
	.w2(32'h3c4a4333),
	.w3(32'h3d02ab49),
	.w4(32'h3ca210b0),
	.w5(32'h3c6313c7),
	.w6(32'h3ca4a588),
	.w7(32'h3c76b2e1),
	.w8(32'h3c1011b0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c487fc2),
	.w1(32'h3bcee9cb),
	.w2(32'h3b9b9b0c),
	.w3(32'h3c0d86a6),
	.w4(32'h3b89ee88),
	.w5(32'h3b49f760),
	.w6(32'h3b81ef30),
	.w7(32'h3b53b80a),
	.w8(32'h3b372949),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a3934),
	.w1(32'h3bc06e16),
	.w2(32'h381a145a),
	.w3(32'hb9d7e54e),
	.w4(32'h3b513a31),
	.w5(32'hb988d5ce),
	.w6(32'hbaf76046),
	.w7(32'h3b65e95e),
	.w8(32'h3a8fec83),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e40b9),
	.w1(32'h39ae4712),
	.w2(32'h3bd353cc),
	.w3(32'hbb2a6657),
	.w4(32'hba0e728a),
	.w5(32'h3c3959c7),
	.w6(32'h3a66b93e),
	.w7(32'h3b09e706),
	.w8(32'h3c1504e6),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc101cec),
	.w1(32'hbc264024),
	.w2(32'hbb85b10d),
	.w3(32'h399844ee),
	.w4(32'hbc3465db),
	.w5(32'hbafb6a61),
	.w6(32'h3c67caac),
	.w7(32'hbb94b5e4),
	.w8(32'hbabab83e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10fdad),
	.w1(32'h3a52ba87),
	.w2(32'hbc509526),
	.w3(32'h3bc3361c),
	.w4(32'h3b669f66),
	.w5(32'hbce6e976),
	.w6(32'h3b073a4d),
	.w7(32'hba968a49),
	.w8(32'hbcbcc0c2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd038000),
	.w1(32'hbcca0b14),
	.w2(32'hbd00546e),
	.w3(32'hbd405ade),
	.w4(32'hbce88093),
	.w5(32'hbd3c0a65),
	.w6(32'hbd00ec8e),
	.w7(32'hbce3fdd6),
	.w8(32'hbd238299),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3b7fe3),
	.w1(32'hbd20364d),
	.w2(32'hbcf5c174),
	.w3(32'hbd99807f),
	.w4(32'hbd5f912e),
	.w5(32'hbd37f701),
	.w6(32'hbd54ba09),
	.w7(32'hbd07d44d),
	.w8(32'hbd05b33c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3b696c),
	.w1(32'hbcf96e93),
	.w2(32'h3b85ccd7),
	.w3(32'hbd787e50),
	.w4(32'hbd20315d),
	.w5(32'hbaa12fc9),
	.w6(32'hbd2654d3),
	.w7(32'hbcb8458d),
	.w8(32'h3bb1d17e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule