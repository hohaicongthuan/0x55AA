module layer_10_featuremap_373(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b972e44),
	.w1(32'h3b9acd91),
	.w2(32'h3be82686),
	.w3(32'hbb47325f),
	.w4(32'h39c1d2ca),
	.w5(32'h3bc40520),
	.w6(32'hbbd9938d),
	.w7(32'h3c0f8fa0),
	.w8(32'hb93903da),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a8f51),
	.w1(32'h3c3e2200),
	.w2(32'hbc3abe7c),
	.w3(32'hbb2cbea5),
	.w4(32'hbc8f7b6f),
	.w5(32'hb9303011),
	.w6(32'h3c31eecd),
	.w7(32'hbbf8f748),
	.w8(32'h3bfbc48b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2485e5),
	.w1(32'hbb1cb8ce),
	.w2(32'h3b0725b6),
	.w3(32'h3bf58cb3),
	.w4(32'hbc20a695),
	.w5(32'h3bfd1243),
	.w6(32'hbbce39cc),
	.w7(32'hbc323a6d),
	.w8(32'h3be9d5a4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e5fdc),
	.w1(32'hbcf33e18),
	.w2(32'h39381cf3),
	.w3(32'hbc676505),
	.w4(32'h3d06cb54),
	.w5(32'h3c815338),
	.w6(32'h3ba927bc),
	.w7(32'hbc6636ce),
	.w8(32'hbc0b31e3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba354c0),
	.w1(32'hbc744a1c),
	.w2(32'hbb46ef99),
	.w3(32'h3c620c00),
	.w4(32'hbc181ec0),
	.w5(32'h3a47f74d),
	.w6(32'hbc873e20),
	.w7(32'hbc45dad0),
	.w8(32'h3beac7ca),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf59cc0),
	.w1(32'hba965de7),
	.w2(32'hbc18e498),
	.w3(32'hbaf4d01d),
	.w4(32'h3a8f60e9),
	.w5(32'h3c872ecb),
	.w6(32'hbb67e1cd),
	.w7(32'h3b0e5a4b),
	.w8(32'h3b1d007a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bbc75),
	.w1(32'hbc1563e7),
	.w2(32'hbb3cb5ce),
	.w3(32'h3c4355c9),
	.w4(32'h3b8a7718),
	.w5(32'hbb241668),
	.w6(32'h3cb36a9c),
	.w7(32'hbc1f9805),
	.w8(32'h3c036ea6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73140),
	.w1(32'hbb961323),
	.w2(32'h3bed8cd1),
	.w3(32'hbbf86bb7),
	.w4(32'h3c0b80d5),
	.w5(32'hb906af49),
	.w6(32'hbb90f340),
	.w7(32'h3ba2e909),
	.w8(32'h3c01dd90),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75cb91),
	.w1(32'hbb713358),
	.w2(32'h3c06551b),
	.w3(32'hbb83db07),
	.w4(32'hbc7d1fbb),
	.w5(32'hbba82f98),
	.w6(32'h3bee18d9),
	.w7(32'h3c247182),
	.w8(32'hbabe24bd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f39a2),
	.w1(32'h39c535b2),
	.w2(32'h3c3f45e1),
	.w3(32'h3b888da9),
	.w4(32'h3d29e7ce),
	.w5(32'h3b7b2824),
	.w6(32'hbc428f40),
	.w7(32'hbb90559e),
	.w8(32'h3b53595c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70979f),
	.w1(32'hbba7c7ce),
	.w2(32'hba91699c),
	.w3(32'hbc828db3),
	.w4(32'hbb595af0),
	.w5(32'hbbad808b),
	.w6(32'hbb83e1d8),
	.w7(32'h3bb3a7aa),
	.w8(32'hbc441a10),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c47b3),
	.w1(32'h38b4c172),
	.w2(32'hbc3ae464),
	.w3(32'h3c39dce8),
	.w4(32'h3b24b17d),
	.w5(32'hbadf1e9a),
	.w6(32'hbb358600),
	.w7(32'hb93f0000),
	.w8(32'hbccb5322),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fd243),
	.w1(32'h3b8da3f8),
	.w2(32'hbb90f181),
	.w3(32'h3bbfb94d),
	.w4(32'hbc2b3d23),
	.w5(32'h3bc6f516),
	.w6(32'hbb1c88ca),
	.w7(32'hbc3e3a30),
	.w8(32'hba149265),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c0776),
	.w1(32'hbaf63e82),
	.w2(32'hbc671d8b),
	.w3(32'hbc245d9b),
	.w4(32'h39f02735),
	.w5(32'h3c7d66bc),
	.w6(32'h3ad2154f),
	.w7(32'hba9b8e54),
	.w8(32'h3bd5afba),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca104dd),
	.w1(32'hbb450504),
	.w2(32'hbae8b695),
	.w3(32'hb7da86e8),
	.w4(32'h3c25ddfa),
	.w5(32'h3b6401b9),
	.w6(32'h3c14e452),
	.w7(32'hbc8c690a),
	.w8(32'hbba2e9a4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaff73e),
	.w1(32'hbb67b0bf),
	.w2(32'h3c6c226d),
	.w3(32'h3bd722f2),
	.w4(32'h3bb2edf7),
	.w5(32'h3c66c43f),
	.w6(32'h3cbc3c1a),
	.w7(32'h3c182c11),
	.w8(32'hba86abdd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195576),
	.w1(32'hbb8711ca),
	.w2(32'hbb579c77),
	.w3(32'hbbb81312),
	.w4(32'h3959a0e4),
	.w5(32'hbbdad135),
	.w6(32'h3b29f80e),
	.w7(32'h39d033c5),
	.w8(32'hbc0cf394),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4fb7e),
	.w1(32'h3c004ed2),
	.w2(32'hbba67482),
	.w3(32'hbc234c3a),
	.w4(32'h3c5df16b),
	.w5(32'hba991922),
	.w6(32'hbc92a717),
	.w7(32'h3c1471b9),
	.w8(32'hbb8253e9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd656e),
	.w1(32'h3bb98840),
	.w2(32'hbc1db5f3),
	.w3(32'hbba43a1f),
	.w4(32'h3a39e60b),
	.w5(32'hbc741acc),
	.w6(32'hbca1d252),
	.w7(32'hbc3d808b),
	.w8(32'hbbb45105),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec6f5a),
	.w1(32'hba06d211),
	.w2(32'hbb871df8),
	.w3(32'h3c8741ef),
	.w4(32'hbbbc6ab5),
	.w5(32'h3aca5ec0),
	.w6(32'h3c3ad4d7),
	.w7(32'h3b9e2eca),
	.w8(32'h39fb9698),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c75f3),
	.w1(32'h39acd580),
	.w2(32'h3b14d524),
	.w3(32'hbc2f155e),
	.w4(32'h3ca8d5a2),
	.w5(32'h3bf51809),
	.w6(32'hbbad53ea),
	.w7(32'hb9dcadd5),
	.w8(32'h3c2bc529),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd05b00),
	.w1(32'h3c91001e),
	.w2(32'hbaf3f281),
	.w3(32'hbb763402),
	.w4(32'hbb0eac47),
	.w5(32'hbc9bb603),
	.w6(32'hbc1c7d6e),
	.w7(32'h3a94a08e),
	.w8(32'h3c95a892),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10e38e),
	.w1(32'h3abda7a5),
	.w2(32'h3bac36f5),
	.w3(32'h3bb25c81),
	.w4(32'hbb3bb475),
	.w5(32'hbc3d5c12),
	.w6(32'h3b4de4e2),
	.w7(32'hbc241e80),
	.w8(32'h3b903f0a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c0154),
	.w1(32'h3a917b64),
	.w2(32'h3b902561),
	.w3(32'h3ccb3a41),
	.w4(32'hbc0c7ac2),
	.w5(32'hbac49628),
	.w6(32'hbc4d837e),
	.w7(32'hbbc651f2),
	.w8(32'h3c7e9cda),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e57dd),
	.w1(32'hbc9c2eec),
	.w2(32'h3a76b200),
	.w3(32'h3c8cde5a),
	.w4(32'h3cc71344),
	.w5(32'h3b543978),
	.w6(32'h3aa9bfe0),
	.w7(32'hbc81e27a),
	.w8(32'h3c0c473e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c167ac3),
	.w1(32'h3b701600),
	.w2(32'hbab5b2a9),
	.w3(32'h3c8a5741),
	.w4(32'hbc59f129),
	.w5(32'h3c92bfd5),
	.w6(32'hba9de9e5),
	.w7(32'hbb8b44a1),
	.w8(32'hbc6f75b3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8f8b2),
	.w1(32'hbc3b8155),
	.w2(32'hbbb6fb05),
	.w3(32'h3a1f9cfa),
	.w4(32'hbb1a740b),
	.w5(32'hbb87814b),
	.w6(32'h3b55c0f2),
	.w7(32'h3a83b7b6),
	.w8(32'h3c879654),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b50ec),
	.w1(32'h3c5d45a9),
	.w2(32'hbc4c1906),
	.w3(32'hbb3e8bc6),
	.w4(32'hbc027703),
	.w5(32'hbb741530),
	.w6(32'h3aa9d02d),
	.w7(32'h3b61c25d),
	.w8(32'h3be24142),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc818a),
	.w1(32'h3c89e040),
	.w2(32'hbb872721),
	.w3(32'hbbe03d0d),
	.w4(32'hbb5fc005),
	.w5(32'h3a9a81cb),
	.w6(32'hbaba0f78),
	.w7(32'hbbc1915c),
	.w8(32'h3c70d628),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84699d),
	.w1(32'hbb763ba6),
	.w2(32'hbaaa68e0),
	.w3(32'h3cabed6f),
	.w4(32'hbb964b7a),
	.w5(32'h3c2562f3),
	.w6(32'h3a81786d),
	.w7(32'hbc221a61),
	.w8(32'hbc2689d4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85c6d6),
	.w1(32'hbc22bf7b),
	.w2(32'h3b320103),
	.w3(32'hbab98eec),
	.w4(32'h3b97aa3a),
	.w5(32'h3ba03446),
	.w6(32'h3c82ecc4),
	.w7(32'hb96c20b4),
	.w8(32'h3b9800a3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d0151),
	.w1(32'hbc35eb89),
	.w2(32'hb9a9d451),
	.w3(32'hbbbdb657),
	.w4(32'hbc437f5b),
	.w5(32'hbc30d5da),
	.w6(32'hbc017a02),
	.w7(32'hb7bb0d00),
	.w8(32'h3c7bd25b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2ab45),
	.w1(32'hba3ddc1d),
	.w2(32'h3c5bb070),
	.w3(32'hbbfe173d),
	.w4(32'hb9bbc922),
	.w5(32'h3c7bd6c0),
	.w6(32'hbbf77fdf),
	.w7(32'h3ca23062),
	.w8(32'h3a38fd79),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7183),
	.w1(32'h3b6fb974),
	.w2(32'h3b91585c),
	.w3(32'h3b2fcd5e),
	.w4(32'h3c0e8b3d),
	.w5(32'h3c4c810f),
	.w6(32'h38683ad6),
	.w7(32'h3b16fc6a),
	.w8(32'hba538ebd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c9e48),
	.w1(32'h3b58a250),
	.w2(32'h3c2e9c63),
	.w3(32'hba8893bd),
	.w4(32'hbc1c787e),
	.w5(32'hbb1d7991),
	.w6(32'h3cc5a079),
	.w7(32'hbb8bd79d),
	.w8(32'h3c51175d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4aec1),
	.w1(32'h3bf6e362),
	.w2(32'h3ad15025),
	.w3(32'hb9477e33),
	.w4(32'h3af80902),
	.w5(32'h3bc25e11),
	.w6(32'hbb9537c8),
	.w7(32'h3d904765),
	.w8(32'hbbcc2fe5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf67e8a),
	.w1(32'h3ba8e6c7),
	.w2(32'hbb14fa35),
	.w3(32'hbb6c6783),
	.w4(32'h3c0fe26c),
	.w5(32'h3c1f62f3),
	.w6(32'hbb162415),
	.w7(32'hbba097c4),
	.w8(32'hbc7ac939),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb996454),
	.w1(32'h3874053b),
	.w2(32'hba813fd9),
	.w3(32'hbc5266b6),
	.w4(32'h3abe3c0f),
	.w5(32'h3adf47c0),
	.w6(32'hbc390102),
	.w7(32'hb8e6f388),
	.w8(32'h3c97a23a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92887d),
	.w1(32'hbb420305),
	.w2(32'hbb9df2c0),
	.w3(32'hbbbee838),
	.w4(32'hbc408728),
	.w5(32'hbbff775a),
	.w6(32'hbb8c191d),
	.w7(32'h3ba3541b),
	.w8(32'hba979223),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc016e05),
	.w1(32'h3b7baf8a),
	.w2(32'h3b4c101d),
	.w3(32'hbbccd2bf),
	.w4(32'h3ab3bed7),
	.w5(32'h3bab4c82),
	.w6(32'hbbd3946d),
	.w7(32'hbb9e5ad6),
	.w8(32'h3bda286b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a13ecf),
	.w1(32'hbcc63429),
	.w2(32'h3caff451),
	.w3(32'h3b91095c),
	.w4(32'h3c1a31df),
	.w5(32'h3b9144b8),
	.w6(32'h3a9fedde),
	.w7(32'h3b7fa190),
	.w8(32'h3b9ed76b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a9734),
	.w1(32'h3c374029),
	.w2(32'h399879e3),
	.w3(32'h3ba098d4),
	.w4(32'h39b52b58),
	.w5(32'hbc30589b),
	.w6(32'h3bc72765),
	.w7(32'hba9df02b),
	.w8(32'h3c342641),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec1b39),
	.w1(32'hbacebea9),
	.w2(32'h3a956b03),
	.w3(32'hbb965e2e),
	.w4(32'hbc9e5687),
	.w5(32'hbbb9aef7),
	.w6(32'h3aa7c8e5),
	.w7(32'h3ca4a23e),
	.w8(32'hbbdce6e7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d03a35),
	.w1(32'h3b04cb48),
	.w2(32'hba798633),
	.w3(32'h3b8918a9),
	.w4(32'hbbd34ee0),
	.w5(32'h3b10c5a3),
	.w6(32'hbc28df87),
	.w7(32'h3a918aba),
	.w8(32'hbb81db1f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a480503),
	.w1(32'h3996b766),
	.w2(32'hbc08d47a),
	.w3(32'hbc12c53b),
	.w4(32'hbc27f0f5),
	.w5(32'h3b3cf185),
	.w6(32'h3b854932),
	.w7(32'h3bcaeca5),
	.w8(32'h3a487209),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e38c2),
	.w1(32'h3ae03bcc),
	.w2(32'h3c083e89),
	.w3(32'h3b7ff916),
	.w4(32'h3c1fd3e1),
	.w5(32'h3c0c9129),
	.w6(32'hbb177234),
	.w7(32'hbc43cfcf),
	.w8(32'hbb8e5ef7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c614358),
	.w1(32'h3c136094),
	.w2(32'h3ba954b3),
	.w3(32'h3a1e0bee),
	.w4(32'h3ba74914),
	.w5(32'hbaed5a4a),
	.w6(32'hbb78024f),
	.w7(32'hbc0e9731),
	.w8(32'hbc028d09),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28260b),
	.w1(32'h3c8ff976),
	.w2(32'h3b5313fc),
	.w3(32'h3bc8e779),
	.w4(32'hbc32f4a8),
	.w5(32'hbb7208f0),
	.w6(32'hbc28d412),
	.w7(32'hbb501176),
	.w8(32'hbbe4c3ae),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a2de6),
	.w1(32'h3c179fb7),
	.w2(32'h3a98b416),
	.w3(32'h3a908638),
	.w4(32'hbc23564d),
	.w5(32'h3b9c93e2),
	.w6(32'h3be247ac),
	.w7(32'h3bfaf670),
	.w8(32'hbb4af272),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a035a),
	.w1(32'hbbb6a94e),
	.w2(32'hbbba8951),
	.w3(32'hbb1802bb),
	.w4(32'hbc0fa08d),
	.w5(32'h3c52203c),
	.w6(32'hbc02be0c),
	.w7(32'hbb80449d),
	.w8(32'h3b59f937),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9c61),
	.w1(32'h3c475341),
	.w2(32'h3bdcabef),
	.w3(32'hba0e55ec),
	.w4(32'hbb5d8ff9),
	.w5(32'h3a33a712),
	.w6(32'hbc902930),
	.w7(32'hbc2826de),
	.w8(32'h3b4c9976),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6fc38),
	.w1(32'h3ce066f2),
	.w2(32'hbb8beafc),
	.w3(32'hbc1afa8f),
	.w4(32'hba7282a0),
	.w5(32'hbc39ee09),
	.w6(32'hbca5487d),
	.w7(32'hbc00124f),
	.w8(32'hbbca3f83),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc238565),
	.w1(32'hbb117db7),
	.w2(32'hbc03b41d),
	.w3(32'hbb3cf0aa),
	.w4(32'hbc1826ea),
	.w5(32'h3b77abd3),
	.w6(32'hbb892b10),
	.w7(32'hbc25cd04),
	.w8(32'hbc5b0618),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ec8d7),
	.w1(32'hbc800379),
	.w2(32'h3aa8f7cd),
	.w3(32'h3c3488ad),
	.w4(32'hbb2a69ce),
	.w5(32'hbc2fbc22),
	.w6(32'h3baca00d),
	.w7(32'h3c8ce6e6),
	.w8(32'hbc0e62b9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ea31d),
	.w1(32'hbaf946e0),
	.w2(32'hbb270d03),
	.w3(32'hbc9a47a1),
	.w4(32'h3c2d7884),
	.w5(32'h38e92309),
	.w6(32'h3b4ff63d),
	.w7(32'hbc278097),
	.w8(32'h3c016d83),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b98f5),
	.w1(32'hbc0e2d4a),
	.w2(32'hbbe9543f),
	.w3(32'h3a478bce),
	.w4(32'h3bf6541b),
	.w5(32'hba72bee3),
	.w6(32'hbaf6a058),
	.w7(32'hbaa8263e),
	.w8(32'h3bfeec42),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a3f89),
	.w1(32'hba7b8f4f),
	.w2(32'hbc1f5a01),
	.w3(32'hbbdad58c),
	.w4(32'h3b7cddfe),
	.w5(32'h3bab8f91),
	.w6(32'h3c1985d0),
	.w7(32'h3c08336e),
	.w8(32'hbc1b6684),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9d017),
	.w1(32'hbb2ed1f7),
	.w2(32'h3c65b129),
	.w3(32'hbcab4457),
	.w4(32'h3b73a719),
	.w5(32'h3b3aa7c1),
	.w6(32'h3bc2b574),
	.w7(32'h3c01c531),
	.w8(32'hbb264c44),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc928c69),
	.w1(32'h3ba57511),
	.w2(32'h3c138dca),
	.w3(32'h3bc0a9b6),
	.w4(32'h3bf9056c),
	.w5(32'h3bf1bd6a),
	.w6(32'h3c295941),
	.w7(32'hbc2f58ac),
	.w8(32'hbc099107),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6c45b),
	.w1(32'h3d99a645),
	.w2(32'h3af35f10),
	.w3(32'hbc08b519),
	.w4(32'h3c3c1af5),
	.w5(32'h3c2e4c26),
	.w6(32'h3c1ba50f),
	.w7(32'hbbe3e599),
	.w8(32'h3bbefc41),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c171c53),
	.w1(32'h3c09ff8c),
	.w2(32'hbab81a9c),
	.w3(32'h3c0a664f),
	.w4(32'h3b5b1eb9),
	.w5(32'h3d079be0),
	.w6(32'hbb34991d),
	.w7(32'h3c1e0740),
	.w8(32'h3c67ae71),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc258cd5),
	.w1(32'hbc37ab68),
	.w2(32'hbad4c6d9),
	.w3(32'hbc84e88a),
	.w4(32'hbb3bd619),
	.w5(32'hbbb3f50b),
	.w6(32'hbc0723c8),
	.w7(32'h3be1bfbf),
	.w8(32'h3acf3248),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b587e98),
	.w1(32'hbbf03284),
	.w2(32'hbb96e769),
	.w3(32'h3c89a0fc),
	.w4(32'hbc25add7),
	.w5(32'hbb52c264),
	.w6(32'h3b65032c),
	.w7(32'h3bd66476),
	.w8(32'h3c543b63),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a657694),
	.w1(32'hbb42b459),
	.w2(32'hbc9c473e),
	.w3(32'h3c37fe1e),
	.w4(32'h3bee1565),
	.w5(32'hbcc319b2),
	.w6(32'hbc346ce1),
	.w7(32'hb96d32af),
	.w8(32'h3b980ed6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b61d),
	.w1(32'hbb113752),
	.w2(32'h3bc4a1bc),
	.w3(32'hbb441fd6),
	.w4(32'hbb75b641),
	.w5(32'h3a83ea13),
	.w6(32'h3b6c7fb6),
	.w7(32'hba78decc),
	.w8(32'h3b8f8851),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba97464),
	.w1(32'hbb12c374),
	.w2(32'h3bf1f8a6),
	.w3(32'h3c0f7a90),
	.w4(32'hb9576195),
	.w5(32'hbb83a5c9),
	.w6(32'hbcb79109),
	.w7(32'h3c97baa1),
	.w8(32'h3b384ee5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc770f13),
	.w1(32'hba938c58),
	.w2(32'h3c0d13f4),
	.w3(32'h3c848174),
	.w4(32'h3b31f4be),
	.w5(32'h3a152b38),
	.w6(32'h3ae24a97),
	.w7(32'hbb7e55c6),
	.w8(32'hbb262631),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74da0c),
	.w1(32'hbaf40247),
	.w2(32'hbc305b84),
	.w3(32'hbb9f6aae),
	.w4(32'hba884786),
	.w5(32'h3c212d6d),
	.w6(32'h3b5ac496),
	.w7(32'h3c1666c3),
	.w8(32'hbb1071fb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf516d9),
	.w1(32'h3bbd5f1a),
	.w2(32'hbb3b547c),
	.w3(32'h3bc0e53c),
	.w4(32'h3984ba7d),
	.w5(32'h3c95f7d3),
	.w6(32'h3a5c3918),
	.w7(32'h3b7caad8),
	.w8(32'hbc31c03f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc825c4a),
	.w1(32'h3a48abbf),
	.w2(32'hbb916d90),
	.w3(32'hbc1b1554),
	.w4(32'h3b9e32ab),
	.w5(32'h3a680cd2),
	.w6(32'hba9107d1),
	.w7(32'h3c325da1),
	.w8(32'hbbaaed27),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0f8e2),
	.w1(32'h3c45befc),
	.w2(32'h3a9627d3),
	.w3(32'hbc63b94a),
	.w4(32'hbb0729b8),
	.w5(32'hbbab0797),
	.w6(32'hbc3e0fa6),
	.w7(32'h3b541ca1),
	.w8(32'h3c58670d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31f1f3),
	.w1(32'hbb5e0e55),
	.w2(32'h3bd7f5ce),
	.w3(32'hbbee7bf0),
	.w4(32'h3c3701e2),
	.w5(32'h3a1fa604),
	.w6(32'h3c2cdb79),
	.w7(32'h3c456815),
	.w8(32'hbc0cceb8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a4ee5),
	.w1(32'h3b805f3f),
	.w2(32'h3b149369),
	.w3(32'h3b384305),
	.w4(32'hb95e265e),
	.w5(32'h3b890e4f),
	.w6(32'h3b695e70),
	.w7(32'h3c4b469b),
	.w8(32'h3b9a435a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe814a),
	.w1(32'hb9ce00bf),
	.w2(32'h3b8a8159),
	.w3(32'h3b6a5664),
	.w4(32'hbad4ec27),
	.w5(32'h3c477a76),
	.w6(32'hbad856d2),
	.w7(32'hbb67787c),
	.w8(32'hbc82303d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc266978),
	.w1(32'h3c850819),
	.w2(32'hbb1636d4),
	.w3(32'hbbd9288d),
	.w4(32'h3c001759),
	.w5(32'h3c090c21),
	.w6(32'hbc49fd73),
	.w7(32'h3c7b502f),
	.w8(32'hbc1fd8e7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d1476),
	.w1(32'h3bd0be80),
	.w2(32'h3c36fb58),
	.w3(32'hbb8d0a96),
	.w4(32'h3bf99289),
	.w5(32'h3bebc743),
	.w6(32'h3c15ee6d),
	.w7(32'hba21d2f9),
	.w8(32'hbcac4a57),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc374eac),
	.w1(32'hba3510fa),
	.w2(32'hbb8a9c3c),
	.w3(32'hbad2de75),
	.w4(32'h3bf9ae87),
	.w5(32'h38604413),
	.w6(32'h3c3e9b02),
	.w7(32'hbab00220),
	.w8(32'hbc174fc3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71640a),
	.w1(32'hbb2e17ee),
	.w2(32'h3b984c56),
	.w3(32'hbb0d98bc),
	.w4(32'h3bc2a7a1),
	.w5(32'h397e387b),
	.w6(32'hb855b11b),
	.w7(32'h3bf6ed62),
	.w8(32'hb7dcb8f3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900e5f4),
	.w1(32'hbb3c376f),
	.w2(32'h3c546d4d),
	.w3(32'hbaaefca4),
	.w4(32'h368b02ce),
	.w5(32'hbb3b5d4b),
	.w6(32'h3c3fb07e),
	.w7(32'h3a3b7d59),
	.w8(32'hbbf86c9b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbab2ce),
	.w1(32'hbaf7f2e3),
	.w2(32'h3d16bfb3),
	.w3(32'hbada2301),
	.w4(32'hbc1802d8),
	.w5(32'h3b1169c7),
	.w6(32'hbac5afa9),
	.w7(32'hba9299ad),
	.w8(32'hbbbce58d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed75e),
	.w1(32'h3c557583),
	.w2(32'h3c120e55),
	.w3(32'h3bfb0f8c),
	.w4(32'h3b9d6c4b),
	.w5(32'hbb103bad),
	.w6(32'hbbbfae5b),
	.w7(32'h3c51d7d1),
	.w8(32'h3c80d667),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c141bb8),
	.w1(32'hbbcf0b4a),
	.w2(32'h3b4f90da),
	.w3(32'hbbb3d008),
	.w4(32'h3ad38293),
	.w5(32'hb9dc7f87),
	.w6(32'hbb334f2c),
	.w7(32'hbc2f6c22),
	.w8(32'h3d05057d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d6108),
	.w1(32'hbb2a0dfd),
	.w2(32'h3bfab394),
	.w3(32'hbb4970db),
	.w4(32'h3b54f750),
	.w5(32'h3c5a9194),
	.w6(32'h3b87d2a0),
	.w7(32'hbb449234),
	.w8(32'hbbde74fd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad16d),
	.w1(32'hb9a70d7a),
	.w2(32'hbae817dc),
	.w3(32'h3c817243),
	.w4(32'h3bb40d37),
	.w5(32'hbbc70274),
	.w6(32'hbc57f59e),
	.w7(32'h3b28dc17),
	.w8(32'hbc764e00),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8d18c),
	.w1(32'hba6c5035),
	.w2(32'hbb50dd34),
	.w3(32'hbb996068),
	.w4(32'hbcaed244),
	.w5(32'h3b6d6732),
	.w6(32'h3bed6306),
	.w7(32'hbd2e9e20),
	.w8(32'h3bcccad2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42c31e),
	.w1(32'hbc96210f),
	.w2(32'h3b450ef8),
	.w3(32'hbc0f8004),
	.w4(32'hbbc583fb),
	.w5(32'h3c15720e),
	.w6(32'hbc34b7cc),
	.w7(32'h3bbdfda8),
	.w8(32'h3c703b2c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc284a),
	.w1(32'h3b0f1b69),
	.w2(32'h3ba0a7ca),
	.w3(32'hbca62bdb),
	.w4(32'h3aeb218a),
	.w5(32'h3abe7bf9),
	.w6(32'h3ada7b02),
	.w7(32'h3bbbf162),
	.w8(32'hbb0d8705),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9c365),
	.w1(32'h3bb8926c),
	.w2(32'hbc57c0f6),
	.w3(32'h3b85a09d),
	.w4(32'hbc452919),
	.w5(32'hbbaf4de7),
	.w6(32'hbb363721),
	.w7(32'hbc018cd1),
	.w8(32'hbc53e058),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8014d8),
	.w1(32'hbbf60a1c),
	.w2(32'h3d03d82a),
	.w3(32'hba1b7369),
	.w4(32'h3bc8e04a),
	.w5(32'hbc80d4c9),
	.w6(32'hbc2022b0),
	.w7(32'hbc7be08d),
	.w8(32'hbc1bdd34),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac9ca5),
	.w1(32'h3b6247c6),
	.w2(32'h3b17c4ce),
	.w3(32'hba489e28),
	.w4(32'hbbbcc61d),
	.w5(32'h3b40dded),
	.w6(32'hbb152e59),
	.w7(32'h3d030da9),
	.w8(32'h39338bbc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67c477),
	.w1(32'h3c316e4e),
	.w2(32'hbc61ebd4),
	.w3(32'h38b38fa4),
	.w4(32'h3b6417c6),
	.w5(32'hbb3f7dd7),
	.w6(32'h3c69f8aa),
	.w7(32'h3d1061ed),
	.w8(32'h39e0a732),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafbfce),
	.w1(32'hbb15b15d),
	.w2(32'h3c86f12e),
	.w3(32'hbbe4cd4a),
	.w4(32'h3c8b0f29),
	.w5(32'h3bd4ef0d),
	.w6(32'h3c581933),
	.w7(32'h3d221be6),
	.w8(32'hb99ceb08),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16e8ec),
	.w1(32'h3b64fe72),
	.w2(32'hbb556d64),
	.w3(32'h3c15b45c),
	.w4(32'hbb0fe9d9),
	.w5(32'h3b97f4f4),
	.w6(32'hba867880),
	.w7(32'h3c32a16f),
	.w8(32'h3ba7619a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd612b9),
	.w1(32'hbbb8ee2e),
	.w2(32'hbb697047),
	.w3(32'h3b24035a),
	.w4(32'h3ba0ccaf),
	.w5(32'hbc871ac3),
	.w6(32'h3743d234),
	.w7(32'hbb5ab2e6),
	.w8(32'h3bcf3f84),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf0f96),
	.w1(32'hbc2ffa19),
	.w2(32'hbab3b8cc),
	.w3(32'hbc4c8b8b),
	.w4(32'h3b98fdbf),
	.w5(32'h3c4b8d0c),
	.w6(32'hbba1e9c5),
	.w7(32'hbc25de94),
	.w8(32'hbc409e72),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe18b5),
	.w1(32'h3b35ffa1),
	.w2(32'hbc1d1653),
	.w3(32'hbb9b8aa6),
	.w4(32'hbc0905cb),
	.w5(32'h3bedf960),
	.w6(32'hba1ef857),
	.w7(32'hb9a40332),
	.w8(32'hbbbb817c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7b2d7),
	.w1(32'hbc0c326b),
	.w2(32'hbbdff339),
	.w3(32'hbaa9daae),
	.w4(32'hbbb3a930),
	.w5(32'hbb84675c),
	.w6(32'hba282c77),
	.w7(32'h3ae7fe07),
	.w8(32'hba38171d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55820f),
	.w1(32'h3cba4c6c),
	.w2(32'h3bbe983d),
	.w3(32'h38bdd7a2),
	.w4(32'hbb9741b1),
	.w5(32'h3b0a7e1e),
	.w6(32'hbd3896a0),
	.w7(32'hbb808117),
	.w8(32'h3c4b0412),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac06ac5),
	.w1(32'hbafcbd1c),
	.w2(32'hbbc0e216),
	.w3(32'hbc2d6eaf),
	.w4(32'hbb895c7d),
	.w5(32'hbb9be737),
	.w6(32'hbbb94ec0),
	.w7(32'hbc634732),
	.w8(32'hba2d2547),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49e17c),
	.w1(32'hbc10fb9c),
	.w2(32'hbc5bbd68),
	.w3(32'hbc0289ab),
	.w4(32'h3cb681f6),
	.w5(32'hbbf928e9),
	.w6(32'hbbf762b8),
	.w7(32'h3cf22e8a),
	.w8(32'hb9b1152e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55315e),
	.w1(32'hbc9a874f),
	.w2(32'hbb077e15),
	.w3(32'hbb1aabf8),
	.w4(32'h3ad8d46d),
	.w5(32'h3926fc8d),
	.w6(32'hbaed4ef8),
	.w7(32'h3ca5288a),
	.w8(32'hbc4f16b3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a141),
	.w1(32'hbb033abb),
	.w2(32'hbc251f00),
	.w3(32'hbc307a96),
	.w4(32'h3b97e735),
	.w5(32'h3a433008),
	.w6(32'h3c3cf811),
	.w7(32'hbba71427),
	.w8(32'h3b94eef5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11b403),
	.w1(32'hba94a3a4),
	.w2(32'h3c50dc75),
	.w3(32'hbb423787),
	.w4(32'hba452b69),
	.w5(32'h3bdadba1),
	.w6(32'h3aa534d0),
	.w7(32'hbbf66799),
	.w8(32'hbc3292c5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc373271),
	.w1(32'h3b4c103b),
	.w2(32'hbc27c6ee),
	.w3(32'hbc39e84d),
	.w4(32'hbc1a9c70),
	.w5(32'h3ab0a1e8),
	.w6(32'h3b1ec532),
	.w7(32'hbba6b8b0),
	.w8(32'h3c7fe3d5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dbf27),
	.w1(32'h3bcc985c),
	.w2(32'h39bf6d7d),
	.w3(32'hbaad02e9),
	.w4(32'h3cb6b58d),
	.w5(32'hbcbb8d7b),
	.w6(32'hbc49c238),
	.w7(32'hbc16272d),
	.w8(32'hbb59213e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e3de0),
	.w1(32'hbb76852b),
	.w2(32'h3b830b21),
	.w3(32'hbaf5a71a),
	.w4(32'hbb1dcb7b),
	.w5(32'h3c55da15),
	.w6(32'h3cd79171),
	.w7(32'h3c32a061),
	.w8(32'h3c14e3af),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3deba),
	.w1(32'hbc3fafff),
	.w2(32'hba4f41f1),
	.w3(32'h3c9dbe8d),
	.w4(32'hbbc8de96),
	.w5(32'h3a57ace0),
	.w6(32'hbb922de1),
	.w7(32'hb9b361e1),
	.w8(32'h39fb269e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3979af),
	.w1(32'hbbd16244),
	.w2(32'h3a2aeafd),
	.w3(32'hbab0bf45),
	.w4(32'hbaeda05c),
	.w5(32'h3be2265d),
	.w6(32'hbab9f27c),
	.w7(32'h3aac28c3),
	.w8(32'h3ac01714),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca69d8a),
	.w1(32'h39343169),
	.w2(32'hbb8001ab),
	.w3(32'hbc3b54d7),
	.w4(32'h3b6da6e8),
	.w5(32'hbc33910d),
	.w6(32'h3ae293a9),
	.w7(32'hbc635ec9),
	.w8(32'hbbad3060),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedc056),
	.w1(32'h3c425a9c),
	.w2(32'h3c39b13d),
	.w3(32'hbb98a5cc),
	.w4(32'hbcdab57b),
	.w5(32'hbb400abc),
	.w6(32'h3ba8ab73),
	.w7(32'hbc16d9f7),
	.w8(32'hbc28bc00),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10b6bf),
	.w1(32'h3cd54179),
	.w2(32'hbc1d4129),
	.w3(32'hbba3f132),
	.w4(32'hbbe14fb2),
	.w5(32'h3b84e5eb),
	.w6(32'h3ae3ebb0),
	.w7(32'hbb2f519e),
	.w8(32'h3c021cba),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c96e7),
	.w1(32'hbc591c39),
	.w2(32'hbbeb0b90),
	.w3(32'hbb0ad2c4),
	.w4(32'hbc33824c),
	.w5(32'hb7edbb50),
	.w6(32'h3a8f0dc3),
	.w7(32'h3bc10abb),
	.w8(32'hbc2fb5ef),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8e3bd),
	.w1(32'hbc0945c3),
	.w2(32'hbc33338f),
	.w3(32'hbb823e70),
	.w4(32'hbc37a0fb),
	.w5(32'hbb224be0),
	.w6(32'hbb1192ef),
	.w7(32'hbb1f07f8),
	.w8(32'h3c66cba7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35cd6c),
	.w1(32'hbb8a45d3),
	.w2(32'hbbce3888),
	.w3(32'h3b163d12),
	.w4(32'hbb48c47d),
	.w5(32'hbbee2e0b),
	.w6(32'h3c186d21),
	.w7(32'hbc0b3ca1),
	.w8(32'hbb675d7f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac60f09),
	.w1(32'hbc6b0f59),
	.w2(32'hbade9ca7),
	.w3(32'hbc8f47a6),
	.w4(32'h3cb1101d),
	.w5(32'h39133b2c),
	.w6(32'hbc90e340),
	.w7(32'h3c67f54b),
	.w8(32'hbc489a21),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b7f6f),
	.w1(32'hbc8b02cb),
	.w2(32'hbbad671c),
	.w3(32'h3a9bae61),
	.w4(32'hbbdc4277),
	.w5(32'h3b852b88),
	.w6(32'h3afd2a0d),
	.w7(32'hbabe4e03),
	.w8(32'hbbdd9fa6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fe950),
	.w1(32'h3b71b6cd),
	.w2(32'hbbd7bf4c),
	.w3(32'hbb60651a),
	.w4(32'h3b787aa9),
	.w5(32'hbc6bafe2),
	.w6(32'hbc76af5f),
	.w7(32'h3a138f92),
	.w8(32'hbc7cec70),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc035482),
	.w1(32'hbb0cf537),
	.w2(32'h3b2ef7a7),
	.w3(32'hbc2ed8df),
	.w4(32'h3cb93aef),
	.w5(32'hbb322468),
	.w6(32'hbbb68999),
	.w7(32'hbb0ca96e),
	.w8(32'hbc9b6828),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5da5),
	.w1(32'hbaa1df27),
	.w2(32'hb916dcfb),
	.w3(32'hbb7eebf0),
	.w4(32'h3b02bfd1),
	.w5(32'hbbf1a57b),
	.w6(32'h3c4c9dfc),
	.w7(32'h3a5706cf),
	.w8(32'hbc3204b9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c8992),
	.w1(32'hbc23b4a3),
	.w2(32'hbcbf9402),
	.w3(32'hba01abd2),
	.w4(32'hbb9e4a92),
	.w5(32'hbcb35cea),
	.w6(32'hbb847e49),
	.w7(32'h3d14a70b),
	.w8(32'h3d21bb18),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c707f0c),
	.w1(32'hbc84faad),
	.w2(32'h3bfa656f),
	.w3(32'hbc4ab3ef),
	.w4(32'h3cb35a39),
	.w5(32'h3be9c2b7),
	.w6(32'hbc0e4e27),
	.w7(32'h3bc6ad48),
	.w8(32'h3b90eb6d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86f1f9),
	.w1(32'hbb4007fe),
	.w2(32'hbca4641c),
	.w3(32'h3c0d2cf4),
	.w4(32'hbbdb8327),
	.w5(32'h3b0d72fb),
	.w6(32'hbb1c7b9a),
	.w7(32'hbb4927df),
	.w8(32'h3ab619ea),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e913f),
	.w1(32'h3af02c56),
	.w2(32'hb9406be9),
	.w3(32'hbcec5fba),
	.w4(32'hbca705b3),
	.w5(32'hbb1066d6),
	.w6(32'hbaf9ec8b),
	.w7(32'hbcc8b32e),
	.w8(32'h3c3b7b38),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbdc924),
	.w1(32'hbc8c5a23),
	.w2(32'h3c0af1e6),
	.w3(32'hbb72720d),
	.w4(32'hbc915990),
	.w5(32'hbc90fb35),
	.w6(32'hbcc37dbf),
	.w7(32'h3b95f74f),
	.w8(32'hbbc33b91),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc514100),
	.w1(32'hbc1b1a42),
	.w2(32'hbc7ebbdf),
	.w3(32'hbc655132),
	.w4(32'hba72f444),
	.w5(32'hbc85cdf0),
	.w6(32'hbbed9b23),
	.w7(32'h3b2abde9),
	.w8(32'hbc7f6d76),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba624b3f),
	.w1(32'h3806d98b),
	.w2(32'hbb4b2354),
	.w3(32'h3bae0490),
	.w4(32'hbb8352db),
	.w5(32'hbb8bcd80),
	.w6(32'h3bc06a29),
	.w7(32'h3b32d5eb),
	.w8(32'hbc18623a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba39f87),
	.w1(32'hba2b7d20),
	.w2(32'hbad61ca0),
	.w3(32'h3bbbb9e9),
	.w4(32'hbb7a64e4),
	.w5(32'hbbf7dbb5),
	.w6(32'hbbe2f6e7),
	.w7(32'h3d209e71),
	.w8(32'h3bf8d7ba),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2812cd),
	.w1(32'h3a32c3eb),
	.w2(32'h3d1d293c),
	.w3(32'hbcbb3d93),
	.w4(32'hbcd9a069),
	.w5(32'hbc855f71),
	.w6(32'h3b0ec457),
	.w7(32'hbba2fb45),
	.w8(32'h3d280751),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af10369),
	.w1(32'hbbf5876a),
	.w2(32'h39ad6102),
	.w3(32'h3c95b382),
	.w4(32'h3b629613),
	.w5(32'h3b1f2042),
	.w6(32'h3b8350c2),
	.w7(32'hbbf43cb7),
	.w8(32'hbb210726),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e9272),
	.w1(32'hbc970090),
	.w2(32'h3c0304af),
	.w3(32'hbc0b5b0d),
	.w4(32'h3ba4410b),
	.w5(32'hb9b01306),
	.w6(32'h3aac2ba0),
	.w7(32'hbc18c70b),
	.w8(32'h398503c8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1fe42),
	.w1(32'hbb6ff66a),
	.w2(32'hbbdd6107),
	.w3(32'hba55fdc7),
	.w4(32'hbb92581f),
	.w5(32'h3b4933db),
	.w6(32'hb9a531a9),
	.w7(32'hbb8d9118),
	.w8(32'hbb271ad0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56aeaf),
	.w1(32'hbb97bd35),
	.w2(32'hbb863ba7),
	.w3(32'hbb4a8f73),
	.w4(32'hbca31738),
	.w5(32'h3cebc019),
	.w6(32'hbcc245f9),
	.w7(32'h3bb7aeb3),
	.w8(32'hbce87455),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c531744),
	.w1(32'hbbecc011),
	.w2(32'hb9a60402),
	.w3(32'hbc35c46c),
	.w4(32'h3c778c8d),
	.w5(32'h3b6116f9),
	.w6(32'hbcaac93d),
	.w7(32'h3a6b64cd),
	.w8(32'hbd1187f0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03a4af),
	.w1(32'hbc99a76e),
	.w2(32'h3c1a9c51),
	.w3(32'h3b40dffa),
	.w4(32'hbbadf89e),
	.w5(32'h3c44d637),
	.w6(32'h3c00bf3e),
	.w7(32'h3a0673d0),
	.w8(32'h3c9cc90a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e734f),
	.w1(32'hbb301175),
	.w2(32'h3ce64dad),
	.w3(32'hbaa6bfec),
	.w4(32'hb9a97c77),
	.w5(32'hbd09ef36),
	.w6(32'h3d10a55f),
	.w7(32'h3b7a587c),
	.w8(32'h3b11f45c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4171c8),
	.w1(32'hba08fb40),
	.w2(32'h3ce2412d),
	.w3(32'h3cf6164b),
	.w4(32'hbb7c863c),
	.w5(32'hb8ede919),
	.w6(32'hb92fe8c4),
	.w7(32'hbb89f352),
	.w8(32'h3c075d17),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace2a7b),
	.w1(32'hba94b31e),
	.w2(32'hbb818697),
	.w3(32'hba6020ed),
	.w4(32'h3b5f7c42),
	.w5(32'hbc373931),
	.w6(32'hbbfc958f),
	.w7(32'hbac93745),
	.w8(32'hbb55f3bc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2936f),
	.w1(32'hb73bfae1),
	.w2(32'hbbb4ab3f),
	.w3(32'h3b8d1f19),
	.w4(32'hbc9c383e),
	.w5(32'hbc2104c7),
	.w6(32'hbccc4607),
	.w7(32'h3b81be01),
	.w8(32'h3bdd2853),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc187e7),
	.w1(32'h3a71b9d9),
	.w2(32'hbb9be809),
	.w3(32'hbc1575a8),
	.w4(32'h3bfabf1d),
	.w5(32'h3c7ba969),
	.w6(32'hbb94fe29),
	.w7(32'h3c8e89d3),
	.w8(32'hbc747d41),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1443b7),
	.w1(32'hbb9b1bb2),
	.w2(32'h3bd7dc90),
	.w3(32'hbcb58538),
	.w4(32'h3c183188),
	.w5(32'h3a863659),
	.w6(32'hbc4ab104),
	.w7(32'h3a99e3d1),
	.w8(32'h3b805701),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8411a3),
	.w1(32'hbbd7fb96),
	.w2(32'h3bb0c437),
	.w3(32'hbc0fa106),
	.w4(32'hbc08736c),
	.w5(32'h3a4f9efa),
	.w6(32'hbc0ecc5e),
	.w7(32'h37ebc232),
	.w8(32'h3c10c4f0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8740bf),
	.w1(32'hbc9831c1),
	.w2(32'hbb052dbb),
	.w3(32'h3d064a51),
	.w4(32'h3b14fbb5),
	.w5(32'hb999b77f),
	.w6(32'hbbbd7004),
	.w7(32'h3c1ac84a),
	.w8(32'h3c94d47f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49129a),
	.w1(32'hbb0090b5),
	.w2(32'hbb7e0357),
	.w3(32'h3ac76bdd),
	.w4(32'h3bad1929),
	.w5(32'h3a1c9dd9),
	.w6(32'h3c8a4511),
	.w7(32'hbbfeb31f),
	.w8(32'h3c148dac),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7018bb),
	.w1(32'hbae82728),
	.w2(32'hbc1c112f),
	.w3(32'hbbda0ec6),
	.w4(32'hbc119341),
	.w5(32'hbbcb3bae),
	.w6(32'h3bba9362),
	.w7(32'h3b4d1d91),
	.w8(32'hbc742128),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248a53),
	.w1(32'hbbbca37d),
	.w2(32'hbc3170f9),
	.w3(32'hbc12500a),
	.w4(32'hbca6e236),
	.w5(32'hbc1a4621),
	.w6(32'h3b5dba43),
	.w7(32'h3bc593bc),
	.w8(32'h3bf023c2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd75c2),
	.w1(32'hbc43471b),
	.w2(32'hbb906bc6),
	.w3(32'hbbe7f26c),
	.w4(32'hbb57d9f9),
	.w5(32'h3bdaaff9),
	.w6(32'h3d1bf933),
	.w7(32'hbc4c7355),
	.w8(32'hbc08b7c5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6bef7),
	.w1(32'hba2f629c),
	.w2(32'h3d10d4fa),
	.w3(32'hbbc4da88),
	.w4(32'hbb630fc3),
	.w5(32'hbbafda3f),
	.w6(32'h3bdd19ef),
	.w7(32'h3bc40948),
	.w8(32'hbb545bad),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab39512),
	.w1(32'hbbba6cb1),
	.w2(32'hbb8fe148),
	.w3(32'h3c290347),
	.w4(32'hbb97f103),
	.w5(32'hbc17aa97),
	.w6(32'hbc042b74),
	.w7(32'h3c126f33),
	.w8(32'h3c35d636),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2ce2a),
	.w1(32'h39f11312),
	.w2(32'hbbabb27c),
	.w3(32'hbb77f8fa),
	.w4(32'h3b767119),
	.w5(32'hbaa22c4f),
	.w6(32'h3c05a6c6),
	.w7(32'h3c45cb72),
	.w8(32'h3b9bfecf),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad19db7),
	.w1(32'hb89fa9c1),
	.w2(32'hbc234b1c),
	.w3(32'hbbd9d192),
	.w4(32'hbbbbf91c),
	.w5(32'hbc3be34b),
	.w6(32'h3a53c7ac),
	.w7(32'h3b6202da),
	.w8(32'h3b9dc841),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ad8e4),
	.w1(32'hbbcf467b),
	.w2(32'h3bd409f3),
	.w3(32'h3b2c36a1),
	.w4(32'hbb0cc5b3),
	.w5(32'hbb9804f4),
	.w6(32'h3c408563),
	.w7(32'hbbddbe40),
	.w8(32'h39a79e8d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed4be1),
	.w1(32'h3c54d5a6),
	.w2(32'h3bab4b20),
	.w3(32'hbb37d53d),
	.w4(32'hbb638750),
	.w5(32'hbc1af5fc),
	.w6(32'hbb14fab0),
	.w7(32'hbb328fac),
	.w8(32'h3d82171f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b721a4c),
	.w1(32'h393b7ea0),
	.w2(32'h3b20bea5),
	.w3(32'hb9ff061e),
	.w4(32'h3c291d75),
	.w5(32'hbbf58842),
	.w6(32'hbc707821),
	.w7(32'h3b86fc82),
	.w8(32'h38bba3bb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb577d1c),
	.w1(32'hba7bccae),
	.w2(32'h3acf1d6a),
	.w3(32'hbd1450f3),
	.w4(32'hba5dd743),
	.w5(32'h391e6262),
	.w6(32'h3b5a57f5),
	.w7(32'hbb06392d),
	.w8(32'h3bcedbc0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ab105),
	.w1(32'h3b3b4d5c),
	.w2(32'h3c1ad7e1),
	.w3(32'hbcb3be30),
	.w4(32'hbb8474cf),
	.w5(32'hba939b7a),
	.w6(32'hbd439e7b),
	.w7(32'h3b199b44),
	.w8(32'hbbf07694),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb103da9),
	.w1(32'hbb27797c),
	.w2(32'hbc343266),
	.w3(32'hbbb2708b),
	.w4(32'hbb06056d),
	.w5(32'h3b32b1d7),
	.w6(32'hbcacc6dc),
	.w7(32'h3bc9c4ac),
	.w8(32'h3c181bf2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62bbd0),
	.w1(32'h3786b257),
	.w2(32'h3992fc65),
	.w3(32'h395ed55c),
	.w4(32'hbbcb1eea),
	.w5(32'hbb24405a),
	.w6(32'h3c3a634d),
	.w7(32'hbbf99425),
	.w8(32'hbb8e649b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9202ab),
	.w1(32'hbba2efbb),
	.w2(32'h39f3e2b0),
	.w3(32'h396a1702),
	.w4(32'hbbe656db),
	.w5(32'hbbc50101),
	.w6(32'hbc0573f3),
	.w7(32'h3ba2e2ba),
	.w8(32'h3aee5164),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cb9e4),
	.w1(32'h3cf9350d),
	.w2(32'h37454780),
	.w3(32'hbc2afac6),
	.w4(32'hbaece6c3),
	.w5(32'h3ad3d774),
	.w6(32'hbb9945ae),
	.w7(32'h3b018999),
	.w8(32'h3a716630),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7d76b),
	.w1(32'hbc3352f0),
	.w2(32'h3acd5fa2),
	.w3(32'h3a645731),
	.w4(32'hbc8057f3),
	.w5(32'h3c2bce96),
	.w6(32'h3a0d4e30),
	.w7(32'hbc44279d),
	.w8(32'hbb0305b9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8888fd),
	.w1(32'h3acc9a23),
	.w2(32'hbc439292),
	.w3(32'h3acc429b),
	.w4(32'hbbb50ca8),
	.w5(32'hbbf60d57),
	.w6(32'h3c177e53),
	.w7(32'hbb9f90a5),
	.w8(32'hbb24e5e2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4caf8),
	.w1(32'hbc8986fd),
	.w2(32'hbb714fa6),
	.w3(32'hb9b18970),
	.w4(32'h3b0407ca),
	.w5(32'hbbb13580),
	.w6(32'h3b3445b8),
	.w7(32'hbb9cea42),
	.w8(32'h3c30574b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35b040),
	.w1(32'h3b858d84),
	.w2(32'h395c03df),
	.w3(32'hbaf0f59f),
	.w4(32'h3c302255),
	.w5(32'hbb33f4f5),
	.w6(32'hbc29bd93),
	.w7(32'h3bed6981),
	.w8(32'hbcfbb63f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc20436),
	.w1(32'h3bb61832),
	.w2(32'hbb1c4917),
	.w3(32'h3bc0fdd5),
	.w4(32'hbb7f0d12),
	.w5(32'h3b354348),
	.w6(32'hbc4ea93c),
	.w7(32'h3b2e1a93),
	.w8(32'hbb056618),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d9744),
	.w1(32'hbb4d1427),
	.w2(32'h3b935434),
	.w3(32'hbbb30832),
	.w4(32'hbb18d2a2),
	.w5(32'hba5e105f),
	.w6(32'h3b1fa3e5),
	.w7(32'h3820f8dc),
	.w8(32'h3a557034),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f38ff),
	.w1(32'h3c17a1ac),
	.w2(32'h3c745c20),
	.w3(32'hbc5d3fa6),
	.w4(32'h3be25e72),
	.w5(32'hbc9fae2e),
	.w6(32'hbbb36996),
	.w7(32'hbbffd047),
	.w8(32'hbabf9cbd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc014bd6),
	.w1(32'h3b4abfc3),
	.w2(32'h3b870ce2),
	.w3(32'hbbb60a8c),
	.w4(32'h3acfaebe),
	.w5(32'hbb8c2630),
	.w6(32'h3baa504c),
	.w7(32'hbb409d55),
	.w8(32'hbb97ef55),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e01c5),
	.w1(32'hbb28449e),
	.w2(32'h3c3c47b4),
	.w3(32'h3ba9c6a3),
	.w4(32'h3b0f3d2a),
	.w5(32'hba5be15c),
	.w6(32'h3c8ab2c2),
	.w7(32'hbc831bc2),
	.w8(32'h3a724fe3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3562b),
	.w1(32'h3b8318d4),
	.w2(32'hbc2e9165),
	.w3(32'hbbd3341f),
	.w4(32'hbba591fa),
	.w5(32'h3bba7473),
	.w6(32'hbc12a135),
	.w7(32'hbc0af950),
	.w8(32'hbc6c86d5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d34e2),
	.w1(32'hbba6497b),
	.w2(32'hbac14a42),
	.w3(32'h39171cd9),
	.w4(32'h3b9949f0),
	.w5(32'h3c8f1f59),
	.w6(32'h399f2968),
	.w7(32'hbb36a730),
	.w8(32'hbcc5ae90),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1480c9),
	.w1(32'hbb661cbf),
	.w2(32'hbae7faa8),
	.w3(32'hba4a9717),
	.w4(32'hbbae073e),
	.w5(32'hbbb52ac4),
	.w6(32'hbc1069cb),
	.w7(32'hbbe0d74e),
	.w8(32'h3bcfb55e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc198a22),
	.w1(32'hbb4b86f3),
	.w2(32'h3a4b6f5f),
	.w3(32'hbbfcccb9),
	.w4(32'hbbbdb421),
	.w5(32'hba9a1c84),
	.w6(32'hbbbe1371),
	.w7(32'hbb3e6769),
	.w8(32'hbbc2313b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc198496),
	.w1(32'h3b9daa3f),
	.w2(32'hba84cea6),
	.w3(32'hbb8fec18),
	.w4(32'hbae54c7a),
	.w5(32'h3b0ddea7),
	.w6(32'h3c15ad6c),
	.w7(32'hbbf25b1c),
	.w8(32'hbc6e4d08),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba069dd8),
	.w1(32'h3b76bab0),
	.w2(32'hbc7ec1f5),
	.w3(32'h3c018f4a),
	.w4(32'hbac29140),
	.w5(32'h3a458177),
	.w6(32'hbc0759b3),
	.w7(32'h3afc5518),
	.w8(32'h38db2e25),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa33a7),
	.w1(32'h3b7a201c),
	.w2(32'h3b82e7ae),
	.w3(32'hbc8c8d54),
	.w4(32'hbb4d677b),
	.w5(32'h3b5d04df),
	.w6(32'hbc244381),
	.w7(32'h3c11f3a3),
	.w8(32'h3b6ad69f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9c88a),
	.w1(32'hb8817cac),
	.w2(32'hbb89afee),
	.w3(32'hbc915574),
	.w4(32'h3a10f90f),
	.w5(32'hbb87bd0f),
	.w6(32'hbc2d5bb6),
	.w7(32'h3bc4fa61),
	.w8(32'hba4dba7c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d8c9c),
	.w1(32'hbc225dce),
	.w2(32'h3b94564e),
	.w3(32'h3b41a843),
	.w4(32'h3b04bce8),
	.w5(32'h3abe0cdb),
	.w6(32'hbbe0af0e),
	.w7(32'hbb18e097),
	.w8(32'hbbe0dba5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d00325),
	.w1(32'h3c1b8087),
	.w2(32'hbc074ddd),
	.w3(32'hbbf31390),
	.w4(32'h3ade5a91),
	.w5(32'hbbf7dcad),
	.w6(32'h3b86321b),
	.w7(32'h3bde4289),
	.w8(32'hbb965477),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fa596),
	.w1(32'hbb0c45fa),
	.w2(32'h3c268a6e),
	.w3(32'hbc01df09),
	.w4(32'hbbd167dd),
	.w5(32'h3b5a55a3),
	.w6(32'h3b0405b8),
	.w7(32'h3c8e4360),
	.w8(32'hbb4077da),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c722),
	.w1(32'hbc8e9326),
	.w2(32'hbc0089dc),
	.w3(32'h3b2f25bf),
	.w4(32'hbc2e9aa7),
	.w5(32'h39a6f826),
	.w6(32'hbb5489f8),
	.w7(32'h3a4e0e24),
	.w8(32'hbafeae87),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59863d),
	.w1(32'hbd386690),
	.w2(32'hbbd901d7),
	.w3(32'hbbc3214c),
	.w4(32'hbb8a51ec),
	.w5(32'h3c150a69),
	.w6(32'hbb3c0958),
	.w7(32'h3bd0aeb1),
	.w8(32'h3b97c4a3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba944237),
	.w1(32'h3abdc42e),
	.w2(32'h3b6c9f58),
	.w3(32'hbba6f7fb),
	.w4(32'h3c19489e),
	.w5(32'hba7469db),
	.w6(32'hbb7caaca),
	.w7(32'h3c2ae6f2),
	.w8(32'hbb44c8a3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9d4ee),
	.w1(32'h3c022f3a),
	.w2(32'h3d07fcce),
	.w3(32'h3b735e31),
	.w4(32'hba9d0ebc),
	.w5(32'hbb269ff6),
	.w6(32'hb933514d),
	.w7(32'hbc8f76b9),
	.w8(32'hbb8d5538),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfabc0),
	.w1(32'h3bf306e3),
	.w2(32'h3c3d1a23),
	.w3(32'h3b0df806),
	.w4(32'h3a66c256),
	.w5(32'hbb2c8093),
	.w6(32'h3c2452e7),
	.w7(32'h3b4bef14),
	.w8(32'hbb87ef1a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc68825),
	.w1(32'h3c0b5d94),
	.w2(32'hbc521cd3),
	.w3(32'h3bb83d92),
	.w4(32'h3be44db8),
	.w5(32'h3ac835f8),
	.w6(32'h3ba36dd1),
	.w7(32'hbc0b00e8),
	.w8(32'hbc708dd7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d38bf),
	.w1(32'hbad590aa),
	.w2(32'h3affeeb2),
	.w3(32'hba4c0132),
	.w4(32'hbafb4e92),
	.w5(32'hbb3d83d6),
	.w6(32'h3afec560),
	.w7(32'h3abddfad),
	.w8(32'hbbc75313),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f7f7d),
	.w1(32'hbba7fe66),
	.w2(32'hb960dde9),
	.w3(32'hbbaded6b),
	.w4(32'h3860d514),
	.w5(32'hbbe3b7a5),
	.w6(32'hbb5faedc),
	.w7(32'h3bbb0f21),
	.w8(32'hbb7fda81),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5accdf),
	.w1(32'hbbb50bbb),
	.w2(32'h3c4080d5),
	.w3(32'h39e4c724),
	.w4(32'hbaab5bee),
	.w5(32'hbabfc926),
	.w6(32'hbb11a042),
	.w7(32'h3b6de3fc),
	.w8(32'hbc70d550),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd112c),
	.w1(32'h3bbc1752),
	.w2(32'h3b65ce2b),
	.w3(32'hb9a590bf),
	.w4(32'hbaafb780),
	.w5(32'hbc342df3),
	.w6(32'h3b0b88d6),
	.w7(32'hbb0ebffd),
	.w8(32'h3a8ad9e9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c367880),
	.w1(32'h3aaedb51),
	.w2(32'h3a37f4a7),
	.w3(32'hbbb4736a),
	.w4(32'hbbf20a75),
	.w5(32'hb94922f6),
	.w6(32'h3c22a09f),
	.w7(32'hbaa16931),
	.w8(32'h3ad49f43),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9766a8),
	.w1(32'hbc0d6758),
	.w2(32'h3b8961c2),
	.w3(32'hbc6628b2),
	.w4(32'hb8ee5189),
	.w5(32'hbb9e9c4f),
	.w6(32'h3bc4e5e6),
	.w7(32'h3bc020fa),
	.w8(32'hbb03e151),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10900a),
	.w1(32'hbc6e4845),
	.w2(32'h3c0f1913),
	.w3(32'hbb0ed1e6),
	.w4(32'h3c3c2206),
	.w5(32'h3a4664dd),
	.w6(32'hbb974f13),
	.w7(32'h3ac09a91),
	.w8(32'h3911242a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073dc6),
	.w1(32'hbbd9c2f2),
	.w2(32'h39f48e9d),
	.w3(32'hbab21bfa),
	.w4(32'hbc0966cb),
	.w5(32'hbbd3ec3f),
	.w6(32'h3af9b63f),
	.w7(32'h3c054042),
	.w8(32'hba39f2f3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b48e7),
	.w1(32'h3a9c9ce4),
	.w2(32'hbb903d23),
	.w3(32'h3b67cd1d),
	.w4(32'hbc5ac107),
	.w5(32'hbb7e766f),
	.w6(32'hbbb97e0d),
	.w7(32'hbae0e7c1),
	.w8(32'hbaf6a6c3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba615317),
	.w1(32'hbc422a5c),
	.w2(32'hbbceca40),
	.w3(32'hbb918781),
	.w4(32'hbc50c2d1),
	.w5(32'hbbfe4bb8),
	.w6(32'hbc17e3bf),
	.w7(32'hba4c1d4b),
	.w8(32'h3ab3b608),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4e1b5),
	.w1(32'h3b18613b),
	.w2(32'hbc206645),
	.w3(32'hbcc44f3b),
	.w4(32'h3bbcbda4),
	.w5(32'hbbb7f6d2),
	.w6(32'hbb408173),
	.w7(32'hbc641a70),
	.w8(32'hbb328430),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbc0ed),
	.w1(32'h3c19e352),
	.w2(32'h3c23e1c4),
	.w3(32'hbc97e398),
	.w4(32'hbb3b27c7),
	.w5(32'hba500a6b),
	.w6(32'hbc6df481),
	.w7(32'hbc2771ea),
	.w8(32'h3b188635),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94642c),
	.w1(32'h3c9375d7),
	.w2(32'h3959d7ee),
	.w3(32'h3ae240ae),
	.w4(32'h3b16afc0),
	.w5(32'h3c5ffbbf),
	.w6(32'h3c22ba41),
	.w7(32'h3ac08036),
	.w8(32'hbc00591e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75e4ff),
	.w1(32'hbc502905),
	.w2(32'h3a82f495),
	.w3(32'hbc0b8a36),
	.w4(32'hbc0328d8),
	.w5(32'h3d01d198),
	.w6(32'hbcb5d9d2),
	.w7(32'h3a2fac02),
	.w8(32'h3d3e62b8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c595c68),
	.w1(32'h3c40a71a),
	.w2(32'hbc46e204),
	.w3(32'hbb005971),
	.w4(32'hbc1e353e),
	.w5(32'h3bc3497e),
	.w6(32'h3b0915fc),
	.w7(32'h3c13a938),
	.w8(32'h3a84140c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bd346),
	.w1(32'hbc16d68c),
	.w2(32'hbc635091),
	.w3(32'hbbef8cbc),
	.w4(32'hbba09b3e),
	.w5(32'hbb7b2704),
	.w6(32'h3a693bce),
	.w7(32'h3c1e4789),
	.w8(32'h3a2eeebc),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fdb98),
	.w1(32'h3be23af8),
	.w2(32'h3abf07b2),
	.w3(32'h3a63f2e5),
	.w4(32'hbacf1ae6),
	.w5(32'h3a9e0812),
	.w6(32'h37dbcd1d),
	.w7(32'hbbe8ce36),
	.w8(32'hbc1c0360),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8adb6),
	.w1(32'hbce29d88),
	.w2(32'hbc183b72),
	.w3(32'hb97d1e56),
	.w4(32'h3c0b6425),
	.w5(32'hbc498606),
	.w6(32'h3cdce420),
	.w7(32'hbc3e1a1b),
	.w8(32'hbc5b6450),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bc321),
	.w1(32'h3b1736d9),
	.w2(32'hbb71e51b),
	.w3(32'h3b6f6188),
	.w4(32'hbb118869),
	.w5(32'hbbeb8f35),
	.w6(32'hba35270a),
	.w7(32'hbc0a975f),
	.w8(32'h39289593),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb453a8b),
	.w1(32'h3a14df45),
	.w2(32'h3b093014),
	.w3(32'h3d01ff9f),
	.w4(32'h3cc483e6),
	.w5(32'hbbd08aaf),
	.w6(32'h3adb088b),
	.w7(32'hba9a9279),
	.w8(32'h3c6df472),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fc0ca),
	.w1(32'hbc631bb1),
	.w2(32'h3b4b4ed7),
	.w3(32'h3adada91),
	.w4(32'hbba5f5ba),
	.w5(32'hbbf299aa),
	.w6(32'hbcce0448),
	.w7(32'h3c9592d5),
	.w8(32'h3c730c10),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ab473),
	.w1(32'h3b1a11ec),
	.w2(32'h3b1467c9),
	.w3(32'hbc8bd973),
	.w4(32'h3c1a5f9c),
	.w5(32'h3b406a16),
	.w6(32'h3cc55d99),
	.w7(32'h3c5e88b0),
	.w8(32'hbb4f2f28),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88e2e),
	.w1(32'hbbf3a7ca),
	.w2(32'hbb4ee0c7),
	.w3(32'hbb97e1d7),
	.w4(32'h3c43706a),
	.w5(32'hbb8edc07),
	.w6(32'hbc7e5967),
	.w7(32'hbcaf1947),
	.w8(32'hbb95c6a0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1c141),
	.w1(32'h3c0503f2),
	.w2(32'hbc0ec511),
	.w3(32'hbc07aec1),
	.w4(32'hba6f1009),
	.w5(32'h3c1d469a),
	.w6(32'hbbcdce70),
	.w7(32'hb9892839),
	.w8(32'hbab0a68e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7c83d),
	.w1(32'hbbcc42b2),
	.w2(32'hbc138f23),
	.w3(32'hbb8246ae),
	.w4(32'hba99129a),
	.w5(32'hbbce87c7),
	.w6(32'h3c3da347),
	.w7(32'h3bb359f3),
	.w8(32'h3ae342b3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc459c4),
	.w1(32'hbbafb77f),
	.w2(32'hb9c62d8e),
	.w3(32'h3b277ed0),
	.w4(32'h3c9d2aca),
	.w5(32'h3c447b19),
	.w6(32'h3c2e7468),
	.w7(32'hbb86af3b),
	.w8(32'h3a76b9ea),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0a77d),
	.w1(32'hbaebd725),
	.w2(32'hbb25bd88),
	.w3(32'hbc004b83),
	.w4(32'hbba52fea),
	.w5(32'h3c34e059),
	.w6(32'hbb81b0f0),
	.w7(32'h3b94f51d),
	.w8(32'hbcee3962),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f6138),
	.w1(32'h3d04f189),
	.w2(32'h3baccb12),
	.w3(32'hbbcb53d6),
	.w4(32'hbc0e6b0e),
	.w5(32'h3a1879a8),
	.w6(32'hba08f8ae),
	.w7(32'hbbb9e07f),
	.w8(32'h3c6904dc),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b1e0f),
	.w1(32'hbaf5d62b),
	.w2(32'hba18c970),
	.w3(32'h3cb024c1),
	.w4(32'hbba3b441),
	.w5(32'h3bd61cf6),
	.w6(32'h3b85d2b6),
	.w7(32'hbc17c838),
	.w8(32'hbbb945a7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36cf66),
	.w1(32'hbc6c4224),
	.w2(32'hbbe970b7),
	.w3(32'hbc896cbc),
	.w4(32'h3bddc51e),
	.w5(32'hbc304333),
	.w6(32'h3be58c35),
	.w7(32'h3a60a56d),
	.w8(32'h3aeb787f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc358439),
	.w1(32'h3c095ca2),
	.w2(32'h38c216b8),
	.w3(32'hbc8285db),
	.w4(32'h3b9f9b8b),
	.w5(32'h3bef1bdf),
	.w6(32'h3c06775b),
	.w7(32'h39417511),
	.w8(32'h3b08e4ee),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5302fd),
	.w1(32'h3c949fc4),
	.w2(32'h3b20673d),
	.w3(32'hbaeabb35),
	.w4(32'hbb2f1fcd),
	.w5(32'hbc1a14b7),
	.w6(32'hbb1c95c6),
	.w7(32'hbc13afda),
	.w8(32'h3a9f06f8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c005b),
	.w1(32'hbb90ffb0),
	.w2(32'hbab58c1b),
	.w3(32'hbb823dec),
	.w4(32'hbb8f7cc1),
	.w5(32'h3bcfdfee),
	.w6(32'h3c16981b),
	.w7(32'hbc91d1c4),
	.w8(32'hbd08c76b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c692ef6),
	.w1(32'hbaa66082),
	.w2(32'hba75d760),
	.w3(32'h3be4229c),
	.w4(32'hbcba988b),
	.w5(32'hbc678a4b),
	.w6(32'h3b83dd29),
	.w7(32'hb9cf305f),
	.w8(32'h3ab625a0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d85e),
	.w1(32'h3c17bc44),
	.w2(32'hbb8379e7),
	.w3(32'h3c5cd0ee),
	.w4(32'hbb6af6dc),
	.w5(32'hbb25ad0f),
	.w6(32'h39b197c6),
	.w7(32'hbc5d8bd3),
	.w8(32'hbc236638),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8b177),
	.w1(32'h3bf3a20d),
	.w2(32'h3a924fc9),
	.w3(32'hbc5399ee),
	.w4(32'h3c110ff9),
	.w5(32'h3a5a7668),
	.w6(32'h3b9f335e),
	.w7(32'h3a35a784),
	.w8(32'hbcb705b3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a5622),
	.w1(32'h3b97378f),
	.w2(32'h3c4fe728),
	.w3(32'h3c12d475),
	.w4(32'h3a99c932),
	.w5(32'hbc4cde73),
	.w6(32'hbc819ecb),
	.w7(32'h3b669663),
	.w8(32'hbbdbc37c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad89c29),
	.w1(32'hb8e48a6b),
	.w2(32'hbc2b25c5),
	.w3(32'hbc9f0f9e),
	.w4(32'h3bbf7425),
	.w5(32'h3b313d28),
	.w6(32'hbbfb5a71),
	.w7(32'hbb7084ba),
	.w8(32'hbc1691c2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedb0bb),
	.w1(32'hbbfb7a4c),
	.w2(32'h3b76d292),
	.w3(32'h3a607876),
	.w4(32'hbb8c2567),
	.w5(32'hbb774f18),
	.w6(32'hbbaa0d0d),
	.w7(32'hbb2f2f04),
	.w8(32'hbaf5588e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea92de),
	.w1(32'h3acb6271),
	.w2(32'hbbb58227),
	.w3(32'hbb309019),
	.w4(32'hbc92f0c7),
	.w5(32'h3bd4d95f),
	.w6(32'hbc57daa7),
	.w7(32'hbbe0b744),
	.w8(32'hbb0759a6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117032),
	.w1(32'h3a798c73),
	.w2(32'h3bb7a896),
	.w3(32'h3ba2f203),
	.w4(32'h3c9a596a),
	.w5(32'hbbc9a3d5),
	.w6(32'h3b7450e2),
	.w7(32'hb9857e42),
	.w8(32'hbb61dcc1),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eaa13),
	.w1(32'hb9da4079),
	.w2(32'hbc86b1bd),
	.w3(32'hbacf64fe),
	.w4(32'hbc277381),
	.w5(32'h3cbfbe89),
	.w6(32'hbc1f31da),
	.w7(32'h3c4e2b5f),
	.w8(32'hba2385fe),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb606074),
	.w1(32'hbbcd453c),
	.w2(32'hbb78cb80),
	.w3(32'hbbbf4ef4),
	.w4(32'h3c250b12),
	.w5(32'hbbca854e),
	.w6(32'h3a407779),
	.w7(32'h3aa45483),
	.w8(32'h3c41fa40),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc6561),
	.w1(32'h3b8abec7),
	.w2(32'h3b655bf3),
	.w3(32'hbc188e31),
	.w4(32'hbb1eb0f6),
	.w5(32'hbc2d4252),
	.w6(32'hbc3bcedb),
	.w7(32'h3b745ce5),
	.w8(32'hbbf9fc0c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83a6af),
	.w1(32'h3bc5dd95),
	.w2(32'hbc2c59d2),
	.w3(32'h3b2fecbc),
	.w4(32'hbbc55ef5),
	.w5(32'hbc223cc4),
	.w6(32'h3be1b08f),
	.w7(32'hbc02243e),
	.w8(32'h3be4cc77),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a828e),
	.w1(32'h3baeecdc),
	.w2(32'hba784a87),
	.w3(32'hbc9298bc),
	.w4(32'hbc20ff2f),
	.w5(32'hbc3676c0),
	.w6(32'hbc1ad179),
	.w7(32'hbbec61f4),
	.w8(32'hbd9d99e3),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06902c),
	.w1(32'h3bc05681),
	.w2(32'hbcbfb6e6),
	.w3(32'h3b54731d),
	.w4(32'h3c75498f),
	.w5(32'hbc36a157),
	.w6(32'hbc2c8eb0),
	.w7(32'hbc2c180a),
	.w8(32'hba4da03a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24bbcf),
	.w1(32'h3ad489a6),
	.w2(32'hbc0a3585),
	.w3(32'hbbad4494),
	.w4(32'hbcab33e2),
	.w5(32'h3c2ed3e2),
	.w6(32'hbc148523),
	.w7(32'h3a608c12),
	.w8(32'hbbac39af),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab74a48),
	.w1(32'h3b35c8f9),
	.w2(32'hbb71be9c),
	.w3(32'h3bff1cf3),
	.w4(32'hbc6345cd),
	.w5(32'h398e6e40),
	.w6(32'h3a9d5df8),
	.w7(32'h3a66ef80),
	.w8(32'h3bffae29),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9c627),
	.w1(32'h3b38311e),
	.w2(32'hbbbffdda),
	.w3(32'h3c0bb12a),
	.w4(32'hba8dd021),
	.w5(32'h39c557ce),
	.w6(32'hbc1b271d),
	.w7(32'h3c822222),
	.w8(32'h3c075677),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d2356),
	.w1(32'h396a573b),
	.w2(32'h3c23b5bb),
	.w3(32'h3c620072),
	.w4(32'h3b18e99a),
	.w5(32'hbc9f24f1),
	.w6(32'hba8db656),
	.w7(32'hbbfb31db),
	.w8(32'h3c9c775e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af529a4),
	.w1(32'hbc07aa4a),
	.w2(32'h3b8117e8),
	.w3(32'hbc0a38f7),
	.w4(32'h3ba2791c),
	.w5(32'hbd57f23a),
	.w6(32'hbc93c223),
	.w7(32'hbadf5267),
	.w8(32'h3b9e5f25),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7157a3),
	.w1(32'hbb5d167b),
	.w2(32'h3afeafcc),
	.w3(32'hbc08da61),
	.w4(32'hbbc5b427),
	.w5(32'h3b8be2c0),
	.w6(32'hbc9cae44),
	.w7(32'h3ae3dda8),
	.w8(32'hbc89913d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc301f6d),
	.w1(32'hbba55413),
	.w2(32'hba113a50),
	.w3(32'h3b84c1e6),
	.w4(32'hbb8cbb43),
	.w5(32'hb9b127db),
	.w6(32'hbb6c3c6a),
	.w7(32'hbb0b5e2c),
	.w8(32'h3b3c5cdf),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8314e),
	.w1(32'h3ac7ced9),
	.w2(32'h3b2f0570),
	.w3(32'hb99f5d7e),
	.w4(32'hbc11d495),
	.w5(32'h3b767482),
	.w6(32'h3b273800),
	.w7(32'hbbd656b8),
	.w8(32'hbc36e0b7),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ea3d5),
	.w1(32'h3c19859c),
	.w2(32'hbc3681d3),
	.w3(32'hbb784f68),
	.w4(32'h39555f14),
	.w5(32'hbc62c873),
	.w6(32'h3c070c22),
	.w7(32'h3bb0b5ba),
	.w8(32'h3b68955c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86df20),
	.w1(32'hbbb7808e),
	.w2(32'hba1bfd9e),
	.w3(32'h3c0c5cd3),
	.w4(32'hbba04812),
	.w5(32'h3c1b38dc),
	.w6(32'hbbf9f4bc),
	.w7(32'h3b6056b5),
	.w8(32'h3b2a3dda),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b928a03),
	.w1(32'h3b0dac4a),
	.w2(32'hba6242ec),
	.w3(32'hba1c905e),
	.w4(32'h3b0f3018),
	.w5(32'h3ba79855),
	.w6(32'h3bd8026e),
	.w7(32'h3af31769),
	.w8(32'hbb5ea816),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b857b34),
	.w1(32'h39a407fa),
	.w2(32'h3bb00d74),
	.w3(32'hbad59af6),
	.w4(32'hbbe3a8c1),
	.w5(32'h3c202df8),
	.w6(32'h3c041967),
	.w7(32'h3b4df94c),
	.w8(32'h3c3bdc9d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a19a03),
	.w1(32'h39d8bfef),
	.w2(32'hbba57a06),
	.w3(32'hbb9b20eb),
	.w4(32'hbbeb740f),
	.w5(32'hbbe5eafb),
	.w6(32'hbbb513f4),
	.w7(32'h3c0e4cd4),
	.w8(32'hbc1b63ef),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc373962),
	.w1(32'hbaee94fa),
	.w2(32'h3c1b0a23),
	.w3(32'h3b6a2325),
	.w4(32'hba5dd19c),
	.w5(32'hbbaf5522),
	.w6(32'h3a011b19),
	.w7(32'h3b5ec50d),
	.w8(32'hbabcae49),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95eaee),
	.w1(32'hbce96b06),
	.w2(32'hbba8802f),
	.w3(32'hbcaa7488),
	.w4(32'h3a249980),
	.w5(32'h3b76ce08),
	.w6(32'hbc5837c9),
	.w7(32'hbb3fc9c9),
	.w8(32'h3988db3c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc5444),
	.w1(32'h3b819ec4),
	.w2(32'hbc0d3793),
	.w3(32'h3a22b40e),
	.w4(32'hbac67fe8),
	.w5(32'hbb82778a),
	.w6(32'h3c32d6d4),
	.w7(32'h3bbeab15),
	.w8(32'hbb6350d4),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35d039),
	.w1(32'h3c9a454b),
	.w2(32'hbb3ca48a),
	.w3(32'hbb8834b3),
	.w4(32'hbc18d86e),
	.w5(32'hbb9e2d05),
	.w6(32'hbaada794),
	.w7(32'h3b14efee),
	.w8(32'h3c8002c4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba069329),
	.w1(32'h3ba5bfc0),
	.w2(32'hb994bae8),
	.w3(32'hbaac9125),
	.w4(32'hbbbc4256),
	.w5(32'h3acb74e8),
	.w6(32'h3bc95e3f),
	.w7(32'h3be9a45d),
	.w8(32'hb9c49971),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ec8c47),
	.w1(32'h382956d7),
	.w2(32'hbba62c54),
	.w3(32'h3bf00575),
	.w4(32'hbcd41695),
	.w5(32'h3bf2c1a4),
	.w6(32'hbce89955),
	.w7(32'hbc8e261a),
	.w8(32'h3a4fd2cd),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10885a),
	.w1(32'h3ab5056a),
	.w2(32'hbb141c33),
	.w3(32'hbb9d9fec),
	.w4(32'hbb319359),
	.w5(32'hbbfc32a1),
	.w6(32'hbcae523a),
	.w7(32'h3afbbfb7),
	.w8(32'hbb28c9c7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65d40a),
	.w1(32'hbbe46d32),
	.w2(32'hbc46b7a0),
	.w3(32'hbb2abcc7),
	.w4(32'hba80b366),
	.w5(32'hbb864c33),
	.w6(32'h3b848db7),
	.w7(32'hbb867b41),
	.w8(32'h3c594869),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91a655),
	.w1(32'hbb15500c),
	.w2(32'h3ba44322),
	.w3(32'hbc96e257),
	.w4(32'h3b8420a3),
	.w5(32'hbc4fe3ab),
	.w6(32'h3b86a271),
	.w7(32'h3cb764c4),
	.w8(32'h399ce6c0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ddcd),
	.w1(32'h3b7e95e5),
	.w2(32'hbb172939),
	.w3(32'hbad6a22c),
	.w4(32'h3a84a6e8),
	.w5(32'h3b8fe4c1),
	.w6(32'hbb5f1220),
	.w7(32'h3c1d29a0),
	.w8(32'hbc22f132),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35965e),
	.w1(32'h3b2186b8),
	.w2(32'h3bc83a13),
	.w3(32'hbb100e9b),
	.w4(32'hbb828031),
	.w5(32'hbc27b21a),
	.w6(32'hbb55f1a4),
	.w7(32'hb9f712e7),
	.w8(32'h3b7c63a0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule