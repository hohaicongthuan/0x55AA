module layer_10_featuremap_98(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31976e),
	.w1(32'hbc11535f),
	.w2(32'h3c7d1879),
	.w3(32'hb9a3dd0f),
	.w4(32'hbc304619),
	.w5(32'h3a34c730),
	.w6(32'hb8c164a6),
	.w7(32'h3b8af8da),
	.w8(32'hbc90a69e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74b0bb),
	.w1(32'hbd2d2ad9),
	.w2(32'h3b8e58d8),
	.w3(32'hbac1c77f),
	.w4(32'hbc3a03c4),
	.w5(32'hbaaebbd6),
	.w6(32'hbc826d40),
	.w7(32'h3c1d9b73),
	.w8(32'h3c7bbf67),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d23d306),
	.w1(32'hbcdd2c5e),
	.w2(32'hba677bcc),
	.w3(32'h3c291cfa),
	.w4(32'hbbd03a9c),
	.w5(32'hba9e89c8),
	.w6(32'hbc7538f5),
	.w7(32'h3bc1e450),
	.w8(32'h3c57c09a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1d763),
	.w1(32'h3b3678f2),
	.w2(32'h3bc584f2),
	.w3(32'h3b3e91a3),
	.w4(32'h3b43bd76),
	.w5(32'h3baa1cc1),
	.w6(32'h39382c8c),
	.w7(32'h3be01254),
	.w8(32'h3bff5935),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1c735),
	.w1(32'h3c4d67ac),
	.w2(32'hbc927c7b),
	.w3(32'h3becd31a),
	.w4(32'h3bd75242),
	.w5(32'hba82195f),
	.w6(32'hbb3e4bb9),
	.w7(32'hbc0f4496),
	.w8(32'hbabbc393),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ba166),
	.w1(32'h3b323eee),
	.w2(32'h3a85e236),
	.w3(32'hbb8de576),
	.w4(32'hbbc1ee07),
	.w5(32'h3bc37dd7),
	.w6(32'h3ab0db57),
	.w7(32'h3b02cb1c),
	.w8(32'h3c0d5eba),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cee24),
	.w1(32'hbd253286),
	.w2(32'hbbc2d1d0),
	.w3(32'h3c66b693),
	.w4(32'hbc5382c9),
	.w5(32'hbc34c188),
	.w6(32'hbca0e1d1),
	.w7(32'h3bcc14a4),
	.w8(32'h3c567f58),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a91f1),
	.w1(32'h3c69a2e2),
	.w2(32'hb9a9eb65),
	.w3(32'h3b058f0e),
	.w4(32'hbc056ff0),
	.w5(32'hba24deb8),
	.w6(32'h3b5a6389),
	.w7(32'hbc31f899),
	.w8(32'hbbb6e5df),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca03277),
	.w1(32'hbb2599a1),
	.w2(32'hbc25d524),
	.w3(32'hbacb28a4),
	.w4(32'hbc1177e7),
	.w5(32'hbbd31cac),
	.w6(32'hbc1e6ce4),
	.w7(32'hbc413464),
	.w8(32'h3b1813b1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93025),
	.w1(32'hbd204fbd),
	.w2(32'hbc01436d),
	.w3(32'h3bc84a8e),
	.w4(32'h3bf4f27d),
	.w5(32'hbbdb03a3),
	.w6(32'hbc4f3ebb),
	.w7(32'h3c16d5da),
	.w8(32'h3cb62b47),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6f28c8),
	.w1(32'h340865d7),
	.w2(32'h3bb9cd23),
	.w3(32'h3c64b45d),
	.w4(32'hbc762041),
	.w5(32'hba8cc123),
	.w6(32'h3b0fe93c),
	.w7(32'h3c33770a),
	.w8(32'h3af7f876),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64b87d),
	.w1(32'h3b02c8b4),
	.w2(32'hbbcb8202),
	.w3(32'h3a8bf4c7),
	.w4(32'hbb52502d),
	.w5(32'hbad877d4),
	.w6(32'h3a304d0f),
	.w7(32'hbb4caf07),
	.w8(32'hbbd75786),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdc5d3),
	.w1(32'hbb858935),
	.w2(32'hbb8ef0d0),
	.w3(32'h3aa2b610),
	.w4(32'hbc1d7963),
	.w5(32'hbbb39bb7),
	.w6(32'hbb622502),
	.w7(32'hbbacc6b7),
	.w8(32'hbaa50ca1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc54a60),
	.w1(32'h3d219e46),
	.w2(32'h3c1990a7),
	.w3(32'hbb27c9d3),
	.w4(32'hba9922e8),
	.w5(32'h3bb201af),
	.w6(32'h3cab7875),
	.w7(32'hbb6760a8),
	.w8(32'h3a749f7b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcde6c48),
	.w1(32'h39f9b91e),
	.w2(32'hbc410a2a),
	.w3(32'hba4494cb),
	.w4(32'h3a4a1650),
	.w5(32'h3bb7fb92),
	.w6(32'hbb3b53c8),
	.w7(32'hbb5695dd),
	.w8(32'hbbab55c9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbe56e),
	.w1(32'hbbedb81d),
	.w2(32'hbbebc475),
	.w3(32'hbbdc5f41),
	.w4(32'hbc3e5451),
	.w5(32'hbb76ab89),
	.w6(32'hbc095daf),
	.w7(32'hbc0a2adf),
	.w8(32'h3b63b62d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb131daf),
	.w1(32'h3b15e38a),
	.w2(32'h3bb6cc25),
	.w3(32'h3bbf42e5),
	.w4(32'h3b73d992),
	.w5(32'h3bd111c6),
	.w6(32'h3bc97634),
	.w7(32'h3b912a60),
	.w8(32'h3b1c82f7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91107b),
	.w1(32'hbd494d78),
	.w2(32'hba5f771d),
	.w3(32'hbaa02e4d),
	.w4(32'hbbd7c4bf),
	.w5(32'hbbb48cc3),
	.w6(32'hbccf659d),
	.w7(32'h3c41a2d0),
	.w8(32'h3cb7f2d5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d779692),
	.w1(32'hbcb48eb7),
	.w2(32'hbb193a62),
	.w3(32'h3c6b0754),
	.w4(32'hbba1e87a),
	.w5(32'hbbc384d0),
	.w6(32'hbbf4290a),
	.w7(32'h3b26e90e),
	.w8(32'h3b6f967c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48e0b0),
	.w1(32'hbb8a8d45),
	.w2(32'hbc1ef1f9),
	.w3(32'hbb3f7b4c),
	.w4(32'hbbdba758),
	.w5(32'hbbc8bdb9),
	.w6(32'hbbdf141a),
	.w7(32'hbc10a063),
	.w8(32'h3b7ec240),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc8e95),
	.w1(32'h39c2e1fa),
	.w2(32'hbc03713b),
	.w3(32'h3b59c383),
	.w4(32'hbc0d1240),
	.w5(32'hbc13b4fa),
	.w6(32'hbc14380e),
	.w7(32'hbc845af8),
	.w8(32'hbba79ca0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd114d2),
	.w1(32'h3b3c861d),
	.w2(32'h3b806dd3),
	.w3(32'h3a3de34f),
	.w4(32'hbc47302d),
	.w5(32'h3ab735de),
	.w6(32'h39b9ae74),
	.w7(32'h3b9b62d3),
	.w8(32'h3c229e51),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1954ee),
	.w1(32'hbc581e86),
	.w2(32'hbc153810),
	.w3(32'hbb7e5302),
	.w4(32'hba7e729b),
	.w5(32'h3a423d8e),
	.w6(32'hbc45dd60),
	.w7(32'hbad427bd),
	.w8(32'h3a490f20),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0cf1e),
	.w1(32'h3c222219),
	.w2(32'h3adf7f41),
	.w3(32'h3b0628ad),
	.w4(32'hbc483631),
	.w5(32'hbb0a8ceb),
	.w6(32'h3b2a6fef),
	.w7(32'hbbff804d),
	.w8(32'hbb0e704b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e7d6c),
	.w1(32'hbc2e2210),
	.w2(32'h3b568dba),
	.w3(32'hba952eb8),
	.w4(32'hbaedadac),
	.w5(32'hbb87c402),
	.w6(32'h3b01c6e6),
	.w7(32'h3bd19f8a),
	.w8(32'h3bacb4a4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3efbb),
	.w1(32'hbb4f6b85),
	.w2(32'h3a98effd),
	.w3(32'hbb2ab2f0),
	.w4(32'h3b9cb6a8),
	.w5(32'h3ba1d6c5),
	.w6(32'hbac06a74),
	.w7(32'h3a4cb1ea),
	.w8(32'hb964cd32),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86a70a),
	.w1(32'hbc430abf),
	.w2(32'hbbd3a250),
	.w3(32'h3b449aa9),
	.w4(32'hbc768bf9),
	.w5(32'hbbd89b1f),
	.w6(32'hbc458752),
	.w7(32'hbc05f4f7),
	.w8(32'h3981dd8f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb314e77),
	.w1(32'hbc491b32),
	.w2(32'h3baeda24),
	.w3(32'h3ab43801),
	.w4(32'hbb55a52f),
	.w5(32'h381a229e),
	.w6(32'h3b41f59d),
	.w7(32'h3ba20317),
	.w8(32'h3b6d66a0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad54a43),
	.w1(32'hbcd7f5c4),
	.w2(32'hbc831d32),
	.w3(32'hbb4e47ed),
	.w4(32'hbcbe1e03),
	.w5(32'hbc054096),
	.w6(32'hbc884314),
	.w7(32'hbc0ec0c0),
	.w8(32'h3b7ccade),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b093d),
	.w1(32'h3af6c85f),
	.w2(32'hbaf339c1),
	.w3(32'h3b46faa7),
	.w4(32'h3b22f4a9),
	.w5(32'h3aa0ea79),
	.w6(32'h3b66de5d),
	.w7(32'hbbc94e67),
	.w8(32'hbbb20142),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb545cba),
	.w1(32'hbbd5a9a6),
	.w2(32'hbba6a465),
	.w3(32'h3b46ffd4),
	.w4(32'hbc264422),
	.w5(32'hbb951d1f),
	.w6(32'hbc15a1f7),
	.w7(32'hbc0b3ef6),
	.w8(32'hbb2308d3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7556),
	.w1(32'hbc1ff702),
	.w2(32'hbbc80d7a),
	.w3(32'h3a4959de),
	.w4(32'hbc751bce),
	.w5(32'hbc17c9da),
	.w6(32'hbc0ca046),
	.w7(32'hbbe98740),
	.w8(32'hbb65a135),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6cc0d),
	.w1(32'hbae53856),
	.w2(32'hbcd839f9),
	.w3(32'hbafc291c),
	.w4(32'hbb1be2f6),
	.w5(32'hbc9131af),
	.w6(32'hb89068a2),
	.w7(32'hbc81efee),
	.w8(32'hbbad82e6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a954b),
	.w1(32'hbcb57e5a),
	.w2(32'hbce6bb15),
	.w3(32'hbc295495),
	.w4(32'hbba72dd7),
	.w5(32'hbc8353b9),
	.w6(32'hbc36ea36),
	.w7(32'hbc5cb988),
	.w8(32'hbc5a5f11),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb7f47),
	.w1(32'hbd49bda6),
	.w2(32'hbbd34c53),
	.w3(32'hbc1dccf6),
	.w4(32'hbc184459),
	.w5(32'hbc374a38),
	.w6(32'hbcd3835a),
	.w7(32'h3b801b8e),
	.w8(32'h3c926963),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d53c41e),
	.w1(32'hbc236630),
	.w2(32'hbb8af008),
	.w3(32'h3c33d52d),
	.w4(32'hbc4257f0),
	.w5(32'hbb480e6f),
	.w6(32'hbc028dad),
	.w7(32'hbbc9d145),
	.w8(32'hbb43278f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917345),
	.w1(32'hbd1f3c61),
	.w2(32'hbc1df39d),
	.w3(32'h3c021d7b),
	.w4(32'h3b4b0bd9),
	.w5(32'hbb44112f),
	.w6(32'hbc3d2f12),
	.w7(32'h3bcdc6dc),
	.w8(32'h3c726bfe),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e8bbb),
	.w1(32'hbd1cbe55),
	.w2(32'h3b828ef3),
	.w3(32'h3c2b644b),
	.w4(32'hbc1167ce),
	.w5(32'hba2d71fa),
	.w6(32'hbc765288),
	.w7(32'h3c26b8b2),
	.w8(32'h3c671a1a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d279e38),
	.w1(32'h3bd6ff3f),
	.w2(32'h3b3bebdd),
	.w3(32'h3c5c93bf),
	.w4(32'hbc6094a4),
	.w5(32'hbb919272),
	.w6(32'h3adf3e48),
	.w7(32'hbbd5329b),
	.w8(32'hbb0d28d9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26a081),
	.w1(32'hbceb70da),
	.w2(32'hbbafb0f4),
	.w3(32'h39ee0801),
	.w4(32'hbb7be6d6),
	.w5(32'hbbd70163),
	.w6(32'hbc43d515),
	.w7(32'h3b6313aa),
	.w8(32'h3bebfcc5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccdc2f1),
	.w1(32'hbb144361),
	.w2(32'hbb726510),
	.w3(32'h3b844ce6),
	.w4(32'h3aa8e3dd),
	.w5(32'h3a92aa09),
	.w6(32'hbb47bafb),
	.w7(32'hbbe9d849),
	.w8(32'hbc49b739),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e1432),
	.w1(32'hbcb9120c),
	.w2(32'hbb482911),
	.w3(32'hba94b3d8),
	.w4(32'hbb218cc2),
	.w5(32'hbb26413e),
	.w6(32'hbbfe8853),
	.w7(32'h3bee6997),
	.w8(32'h3c31bcad),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd4f80f),
	.w1(32'hbc09864e),
	.w2(32'hbc1adb68),
	.w3(32'h3c3952f6),
	.w4(32'hbc516f6f),
	.w5(32'hbc28613b),
	.w6(32'hbbf1a3f3),
	.w7(32'hbc04b980),
	.w8(32'hbb80a8f1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd1bec),
	.w1(32'hbcb1573a),
	.w2(32'h3956f946),
	.w3(32'hbb2746a2),
	.w4(32'h3cabb027),
	.w5(32'hbaf46ab0),
	.w6(32'h3b4c24a0),
	.w7(32'h3c63dee1),
	.w8(32'h3cc28a60),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d81a494),
	.w1(32'hbc90654b),
	.w2(32'hbbcb7e52),
	.w3(32'h3c8a0356),
	.w4(32'hbb0fb4a2),
	.w5(32'hbae5ce12),
	.w6(32'hbc3fc2de),
	.w7(32'h3b6d43a9),
	.w8(32'h3b96b869),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93e581),
	.w1(32'hbcb74bc2),
	.w2(32'hba86d803),
	.w3(32'h3adf051a),
	.w4(32'hbc355681),
	.w5(32'hbc29fb15),
	.w6(32'hbc57378e),
	.w7(32'h3ad9847e),
	.w8(32'h3c3e34ad),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c6d93),
	.w1(32'h3bba84a6),
	.w2(32'hbbe454d8),
	.w3(32'h3b3ae703),
	.w4(32'h3bacf5e9),
	.w5(32'h3b8601d4),
	.w6(32'hb9bf65b0),
	.w7(32'hbbb780bf),
	.w8(32'h39b42e0c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c56ba8),
	.w1(32'hbbd90fec),
	.w2(32'hbc166f1a),
	.w3(32'hbaf15500),
	.w4(32'h3b2bdf79),
	.w5(32'h3ac2d64a),
	.w6(32'h3a98fcac),
	.w7(32'hbbddab73),
	.w8(32'hb9a3c303),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83d2d1),
	.w1(32'hbc3cd2cf),
	.w2(32'hbc27fab2),
	.w3(32'h3b9597e1),
	.w4(32'hbc5a5c91),
	.w5(32'hbc10df40),
	.w6(32'hbc0149d7),
	.w7(32'hbbedafe0),
	.w8(32'hba39ba2a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6c8b3),
	.w1(32'h3c97b7c1),
	.w2(32'h3bf02776),
	.w3(32'hbb289cce),
	.w4(32'hbba9ac1c),
	.w5(32'h3b0c339d),
	.w6(32'h3c10486f),
	.w7(32'hbb3b04f1),
	.w8(32'hba2a2ad0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc782543),
	.w1(32'hbcd7a9da),
	.w2(32'hb9ecccd8),
	.w3(32'hbad47774),
	.w4(32'hbbe33f85),
	.w5(32'hbb96054c),
	.w6(32'hbc336f76),
	.w7(32'h3b96d4f7),
	.w8(32'h3c1a48b4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97ec2f),
	.w1(32'h3b922a42),
	.w2(32'h3c44eeb7),
	.w3(32'hb9cea2cc),
	.w4(32'h3a379719),
	.w5(32'hbc0c010a),
	.w6(32'h3c8c903e),
	.w7(32'h3bd21e48),
	.w8(32'hbb9f4be3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0806b8),
	.w1(32'hbc68788f),
	.w2(32'h3b5d6e5f),
	.w3(32'hbba4eaaa),
	.w4(32'hbc4dd0f3),
	.w5(32'h3b44a824),
	.w6(32'hbbf1b55b),
	.w7(32'h3b1156e6),
	.w8(32'h3be4b492),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b807ba7),
	.w1(32'hbaede66d),
	.w2(32'hbc90f33b),
	.w3(32'h3bf59094),
	.w4(32'h3b942c8e),
	.w5(32'hbba3c7f2),
	.w6(32'hbb41d0db),
	.w7(32'hbbce13a8),
	.w8(32'hbac85997),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4153ca),
	.w1(32'hbc551f5c),
	.w2(32'hb8988649),
	.w3(32'hbb7b0658),
	.w4(32'h3a088f10),
	.w5(32'hbaab1b11),
	.w6(32'hbb309a36),
	.w7(32'h3b284a9b),
	.w8(32'h3b3bc50d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be30248),
	.w1(32'hbc309fe6),
	.w2(32'h3b928943),
	.w3(32'hbb047d06),
	.w4(32'hbb97c83a),
	.w5(32'h3b914afa),
	.w6(32'hbc46f3da),
	.w7(32'hbb9fda2c),
	.w8(32'hbc1ebef2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02f72f),
	.w1(32'hbc2aadea),
	.w2(32'h3adf0904),
	.w3(32'hbb3830c4),
	.w4(32'hba04db60),
	.w5(32'hbac02700),
	.w6(32'hb8e89fe8),
	.w7(32'h3b4bf0e0),
	.w8(32'h3bba7109),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c667aec),
	.w1(32'h3ac6e5a4),
	.w2(32'h3c21c071),
	.w3(32'h3c1249b4),
	.w4(32'hbb4e83a2),
	.w5(32'h3a25590e),
	.w6(32'h39a6d146),
	.w7(32'h3b1d02a4),
	.w8(32'hbc70c21f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54f360),
	.w1(32'hbd264472),
	.w2(32'h3c21d54e),
	.w3(32'hbbbfc88c),
	.w4(32'hbc66e57e),
	.w5(32'h3af3e06e),
	.w6(32'hbc935a14),
	.w7(32'h3c5374e3),
	.w8(32'h3c1a9ac7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d185aac),
	.w1(32'h3bc853fd),
	.w2(32'h39503486),
	.w3(32'h3c2d7710),
	.w4(32'hbc4b4752),
	.w5(32'hbb90a125),
	.w6(32'h39d035cb),
	.w7(32'hbbd22ddc),
	.w8(32'hb9d8edf2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5393de),
	.w1(32'hbd0b8e8c),
	.w2(32'hbbcb7243),
	.w3(32'hbb0b6b02),
	.w4(32'hbbad20de),
	.w5(32'hbb7d0b98),
	.w6(32'hbc7d637d),
	.w7(32'h3bffc7e3),
	.w8(32'h3c8c42d6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d13ec10),
	.w1(32'h3bd8848e),
	.w2(32'hbb3ace6d),
	.w3(32'h3a94571b),
	.w4(32'hbb6e4a35),
	.w5(32'h39a36b17),
	.w6(32'hb7c7e4dc),
	.w7(32'hbbd73b6c),
	.w8(32'hbaa343f7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc190474),
	.w1(32'h38c5a6b7),
	.w2(32'hbd1c7b29),
	.w3(32'hbacf13dd),
	.w4(32'h3beb837a),
	.w5(32'hbc1743c5),
	.w6(32'hbc0b6eab),
	.w7(32'hbc81030b),
	.w8(32'h3b8b00f9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e89df),
	.w1(32'hbca76fe4),
	.w2(32'hbb121ee0),
	.w3(32'h3b1b727d),
	.w4(32'h3c314816),
	.w5(32'hbb9d616a),
	.w6(32'hba59b1ce),
	.w7(32'h3c1d5469),
	.w8(32'h3c88744d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3c1c89),
	.w1(32'hbc91f116),
	.w2(32'hbc4b817b),
	.w3(32'h3c32000e),
	.w4(32'hbbb227f3),
	.w5(32'hbc03c376),
	.w6(32'hbc34a815),
	.w7(32'hbb192ed8),
	.w8(32'h3c1a3e36),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c835951),
	.w1(32'h3c40044b),
	.w2(32'hbb97794b),
	.w3(32'hba2965e1),
	.w4(32'h3a248b96),
	.w5(32'hbbde0b07),
	.w6(32'h3be9c6d6),
	.w7(32'hbba3ea7e),
	.w8(32'hbb5bdf6d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe942bb),
	.w1(32'hbba7a9ec),
	.w2(32'hbb92d0e9),
	.w3(32'hbb3b4628),
	.w4(32'h3bbfbb3d),
	.w5(32'h3bae7abf),
	.w6(32'hbb976e24),
	.w7(32'hbbb2f7f5),
	.w8(32'hbc251092),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf553b),
	.w1(32'hbc521be0),
	.w2(32'hbab92065),
	.w3(32'h3a95f235),
	.w4(32'hbbace909),
	.w5(32'h3b6058ad),
	.w6(32'hbc224cee),
	.w7(32'hbb42a2bd),
	.w8(32'hbc02059f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94ed80),
	.w1(32'hbbe30556),
	.w2(32'h3b72a744),
	.w3(32'h3b084817),
	.w4(32'hbc8206a7),
	.w5(32'hbb34ece1),
	.w6(32'hbbed368e),
	.w7(32'hbaa7656d),
	.w8(32'h3b51ee81),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6de701),
	.w1(32'h3c010104),
	.w2(32'h3b89aa89),
	.w3(32'h3bdb4177),
	.w4(32'h3c0141ba),
	.w5(32'hbbf3d097),
	.w6(32'h3beabe47),
	.w7(32'hbad1c6a2),
	.w8(32'h3981f312),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12df45),
	.w1(32'hbd222522),
	.w2(32'h3bf41158),
	.w3(32'hbb8af364),
	.w4(32'hbc2c62ee),
	.w5(32'h3a16699b),
	.w6(32'hbc87e421),
	.w7(32'h3c5bb7ce),
	.w8(32'h3c803fb6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3d91bd),
	.w1(32'h3aaa7d9a),
	.w2(32'h3bb511c2),
	.w3(32'h3c7598e2),
	.w4(32'hbc60022d),
	.w5(32'hbae5045e),
	.w6(32'hbb8c48e7),
	.w7(32'hbb25b99c),
	.w8(32'h3a31fcb8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedf3b0),
	.w1(32'h3b9b49c3),
	.w2(32'h3b1154e3),
	.w3(32'h3a8fd14f),
	.w4(32'hbc4539b5),
	.w5(32'hbb49f77d),
	.w6(32'hb988b691),
	.w7(32'hbba1ac63),
	.w8(32'hb9f460a4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1777c9),
	.w1(32'hbc5d87c0),
	.w2(32'hbbd2bed5),
	.w3(32'h3aa7c543),
	.w4(32'hbca0d49e),
	.w5(32'hbc0a5ef3),
	.w6(32'hbc0ee18c),
	.w7(32'hbbd1e333),
	.w8(32'hba84a2b1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfabc2),
	.w1(32'hbd00de53),
	.w2(32'h3bec79ec),
	.w3(32'h3a9bc3ba),
	.w4(32'hbbd07664),
	.w5(32'hb9d6c548),
	.w6(32'hbc31d2ba),
	.w7(32'h3c3bcd8b),
	.w8(32'h3c524baf),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cff86b7),
	.w1(32'hbba0b604),
	.w2(32'h3b1bc1de),
	.w3(32'h3ba2ee68),
	.w4(32'h3b0551cc),
	.w5(32'hba962ffe),
	.w6(32'h3b5a238f),
	.w7(32'hba567d36),
	.w8(32'hbba93f1d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3865d),
	.w1(32'h3d13fbf6),
	.w2(32'h3acec11f),
	.w3(32'h3c3a2e11),
	.w4(32'hbac2c08b),
	.w5(32'h3a3c2ed1),
	.w6(32'h3c4f2b38),
	.w7(32'hbc5505b5),
	.w8(32'hbbb9b79b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceb91b4),
	.w1(32'hbcbc6312),
	.w2(32'hbb75821e),
	.w3(32'hbb158e25),
	.w4(32'h3b8f58cd),
	.w5(32'h3b9cc084),
	.w6(32'hbbcc7c81),
	.w7(32'h3c356f36),
	.w8(32'h3c2e384f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf8a785),
	.w1(32'h3ba04830),
	.w2(32'h3b70827c),
	.w3(32'h3ba59e85),
	.w4(32'h3bf8c45d),
	.w5(32'h3b5f4696),
	.w6(32'h3b9425f8),
	.w7(32'hbb000ef9),
	.w8(32'hb9bfda54),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d4cfb),
	.w1(32'hbc057ab7),
	.w2(32'hbc4eeaa3),
	.w3(32'hbb2888ca),
	.w4(32'hbc89ff35),
	.w5(32'hbc3da873),
	.w6(32'hbc76e243),
	.w7(32'hbc95d71c),
	.w8(32'hbb865610),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed8382),
	.w1(32'hbc766603),
	.w2(32'hbb0275ad),
	.w3(32'h39ffe1f8),
	.w4(32'hbbec4235),
	.w5(32'h3b1a922c),
	.w6(32'hbc31439f),
	.w7(32'hbba3294c),
	.w8(32'hbbca7ecb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb797338),
	.w1(32'hbcc127dc),
	.w2(32'hbafb687e),
	.w3(32'h3b1f5cf6),
	.w4(32'hba5f26b0),
	.w5(32'h38c67d20),
	.w6(32'hbbcb9fd7),
	.w7(32'h3c05db18),
	.w8(32'h3c6d9a97),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d11cf82),
	.w1(32'hbbe23db6),
	.w2(32'h3b04fca4),
	.w3(32'h3c6943aa),
	.w4(32'hb9bec729),
	.w5(32'hbaa9e9b8),
	.w6(32'hbb3ebfda),
	.w7(32'h3aecfc14),
	.w8(32'h381f6288),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b397aab),
	.w1(32'hbccf9187),
	.w2(32'h3b7b6541),
	.w3(32'h39752bef),
	.w4(32'hbbaadd80),
	.w5(32'h3b0a9daa),
	.w6(32'hbc344db8),
	.w7(32'h3bf501e2),
	.w8(32'h3c316cb4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09c0c1),
	.w1(32'hbbdd5819),
	.w2(32'hbbc9adcd),
	.w3(32'h3c2a1b23),
	.w4(32'hbc3c99fb),
	.w5(32'hbb0d9323),
	.w6(32'h3bd6e0da),
	.w7(32'h3bbfe495),
	.w8(32'hba82af55),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf6a2b),
	.w1(32'hbc2aa21b),
	.w2(32'h3c09ac54),
	.w3(32'h39d6e055),
	.w4(32'h3b981970),
	.w5(32'h3be0afb4),
	.w6(32'hb99961c2),
	.w7(32'h3bcddf3f),
	.w8(32'h3afeeb48),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c33d2),
	.w1(32'hbb762cae),
	.w2(32'h3bf0d8f0),
	.w3(32'h3b80dc4e),
	.w4(32'h3b1d7a8d),
	.w5(32'hba0c8f7a),
	.w6(32'h3bf18009),
	.w7(32'h3b848cdc),
	.w8(32'hbb830de2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa34227),
	.w1(32'hbbaf3b16),
	.w2(32'hbb8d4cec),
	.w3(32'h3b7b2348),
	.w4(32'hbc23460d),
	.w5(32'hbba64407),
	.w6(32'hbc030d7d),
	.w7(32'hbbf68484),
	.w8(32'hbb227c12),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd4346),
	.w1(32'hbc70e26a),
	.w2(32'h3adf8dad),
	.w3(32'hb8fe8de1),
	.w4(32'hba79ed6e),
	.w5(32'hbaab88bb),
	.w6(32'hbb151416),
	.w7(32'h3b63c7e9),
	.w8(32'h3b576167),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23157f),
	.w1(32'hbc01aef5),
	.w2(32'hbc4029e8),
	.w3(32'hbb420ee7),
	.w4(32'hbc7bcbaa),
	.w5(32'hbc3d1d82),
	.w6(32'hbc860e10),
	.w7(32'hbc9ac022),
	.w8(32'hbbefeeb3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c5753),
	.w1(32'hbb9c3fe4),
	.w2(32'hbade6cea),
	.w3(32'hba383d01),
	.w4(32'hbc1a6bbf),
	.w5(32'hbb6504d1),
	.w6(32'hba9a0377),
	.w7(32'hbaf3fe0d),
	.w8(32'hba8c67ba),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0dc42),
	.w1(32'hbd04523b),
	.w2(32'hbbcb634b),
	.w3(32'h3aea90a6),
	.w4(32'h3a341323),
	.w5(32'hbb8bf4fc),
	.w6(32'hbc70861b),
	.w7(32'h3c054222),
	.w8(32'h3c871e9e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3b9167),
	.w1(32'hbc9dbd93),
	.w2(32'h3bd40eff),
	.w3(32'h3c3df1ae),
	.w4(32'hbb0996a9),
	.w5(32'h3b9d4604),
	.w6(32'hbbaa76d8),
	.w7(32'h3bfc44b5),
	.w8(32'h3c90818f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1e02ab),
	.w1(32'hbc8542ce),
	.w2(32'hbc13e7c2),
	.w3(32'h3c99e589),
	.w4(32'hbc14577d),
	.w5(32'hbb6fae59),
	.w6(32'hbc6315b1),
	.w7(32'hbc2e0a1d),
	.w8(32'hbbd50e3e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdb2b2),
	.w1(32'hbcd4e8d7),
	.w2(32'h3a74de67),
	.w3(32'h3b00709f),
	.w4(32'hbc03e424),
	.w5(32'hbb74a3de),
	.w6(32'hbc81e425),
	.w7(32'h3b2b40b4),
	.w8(32'h3bf69bc8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9ecb0),
	.w1(32'hb9fe722b),
	.w2(32'h3b617ed9),
	.w3(32'h3be60a87),
	.w4(32'hbc074618),
	.w5(32'hb9089ceb),
	.w6(32'h3b8422db),
	.w7(32'h3b6a48e3),
	.w8(32'h3b85d39a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb712bb),
	.w1(32'hbc03af5b),
	.w2(32'hb924936e),
	.w3(32'h3c25e3ff),
	.w4(32'h3b372b74),
	.w5(32'h3b971b68),
	.w6(32'hbc3ae643),
	.w7(32'hbb66e866),
	.w8(32'h39dd3839),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b1443),
	.w1(32'hbc8c49bf),
	.w2(32'hbc8238c6),
	.w3(32'hbb5490bc),
	.w4(32'hbc9d2338),
	.w5(32'hbc9a14f7),
	.w6(32'hbc088dcd),
	.w7(32'hbc2b6736),
	.w8(32'hbc23a8d4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d8dd),
	.w1(32'hbd18319d),
	.w2(32'hbc327005),
	.w3(32'hbb9e4caa),
	.w4(32'hbbcf0e3c),
	.w5(32'hbbcfee78),
	.w6(32'hbc82abf7),
	.w7(32'h3bdd78bf),
	.w8(32'h3c515a63),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07d13b),
	.w1(32'hbc477598),
	.w2(32'h3b1e2d04),
	.w3(32'h3bd12b65),
	.w4(32'h3b6100c8),
	.w5(32'h3bc31efb),
	.w6(32'hbb3157c2),
	.w7(32'h3b820386),
	.w8(32'h3bc3ac2e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51a4c6),
	.w1(32'h3b377c02),
	.w2(32'hbcad66f6),
	.w3(32'h3c16358b),
	.w4(32'h3c0f46e0),
	.w5(32'hbc8d41e7),
	.w6(32'h3b2d5f27),
	.w7(32'hbbc46c95),
	.w8(32'hbb63a498),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe6652),
	.w1(32'h3c71aac9),
	.w2(32'hbb6f95b8),
	.w3(32'hbc141df5),
	.w4(32'h3bc4e1a1),
	.w5(32'hbb9c47cf),
	.w6(32'h3c065a0d),
	.w7(32'h3b8dcb96),
	.w8(32'h3ba518d3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144ce7),
	.w1(32'h3d64bde3),
	.w2(32'h3b412e1c),
	.w3(32'hbb6f9270),
	.w4(32'h3b2205da),
	.w5(32'h3b17235b),
	.w6(32'h3cc34e77),
	.w7(32'hbc730c24),
	.w8(32'hbbf4c999),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2c30ee),
	.w1(32'hbb68e3b7),
	.w2(32'h3baea34b),
	.w3(32'hbb4ada0b),
	.w4(32'hbc85cad5),
	.w5(32'h3a666d5d),
	.w6(32'hbc196b1a),
	.w7(32'hbb10208e),
	.w8(32'h3ac0666a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef2337),
	.w1(32'h3cd18e98),
	.w2(32'hba43d513),
	.w3(32'h3afd2bca),
	.w4(32'hba788a2b),
	.w5(32'h3942dcd5),
	.w6(32'h3c2be202),
	.w7(32'hbc14a4fe),
	.w8(32'hbbbf9f4e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1e26e),
	.w1(32'hbbd5c0ca),
	.w2(32'hbc37e474),
	.w3(32'h39127610),
	.w4(32'hbc2447f4),
	.w5(32'hbc0bc67a),
	.w6(32'hbc006e87),
	.w7(32'hbc565551),
	.w8(32'hbb2e7e60),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdca0c4),
	.w1(32'hbcd31a5f),
	.w2(32'hbb3766eb),
	.w3(32'h39497a6c),
	.w4(32'hbbc9c942),
	.w5(32'hba47f86d),
	.w6(32'hbc8b35ac),
	.w7(32'h3a97c525),
	.w8(32'h3c1f3163),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05a484),
	.w1(32'hbb809899),
	.w2(32'hbb1e9727),
	.w3(32'h3c1164a7),
	.w4(32'hbc0c2be2),
	.w5(32'hbb3be5c3),
	.w6(32'hbb9b022d),
	.w7(32'hbbb36028),
	.w8(32'hbb123c6c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d3473),
	.w1(32'h3cf0656b),
	.w2(32'h3b14dcae),
	.w3(32'h3b49f6c8),
	.w4(32'h3a7c3665),
	.w5(32'h3ac5b71a),
	.w6(32'h3c4918ed),
	.w7(32'hbc0ef935),
	.w8(32'hbb586f1a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb507e2),
	.w1(32'hbcd1b698),
	.w2(32'h3b0ace64),
	.w3(32'hba8da3e8),
	.w4(32'h3af04405),
	.w5(32'h3b34bbe9),
	.w6(32'hbc13e0b1),
	.w7(32'h3bc4dc07),
	.w8(32'h3c131bcf),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfb2ebd),
	.w1(32'hbb0edeec),
	.w2(32'hbac77681),
	.w3(32'h3be1b5b7),
	.w4(32'hbc53071a),
	.w5(32'hbbe06ad3),
	.w6(32'hbaec392c),
	.w7(32'hbbb00857),
	.w8(32'h3a86077a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec2c30),
	.w1(32'h3c55ef2c),
	.w2(32'hbcb4cb2e),
	.w3(32'h3b55ef6f),
	.w4(32'h3c53169d),
	.w5(32'hbbc5921f),
	.w6(32'h3b19f5a3),
	.w7(32'hbbc9b4aa),
	.w8(32'hba541c7e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefa60f),
	.w1(32'hbb99cb6b),
	.w2(32'h3aa5b9e0),
	.w3(32'hbc0cbdf3),
	.w4(32'hbc78b450),
	.w5(32'hbb849b25),
	.w6(32'hbb7f0d31),
	.w7(32'hbb53dda9),
	.w8(32'h3b059dad),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5e341),
	.w1(32'hbd1024e4),
	.w2(32'h3b2b03f6),
	.w3(32'h3b7192e3),
	.w4(32'hbc5793e7),
	.w5(32'hbb1f732d),
	.w6(32'hbc4e3b93),
	.w7(32'h3bf67494),
	.w8(32'h3adf9ee9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab6f50),
	.w1(32'h3b54f59d),
	.w2(32'h3abb632a),
	.w3(32'hba674017),
	.w4(32'hbb936124),
	.w5(32'h3b8f2f7a),
	.w6(32'hba44d0d6),
	.w7(32'hbb6c634d),
	.w8(32'h3bfac4ae),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4864f6),
	.w1(32'h3d28145b),
	.w2(32'h3b32a108),
	.w3(32'h3ba5261b),
	.w4(32'h39b1a09a),
	.w5(32'h3aa26537),
	.w6(32'h3c89b427),
	.w7(32'hbc4359fd),
	.w8(32'hbb95faa1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd009366),
	.w1(32'h3c5663bf),
	.w2(32'h3ac8e2d5),
	.w3(32'hbb41e587),
	.w4(32'hbc02d071),
	.w5(32'hbab1572e),
	.w6(32'h3b77db11),
	.w7(32'hbbb13e10),
	.w8(32'hbb82508d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc669370),
	.w1(32'h3c86b8ac),
	.w2(32'h39a0d8b9),
	.w3(32'hba53a87c),
	.w4(32'hbbda896d),
	.w5(32'hba96e20d),
	.w6(32'h3ba96f29),
	.w7(32'hbbdf49db),
	.w8(32'hbaec3f36),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70d367),
	.w1(32'h3be8466b),
	.w2(32'hbb1965de),
	.w3(32'h3a9a72fb),
	.w4(32'h3a2c1bbd),
	.w5(32'hbb547787),
	.w6(32'h3b19d1ec),
	.w7(32'hb99c8c44),
	.w8(32'hba893b08),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc58dd3),
	.w1(32'hbcb4fdfa),
	.w2(32'hbb7293b0),
	.w3(32'hbbe919fa),
	.w4(32'hbb8c64dd),
	.w5(32'hbc607f7d),
	.w6(32'hba1b87f2),
	.w7(32'h3a2a5c50),
	.w8(32'hbb58906f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fa6c2),
	.w1(32'hbc42a2b3),
	.w2(32'h39ef4de2),
	.w3(32'hbc9cc32c),
	.w4(32'hbc65229f),
	.w5(32'h39a8c1f4),
	.w6(32'hbc11ea54),
	.w7(32'h3bbd9e28),
	.w8(32'h3c0d33d9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b9ec2),
	.w1(32'hbbafecb5),
	.w2(32'hba1ac56f),
	.w3(32'h3be55242),
	.w4(32'hbbae3917),
	.w5(32'hba934a7a),
	.w6(32'hbb461cbd),
	.w7(32'hba613a64),
	.w8(32'h3bd1599a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9754),
	.w1(32'h3bffc63c),
	.w2(32'h3a91f813),
	.w3(32'h3bd788de),
	.w4(32'hbc5baa83),
	.w5(32'hbb5fc51c),
	.w6(32'h3b33f93c),
	.w7(32'hbbe9a23f),
	.w8(32'hbafccb7f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78725f),
	.w1(32'hbaa4877c),
	.w2(32'hbbd6a37d),
	.w3(32'hbac187a0),
	.w4(32'h3bc7df61),
	.w5(32'hba245f11),
	.w6(32'hbc3afadd),
	.w7(32'h38c220bc),
	.w8(32'h3b57375f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c4f8e),
	.w1(32'hbc6fbadc),
	.w2(32'h3b85f59e),
	.w3(32'hbbb63a49),
	.w4(32'hbc4ed938),
	.w5(32'h3c33d86e),
	.w6(32'hbba6bf2c),
	.w7(32'h3bf55ec9),
	.w8(32'h3c83b906),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8322f9),
	.w1(32'hbc2bbb61),
	.w2(32'hbbe0cdb5),
	.w3(32'h3c91fe78),
	.w4(32'hbc84aabd),
	.w5(32'hbbc9bf37),
	.w6(32'hbc541bc3),
	.w7(32'hbc16a777),
	.w8(32'hba54d7aa),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaed64b),
	.w1(32'hb88279dc),
	.w2(32'hb9b7402d),
	.w3(32'h3ad79d08),
	.w4(32'h39536fdf),
	.w5(32'hb9b0d386),
	.w6(32'h391af744),
	.w7(32'h37bdac10),
	.w8(32'hb9cd86d7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51699a),
	.w1(32'hba096e90),
	.w2(32'hbaf7bc70),
	.w3(32'h3a5fa785),
	.w4(32'hba986111),
	.w5(32'hbae0633e),
	.w6(32'hbabafb25),
	.w7(32'hbafb1023),
	.w8(32'hba9dcb2f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8e5b4),
	.w1(32'h3a54a412),
	.w2(32'hb8837f5b),
	.w3(32'h3a196348),
	.w4(32'hba8f82b4),
	.w5(32'hb9cf13a4),
	.w6(32'h3ab7e723),
	.w7(32'h39270e24),
	.w8(32'h3a4b31ce),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a916cb9),
	.w1(32'hba1f4f66),
	.w2(32'hba985eb6),
	.w3(32'h385a75b2),
	.w4(32'hba21ada2),
	.w5(32'hba6fa269),
	.w6(32'hb9f93095),
	.w7(32'hba609274),
	.w8(32'hba7e502e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84bb10),
	.w1(32'hba9f710c),
	.w2(32'hba9028ed),
	.w3(32'hba6701ce),
	.w4(32'hba18c90c),
	.w5(32'hba1cf9bc),
	.w6(32'hba877c21),
	.w7(32'hba6974db),
	.w8(32'hba3367f9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba419f79),
	.w1(32'hb9b5bf59),
	.w2(32'hb8edfefb),
	.w3(32'hb9b49f8b),
	.w4(32'h3891e295),
	.w5(32'h376dd68c),
	.w6(32'hba11be93),
	.w7(32'hba811272),
	.w8(32'hb9e782c1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba090483),
	.w1(32'hba02ee13),
	.w2(32'hba1866e6),
	.w3(32'h37630bcd),
	.w4(32'hb92ff80f),
	.w5(32'h399c59f7),
	.w6(32'hb97d5db0),
	.w7(32'hb875ef4c),
	.w8(32'hb8d2d90b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b7f90),
	.w1(32'hbaa258a2),
	.w2(32'hba89a576),
	.w3(32'hb9ecfbec),
	.w4(32'hb9a26488),
	.w5(32'h3a578417),
	.w6(32'hb985f1e8),
	.w7(32'hb8dbbec2),
	.w8(32'h3a7032fb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b2ced),
	.w1(32'hb983e6b3),
	.w2(32'hbb232918),
	.w3(32'h3a3fb4c1),
	.w4(32'hb9986ce0),
	.w5(32'hba76265b),
	.w6(32'hbaa96f55),
	.w7(32'hbb0f243f),
	.w8(32'hbabd3d76),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba796e4c),
	.w1(32'hb96a507f),
	.w2(32'h39f34479),
	.w3(32'h3797dab5),
	.w4(32'h3a6b9114),
	.w5(32'h3a77d5f6),
	.w6(32'h3a8308b3),
	.w7(32'h3a034830),
	.w8(32'h3a60bd1f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c2375),
	.w1(32'hba3ce148),
	.w2(32'hbacc2bcd),
	.w3(32'h3a8312e9),
	.w4(32'hb9316cb6),
	.w5(32'hba7a6125),
	.w6(32'hb9c75b43),
	.w7(32'hb897018e),
	.w8(32'hba50a847),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e4c00),
	.w1(32'h39938562),
	.w2(32'hbaa6e5a0),
	.w3(32'h3a3660ec),
	.w4(32'h395f2bf8),
	.w5(32'hb9120c16),
	.w6(32'hba6224c0),
	.w7(32'hba7c419b),
	.w8(32'hba089c0a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e42af),
	.w1(32'hba94e737),
	.w2(32'hb921290f),
	.w3(32'hb96ea2a7),
	.w4(32'h38e6a7ca),
	.w5(32'h37cd9872),
	.w6(32'hba6d7c70),
	.w7(32'hba2fdf18),
	.w8(32'h39deafdd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee3d01),
	.w1(32'hb7ed8e7d),
	.w2(32'hb80df2df),
	.w3(32'h3a89a8c6),
	.w4(32'h3a3bc901),
	.w5(32'hb672f83d),
	.w6(32'h39e2aed6),
	.w7(32'h39243d20),
	.w8(32'hb93b82c7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39156307),
	.w1(32'hb98dbb11),
	.w2(32'hb8b685ea),
	.w3(32'h39555d50),
	.w4(32'h388fa926),
	.w5(32'h397c299d),
	.w6(32'hb8610e6a),
	.w7(32'hb958ca72),
	.w8(32'h38b3d89a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a057eed),
	.w1(32'hba9fb82c),
	.w2(32'h3a5afd5f),
	.w3(32'h3a8b2e00),
	.w4(32'h39879d6f),
	.w5(32'h3a6f6f18),
	.w6(32'h3b229877),
	.w7(32'hba3f4d31),
	.w8(32'h3a118ecd),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ded97),
	.w1(32'hba0e869e),
	.w2(32'h398a0533),
	.w3(32'h3a79fa2e),
	.w4(32'hba699453),
	.w5(32'hba64fe91),
	.w6(32'hba2a8c4a),
	.w7(32'hba5d1a64),
	.w8(32'hba4a7914),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de0477),
	.w1(32'hba20a430),
	.w2(32'hba32e3a7),
	.w3(32'hb9532dec),
	.w4(32'hb9a10194),
	.w5(32'hb99e462c),
	.w6(32'hb99f271c),
	.w7(32'hb9c11448),
	.w8(32'hb99fc44d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9baebaa),
	.w1(32'h382ffec4),
	.w2(32'h39b6f635),
	.w3(32'hb98eb643),
	.w4(32'h384b6662),
	.w5(32'h395dbeac),
	.w6(32'hb91cb98c),
	.w7(32'h390f5f42),
	.w8(32'h3882a6ac),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4518e),
	.w1(32'hba55f45c),
	.w2(32'hba548b85),
	.w3(32'h39536899),
	.w4(32'hba5aaa31),
	.w5(32'hba32fb14),
	.w6(32'hb9eb96c7),
	.w7(32'hba750a1c),
	.w8(32'hba8fe955),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad297b8),
	.w1(32'hba158138),
	.w2(32'h39061a2d),
	.w3(32'hba4d637b),
	.w4(32'h3a35301a),
	.w5(32'h3a689877),
	.w6(32'h38d2775e),
	.w7(32'h36ec071f),
	.w8(32'hb970eaae),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba879a2b),
	.w1(32'hba9a01d9),
	.w2(32'h39f38594),
	.w3(32'hb987e23a),
	.w4(32'hba11297e),
	.w5(32'h3a60d7e4),
	.w6(32'hba029d54),
	.w7(32'hba3b2539),
	.w8(32'h3a5d7282),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7c7ed),
	.w1(32'hb97c22a1),
	.w2(32'hb9850bb1),
	.w3(32'hb71144ff),
	.w4(32'hb981e26f),
	.w5(32'hb95b1176),
	.w6(32'hb97135c6),
	.w7(32'hb97ab391),
	.w8(32'hb9d46229),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f131c),
	.w1(32'hb9e0e106),
	.w2(32'h3a900df3),
	.w3(32'h3a12509d),
	.w4(32'h390148ee),
	.w5(32'h3a11b7d7),
	.w6(32'h3a22b579),
	.w7(32'hba4be0cb),
	.w8(32'h3a01b857),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2ff7c),
	.w1(32'hba9e3c06),
	.w2(32'hb9e0769c),
	.w3(32'h39211713),
	.w4(32'hba2af590),
	.w5(32'hb88a481e),
	.w6(32'hb92fcba6),
	.w7(32'hba0d9379),
	.w8(32'h381b1c98),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02e0fa),
	.w1(32'hb8ba00d0),
	.w2(32'hbabcde51),
	.w3(32'h39cc93ea),
	.w4(32'h3a0359f3),
	.w5(32'hb95af421),
	.w6(32'h3897a065),
	.w7(32'hba3ab705),
	.w8(32'hba36255e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a532d69),
	.w1(32'hbaae5310),
	.w2(32'h3a369c36),
	.w3(32'h3ae552bd),
	.w4(32'hba0a8ce3),
	.w5(32'h3a261c2e),
	.w6(32'h3aaf18d8),
	.w7(32'hbb05acc8),
	.w8(32'hb98660fb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ec545),
	.w1(32'h3a34df3e),
	.w2(32'h39f87dc1),
	.w3(32'h3934bdad),
	.w4(32'h3a23f2b2),
	.w5(32'h39ba58ab),
	.w6(32'h3a702ddd),
	.w7(32'h3a0d59b7),
	.w8(32'hb7f5b8b5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaa444),
	.w1(32'h3a8488a0),
	.w2(32'h3a1e3499),
	.w3(32'h3ac18ae2),
	.w4(32'h3a39a4ae),
	.w5(32'h384b55e8),
	.w6(32'h3a34c1a8),
	.w7(32'h39bcb546),
	.w8(32'h39680555),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9758ae6),
	.w1(32'hba2c49f3),
	.w2(32'h389d34c7),
	.w3(32'h3a810ede),
	.w4(32'h3a10672b),
	.w5(32'h3a2d395b),
	.w6(32'h3a189bb4),
	.w7(32'h37ec7f07),
	.w8(32'hb8ae1d8d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d8d8),
	.w1(32'hbaa05c6d),
	.w2(32'hba885567),
	.w3(32'hb9aaff0b),
	.w4(32'hba056872),
	.w5(32'hb9e1ac7d),
	.w6(32'h37994463),
	.w7(32'hb98a0c15),
	.w8(32'hba65c2ca),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9f277),
	.w1(32'hb8890cf5),
	.w2(32'h39c7f972),
	.w3(32'hb9dba800),
	.w4(32'hb8f7e9f7),
	.w5(32'hb7f680d4),
	.w6(32'h37eef2eb),
	.w7(32'h392f6be5),
	.w8(32'h39211d31),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd20f1),
	.w1(32'h3904b3fb),
	.w2(32'hb9a34b32),
	.w3(32'h3819760a),
	.w4(32'h389d914f),
	.w5(32'hb8fc94c2),
	.w6(32'hb9dfa7fa),
	.w7(32'hba0248b0),
	.w8(32'hba0549b6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922133f),
	.w1(32'hb8773014),
	.w2(32'hb95a1726),
	.w3(32'hb8b20296),
	.w4(32'h38b79160),
	.w5(32'hb834ecea),
	.w6(32'hb907ce10),
	.w7(32'h36aadf30),
	.w8(32'hb92043c2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39088205),
	.w1(32'h398ca5d7),
	.w2(32'hba489b28),
	.w3(32'h3a02147a),
	.w4(32'h3a182f18),
	.w5(32'h390dda37),
	.w6(32'hb90844d5),
	.w7(32'hb99adca2),
	.w8(32'h3883a8f4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79f625),
	.w1(32'h3a11ac15),
	.w2(32'hb8c55e31),
	.w3(32'h3a4200cd),
	.w4(32'h3889d846),
	.w5(32'hb94c215a),
	.w6(32'h39d3916e),
	.w7(32'h39109657),
	.w8(32'hb953482c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dbbec),
	.w1(32'hba9037cf),
	.w2(32'hb99d9a79),
	.w3(32'h3a1a5397),
	.w4(32'hb9171410),
	.w5(32'h3882392d),
	.w6(32'h382341c3),
	.w7(32'hba26af5e),
	.w8(32'hb84e6c63),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cef2f),
	.w1(32'hb84e2783),
	.w2(32'hb9a7e3cb),
	.w3(32'hb9b7de50),
	.w4(32'h389b37dd),
	.w5(32'hb761d969),
	.w6(32'h38194776),
	.w7(32'h39208cf5),
	.w8(32'h38c78c83),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d4a5c),
	.w1(32'hba1034d5),
	.w2(32'hba83031c),
	.w3(32'hb9a6fa6a),
	.w4(32'hbaca88e7),
	.w5(32'hbaae78b8),
	.w6(32'hba9163cf),
	.w7(32'hbae31e54),
	.w8(32'hbac0abc5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba761918),
	.w1(32'hb9cb1021),
	.w2(32'hb9f1d5e2),
	.w3(32'hba120dec),
	.w4(32'hba063263),
	.w5(32'hba030819),
	.w6(32'hb9f800e2),
	.w7(32'hb9d7189e),
	.w8(32'hb9c2ea9b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcae89),
	.w1(32'h37df9b17),
	.w2(32'hb940e8b5),
	.w3(32'hba47b8b2),
	.w4(32'h38ffd510),
	.w5(32'hb891ebfc),
	.w6(32'h38e62f8c),
	.w7(32'h37a8d7c1),
	.w8(32'hb8c13b58),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8912429),
	.w1(32'hb9dd62f0),
	.w2(32'hb943c26e),
	.w3(32'h3a9fa235),
	.w4(32'h3a61fed5),
	.w5(32'h39441aa9),
	.w6(32'h3a59ae56),
	.w7(32'h39ccf38f),
	.w8(32'hba3eb48b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ed4a4),
	.w1(32'hb931b4ac),
	.w2(32'h3a1d0028),
	.w3(32'h3a821ed9),
	.w4(32'h3a0b18b6),
	.w5(32'h3a2371b8),
	.w6(32'hba9e0925),
	.w7(32'hb9f1cc1a),
	.w8(32'hba7315e9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39240e7a),
	.w1(32'hb962e986),
	.w2(32'hba6b2009),
	.w3(32'h38c54b71),
	.w4(32'h376de130),
	.w5(32'hba57239f),
	.w6(32'h36c63d58),
	.w7(32'hb92746cb),
	.w8(32'hb9ba52c7),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9585fb0),
	.w1(32'hb9c27124),
	.w2(32'h39146b73),
	.w3(32'h39d84ec5),
	.w4(32'h3a00ebcf),
	.w5(32'h3a3ab202),
	.w6(32'h3a95875b),
	.w7(32'h3a0dcba2),
	.w8(32'h39abc491),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e59a79),
	.w1(32'h3911dc7b),
	.w2(32'hb9ba0cfe),
	.w3(32'h39a734cd),
	.w4(32'hb979c41e),
	.w5(32'hb984138f),
	.w6(32'h3a60de78),
	.w7(32'hb87bda92),
	.w8(32'h39c31d24),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fd61c),
	.w1(32'hb97b5e97),
	.w2(32'hba9a820e),
	.w3(32'h3a58401a),
	.w4(32'h395b9927),
	.w5(32'h3a0f1d11),
	.w6(32'h39b2dbc1),
	.w7(32'hba8734f1),
	.w8(32'h398ec008),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9033056),
	.w1(32'hba81750c),
	.w2(32'hbacbdd17),
	.w3(32'h38fc0efc),
	.w4(32'hb9dd252f),
	.w5(32'hba210576),
	.w6(32'hba074b69),
	.w7(32'hba610383),
	.w8(32'hba2b055f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389665cc),
	.w1(32'h3a5aab79),
	.w2(32'h3a927736),
	.w3(32'h389eae1e),
	.w4(32'h39ad85e7),
	.w5(32'h3a3f3555),
	.w6(32'hb941b9d3),
	.w7(32'hba3cc8e5),
	.w8(32'h39b90453),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a984768),
	.w1(32'hba594a88),
	.w2(32'hba0de47f),
	.w3(32'h3a506cdb),
	.w4(32'hb9de977b),
	.w5(32'hb9efa0e5),
	.w6(32'hb9f8c412),
	.w7(32'hb9b6d365),
	.w8(32'hb9d84db0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20b336),
	.w1(32'hba933c17),
	.w2(32'hba5dfa3a),
	.w3(32'hb9ef279a),
	.w4(32'hb99232e8),
	.w5(32'h39bb7edf),
	.w6(32'h39488af3),
	.w7(32'h3832f4fc),
	.w8(32'hb91f81fa),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37994a68),
	.w1(32'h398f6b50),
	.w2(32'hb7b69279),
	.w3(32'h392d29b5),
	.w4(32'h39e081c4),
	.w5(32'h39b23372),
	.w6(32'h3a0d50ce),
	.w7(32'h39a3118b),
	.w8(32'h39d3d7c5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39929fa2),
	.w1(32'h391b4a3f),
	.w2(32'hb8501584),
	.w3(32'h39abe08c),
	.w4(32'hb8ac7050),
	.w5(32'hb52c9448),
	.w6(32'h3782c3f0),
	.w7(32'h38f66269),
	.w8(32'h398edd59),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7741004),
	.w1(32'h384746cd),
	.w2(32'hba43afa6),
	.w3(32'hb9c293fb),
	.w4(32'h3a458b64),
	.w5(32'hb8fe28fb),
	.w6(32'hb91a0a46),
	.w7(32'h38f0f1ff),
	.w8(32'h3a358e8c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5d372),
	.w1(32'hbafd9a2a),
	.w2(32'hbb1fae8d),
	.w3(32'hb8c2981b),
	.w4(32'hbaa1a389),
	.w5(32'hba66fbfd),
	.w6(32'hba7be4ea),
	.w7(32'hbaada771),
	.w8(32'hb9562143),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3e6f6),
	.w1(32'h39a084e5),
	.w2(32'h39548c2c),
	.w3(32'hb9837c84),
	.w4(32'hb8518768),
	.w5(32'h39574886),
	.w6(32'hb965212b),
	.w7(32'h39d5e6ac),
	.w8(32'h38b194a1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c733d9),
	.w1(32'h39050577),
	.w2(32'hb824158b),
	.w3(32'hb8b03a9a),
	.w4(32'hb89b152c),
	.w5(32'hb94f5287),
	.w6(32'h38af7d68),
	.w7(32'hb8bc1061),
	.w8(32'hb9e32ed7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9213bca),
	.w1(32'hba86cd70),
	.w2(32'h39416654),
	.w3(32'hb94d4635),
	.w4(32'hb99b3879),
	.w5(32'h398ffa90),
	.w6(32'hb9d35731),
	.w7(32'hba0f2ff2),
	.w8(32'h39e1c888),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e343a),
	.w1(32'hba4fc764),
	.w2(32'hbae113eb),
	.w3(32'h3adc1f50),
	.w4(32'h39f4da3b),
	.w5(32'hb96ca724),
	.w6(32'h3a870a2a),
	.w7(32'hb9b84b38),
	.w8(32'hba03b922),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7181e7),
	.w1(32'hb86a5ed2),
	.w2(32'h39fb8d4b),
	.w3(32'hb9022912),
	.w4(32'h39642132),
	.w5(32'h39c5fe06),
	.w6(32'hb9000016),
	.w7(32'h39b63c90),
	.w8(32'hb9a7a805),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941db53),
	.w1(32'hba017bfb),
	.w2(32'hba621b3f),
	.w3(32'hb99612e1),
	.w4(32'hb9c8fb03),
	.w5(32'hba4ddbf0),
	.w6(32'hba1cdfc7),
	.w7(32'hba30c22c),
	.w8(32'hb971109a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb27ba),
	.w1(32'hba39fc00),
	.w2(32'h3a15c610),
	.w3(32'h3a7af54f),
	.w4(32'hb9bee7a4),
	.w5(32'h3ae91629),
	.w6(32'hb9d5103c),
	.w7(32'hba884064),
	.w8(32'h3afbb177),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a821f6d),
	.w1(32'hba8bc311),
	.w2(32'hba59f1bf),
	.w3(32'h3b0360e2),
	.w4(32'h3a139ee7),
	.w5(32'h3a1458f3),
	.w6(32'h3b184fcd),
	.w7(32'hb8a38b7a),
	.w8(32'h37984c17),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3a570),
	.w1(32'h3a13e8c6),
	.w2(32'hb896581e),
	.w3(32'h399bd6a7),
	.w4(32'h39c486aa),
	.w5(32'h385a18b7),
	.w6(32'h3a6ce4c5),
	.w7(32'hb7cda861),
	.w8(32'hb9dbb498),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bcd61),
	.w1(32'h38c4ec51),
	.w2(32'hb9c34ab7),
	.w3(32'h398d6119),
	.w4(32'hb988a8cc),
	.w5(32'hba2aef44),
	.w6(32'h39cb6095),
	.w7(32'hba2a5d7c),
	.w8(32'hb9347b5f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dfad7f),
	.w1(32'hb6ff1cd8),
	.w2(32'hb94253b4),
	.w3(32'h3a13e0a6),
	.w4(32'hb8a721ef),
	.w5(32'hb9ae158e),
	.w6(32'h389c7dda),
	.w7(32'hb7a3945f),
	.w8(32'hb9053471),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4fd43),
	.w1(32'hb9bb5e6c),
	.w2(32'hba20c300),
	.w3(32'hb91d8909),
	.w4(32'hb9d3318f),
	.w5(32'hb9f84ee9),
	.w6(32'hb9a490dd),
	.w7(32'hb9fa9835),
	.w8(32'hb9c2205e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e4327),
	.w1(32'h3a4532f8),
	.w2(32'hba2692e0),
	.w3(32'h3a5cda1b),
	.w4(32'h3a2f9916),
	.w5(32'hba1f88f2),
	.w6(32'h396b31c5),
	.w7(32'hb96cdc85),
	.w8(32'hba42c923),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7cd13),
	.w1(32'h39d223fc),
	.w2(32'h37460380),
	.w3(32'h3a27f431),
	.w4(32'h3a6610e3),
	.w5(32'h39ec2354),
	.w6(32'h39c07705),
	.w7(32'h3a4d53d7),
	.w8(32'h39e96bed),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2909c7),
	.w1(32'hbace9a15),
	.w2(32'h3a2c6f26),
	.w3(32'h39c1810f),
	.w4(32'hb92dff3b),
	.w5(32'h3aade7e8),
	.w6(32'hb93b4e4e),
	.w7(32'h37d289e3),
	.w8(32'h3a7d40f6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76ace2),
	.w1(32'hba2be650),
	.w2(32'hba379d3e),
	.w3(32'hba223ae4),
	.w4(32'hb9747579),
	.w5(32'hb90ab2ec),
	.w6(32'hb97de569),
	.w7(32'hb98facbd),
	.w8(32'h392320c6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fed03a),
	.w1(32'hb8811c64),
	.w2(32'hb9f8ba02),
	.w3(32'h3a566d40),
	.w4(32'h3a207607),
	.w5(32'h38f935f2),
	.w6(32'h3a20915a),
	.w7(32'h39669984),
	.w8(32'h39b3e2c2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a59f6e),
	.w1(32'hba4f113f),
	.w2(32'hba0a0408),
	.w3(32'h3a829751),
	.w4(32'hba095c3c),
	.w5(32'hba3b7f39),
	.w6(32'hb97645b9),
	.w7(32'hb9e7b13b),
	.w8(32'hb9d76144),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba398929),
	.w1(32'hb90bb5d8),
	.w2(32'hb9a07381),
	.w3(32'hba2ed9e1),
	.w4(32'h388bd461),
	.w5(32'hb86b0ae2),
	.w6(32'h36107ad9),
	.w7(32'hb8d33e54),
	.w8(32'h37fef0e0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba516425),
	.w1(32'hbaa06655),
	.w2(32'hbac1f264),
	.w3(32'hb99bf266),
	.w4(32'hba20f140),
	.w5(32'hb9e6149a),
	.w6(32'hb96eefbf),
	.w7(32'hb963b917),
	.w8(32'hb9ce20cf),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb754f78d),
	.w1(32'hb9205826),
	.w2(32'hb9441f07),
	.w3(32'h38f172be),
	.w4(32'hb7d628b1),
	.w5(32'h36df1a44),
	.w6(32'hb9223f8e),
	.w7(32'hb8fe121d),
	.w8(32'hb89012fa),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f0a48),
	.w1(32'hb9d87052),
	.w2(32'hba8fdef4),
	.w3(32'h39eff4d2),
	.w4(32'h3906f0aa),
	.w5(32'hb9a1027f),
	.w6(32'hba5dc3ac),
	.w7(32'hba8d05e7),
	.w8(32'hba5d5767),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5494f3),
	.w1(32'hb992e1b8),
	.w2(32'h3a2ffcbc),
	.w3(32'hb9dbad3b),
	.w4(32'h396a3fe2),
	.w5(32'hba8b520f),
	.w6(32'h3a0d2d62),
	.w7(32'h3a55ed69),
	.w8(32'h39ff44f6),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa0364),
	.w1(32'hb8e65794),
	.w2(32'h38bd6aa7),
	.w3(32'hb8e3e79b),
	.w4(32'h3abbc30c),
	.w5(32'h3a86ebe6),
	.w6(32'h3aae0c43),
	.w7(32'h3a68b4c0),
	.w8(32'h3a81b0e9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c819fd),
	.w1(32'hba4066b8),
	.w2(32'hba90bc2f),
	.w3(32'h3a44eb9f),
	.w4(32'hba693007),
	.w5(32'hbaa688ca),
	.w6(32'hba4a9f3a),
	.w7(32'hba83aec3),
	.w8(32'hba38d399),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec5ab),
	.w1(32'hba773a24),
	.w2(32'hb974f103),
	.w3(32'h39aa0138),
	.w4(32'h3a834d35),
	.w5(32'h3aec499c),
	.w6(32'h3ac875b7),
	.w7(32'h3a3165a1),
	.w8(32'h3a544afe),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f5327e),
	.w1(32'hba58ce1a),
	.w2(32'hba31c818),
	.w3(32'h39940aae),
	.w4(32'hb861d32f),
	.w5(32'h3791cc6d),
	.w6(32'hb9b4d349),
	.w7(32'hb9e1f958),
	.w8(32'hba188211),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa0639),
	.w1(32'hbb0ab72d),
	.w2(32'hb99b1329),
	.w3(32'hb9bc2fa5),
	.w4(32'hbab0bef4),
	.w5(32'h399fae20),
	.w6(32'hba82cc6b),
	.w7(32'hbaa7ed42),
	.w8(32'h394d3bb7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f6b10),
	.w1(32'hb9ee5f54),
	.w2(32'hba4912e2),
	.w3(32'hba142efb),
	.w4(32'hb9e7275b),
	.w5(32'hba200015),
	.w6(32'hb9fac92c),
	.w7(32'hba11cf85),
	.w8(32'hb9e60f93),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba034cde),
	.w1(32'hba415e38),
	.w2(32'hba061f36),
	.w3(32'hba146422),
	.w4(32'hba1429be),
	.w5(32'hb9c7773b),
	.w6(32'hba2c6ad9),
	.w7(32'hba464b93),
	.w8(32'hba0f36c8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fb87f4),
	.w1(32'hb97cf649),
	.w2(32'hb9de9d09),
	.w3(32'h3a82d109),
	.w4(32'hba08225f),
	.w5(32'hbab88b0b),
	.w6(32'hba866acf),
	.w7(32'hba8e3101),
	.w8(32'hba2b88e6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f76e4),
	.w1(32'hbab2cbdd),
	.w2(32'hbaeea446),
	.w3(32'h3a294669),
	.w4(32'h38796717),
	.w5(32'hba890009),
	.w6(32'hbb10f7ec),
	.w7(32'hbb1a05dc),
	.w8(32'hbaf75017),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfccec),
	.w1(32'hba8996a9),
	.w2(32'h3a82b6dd),
	.w3(32'h38c1f853),
	.w4(32'h39d42b37),
	.w5(32'h3a83be89),
	.w6(32'hb912da64),
	.w7(32'h38a4aad6),
	.w8(32'h3a64f512),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d5f66),
	.w1(32'h3a80b0c7),
	.w2(32'hba8e3f23),
	.w3(32'h3ad3be23),
	.w4(32'h3a2092a6),
	.w5(32'hba0a3d75),
	.w6(32'h3ad1762f),
	.w7(32'hb9c1d7ad),
	.w8(32'hbab8fd54),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958dbc4),
	.w1(32'hb9966082),
	.w2(32'hba08fb3a),
	.w3(32'hb7982770),
	.w4(32'hb9b86231),
	.w5(32'hb9ddcc9f),
	.w6(32'hb998c489),
	.w7(32'hb9fd3a9b),
	.w8(32'hb9829ac3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f8045),
	.w1(32'hb9fc7dff),
	.w2(32'hba271242),
	.w3(32'hba17b0ad),
	.w4(32'hba3ddc69),
	.w5(32'hba1c6fcc),
	.w6(32'hb9dd3b03),
	.w7(32'hb9e0f5ea),
	.w8(32'hb9d443b4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2a1c8),
	.w1(32'h3b438921),
	.w2(32'h3955abf3),
	.w3(32'h3ad90789),
	.w4(32'h3a8719d9),
	.w5(32'hb9dad3e6),
	.w6(32'hb9d6c0b3),
	.w7(32'hb8c40a06),
	.w8(32'hba82169f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3765c),
	.w1(32'hba3f4892),
	.w2(32'hba85ad55),
	.w3(32'hb9de9815),
	.w4(32'hba655d2d),
	.w5(32'hb9b71afe),
	.w6(32'hbb103194),
	.w7(32'hbb16adbc),
	.w8(32'hb993fbd6),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f5a12),
	.w1(32'h391aa98d),
	.w2(32'hba728d84),
	.w3(32'h39d31b41),
	.w4(32'hb9ad0f69),
	.w5(32'hba155111),
	.w6(32'hbad5c562),
	.w7(32'hba38138a),
	.w8(32'hbacb2012),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88dd7b8),
	.w1(32'hba4371ff),
	.w2(32'hba231efe),
	.w3(32'hb78e7319),
	.w4(32'hba20b95b),
	.w5(32'hba8a348c),
	.w6(32'hb9bdce35),
	.w7(32'hba87d6da),
	.w8(32'hba692dc5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b78d7),
	.w1(32'hbb14030d),
	.w2(32'hb9fc289e),
	.w3(32'hb8e5ac3c),
	.w4(32'hba084182),
	.w5(32'h3a03a959),
	.w6(32'hb8d4d9e7),
	.w7(32'hb9c2cd7c),
	.w8(32'hb8466fc3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d3152),
	.w1(32'hba0c8318),
	.w2(32'hba04ab84),
	.w3(32'hb9f2fc51),
	.w4(32'hb99e864e),
	.w5(32'hb9a98f73),
	.w6(32'hb9172104),
	.w7(32'hb98ac105),
	.w8(32'hb9bdcb44),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23c152),
	.w1(32'h39ae9a45),
	.w2(32'h39ebbbe3),
	.w3(32'hba11d807),
	.w4(32'hb9dd26c8),
	.w5(32'hba2c04ee),
	.w6(32'h394ede3e),
	.w7(32'h3a2c64a0),
	.w8(32'h3a8a296e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55e907),
	.w1(32'hb9adb0d3),
	.w2(32'hb9756380),
	.w3(32'hb9d8863e),
	.w4(32'hba45944f),
	.w5(32'hba09b252),
	.w6(32'hb98327f3),
	.w7(32'hb9bba0a3),
	.w8(32'hb98e9c96),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9156951),
	.w1(32'hb950ff62),
	.w2(32'hba28250a),
	.w3(32'h3732aadf),
	.w4(32'hb99a1e33),
	.w5(32'hba2ce521),
	.w6(32'h34b049ba),
	.w7(32'hb9bd25b1),
	.w8(32'h3906fd07),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51e026),
	.w1(32'hb8249a2c),
	.w2(32'hba8cd739),
	.w3(32'h3a13cdf1),
	.w4(32'hb9ff6282),
	.w5(32'hbaa77d0e),
	.w6(32'hb9742367),
	.w7(32'hba3cea63),
	.w8(32'hba79bb25),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9888be),
	.w1(32'hbb1e62e3),
	.w2(32'hbb35693b),
	.w3(32'h3916e3c7),
	.w4(32'hbaa0c540),
	.w5(32'hbaf6022f),
	.w6(32'hbaab52fe),
	.w7(32'hbaca59e0),
	.w8(32'hbad0bf85),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c88a2),
	.w1(32'hba320c9f),
	.w2(32'hba08c3ce),
	.w3(32'h3775f882),
	.w4(32'hb980d788),
	.w5(32'hb9837233),
	.w6(32'h3919115d),
	.w7(32'h39e7cb90),
	.w8(32'hb8fe73f4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05cd1e),
	.w1(32'h39237adb),
	.w2(32'h39f097e1),
	.w3(32'hba4df823),
	.w4(32'hb8123599),
	.w5(32'hb9847946),
	.w6(32'hb9bb279c),
	.w7(32'h3939068b),
	.w8(32'h3a1afdbd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac992b5),
	.w1(32'hb925bbed),
	.w2(32'hb9f930e6),
	.w3(32'hba6e2eaa),
	.w4(32'h3934c6e6),
	.w5(32'h3984f3f8),
	.w6(32'hba582738),
	.w7(32'hb94a50dd),
	.w8(32'hba2952da),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57e5a2),
	.w1(32'h39791ff7),
	.w2(32'hb9b57523),
	.w3(32'h3ab52911),
	.w4(32'h391a2c89),
	.w5(32'hb710f2aa),
	.w6(32'hb9d4a260),
	.w7(32'hba2f928c),
	.w8(32'hb8d14de5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4f06d),
	.w1(32'h38f953fc),
	.w2(32'hb780c5d3),
	.w3(32'h381780f8),
	.w4(32'h39e6df18),
	.w5(32'h39bc8fc0),
	.w6(32'h3a0b7602),
	.w7(32'h39a82e3d),
	.w8(32'h3a047f08),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f5b3d),
	.w1(32'hb7931b82),
	.w2(32'hba04adaa),
	.w3(32'h3a5d7745),
	.w4(32'hb9304386),
	.w5(32'hb9f2fa4b),
	.w6(32'hba066410),
	.w7(32'hba07dc89),
	.w8(32'hb9a9a49b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3877b8c7),
	.w1(32'hba0dbfbe),
	.w2(32'hba1a64b6),
	.w3(32'h38a03615),
	.w4(32'hb9f68d8b),
	.w5(32'hba10cf7e),
	.w6(32'hb9816e4c),
	.w7(32'hb9cf40ce),
	.w8(32'hb9bd5725),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ebd03),
	.w1(32'hb935ddc9),
	.w2(32'hb9849271),
	.w3(32'hba1f5fbd),
	.w4(32'hb7dde148),
	.w5(32'hb810a5b7),
	.w6(32'hb94cadb0),
	.w7(32'hb9282be8),
	.w8(32'hb9770504),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9268e81),
	.w1(32'h394690a1),
	.w2(32'h38a789a5),
	.w3(32'hb8644004),
	.w4(32'h3a135cb1),
	.w5(32'h3a02da9c),
	.w6(32'h3a127b9a),
	.w7(32'h39c54d1d),
	.w8(32'h3a113cbc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0212b),
	.w1(32'hb9a1e227),
	.w2(32'hba62bc83),
	.w3(32'h3a1eb024),
	.w4(32'hb9cef146),
	.w5(32'hb9f22e41),
	.w6(32'hb9bf7a15),
	.w7(32'hba398fcf),
	.w8(32'hb9acd502),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9370a),
	.w1(32'h39eec0b4),
	.w2(32'h39389d8d),
	.w3(32'hb99585a2),
	.w4(32'h3a152081),
	.w5(32'h38a80992),
	.w6(32'hb9e455f6),
	.w7(32'hb8c8593a),
	.w8(32'hb864960b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a477f9a),
	.w1(32'h39a4d3ad),
	.w2(32'hbac1f863),
	.w3(32'h3ab231f7),
	.w4(32'h39fac80e),
	.w5(32'h3a4dfc11),
	.w6(32'h3a5c9322),
	.w7(32'hb9d2edaf),
	.w8(32'h38404143),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a739c6b),
	.w1(32'hb9929e01),
	.w2(32'hba04734a),
	.w3(32'h3a9b4382),
	.w4(32'h38a07678),
	.w5(32'h397e13aa),
	.w6(32'hb90bc621),
	.w7(32'hba411ce9),
	.w8(32'h38a1ca0e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7be9192),
	.w1(32'hba3766ac),
	.w2(32'hba969374),
	.w3(32'h39a8da9c),
	.w4(32'h3963f8fa),
	.w5(32'h399d478a),
	.w6(32'hb9fdd45d),
	.w7(32'hba84f4de),
	.w8(32'hba482b3c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b55760),
	.w1(32'h397aa1c2),
	.w2(32'hb6722a17),
	.w3(32'hb99f407d),
	.w4(32'h39fd4b2d),
	.w5(32'h3a0b4375),
	.w6(32'h39ba080f),
	.w7(32'h39fc63c6),
	.w8(32'h39e1130d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b08108),
	.w1(32'h38d0517e),
	.w2(32'hb94cde4c),
	.w3(32'h396824b6),
	.w4(32'h3a3190bc),
	.w5(32'h3a0b7a39),
	.w6(32'h3a409320),
	.w7(32'h39f4dcdb),
	.w8(32'h3a22c491),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c05361),
	.w1(32'hb816614a),
	.w2(32'hb8b62ca3),
	.w3(32'h3a5ccb9e),
	.w4(32'h39abc499),
	.w5(32'h396f1efd),
	.w6(32'h39710f23),
	.w7(32'h39346fc6),
	.w8(32'h399e760c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b3595),
	.w1(32'hb858bc0b),
	.w2(32'hb92d4d82),
	.w3(32'h399e5598),
	.w4(32'h39bf8948),
	.w5(32'h39562b06),
	.w6(32'h39982fa3),
	.w7(32'h391dadc7),
	.w8(32'h39a313f6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39100b89),
	.w1(32'hbaa38634),
	.w2(32'hbae95418),
	.w3(32'h3a0cf09a),
	.w4(32'hba6bc25b),
	.w5(32'hba5a08e8),
	.w6(32'hb91a7d28),
	.w7(32'hba85d05d),
	.w8(32'hb9c8eac0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ef8c5),
	.w1(32'hba3bfbc0),
	.w2(32'hba50182e),
	.w3(32'hb9af2b9e),
	.w4(32'hba6f59ac),
	.w5(32'hba6be196),
	.w6(32'hba29bf99),
	.w7(32'hba4d157c),
	.w8(32'hba9b2674),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22da71),
	.w1(32'hb8ba07a8),
	.w2(32'hba347d67),
	.w3(32'hba81003d),
	.w4(32'h36a63091),
	.w5(32'hba27f439),
	.w6(32'hba0538f5),
	.w7(32'hba154283),
	.w8(32'hba34f955),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a7688),
	.w1(32'hba8f6d9b),
	.w2(32'hbaa981b0),
	.w3(32'hba4ce398),
	.w4(32'hba7cbe98),
	.w5(32'hba653bbf),
	.w6(32'hb99e266b),
	.w7(32'hb994c035),
	.w8(32'hb981d645),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a6743),
	.w1(32'h3999fdd2),
	.w2(32'h38c14bb7),
	.w3(32'hb91328c7),
	.w4(32'h3a103be7),
	.w5(32'h39e8f263),
	.w6(32'h3a0dbd00),
	.w7(32'h39ddec1a),
	.w8(32'h39bf94b3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abdb9a),
	.w1(32'h3a6c76e5),
	.w2(32'h3acd1e31),
	.w3(32'h3a43c0d5),
	.w4(32'hb9f4766c),
	.w5(32'hba34562c),
	.w6(32'h3a396dbf),
	.w7(32'h39a09c60),
	.w8(32'h3a695c4a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97e81a),
	.w1(32'hba8085a7),
	.w2(32'hbad01024),
	.w3(32'hb9d486e8),
	.w4(32'hba61532f),
	.w5(32'hba9b26af),
	.w6(32'hba21fc2e),
	.w7(32'hba3659f8),
	.w8(32'hba0b6845),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9940427),
	.w1(32'hbb0cc9c1),
	.w2(32'hbbab5853),
	.w3(32'hbab579ab),
	.w4(32'hbb00ee0d),
	.w5(32'hba4c3e93),
	.w6(32'hbaecdcb8),
	.w7(32'hbaf7bcc2),
	.w8(32'hb9665b7e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a38e7),
	.w1(32'hb5f74491),
	.w2(32'hb8070d3c),
	.w3(32'hb990099f),
	.w4(32'hb862f453),
	.w5(32'hb897a666),
	.w6(32'hb8224336),
	.w7(32'hb8c8bcf7),
	.w8(32'hb8cd4877),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bce9ad),
	.w1(32'hba041ecc),
	.w2(32'h3a3001bd),
	.w3(32'h38a22436),
	.w4(32'h389e53fe),
	.w5(32'h39853d0f),
	.w6(32'hba852a10),
	.w7(32'hba975021),
	.w8(32'hba0081c0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule