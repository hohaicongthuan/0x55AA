module layer_10_featuremap_460(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9681786),
	.w1(32'hbb973d4f),
	.w2(32'hbab8279a),
	.w3(32'h3b89075a),
	.w4(32'h382c0f67),
	.w5(32'hba9fae90),
	.w6(32'h3a8187ef),
	.w7(32'h3b8aa2d4),
	.w8(32'h3b364052),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a67f18),
	.w1(32'h3c1c7b60),
	.w2(32'hbbb19a5b),
	.w3(32'h3b0e9fb7),
	.w4(32'h3b29d08a),
	.w5(32'h3c485cec),
	.w6(32'h390f95be),
	.w7(32'hbb8ebe6c),
	.w8(32'h3bf916e4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c74ec),
	.w1(32'hbb14ec69),
	.w2(32'hbc03b325),
	.w3(32'hbba20151),
	.w4(32'h3c3aefce),
	.w5(32'hba7f85c2),
	.w6(32'h3b1035aa),
	.w7(32'hba81cb64),
	.w8(32'h3c3e94a3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89af1f),
	.w1(32'hbac69ddb),
	.w2(32'h391f43d7),
	.w3(32'hbc104f53),
	.w4(32'hbbb8a5a6),
	.w5(32'h3bb37bcf),
	.w6(32'hbbe783ea),
	.w7(32'hbb05676d),
	.w8(32'h3acdcac9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b676e),
	.w1(32'hbb7ea6e6),
	.w2(32'hba8ae995),
	.w3(32'h3b4101a3),
	.w4(32'h3b637b46),
	.w5(32'hbb040586),
	.w6(32'h3c148886),
	.w7(32'h3b8c51ae),
	.w8(32'h3ad863fd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55f2c9),
	.w1(32'hba02efc1),
	.w2(32'h3a7b2ea2),
	.w3(32'h3adba4a9),
	.w4(32'h3b4b62cc),
	.w5(32'h3a984ddc),
	.w6(32'hbb6b2598),
	.w7(32'h3af73fdd),
	.w8(32'hb9ce9abb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be992e1),
	.w1(32'h3b8a698a),
	.w2(32'hbafdad34),
	.w3(32'h3bdd06cc),
	.w4(32'hbafed3d3),
	.w5(32'hbb92fb51),
	.w6(32'hbabbbb2c),
	.w7(32'hbbcfb4f7),
	.w8(32'h3c02cc77),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb931b14),
	.w1(32'hbcbe98ba),
	.w2(32'hbbdca2f5),
	.w3(32'hbc39ff0a),
	.w4(32'h3acdec1a),
	.w5(32'hbad69823),
	.w6(32'hbb21aec8),
	.w7(32'hb846b8ca),
	.w8(32'h3b029691),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba412d6),
	.w1(32'h397533f1),
	.w2(32'h3b485214),
	.w3(32'hbc426b61),
	.w4(32'hbb5945e6),
	.w5(32'h3ae7b4d0),
	.w6(32'hbb322c91),
	.w7(32'hbaf43a1f),
	.w8(32'hbbb65379),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dce0d0),
	.w1(32'hba2892f7),
	.w2(32'h3b21c48f),
	.w3(32'h3b6f4f23),
	.w4(32'hbb6eb09d),
	.w5(32'hbc38d6ec),
	.w6(32'hbafe8619),
	.w7(32'hba3f7607),
	.w8(32'hbbcf97ca),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb062bc3),
	.w1(32'hbb307599),
	.w2(32'hbaa4f8dd),
	.w3(32'h3b12ce7c),
	.w4(32'h3ba5db3c),
	.w5(32'h3a8b3f29),
	.w6(32'hbbc6304b),
	.w7(32'h3b4f247a),
	.w8(32'h3a09157f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6c417),
	.w1(32'hbb04a46d),
	.w2(32'h3b28720c),
	.w3(32'h3bf2ff99),
	.w4(32'h3a60de25),
	.w5(32'h3a4b4094),
	.w6(32'hbab0d39f),
	.w7(32'h3b0dcfa3),
	.w8(32'hbaaf918b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eaf6f),
	.w1(32'hb9bf271c),
	.w2(32'hbae1cad2),
	.w3(32'h3b9166b6),
	.w4(32'hbc0ac03c),
	.w5(32'h3b840656),
	.w6(32'h3a41f90b),
	.w7(32'hbbc160fc),
	.w8(32'hbba9c491),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fb24c),
	.w1(32'hbbdccd0c),
	.w2(32'hbb1446eb),
	.w3(32'h3aaa4ff5),
	.w4(32'h3b0b8962),
	.w5(32'hbb1f68f3),
	.w6(32'h39d5cae2),
	.w7(32'h3ad2aedb),
	.w8(32'hbb4db769),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f367b),
	.w1(32'h3b999a60),
	.w2(32'hba69aec2),
	.w3(32'h3b23f40e),
	.w4(32'hbb071ec1),
	.w5(32'h3a913f66),
	.w6(32'h3b0df027),
	.w7(32'hbb0363d3),
	.w8(32'hbb3ed2ef),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa687),
	.w1(32'hb9b507bc),
	.w2(32'hbbcf01b4),
	.w3(32'hba8bb40d),
	.w4(32'hbbf1bf3f),
	.w5(32'hbba418bf),
	.w6(32'hbb63c42e),
	.w7(32'hbbc59ef0),
	.w8(32'hbbca34b9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b497073),
	.w1(32'hbb1dad33),
	.w2(32'hbaa1bee8),
	.w3(32'h3acb5e2d),
	.w4(32'hbb41cdf1),
	.w5(32'hba3727ff),
	.w6(32'hb908c2f9),
	.w7(32'hb9accb60),
	.w8(32'h3a99512b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba922a),
	.w1(32'hbc8a7374),
	.w2(32'hbc0f46fa),
	.w3(32'hbc08030a),
	.w4(32'hbbb8e4b7),
	.w5(32'hbbfb6490),
	.w6(32'hbbc37946),
	.w7(32'h3bb4516c),
	.w8(32'h3af39a39),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29b54e),
	.w1(32'hbbea82b9),
	.w2(32'hbaa4e62d),
	.w3(32'hbb9cac90),
	.w4(32'hbb9dceab),
	.w5(32'hba419e2a),
	.w6(32'hbbdbd288),
	.w7(32'h3a8fd94c),
	.w8(32'h3a5a77e8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db2c10),
	.w1(32'h3ac52b8c),
	.w2(32'h3b2c5a57),
	.w3(32'hbaa1dae3),
	.w4(32'hbbe49679),
	.w5(32'h3bc2f30d),
	.w6(32'h3a83891a),
	.w7(32'hbbb034b7),
	.w8(32'hbc1377e9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3726ce),
	.w1(32'hbabc91cc),
	.w2(32'h3a47df12),
	.w3(32'h394787a2),
	.w4(32'h3b309c43),
	.w5(32'hbabf2550),
	.w6(32'h3ba8e28c),
	.w7(32'h3b3d8885),
	.w8(32'hba85b546),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15cfa8),
	.w1(32'h3a24a285),
	.w2(32'h3b26ab72),
	.w3(32'h3b888ed3),
	.w4(32'hbbb6ccbe),
	.w5(32'h3b25ed54),
	.w6(32'h3ba1f6fb),
	.w7(32'hbbc0fda0),
	.w8(32'hba9e62ca),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba19e3f),
	.w1(32'hbc8a571d),
	.w2(32'h3b605c58),
	.w3(32'hbc938b01),
	.w4(32'hbc0f183d),
	.w5(32'h3b3fda7b),
	.w6(32'hbc7c97cc),
	.w7(32'h3b45d6a6),
	.w8(32'h3a103cd9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24048a),
	.w1(32'hba4ed631),
	.w2(32'hbae7e664),
	.w3(32'h3c0023af),
	.w4(32'hbb4faa19),
	.w5(32'hbbbb360b),
	.w6(32'h3b96c1b3),
	.w7(32'hba8404e4),
	.w8(32'hbbe377a7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b88e3),
	.w1(32'h3b883717),
	.w2(32'hbbc14a95),
	.w3(32'hba8c9555),
	.w4(32'hba2ac657),
	.w5(32'hbc172ab6),
	.w6(32'hbaf33cd9),
	.w7(32'hbc7d9dd5),
	.w8(32'hbc50267a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a154c),
	.w1(32'hbb887023),
	.w2(32'hbb389798),
	.w3(32'hba8543d2),
	.w4(32'h3b3a2c87),
	.w5(32'hbb9aa52b),
	.w6(32'hbb84480e),
	.w7(32'h39cfff11),
	.w8(32'hbb9a18d5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9fa8f),
	.w1(32'hbb83c117),
	.w2(32'hbb3d60ee),
	.w3(32'h3b0910d0),
	.w4(32'hba604ed2),
	.w5(32'hbbc23641),
	.w6(32'hba8e06b6),
	.w7(32'hbadb9118),
	.w8(32'hbaf53d98),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36af99),
	.w1(32'hbadc21d3),
	.w2(32'h3b859e15),
	.w3(32'hbb881bd0),
	.w4(32'hbb88538f),
	.w5(32'hbc0e9de4),
	.w6(32'hb9da1ab9),
	.w7(32'hba607249),
	.w8(32'hbb91b02d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9cd12),
	.w1(32'hbbd130a1),
	.w2(32'hbbcf1e98),
	.w3(32'h3b0f93e2),
	.w4(32'hba00a51c),
	.w5(32'hbba317c7),
	.w6(32'hbb63f13a),
	.w7(32'h3b8bfa82),
	.w8(32'hbaf52682),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a785bad),
	.w1(32'h3bc803ae),
	.w2(32'hba8d23c9),
	.w3(32'h3c31a82c),
	.w4(32'h3b284c94),
	.w5(32'hbc0e746d),
	.w6(32'h3c3b7e83),
	.w7(32'hb9ef7670),
	.w8(32'hbc0d13a5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6127b8),
	.w1(32'hbb978fa8),
	.w2(32'hbb79b96f),
	.w3(32'h3b926d00),
	.w4(32'hbae8fb8f),
	.w5(32'hbb11376f),
	.w6(32'h3b8ac2a1),
	.w7(32'h3bc6db51),
	.w8(32'h3a1d5c89),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4432d5),
	.w1(32'h3ba9f7f6),
	.w2(32'hbba5779e),
	.w3(32'h3b3130b0),
	.w4(32'h3b3901e7),
	.w5(32'h3c3e1f3f),
	.w6(32'h3a6cdaa6),
	.w7(32'hbb92b70d),
	.w8(32'h3c232079),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4c3c5),
	.w1(32'h3bda7be2),
	.w2(32'hbb554462),
	.w3(32'hbc15399b),
	.w4(32'h3b46bde7),
	.w5(32'h3c1a8705),
	.w6(32'hbb2e1dc4),
	.w7(32'hbb317f9b),
	.w8(32'h3c5effc0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7f435),
	.w1(32'h3b4a924f),
	.w2(32'hbb94f1ec),
	.w3(32'hbb74ecc6),
	.w4(32'hbae7980e),
	.w5(32'hbbb6f5d6),
	.w6(32'hbbc98e24),
	.w7(32'hbbb5894d),
	.w8(32'hbab061f2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43a7a6),
	.w1(32'hb992b7ac),
	.w2(32'h39a30008),
	.w3(32'hba93579d),
	.w4(32'h3b9067e7),
	.w5(32'hbbce6d5d),
	.w6(32'hbbcbf1aa),
	.w7(32'h3b4129ec),
	.w8(32'hbc382648),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be89425),
	.w1(32'h3a0bce18),
	.w2(32'hbad570fb),
	.w3(32'hbb0d6485),
	.w4(32'hbb86307b),
	.w5(32'h3b749717),
	.w6(32'hbb06dd56),
	.w7(32'h3ab28312),
	.w8(32'h3a0d057b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07a147),
	.w1(32'hbbd36730),
	.w2(32'hbc05cd12),
	.w3(32'h3c33535d),
	.w4(32'hbb405dd6),
	.w5(32'h3bde5c02),
	.w6(32'h3bb12064),
	.w7(32'hbc202ed1),
	.w8(32'hbafeb969),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e66ef),
	.w1(32'h3cbf3fcf),
	.w2(32'hbc196bc1),
	.w3(32'h3c3d40d0),
	.w4(32'h3ad68382),
	.w5(32'h3c97f303),
	.w6(32'h3bc02114),
	.w7(32'hbc861077),
	.w8(32'h3b9007cc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb6fbc),
	.w1(32'h3b612dc0),
	.w2(32'hbb2d4ee8),
	.w3(32'hbac77a9f),
	.w4(32'h3b67e992),
	.w5(32'hbc6f1977),
	.w6(32'h3c2ff614),
	.w7(32'h3ba96a5e),
	.w8(32'hbc22c77a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb78233),
	.w1(32'h3b12f350),
	.w2(32'h3bc3ff0e),
	.w3(32'h3bf1091b),
	.w4(32'hbb9de476),
	.w5(32'h3c792b02),
	.w6(32'hb9e82d43),
	.w7(32'hbb9eb0a7),
	.w8(32'h3b2602b6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bc3e7),
	.w1(32'hbc001970),
	.w2(32'h3c4e4186),
	.w3(32'hbba7bb22),
	.w4(32'hbbbcb457),
	.w5(32'h3c2c53a0),
	.w6(32'h3bf00052),
	.w7(32'hbb2d68df),
	.w8(32'h3b13878e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36a167),
	.w1(32'h3b1c7e42),
	.w2(32'h3b1d2431),
	.w3(32'hbb99dbcf),
	.w4(32'hbb5d19f0),
	.w5(32'h3bf30b8c),
	.w6(32'h3bfee81f),
	.w7(32'h3a403a91),
	.w8(32'h3ad553cc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8885c2),
	.w1(32'h3bc1f940),
	.w2(32'hbc4eddb3),
	.w3(32'hbba16ffd),
	.w4(32'hbbbab057),
	.w5(32'h3ba7923c),
	.w6(32'hba844406),
	.w7(32'hbc191b94),
	.w8(32'h3b72652b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd889),
	.w1(32'hbb6f290e),
	.w2(32'hba75a3b6),
	.w3(32'hbc2d19b5),
	.w4(32'h3a7eca62),
	.w5(32'hbb634378),
	.w6(32'hbb9ae340),
	.w7(32'h3b86130a),
	.w8(32'h3a8b90f6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54b8b0),
	.w1(32'hba15f8b8),
	.w2(32'hba9aad09),
	.w3(32'hba428860),
	.w4(32'hbaf42508),
	.w5(32'hbbd69ce7),
	.w6(32'h3b12c057),
	.w7(32'hbbbdf8e3),
	.w8(32'hbba5b7eb),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac0df),
	.w1(32'h3b98f8fa),
	.w2(32'hbac3fe7e),
	.w3(32'hbb3ca78f),
	.w4(32'hbb1a78e6),
	.w5(32'hbb5a9095),
	.w6(32'hbb75d569),
	.w7(32'hbbed60d2),
	.w8(32'hbb878ade),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ef4c3),
	.w1(32'hbb0ffd0a),
	.w2(32'h3bb113d4),
	.w3(32'hbbd67777),
	.w4(32'h3b138164),
	.w5(32'hbb8e7dfb),
	.w6(32'hbbb95fe2),
	.w7(32'h3a86ddcf),
	.w8(32'hbb27d607),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2639c),
	.w1(32'hbc4ed517),
	.w2(32'h3acb35aa),
	.w3(32'hbc03f418),
	.w4(32'hbc20d24c),
	.w5(32'h3c195ef0),
	.w6(32'hbbcc2e43),
	.w7(32'hba1b56be),
	.w8(32'h3be467e4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa66469),
	.w1(32'hbbdf8015),
	.w2(32'h3afb101f),
	.w3(32'h3afbee29),
	.w4(32'hbb0cd720),
	.w5(32'hbbaddbaf),
	.w6(32'h3bb6573f),
	.w7(32'h3b8806a4),
	.w8(32'hbb0a6cac),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba42df4),
	.w1(32'hb936fbf8),
	.w2(32'hbb105e10),
	.w3(32'h3aadf4e3),
	.w4(32'hb920974e),
	.w5(32'hbab161f0),
	.w6(32'hb79db39b),
	.w7(32'hba965079),
	.w8(32'hbab93c79),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93377e),
	.w1(32'h3b37bb44),
	.w2(32'hbb019524),
	.w3(32'hbb3a26f0),
	.w4(32'h3b50e0e1),
	.w5(32'hbbd80223),
	.w6(32'h3b309a6a),
	.w7(32'h3b4df910),
	.w8(32'hbb7d3537),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ee37),
	.w1(32'hba7eed68),
	.w2(32'h39a95121),
	.w3(32'hba0775bc),
	.w4(32'h3b10d9ba),
	.w5(32'h3b959641),
	.w6(32'hbb9bcc34),
	.w7(32'hba4b2d0c),
	.w8(32'h3bb2c680),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf1c55),
	.w1(32'hbac28db9),
	.w2(32'hba2a75d7),
	.w3(32'hbbc03cbc),
	.w4(32'hbad914f6),
	.w5(32'hbb659ccb),
	.w6(32'h3a483c0f),
	.w7(32'hbbab40c3),
	.w8(32'h39f95991),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03039a),
	.w1(32'hbbdf4932),
	.w2(32'hbbd49057),
	.w3(32'hbc4d967e),
	.w4(32'hbb9aa396),
	.w5(32'h3bb6b1fb),
	.w6(32'hbbc4d80b),
	.w7(32'hbbbf1f25),
	.w8(32'h3c084f2e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce11a7),
	.w1(32'h3b1cc085),
	.w2(32'hbb7e3a01),
	.w3(32'hbc08bd14),
	.w4(32'hbb923b36),
	.w5(32'h3ca88c2e),
	.w6(32'hbb4b2253),
	.w7(32'hbb961da6),
	.w8(32'h3bd11d6f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aad1c3),
	.w1(32'h3c0a15be),
	.w2(32'hbc42d75d),
	.w3(32'hbbd02c2d),
	.w4(32'h3ae5740b),
	.w5(32'h3cb6ade2),
	.w6(32'h3b6f20db),
	.w7(32'hbbcd4c91),
	.w8(32'h3c83d30b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb319bd1),
	.w1(32'hbb516d67),
	.w2(32'hbb7fe115),
	.w3(32'hbbca9712),
	.w4(32'hba667914),
	.w5(32'hbb5ee34a),
	.w6(32'hbbab8e8a),
	.w7(32'h3a7a2d1c),
	.w8(32'hba87adaf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143e40),
	.w1(32'h3af693b0),
	.w2(32'hbb87f49c),
	.w3(32'hbae555f0),
	.w4(32'hbbb1d1c4),
	.w5(32'hb88071e0),
	.w6(32'hbac3a239),
	.w7(32'hbc1df898),
	.w8(32'hbb4162c8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ebe46),
	.w1(32'h3a616ff0),
	.w2(32'hbc159480),
	.w3(32'h395f224f),
	.w4(32'hbbaad8f9),
	.w5(32'hbbafe13d),
	.w6(32'hbaacc1a7),
	.w7(32'hbc01940e),
	.w8(32'hbb4f6baf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca25f),
	.w1(32'hbba631b9),
	.w2(32'hbb87222c),
	.w3(32'hba4b065a),
	.w4(32'hbbfda2e9),
	.w5(32'hbb136daa),
	.w6(32'hb9ce3185),
	.w7(32'hbb9e8c65),
	.w8(32'hbbd79b79),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18925b),
	.w1(32'hbbfef279),
	.w2(32'hbbd9ca53),
	.w3(32'hbbce46b1),
	.w4(32'h3a168f5c),
	.w5(32'hbb6eec4a),
	.w6(32'h3a17c4bc),
	.w7(32'h3a8fb713),
	.w8(32'hbb71c321),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc311424),
	.w1(32'hbbe576a7),
	.w2(32'h3ba43374),
	.w3(32'hbbdef8d6),
	.w4(32'hbaddb774),
	.w5(32'hb8a773b6),
	.w6(32'hbb0abc57),
	.w7(32'hb932b7ba),
	.w8(32'hbafb1f44),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920608),
	.w1(32'h3beb44f0),
	.w2(32'hbc42fb97),
	.w3(32'h3b4b5c5b),
	.w4(32'h3b3e930f),
	.w5(32'hbbb1c776),
	.w6(32'hb909cd6e),
	.w7(32'h3b3aa1c5),
	.w8(32'h3bf0820f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96eb91),
	.w1(32'h3a17a104),
	.w2(32'h39e349ec),
	.w3(32'hbb88fabc),
	.w4(32'h39056713),
	.w5(32'hbb68cc46),
	.w6(32'hba762b42),
	.w7(32'h3b4383a3),
	.w8(32'hbb23267d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01f69c),
	.w1(32'h3b67a116),
	.w2(32'h3b4fff33),
	.w3(32'hbac514dd),
	.w4(32'h3ba80744),
	.w5(32'h3b27e62f),
	.w6(32'hbb7795b0),
	.w7(32'h3b82db8e),
	.w8(32'h3a80ec5c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a910950),
	.w1(32'hbb4b99c7),
	.w2(32'h3b9b952d),
	.w3(32'h3af0dcdf),
	.w4(32'h3bb0a5d7),
	.w5(32'hba8ed63a),
	.w6(32'h3b141d87),
	.w7(32'h3b960e7f),
	.w8(32'h3a8d51a6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29aeec),
	.w1(32'hbb40a077),
	.w2(32'h3c142d34),
	.w3(32'h3be4f252),
	.w4(32'hbb99f8db),
	.w5(32'h39438055),
	.w6(32'h3a34e65a),
	.w7(32'h3a684edc),
	.w8(32'hb96f3489),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d46da),
	.w1(32'hbac90ef8),
	.w2(32'hbae7acfd),
	.w3(32'h3a87fb2d),
	.w4(32'hbb80cd40),
	.w5(32'hbbbeefc4),
	.w6(32'hbb0c16ec),
	.w7(32'h3b66614f),
	.w8(32'hbbd98d60),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37c7db),
	.w1(32'hbbc34c35),
	.w2(32'hbbeddc3f),
	.w3(32'hbb899593),
	.w4(32'h3b562937),
	.w5(32'h3a4970a0),
	.w6(32'hbb9261cc),
	.w7(32'h3b530156),
	.w8(32'h39b6c8da),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ec2c5),
	.w1(32'h3b0689c9),
	.w2(32'hbc0e72c3),
	.w3(32'h396448ba),
	.w4(32'hba4288bc),
	.w5(32'hbc046c91),
	.w6(32'hbbc5a109),
	.w7(32'hbc2af6c2),
	.w8(32'hbc59f012),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b756b23),
	.w1(32'hbb401c05),
	.w2(32'hb9da300e),
	.w3(32'h3b04f300),
	.w4(32'hbb407c9d),
	.w5(32'h3ad4715d),
	.w6(32'h3ab2124b),
	.w7(32'hbaa627f8),
	.w8(32'h3a0175fc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d02bd),
	.w1(32'hbb2af5e1),
	.w2(32'hbb8ba903),
	.w3(32'h3ab7617a),
	.w4(32'hbbcd41e1),
	.w5(32'hbb8d1cdf),
	.w6(32'hba4da520),
	.w7(32'hbbbd9a28),
	.w8(32'hbba1a97f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34ff5f),
	.w1(32'h3a5d08bb),
	.w2(32'hbace3061),
	.w3(32'hbb3b9123),
	.w4(32'h3b2df490),
	.w5(32'hbaf00d18),
	.w6(32'hba312e6f),
	.w7(32'h3afde5d8),
	.w8(32'hba5d6822),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10f2ae),
	.w1(32'hbad3daed),
	.w2(32'h3978aedb),
	.w3(32'hbc136556),
	.w4(32'h3aea73dd),
	.w5(32'h3acda1b4),
	.w6(32'hbbb4dd3a),
	.w7(32'h3a80f4fb),
	.w8(32'h3a887fee),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f82dd),
	.w1(32'h3b7bec87),
	.w2(32'h3b840fb4),
	.w3(32'h3b7a3783),
	.w4(32'hb42a21de),
	.w5(32'h3b935a2c),
	.w6(32'h3b3030fe),
	.w7(32'h3b177b96),
	.w8(32'h3b03abb9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393feafa),
	.w1(32'hbc315592),
	.w2(32'hbbf0fdd1),
	.w3(32'hbba1b6fb),
	.w4(32'hbbabf285),
	.w5(32'hb95b9732),
	.w6(32'hbab006d9),
	.w7(32'h3c0454ab),
	.w8(32'h3b7f8394),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ddd2a),
	.w1(32'hbc1085d0),
	.w2(32'hbb995236),
	.w3(32'hbb72df90),
	.w4(32'hbc14b372),
	.w5(32'h3b9acd54),
	.w6(32'hbc1fc59c),
	.w7(32'hbafea16b),
	.w8(32'hb998b78e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae35ac2),
	.w1(32'h3b56dbb2),
	.w2(32'h3b94fef0),
	.w3(32'h3b80fb0d),
	.w4(32'h3b98d48e),
	.w5(32'h3be2ba10),
	.w6(32'h3b68db75),
	.w7(32'hbb8ff3e3),
	.w8(32'hbb8f09d5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79e1ec),
	.w1(32'h3a90732b),
	.w2(32'h3c0db730),
	.w3(32'h3c1a885b),
	.w4(32'h3a6df212),
	.w5(32'h3c20ca88),
	.w6(32'h3b9275ac),
	.w7(32'h3b8bedbf),
	.w8(32'h3c0852d3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074838),
	.w1(32'hba89a6de),
	.w2(32'h3bb8b1ea),
	.w3(32'h3c146bed),
	.w4(32'h3b4e0032),
	.w5(32'h3c090301),
	.w6(32'h3bb39c21),
	.w7(32'h3b1ca6ca),
	.w8(32'h3b9f31b8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad389b0),
	.w1(32'h3b90d86b),
	.w2(32'hb9bf5c3b),
	.w3(32'hb93f818e),
	.w4(32'h398bd9f0),
	.w5(32'hbb9c9455),
	.w6(32'hb9a67c6a),
	.w7(32'hb7a48764),
	.w8(32'hbad3d924),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5899e),
	.w1(32'hbc08b94b),
	.w2(32'hbb8b89d1),
	.w3(32'h3a3b4c94),
	.w4(32'hbbe7d065),
	.w5(32'h39964e83),
	.w6(32'h3a7126a2),
	.w7(32'hbb205700),
	.w8(32'h3b480678),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba861964),
	.w1(32'h3aa30234),
	.w2(32'hb753c621),
	.w3(32'h3afa5edb),
	.w4(32'hbaebe692),
	.w5(32'hbaf28702),
	.w6(32'hb9b8c924),
	.w7(32'hba18c89e),
	.w8(32'hbac40ecf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8635a8),
	.w1(32'h3bfac958),
	.w2(32'hba6b2286),
	.w3(32'h3a43db00),
	.w4(32'h3bba12a9),
	.w5(32'hbb3814f5),
	.w6(32'h3a066b73),
	.w7(32'h3abe8e44),
	.w8(32'hbb2e7cab),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad174b4),
	.w1(32'hb99018e8),
	.w2(32'h3b8cd329),
	.w3(32'hba57b6f8),
	.w4(32'hba9193bf),
	.w5(32'h3b4ffc0f),
	.w6(32'hba3b8197),
	.w7(32'hbac76c64),
	.w8(32'h3b245079),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46f136),
	.w1(32'hba576c15),
	.w2(32'hbb896e9e),
	.w3(32'h3b55db6b),
	.w4(32'h3a9d7e8e),
	.w5(32'hbb7bdc3a),
	.w6(32'h3a993fef),
	.w7(32'hb99712fa),
	.w8(32'hbba683e8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74f7a8),
	.w1(32'h3afd86ac),
	.w2(32'h3a3079e3),
	.w3(32'h3b872f41),
	.w4(32'hbb0206e9),
	.w5(32'h3ac63b57),
	.w6(32'hbb7b66ff),
	.w7(32'hbc11dd41),
	.w8(32'hbbea4b92),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ab99a),
	.w1(32'hbb96eba9),
	.w2(32'hbb5fa131),
	.w3(32'hbb2048dd),
	.w4(32'hbae4d24e),
	.w5(32'h3b0e3fed),
	.w6(32'hbb467d78),
	.w7(32'hbbc21c29),
	.w8(32'hbb95c7d4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01119),
	.w1(32'h3a161a1f),
	.w2(32'h3b7f34a1),
	.w3(32'hba909af9),
	.w4(32'h3894f0f9),
	.w5(32'h3adca8e2),
	.w6(32'hbb366f98),
	.w7(32'hbb917795),
	.w8(32'hbab03f78),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf15950),
	.w1(32'hbc734dd8),
	.w2(32'hba845cad),
	.w3(32'hbc510b2f),
	.w4(32'hbbf5f3e3),
	.w5(32'h3c48ad2b),
	.w6(32'hbc25e8d6),
	.w7(32'h3b37565b),
	.w8(32'h3c0bbbd0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9603aa),
	.w1(32'hb9aea700),
	.w2(32'hbb914057),
	.w3(32'hbac2ef20),
	.w4(32'hbaee21b3),
	.w5(32'hbb85c588),
	.w6(32'hbb1a2a8b),
	.w7(32'hbae43e77),
	.w8(32'hbb4e6ae5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b528b9c),
	.w1(32'h39d70274),
	.w2(32'h38ba7cec),
	.w3(32'h3b6240b6),
	.w4(32'hbac049d2),
	.w5(32'hbaecfb09),
	.w6(32'hbadf4442),
	.w7(32'hb9f9a9ae),
	.w8(32'hbb1d1b72),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb166e6),
	.w1(32'hbb096a5f),
	.w2(32'hbb6d3a9e),
	.w3(32'hbac4cb01),
	.w4(32'h3b243f73),
	.w5(32'h3a0966a2),
	.w6(32'hbb7b84e1),
	.w7(32'h3b59af58),
	.w8(32'h3b3ebed6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab481f1),
	.w1(32'h3b19fd9d),
	.w2(32'h3b48f8a3),
	.w3(32'h3a72d13b),
	.w4(32'h3ba25eb0),
	.w5(32'h3b428fbe),
	.w6(32'h3a9a7257),
	.w7(32'h3b290040),
	.w8(32'h39c3c27d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afca8bf),
	.w1(32'h3b16fc70),
	.w2(32'hbb7c6f3c),
	.w3(32'h3ba1eeec),
	.w4(32'hba756141),
	.w5(32'hbbac2498),
	.w6(32'h3b104aba),
	.w7(32'hbbb6574d),
	.w8(32'hbbe75dec),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba938d34),
	.w1(32'h3c12b9b2),
	.w2(32'h3bab081e),
	.w3(32'h3a9e79c1),
	.w4(32'h3c22f65f),
	.w5(32'h3bb81f8d),
	.w6(32'hbaf40060),
	.w7(32'h3b0e04b0),
	.w8(32'h3adeb486),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0fdd1),
	.w1(32'h3a31be7c),
	.w2(32'hba613d33),
	.w3(32'hbb3292c7),
	.w4(32'h3b75394a),
	.w5(32'h3b291593),
	.w6(32'hbb2ace21),
	.w7(32'h396ee7a6),
	.w8(32'hbaa63e4e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf73a7d),
	.w1(32'hbab0bfb8),
	.w2(32'hbb0a97fa),
	.w3(32'hb93176aa),
	.w4(32'hb9c31088),
	.w5(32'hbba9855f),
	.w6(32'hbbae50d3),
	.w7(32'h3aad6a2e),
	.w8(32'hbb392956),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb6d65),
	.w1(32'hbb91c0a4),
	.w2(32'hbb3f145a),
	.w3(32'h3b79d544),
	.w4(32'hbb14483c),
	.w5(32'hbb8e81fa),
	.w6(32'h3a9fef07),
	.w7(32'h3a57f388),
	.w8(32'h3a4038d4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1ebe4),
	.w1(32'hbc9ae0ec),
	.w2(32'hbc1c5e33),
	.w3(32'hbc529cf5),
	.w4(32'hbc65952b),
	.w5(32'h3b9e58cc),
	.w6(32'hbc935731),
	.w7(32'h3a59e455),
	.w8(32'hb85b6688),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818dbc),
	.w1(32'h3bb905bc),
	.w2(32'hbb4d545d),
	.w3(32'h3a9b7b5b),
	.w4(32'hba8aaeab),
	.w5(32'hbbcd7e64),
	.w6(32'h3b4d51de),
	.w7(32'hbbc91746),
	.w8(32'hbc32c28c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b544e6f),
	.w1(32'h3c0bc574),
	.w2(32'h3bfadd67),
	.w3(32'h3c2752d0),
	.w4(32'h3c0cd923),
	.w5(32'h3b9d36a0),
	.w6(32'h3b007aef),
	.w7(32'h39ba3c0f),
	.w8(32'h39724799),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514d73),
	.w1(32'h3b5c9359),
	.w2(32'h39e26102),
	.w3(32'h3bf8c566),
	.w4(32'h3bdc8259),
	.w5(32'h3b3d6f61),
	.w6(32'hbb128c5c),
	.w7(32'h396d0672),
	.w8(32'hbb8a4600),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a0d58),
	.w1(32'hbb0cc867),
	.w2(32'h3bae5b74),
	.w3(32'hbb43668a),
	.w4(32'hbbd42e21),
	.w5(32'h3a89e899),
	.w6(32'hbb1d9dfe),
	.w7(32'hbbf22eb6),
	.w8(32'hbb409792),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6360db),
	.w1(32'hbcb5b3a1),
	.w2(32'hbc983940),
	.w3(32'hbaf5e9eb),
	.w4(32'hbc3f1a0d),
	.w5(32'h3b1a0291),
	.w6(32'hbbc3d54b),
	.w7(32'hbb82cc62),
	.w8(32'hbb0c32c7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45274),
	.w1(32'h3b961fd4),
	.w2(32'hbb6dfcb7),
	.w3(32'h3c01c9b8),
	.w4(32'h3bba7f86),
	.w5(32'hba3ef91b),
	.w6(32'h3a44b3b2),
	.w7(32'h3bf74b82),
	.w8(32'h3bb8c087),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccc013),
	.w1(32'hbad7b02a),
	.w2(32'hbb44ced6),
	.w3(32'h3c023998),
	.w4(32'hbbb91247),
	.w5(32'hbb9f3243),
	.w6(32'h3b8c8223),
	.w7(32'hbb89e18c),
	.w8(32'hbbb6965d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71649f),
	.w1(32'hbaaa9901),
	.w2(32'hbb0f4862),
	.w3(32'hbbf32863),
	.w4(32'hbada7028),
	.w5(32'hbb6f3772),
	.w6(32'hbc0cb9d8),
	.w7(32'hbb53adda),
	.w8(32'hb8f6dd4d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b904827),
	.w1(32'h3a91b346),
	.w2(32'hba942a96),
	.w3(32'h3be169d2),
	.w4(32'h3b5180b4),
	.w5(32'hbaa56179),
	.w6(32'h3b3e3e4b),
	.w7(32'h3b83353b),
	.w8(32'h3b341dd6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ab2ef),
	.w1(32'h3b77a0d4),
	.w2(32'hbb31bd92),
	.w3(32'h3aed0006),
	.w4(32'h3c4ffeff),
	.w5(32'h3aa95e13),
	.w6(32'h3b381aa3),
	.w7(32'h3c16c588),
	.w8(32'h3b971d29),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1acb1),
	.w1(32'h3b1e6d09),
	.w2(32'hbbcb0361),
	.w3(32'h3a6b133e),
	.w4(32'hbb7eaadb),
	.w5(32'hbbf607a9),
	.w6(32'h3b5798f3),
	.w7(32'hbbc689c2),
	.w8(32'hbbb1047c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf04125),
	.w1(32'h3b9951b6),
	.w2(32'h3939f33c),
	.w3(32'hbbc33460),
	.w4(32'h3b43dde4),
	.w5(32'h3b03b08b),
	.w6(32'hbbcdaec5),
	.w7(32'hb9db3d38),
	.w8(32'hbb1a9b56),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91b4d3),
	.w1(32'hb9b5d6dc),
	.w2(32'hbb1a9728),
	.w3(32'hb97821e0),
	.w4(32'h3aaacc13),
	.w5(32'h3b4748a2),
	.w6(32'hbb2c32e1),
	.w7(32'h3b10c3fd),
	.w8(32'hb9a64bf1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab820d7),
	.w1(32'hbc0119ae),
	.w2(32'hbbe79709),
	.w3(32'hbadb12ef),
	.w4(32'hbc247892),
	.w5(32'hbbfc323e),
	.w6(32'hb94d05a2),
	.w7(32'hbba17a68),
	.w8(32'hbbbf1e21),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99f7f6),
	.w1(32'hbb1fa554),
	.w2(32'hbb363cce),
	.w3(32'hbac4cdec),
	.w4(32'hbb536754),
	.w5(32'hbb8ba739),
	.w6(32'hbbbaf929),
	.w7(32'hbb794c03),
	.w8(32'hbb92d14b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae683da),
	.w1(32'h3b3c15ee),
	.w2(32'h3c14f586),
	.w3(32'h3a5133e6),
	.w4(32'h3b5ac663),
	.w5(32'h3c69b19d),
	.w6(32'hb8914a1f),
	.w7(32'h3be2d1cd),
	.w8(32'h3c1f423f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa3adf),
	.w1(32'hbad1486a),
	.w2(32'h3a8888d2),
	.w3(32'h3c45d6a9),
	.w4(32'h3b4e4ed9),
	.w5(32'h3aaacd8b),
	.w6(32'h3befce93),
	.w7(32'h3b815e80),
	.w8(32'h3a36cb0b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae597f0),
	.w1(32'hbb3962d6),
	.w2(32'hbb2f5236),
	.w3(32'hba4f604a),
	.w4(32'h3b9f06a5),
	.w5(32'h3b17cd2b),
	.w6(32'h3ae33c31),
	.w7(32'h3b887430),
	.w8(32'h3b6e1cec),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ffcaf),
	.w1(32'h3bb447ad),
	.w2(32'h3bc5d603),
	.w3(32'h3b7c869f),
	.w4(32'h3c0cf6bf),
	.w5(32'h3c4fde39),
	.w6(32'h3b346bd5),
	.w7(32'hba3c0230),
	.w8(32'h3a87eb40),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb572985),
	.w1(32'hba954466),
	.w2(32'hbbb155cc),
	.w3(32'h3af8d376),
	.w4(32'hbacdd42c),
	.w5(32'hbc2d7d37),
	.w6(32'hb90d14c2),
	.w7(32'hbb4d89d8),
	.w8(32'hbc1d7575),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43cb18),
	.w1(32'h3b9fe3ad),
	.w2(32'h3b834c78),
	.w3(32'hbb9f819d),
	.w4(32'h3bcf4aaa),
	.w5(32'h3ba6e965),
	.w6(32'hbb74c70d),
	.w7(32'h3ba7b93b),
	.w8(32'h3b452f03),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba340b3d),
	.w1(32'hbc0255f2),
	.w2(32'hbb76481b),
	.w3(32'h3aead0bf),
	.w4(32'hbb8bcbdd),
	.w5(32'h3a5d11d8),
	.w6(32'hba8024a1),
	.w7(32'h3b0b6b29),
	.w8(32'h3ab522f5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66f156),
	.w1(32'h3bcb061f),
	.w2(32'hbb8d2b25),
	.w3(32'h3c15ce8a),
	.w4(32'hbb188261),
	.w5(32'hbc1b53e8),
	.w6(32'h3bacc08f),
	.w7(32'hbc1f2f2c),
	.w8(32'hbc5f08f0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc506),
	.w1(32'h3a96d740),
	.w2(32'h39c1706b),
	.w3(32'hbbcf4325),
	.w4(32'hba869f1b),
	.w5(32'hbad669e0),
	.w6(32'hbbd1c82a),
	.w7(32'hba4426cc),
	.w8(32'hbafaf5de),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b8bc5),
	.w1(32'hbb33c38e),
	.w2(32'hbb37033a),
	.w3(32'hbacdd2e3),
	.w4(32'h398f1f93),
	.w5(32'h3a34efb7),
	.w6(32'hbb00ae29),
	.w7(32'hbad84620),
	.w8(32'hbae30d76),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6644b7),
	.w1(32'h3b3ba3c2),
	.w2(32'h3a301220),
	.w3(32'h3908217a),
	.w4(32'h3c0111a2),
	.w5(32'h3c74b34c),
	.w6(32'hba373c06),
	.w7(32'h3bfee6e2),
	.w8(32'h3c477517),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0884ee),
	.w1(32'h3a0aecce),
	.w2(32'h3b3e041a),
	.w3(32'h3c2bb5a2),
	.w4(32'h3b9228af),
	.w5(32'h3ba002d8),
	.w6(32'h3bb47e74),
	.w7(32'hba54b574),
	.w8(32'hba787b16),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29baad),
	.w1(32'h3c2e0c2b),
	.w2(32'h3b8d1ec7),
	.w3(32'h3b8a841a),
	.w4(32'h3ba98393),
	.w5(32'h3a8fbee3),
	.w6(32'hbb8b0ce3),
	.w7(32'hbaa0922b),
	.w8(32'hba7f9491),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98d790),
	.w1(32'hba9cc10a),
	.w2(32'h3a441505),
	.w3(32'hbb7e0906),
	.w4(32'hba2fc216),
	.w5(32'hba5a0137),
	.w6(32'hbb7e4ce1),
	.w7(32'h39f8dcc5),
	.w8(32'h3b093b84),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb747bf9),
	.w1(32'h3696ef74),
	.w2(32'h3a83425d),
	.w3(32'hbb96410f),
	.w4(32'h3b95e427),
	.w5(32'h3ba37955),
	.w6(32'hbb32e817),
	.w7(32'h3b8ee049),
	.w8(32'h3b35486f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e98d3),
	.w1(32'hbbe9291d),
	.w2(32'hbb99f620),
	.w3(32'h3b3227a7),
	.w4(32'h3adcf1c5),
	.w5(32'h3a9e7c71),
	.w6(32'h3a9f7295),
	.w7(32'hbba1e653),
	.w8(32'hbb70883a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9411dde),
	.w1(32'hbb77f8ee),
	.w2(32'h38b190a0),
	.w3(32'hba474fdb),
	.w4(32'hbabd0d69),
	.w5(32'h3bd53941),
	.w6(32'hbb203f4f),
	.w7(32'hbb12c8d8),
	.w8(32'h3ad5c44c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93de44),
	.w1(32'h39c98ebb),
	.w2(32'h3aa3e5aa),
	.w3(32'h3a961e24),
	.w4(32'h39d2f713),
	.w5(32'hb9f78df6),
	.w6(32'hb9ca2766),
	.w7(32'h3a0bccda),
	.w8(32'hba0b4514),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b5038),
	.w1(32'h398473a1),
	.w2(32'h3b9bac0d),
	.w3(32'h3a278cbd),
	.w4(32'hbaefaff3),
	.w5(32'h3a91eb7f),
	.w6(32'h3b0249c1),
	.w7(32'h386b1193),
	.w8(32'h3ad106fa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074806),
	.w1(32'hbc568565),
	.w2(32'hbbc76dcc),
	.w3(32'hbb6cab51),
	.w4(32'hbbca73aa),
	.w5(32'hbb5544cf),
	.w6(32'hbbd93f75),
	.w7(32'hbbd9d1e2),
	.w8(32'hbbb3bbec),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb4c1),
	.w1(32'h3ba16646),
	.w2(32'hbb4560a3),
	.w3(32'hbaf8c188),
	.w4(32'h3b51fac4),
	.w5(32'hba28a889),
	.w6(32'hbb5d03f7),
	.w7(32'hbb9bf7d7),
	.w8(32'hbb850178),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb627069),
	.w1(32'hbb32661f),
	.w2(32'hbaf8e99c),
	.w3(32'h3b10de0d),
	.w4(32'hbac31e45),
	.w5(32'hbb650590),
	.w6(32'hbb883927),
	.w7(32'hba8f333f),
	.w8(32'hbb2b0f7d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4288ba),
	.w1(32'hbbf8725e),
	.w2(32'h39bf66ec),
	.w3(32'h3b2a890d),
	.w4(32'hbb9d275e),
	.w5(32'h3b81fe7d),
	.w6(32'h3a0a1fd4),
	.w7(32'h39f25608),
	.w8(32'h391555d8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8a4d),
	.w1(32'h3c092fe9),
	.w2(32'h3bf2037e),
	.w3(32'hbb173446),
	.w4(32'hbb05b6c1),
	.w5(32'hbb555729),
	.w6(32'hbbadc096),
	.w7(32'hbc2174c8),
	.w8(32'hbc1f9332),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49cd23),
	.w1(32'h3c07b3fe),
	.w2(32'h3c1df70c),
	.w3(32'hbb5bf733),
	.w4(32'h3bddcc9b),
	.w5(32'h3c097b22),
	.w6(32'hbc08734c),
	.w7(32'h3bea43ff),
	.w8(32'h3bdd4b39),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aa3c6),
	.w1(32'hb8facad6),
	.w2(32'h3bdee26a),
	.w3(32'h3bd02eca),
	.w4(32'hba9acfc6),
	.w5(32'h3ca0ea4d),
	.w6(32'h3baba70d),
	.w7(32'h3b418463),
	.w8(32'h3c5e1ec6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31e843),
	.w1(32'hb9f6c57a),
	.w2(32'hbad3128b),
	.w3(32'h3cc1f12a),
	.w4(32'hbb378fb8),
	.w5(32'hbbd5c1cf),
	.w6(32'h3c8d16c5),
	.w7(32'hbbd13dfe),
	.w8(32'hbbde498f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c80b),
	.w1(32'hbb92a82e),
	.w2(32'hbbccd4d4),
	.w3(32'hbbc92b78),
	.w4(32'hb99fe573),
	.w5(32'hbb606d6b),
	.w6(32'hbba26820),
	.w7(32'hbb3b13c2),
	.w8(32'hbb9614d2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4f742),
	.w1(32'h3b070832),
	.w2(32'hbb4427c0),
	.w3(32'hbbe0a3f6),
	.w4(32'h3aa0d9f8),
	.w5(32'hbb1af073),
	.w6(32'hbbf92df6),
	.w7(32'h3b0fae94),
	.w8(32'hbae92528),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b1a35),
	.w1(32'h3b23a738),
	.w2(32'hba815c06),
	.w3(32'hbb65bed0),
	.w4(32'h3aa8d6ea),
	.w5(32'h3ab941bb),
	.w6(32'hbb191ca5),
	.w7(32'hb9f3d661),
	.w8(32'hbb4e0fb4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc073ff3),
	.w1(32'h3aca331e),
	.w2(32'hbac156e9),
	.w3(32'hba431c4c),
	.w4(32'hbaf25f62),
	.w5(32'hbc00391d),
	.w6(32'hba78fdd0),
	.w7(32'hbac38c02),
	.w8(32'hbb812863),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacd610),
	.w1(32'h3ba93591),
	.w2(32'hba8d82c9),
	.w3(32'hbb893ae6),
	.w4(32'hbac52576),
	.w5(32'hba3d3d65),
	.w6(32'hbba2aeba),
	.w7(32'hbbaeca5d),
	.w8(32'hbb4820bd),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a7bd5),
	.w1(32'h3aedec02),
	.w2(32'hbb103b48),
	.w3(32'h3b889909),
	.w4(32'h3bb25253),
	.w5(32'hbacd9e99),
	.w6(32'h3ac6e3cb),
	.w7(32'h3b8c2744),
	.w8(32'h3abae4ce),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3690f539),
	.w1(32'hbb2f22af),
	.w2(32'hbb69bb4e),
	.w3(32'hbb34488b),
	.w4(32'hbba84ced),
	.w5(32'hbbd897ce),
	.w6(32'h3a2e602f),
	.w7(32'hbbb5163b),
	.w8(32'hbbccdc32),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e1c9e),
	.w1(32'hbaa20d8f),
	.w2(32'h39231104),
	.w3(32'h3ac8f4d0),
	.w4(32'hba05af80),
	.w5(32'hbb679e14),
	.w6(32'hbb526878),
	.w7(32'hbb727128),
	.w8(32'hb9d7eeaa),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9728e4),
	.w1(32'hb89acd22),
	.w2(32'h3b72ffa5),
	.w3(32'h3bde8b3f),
	.w4(32'h39af86c8),
	.w5(32'h3afd4bb9),
	.w6(32'h3b9c8a61),
	.w7(32'hbaaaad7e),
	.w8(32'h399c9096),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a943e),
	.w1(32'hbbc781cf),
	.w2(32'hbbc36b32),
	.w3(32'hba36f11f),
	.w4(32'hba775468),
	.w5(32'h3a9e2232),
	.w6(32'hbb02992f),
	.w7(32'hbb0fd9d9),
	.w8(32'hb9646447),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35b767),
	.w1(32'h3ace8188),
	.w2(32'h3b986e6f),
	.w3(32'hba6c0a0c),
	.w4(32'hba207dd5),
	.w5(32'hbaa6ff7d),
	.w6(32'hbb07b795),
	.w7(32'hbb3d3034),
	.w8(32'hbb736048),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6d923),
	.w1(32'h3bef5f2a),
	.w2(32'hbaeb9bb4),
	.w3(32'h3ae869d4),
	.w4(32'h3b10d245),
	.w5(32'hbbbc6ee0),
	.w6(32'h3b868ed6),
	.w7(32'h3aa9689a),
	.w8(32'hbb5ced20),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdccae4),
	.w1(32'h3ac9f80e),
	.w2(32'hba010c66),
	.w3(32'h3b41c192),
	.w4(32'h3a883d41),
	.w5(32'hbae2d94c),
	.w6(32'h3b88cced),
	.w7(32'hbaf46645),
	.w8(32'hbb117b70),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1c6eb),
	.w1(32'h3abfdee6),
	.w2(32'h3a01b1ee),
	.w3(32'h3aba893d),
	.w4(32'h3b0c87a8),
	.w5(32'hbb2d2795),
	.w6(32'h3b262327),
	.w7(32'hbaa23001),
	.w8(32'hbb877514),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba543777),
	.w1(32'h3b8d2aeb),
	.w2(32'h3bf500cb),
	.w3(32'hbab4728a),
	.w4(32'h3b2d2200),
	.w5(32'h3b3fe845),
	.w6(32'hba98fd90),
	.w7(32'hba4fb29c),
	.w8(32'hb91924e4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c303d),
	.w1(32'h39f44691),
	.w2(32'hba447040),
	.w3(32'hba7a8742),
	.w4(32'hb9650a60),
	.w5(32'hba67d01d),
	.w6(32'hbab79df0),
	.w7(32'hba972e08),
	.w8(32'hba8ef897),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac99106),
	.w1(32'hbb4230a8),
	.w2(32'hbab04247),
	.w3(32'hbaa64d40),
	.w4(32'hbacd585a),
	.w5(32'h3b3c3214),
	.w6(32'hbb1fad44),
	.w7(32'h3a7fac5e),
	.w8(32'h3b029f49),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e46eb),
	.w1(32'hbb171294),
	.w2(32'hbb3c320b),
	.w3(32'h3b30d2cf),
	.w4(32'h3a9e62ed),
	.w5(32'hbb1b5274),
	.w6(32'h3b7678a3),
	.w7(32'hbab64443),
	.w8(32'hbb999822),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb473f1c),
	.w1(32'hbb697961),
	.w2(32'h3b9a6ee9),
	.w3(32'hbb31046b),
	.w4(32'hbb89ced6),
	.w5(32'hbb299580),
	.w6(32'hbbc06eb2),
	.w7(32'hbb8abb0d),
	.w8(32'hbba27ccb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f72eae),
	.w1(32'hbb09e8fe),
	.w2(32'h3933fad7),
	.w3(32'hba544d0b),
	.w4(32'h3a26300a),
	.w5(32'h3844459e),
	.w6(32'hbaa27734),
	.w7(32'hbb5e3417),
	.w8(32'hbb4dc2ee),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e1cee),
	.w1(32'h3b339f4f),
	.w2(32'h3abbd474),
	.w3(32'hbb4b5b69),
	.w4(32'hb94d1adb),
	.w5(32'hbb9e0265),
	.w6(32'hbb6905cc),
	.w7(32'hbbafc2df),
	.w8(32'hbc116614),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da1c68),
	.w1(32'hbbb518d7),
	.w2(32'hbb21dab8),
	.w3(32'hbb3f1566),
	.w4(32'hbbb5430f),
	.w5(32'hba5f9650),
	.w6(32'hbbb8027a),
	.w7(32'hbb259cdb),
	.w8(32'hbb3693be),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae95e3),
	.w1(32'hbae98061),
	.w2(32'hbb8444ae),
	.w3(32'hba186413),
	.w4(32'hbb51993d),
	.w5(32'hbc1e49cf),
	.w6(32'hbade4d86),
	.w7(32'hbb6aa719),
	.w8(32'hbbba1861),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f18f5),
	.w1(32'h39af4f78),
	.w2(32'h3a042f2e),
	.w3(32'hba939e64),
	.w4(32'h3b86486e),
	.w5(32'h3bc6f682),
	.w6(32'hba99d4ed),
	.w7(32'h3a99f8f4),
	.w8(32'hba038735),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1500),
	.w1(32'hba42129f),
	.w2(32'hbad4afd8),
	.w3(32'hba26814b),
	.w4(32'h3b0c8e3b),
	.w5(32'hbad7467d),
	.w6(32'hbb673227),
	.w7(32'h3b0b50af),
	.w8(32'h3a91b9ce),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b22af),
	.w1(32'h3afb6e9c),
	.w2(32'hbb65852f),
	.w3(32'hbb135090),
	.w4(32'hb7d9ca2e),
	.w5(32'hbb2dbc8a),
	.w6(32'hbb00a540),
	.w7(32'hbb17706c),
	.w8(32'hbb592669),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c673f),
	.w1(32'h3aa71ea7),
	.w2(32'h3b5e35ad),
	.w3(32'hbad720af),
	.w4(32'h3c1ff209),
	.w5(32'h3c7551d4),
	.w6(32'hbbc0b912),
	.w7(32'h3c10a5eb),
	.w8(32'h3bac2561),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a6a7d),
	.w1(32'h3b818182),
	.w2(32'h39fe3610),
	.w3(32'h3c62826d),
	.w4(32'h3bc4597e),
	.w5(32'h3b08af48),
	.w6(32'h3c56671b),
	.w7(32'hb93d4cef),
	.w8(32'hbaea7375),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aab9b),
	.w1(32'hba3f540a),
	.w2(32'hbad51545),
	.w3(32'hbaab14e1),
	.w4(32'h39187545),
	.w5(32'h3bbaf0bd),
	.w6(32'hbb142e8e),
	.w7(32'hbaee2ecd),
	.w8(32'h39f56820),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f80bf),
	.w1(32'h3b5ce9b0),
	.w2(32'h3a82b441),
	.w3(32'h3b9d613a),
	.w4(32'h3b9aee3e),
	.w5(32'hbb431242),
	.w6(32'h3b106cd5),
	.w7(32'h3b847af8),
	.w8(32'h38e34b46),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2b09e),
	.w1(32'hbb583f4e),
	.w2(32'hbb0fb0b5),
	.w3(32'hbb6f9153),
	.w4(32'hba89fbc8),
	.w5(32'hbb9ca625),
	.w6(32'hbb776c91),
	.w7(32'hba941641),
	.w8(32'hbafa0103),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4f40f),
	.w1(32'h3ac8435b),
	.w2(32'hbb5f7ee7),
	.w3(32'h3a6a6dc7),
	.w4(32'h3b3a4e36),
	.w5(32'hbb9acdd7),
	.w6(32'hba01173c),
	.w7(32'h3b86c868),
	.w8(32'hbb7a6097),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3dc6e),
	.w1(32'hbbd150ac),
	.w2(32'hbba9c4f9),
	.w3(32'hbbd9052b),
	.w4(32'hbbee2e42),
	.w5(32'hbb87b1f5),
	.w6(32'hbba5b9c2),
	.w7(32'hba9b2468),
	.w8(32'hb9c0c10e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c8f3f),
	.w1(32'hbbb1baa9),
	.w2(32'hbba425ce),
	.w3(32'hb9f77211),
	.w4(32'hbb71945c),
	.w5(32'hbb858513),
	.w6(32'hb9059667),
	.w7(32'hbb193296),
	.w8(32'hbba23652),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0545bc),
	.w1(32'hbb297e6f),
	.w2(32'h393ccb6b),
	.w3(32'hbc0a5539),
	.w4(32'hbbcef4fc),
	.w5(32'hbbf9104a),
	.w6(32'hbbff7a23),
	.w7(32'hbb4a7e01),
	.w8(32'hbb6d9db9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21c3ac),
	.w1(32'hbba3213b),
	.w2(32'hbb704a8c),
	.w3(32'hbb43dac8),
	.w4(32'hbbcbf5b3),
	.w5(32'hbbe243d9),
	.w6(32'h3a9609e7),
	.w7(32'hba2e0d8b),
	.w8(32'hbb40572f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8ea6f),
	.w1(32'hbabb2651),
	.w2(32'h3b8b3150),
	.w3(32'hbc3e94a9),
	.w4(32'hbabf590c),
	.w5(32'h3c0454bf),
	.w6(32'hbbe08af4),
	.w7(32'hba1a68dc),
	.w8(32'h3bcbbf72),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bcba2),
	.w1(32'h3ab0b550),
	.w2(32'hbb959fb8),
	.w3(32'h3b777f0c),
	.w4(32'hb9d840dd),
	.w5(32'hbb9dbc5b),
	.w6(32'h399d84f8),
	.w7(32'hbb542147),
	.w8(32'hbb7c32eb),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf3320),
	.w1(32'hbb3a05ee),
	.w2(32'h3851b6b3),
	.w3(32'hbb74ee12),
	.w4(32'hbac90b06),
	.w5(32'hba99218f),
	.w6(32'h373bf870),
	.w7(32'hbb942843),
	.w8(32'hbb82aa4d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49ff65),
	.w1(32'hbac5ca15),
	.w2(32'hbb66d4ce),
	.w3(32'h3a89d293),
	.w4(32'hbb2fd973),
	.w5(32'hbb68e587),
	.w6(32'hba6fdf2e),
	.w7(32'hbbbefd83),
	.w8(32'hbc036a82),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1429ba),
	.w1(32'hbacf576f),
	.w2(32'h3b3bd5fd),
	.w3(32'hba65722f),
	.w4(32'h3b45d046),
	.w5(32'h3c2737fc),
	.w6(32'hbb4683a1),
	.w7(32'h39e102aa),
	.w8(32'h3b9b6f41),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba906779),
	.w1(32'h3b0a3821),
	.w2(32'h3bcebda9),
	.w3(32'h3b5799b4),
	.w4(32'h3baa04e5),
	.w5(32'h3bc81ff9),
	.w6(32'hb81e131a),
	.w7(32'h3b34ffe3),
	.w8(32'hbb15e832),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c3526),
	.w1(32'hbc305026),
	.w2(32'hbb99d4a2),
	.w3(32'h3b8c8c3f),
	.w4(32'hbbdf4493),
	.w5(32'hbba62045),
	.w6(32'h3abd98c1),
	.w7(32'hbc1f5bab),
	.w8(32'hbbfe64b6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39eadf),
	.w1(32'hbb8091bc),
	.w2(32'hbb937b82),
	.w3(32'hba27b90f),
	.w4(32'hb9b7ff33),
	.w5(32'hbb8f1f88),
	.w6(32'hbaf08912),
	.w7(32'hba9c4440),
	.w8(32'hbba3de31),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef3e98),
	.w1(32'h3b518e0e),
	.w2(32'h39cd03f7),
	.w3(32'hbb44b200),
	.w4(32'h3c0f4f0f),
	.w5(32'h3c0bc9b3),
	.w6(32'hbabf6d01),
	.w7(32'h3a62946d),
	.w8(32'h39c5b28c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024847),
	.w1(32'hbc17af89),
	.w2(32'hbc13f125),
	.w3(32'hbb565d28),
	.w4(32'hbc3f63f2),
	.w5(32'hbbbecb7b),
	.w6(32'hbc05d992),
	.w7(32'hbb3a2420),
	.w8(32'hbae1f483),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7cba6),
	.w1(32'h3c6873e2),
	.w2(32'h3bd85bcf),
	.w3(32'h3b81a2aa),
	.w4(32'h3aef5103),
	.w5(32'hbbc18f80),
	.w6(32'h3b942586),
	.w7(32'h39e35f18),
	.w8(32'hb9ab7fe1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb199a2),
	.w1(32'hba784edb),
	.w2(32'hba67330a),
	.w3(32'h3bbbd11a),
	.w4(32'h3c088202),
	.w5(32'h3a5be76b),
	.w6(32'h3b90897e),
	.w7(32'h3b5fbb03),
	.w8(32'hb9d5c7a1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1a3f3),
	.w1(32'h3c02fc99),
	.w2(32'hba333f3e),
	.w3(32'hba952c12),
	.w4(32'h3c0a117d),
	.w5(32'h39d08882),
	.w6(32'hb96b2a42),
	.w7(32'h3b7e536f),
	.w8(32'hbb516314),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985a7c0),
	.w1(32'h3b505505),
	.w2(32'h3b9c3e5f),
	.w3(32'hbaf6c524),
	.w4(32'h3af3e980),
	.w5(32'h3bf60b9d),
	.w6(32'hbaa0748d),
	.w7(32'h3b3c5cbb),
	.w8(32'h3b97f468),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66f10f),
	.w1(32'h3bbef20f),
	.w2(32'h3b1eb6ec),
	.w3(32'h3b9c4ac0),
	.w4(32'h37faa66f),
	.w5(32'hbad985d3),
	.w6(32'h3b307e57),
	.w7(32'h3a872799),
	.w8(32'hba1da0cf),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0efbc7),
	.w1(32'h3a82693c),
	.w2(32'h39b693d8),
	.w3(32'h3bc37aa0),
	.w4(32'h3bb88f96),
	.w5(32'h38e98c85),
	.w6(32'h3b6ca802),
	.w7(32'h3b1fb02c),
	.w8(32'hba7b4637),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8be0f4),
	.w1(32'hbb77ff68),
	.w2(32'hb8956fa3),
	.w3(32'hbb9ad895),
	.w4(32'hb99c2de8),
	.w5(32'h3b56a466),
	.w6(32'hbb81d3d4),
	.w7(32'hbb91f5fb),
	.w8(32'hbb4def88),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd1e87),
	.w1(32'hbbc425ab),
	.w2(32'hb9ac8044),
	.w3(32'h3bc6eee0),
	.w4(32'hba3c0583),
	.w5(32'h3b374aef),
	.w6(32'hbb3cae74),
	.w7(32'hbabad9fa),
	.w8(32'h3b866017),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb697c8c),
	.w1(32'h3b9cb578),
	.w2(32'h39a9fac2),
	.w3(32'hb85ffab1),
	.w4(32'h3c0b158a),
	.w5(32'hba26b7f2),
	.w6(32'hba230d39),
	.w7(32'h3b7e7e29),
	.w8(32'h3a88b0ca),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7033bf),
	.w1(32'h3a56e5db),
	.w2(32'hb9b124c5),
	.w3(32'hbb9353d6),
	.w4(32'h38b1d7f2),
	.w5(32'hbb33caa2),
	.w6(32'hbbf5cb41),
	.w7(32'hba5bdb92),
	.w8(32'hbb13cffc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97c2e1),
	.w1(32'hba701560),
	.w2(32'hbb897f99),
	.w3(32'h3a97667d),
	.w4(32'hbadb1953),
	.w5(32'hbb91be86),
	.w6(32'hba04d000),
	.w7(32'hbb1349d8),
	.w8(32'hbb2cd43f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3718bc44),
	.w1(32'h33bb11a2),
	.w2(32'h3817b367),
	.w3(32'h370f38da),
	.w4(32'hb5fdd8bd),
	.w5(32'h380bd9f5),
	.w6(32'h37f33d6b),
	.w7(32'h375d384a),
	.w8(32'h38209be0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb370d1c),
	.w1(32'hbba76117),
	.w2(32'hbb4adc63),
	.w3(32'hba8b1c0f),
	.w4(32'hbb304df1),
	.w5(32'hbaddb5b6),
	.w6(32'h3a9c2054),
	.w7(32'h3a2bdbe7),
	.w8(32'hbb2797a5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376d4b9b),
	.w1(32'h375531db),
	.w2(32'h3870259b),
	.w3(32'h380535f3),
	.w4(32'hb7984e72),
	.w5(32'h38269f2c),
	.w6(32'h38a80fec),
	.w7(32'h3605ada3),
	.w8(32'h388b4e87),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6fa46),
	.w1(32'hba712a62),
	.w2(32'h388bc31b),
	.w3(32'hbacf1680),
	.w4(32'hb7985a64),
	.w5(32'h3a35ea5d),
	.w6(32'hbb3507fc),
	.w7(32'hb9ba10ad),
	.w8(32'hba70c49f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bbf8b),
	.w1(32'h3b98dc13),
	.w2(32'hba3dd4e1),
	.w3(32'h3a17e6c4),
	.w4(32'h3a12554e),
	.w5(32'hbb01ed90),
	.w6(32'hbadb9825),
	.w7(32'hbb8b421f),
	.w8(32'hbb9dcbdf),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378dc353),
	.w1(32'h3b197492),
	.w2(32'hba7089d1),
	.w3(32'h3ab33ee9),
	.w4(32'h3ab1fcf0),
	.w5(32'hbb14877d),
	.w6(32'h3a1a10fe),
	.w7(32'hb9d9905b),
	.w8(32'hbb208360),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39954b27),
	.w1(32'h3973d3c6),
	.w2(32'hba1aca61),
	.w3(32'hb90823b7),
	.w4(32'hba0a6cc3),
	.w5(32'hba589834),
	.w6(32'hb98abd1f),
	.w7(32'hba162b90),
	.w8(32'hba40dd2f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80e4fe),
	.w1(32'h3b9a43c7),
	.w2(32'hbb3c273b),
	.w3(32'h3b819c3e),
	.w4(32'h3a4c69e6),
	.w5(32'hbb8d7249),
	.w6(32'h3b60b1cf),
	.w7(32'hba690b73),
	.w8(32'hbb453ff1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f221f5),
	.w1(32'hb98dc632),
	.w2(32'h3abf8093),
	.w3(32'hb8f22029),
	.w4(32'hb9c7b28b),
	.w5(32'h3a055605),
	.w6(32'hba2eb5d7),
	.w7(32'h39186374),
	.w8(32'h39e3764a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac96f7),
	.w1(32'h3aa5f51d),
	.w2(32'hbadd6a89),
	.w3(32'h3b4cd904),
	.w4(32'hbac18376),
	.w5(32'hbba7b265),
	.w6(32'h3a06295d),
	.w7(32'hbb1549e3),
	.w8(32'hbb88c079),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb831b775),
	.w1(32'h361263f9),
	.w2(32'h37671a4d),
	.w3(32'h36653680),
	.w4(32'h38764e90),
	.w5(32'h37cd7632),
	.w6(32'h37fb3591),
	.w7(32'h380c9859),
	.w8(32'hb50bbfbe),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c79c46),
	.w1(32'h3817c737),
	.w2(32'h38ae6a28),
	.w3(32'h38cd8eb3),
	.w4(32'hb826c512),
	.w5(32'h360b2d1a),
	.w6(32'h399120f1),
	.w7(32'h3825981d),
	.w8(32'h362fb973),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94e9eb),
	.w1(32'h3b39f366),
	.w2(32'hbb04c178),
	.w3(32'h3b465ece),
	.w4(32'hb9d9c8d4),
	.w5(32'hbb1c05bc),
	.w6(32'hba84f893),
	.w7(32'h3a81ab19),
	.w8(32'hbb042f6c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf1b57),
	.w1(32'hbba063e2),
	.w2(32'hbb827929),
	.w3(32'hbaf3a88b),
	.w4(32'h3afb8d96),
	.w5(32'hbb0a374c),
	.w6(32'hbb6a7c83),
	.w7(32'h3a58f39a),
	.w8(32'hbb8614b2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb889e961),
	.w1(32'h3adb14f5),
	.w2(32'h3b35f5cb),
	.w3(32'h3b162a0c),
	.w4(32'h3a5011d1),
	.w5(32'hbafebd89),
	.w6(32'hb9a7a501),
	.w7(32'hbb3a5c83),
	.w8(32'hbb832ba9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a26bf),
	.w1(32'hb8f62b48),
	.w2(32'h3b6707ab),
	.w3(32'h3c01e8cd),
	.w4(32'h3b25e56a),
	.w5(32'h3a949e55),
	.w6(32'h3ae4c761),
	.w7(32'h3a1d67eb),
	.w8(32'h3a3ccfb4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d89a3),
	.w1(32'h3a224927),
	.w2(32'hb7d5f4ee),
	.w3(32'h39438867),
	.w4(32'h39bd65bd),
	.w5(32'hba17514e),
	.w6(32'hb9845f42),
	.w7(32'hb9b1128c),
	.w8(32'hb96d5974),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397844e9),
	.w1(32'hba642a8f),
	.w2(32'hb964c2db),
	.w3(32'h37179ade),
	.w4(32'hb9a976ed),
	.w5(32'h391e53bc),
	.w6(32'h3a7b59e2),
	.w7(32'h38b3ca50),
	.w8(32'hb9f97a21),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd4986),
	.w1(32'hba302fae),
	.w2(32'h39343a76),
	.w3(32'h3b675778),
	.w4(32'hbb126d0c),
	.w5(32'h3b94de5f),
	.w6(32'hbbf34710),
	.w7(32'hbaefbc52),
	.w8(32'h3afcdf7a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ea135),
	.w1(32'hbbe6c9b2),
	.w2(32'hbb7f851d),
	.w3(32'hbb99f9b9),
	.w4(32'hbb9c764f),
	.w5(32'hbb1e7eeb),
	.w6(32'hbbab2b2d),
	.w7(32'hba69f7f7),
	.w8(32'h3988f2d0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac84cb2),
	.w1(32'hbbd00edf),
	.w2(32'hbb31b318),
	.w3(32'hbafd3912),
	.w4(32'hbbff7811),
	.w5(32'h3aa1e973),
	.w6(32'hbc197f9d),
	.w7(32'hbacd6add),
	.w8(32'h3b68eb1e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba491f4a),
	.w1(32'h3b377856),
	.w2(32'hbab564b0),
	.w3(32'h3a50cc28),
	.w4(32'h39ba9d56),
	.w5(32'hbb2a1772),
	.w6(32'hb8bfadc4),
	.w7(32'hbb414ad7),
	.w8(32'hbb906ff2),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b2b1f),
	.w1(32'h3ba97bc2),
	.w2(32'hba5a148b),
	.w3(32'h3b18f943),
	.w4(32'h3b050050),
	.w5(32'hbb28eb9e),
	.w6(32'h3abca242),
	.w7(32'hbb1e78f3),
	.w8(32'hbb99ca8b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f0c572),
	.w1(32'h37052942),
	.w2(32'h370b5980),
	.w3(32'h37639c94),
	.w4(32'h36300df9),
	.w5(32'h3718dd63),
	.w6(32'h37523659),
	.w7(32'h3606cfc6),
	.w8(32'h3788a934),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37817864),
	.w1(32'h3628eb12),
	.w2(32'h3726a8ca),
	.w3(32'h375b1a96),
	.w4(32'hb6e3fa23),
	.w5(32'h37291a2f),
	.w6(32'h379b4c79),
	.w7(32'h368e27c9),
	.w8(32'h376961c8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1779a),
	.w1(32'h3ade7e66),
	.w2(32'h3a674daa),
	.w3(32'hb6310997),
	.w4(32'h3a8a2afd),
	.w5(32'h3953fad6),
	.w6(32'h38bba7ae),
	.w7(32'h39ea6f9e),
	.w8(32'h3a49aad5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372de4b3),
	.w1(32'hb69c334c),
	.w2(32'h378dc2b2),
	.w3(32'h37ef8ed1),
	.w4(32'h37b0c9eb),
	.w5(32'h37bc1ff6),
	.w6(32'h38321c5a),
	.w7(32'h37a22d60),
	.w8(32'h37fa794d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b593aae),
	.w1(32'h3a91547a),
	.w2(32'hbb1a4831),
	.w3(32'h3b1ab963),
	.w4(32'h3ab733bf),
	.w5(32'hba246878),
	.w6(32'h3a802f94),
	.w7(32'h3adf98be),
	.w8(32'h39cb55c4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae438d1),
	.w1(32'h3a6557f3),
	.w2(32'h38cd0506),
	.w3(32'h3a422a88),
	.w4(32'h39c57823),
	.w5(32'hbb04ac18),
	.w6(32'hbabf701b),
	.w7(32'h398eb502),
	.w8(32'hbb160d1a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d9cfc),
	.w1(32'h3abc3509),
	.w2(32'hbb01672a),
	.w3(32'h3b33682a),
	.w4(32'h3a80cc19),
	.w5(32'hbafeb878),
	.w6(32'h3a2a4fb6),
	.w7(32'hb97aded8),
	.w8(32'hbb513d2b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fbbebc),
	.w1(32'h38318c6d),
	.w2(32'h384d7c8c),
	.w3(32'h380e6a48),
	.w4(32'h3703ede1),
	.w5(32'h3828e24d),
	.w6(32'h37f372a2),
	.w7(32'h35e5f6ae),
	.w8(32'h37e981a3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a590a2a),
	.w1(32'hbc26f220),
	.w2(32'hbbdcd542),
	.w3(32'hbae8c296),
	.w4(32'hbc07277e),
	.w5(32'hba621e72),
	.w6(32'hbbff6a0f),
	.w7(32'hbaf49864),
	.w8(32'h3a70c345),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77d996),
	.w1(32'hbb283b1a),
	.w2(32'hb8f9bc25),
	.w3(32'hbaaa2823),
	.w4(32'hbb10f16c),
	.w5(32'hb8e410ae),
	.w6(32'hbb032b77),
	.w7(32'hba8ece18),
	.w8(32'h39da04c0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7936b1e),
	.w1(32'hb8b23a26),
	.w2(32'hb81063f0),
	.w3(32'h38150850),
	.w4(32'hb88ca7ba),
	.w5(32'hb8859e07),
	.w6(32'h381317ac),
	.w7(32'hb876a6ed),
	.w8(32'hb694b63b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058095),
	.w1(32'hbb56f6b4),
	.w2(32'hb9b4b576),
	.w3(32'hbaf6626e),
	.w4(32'hbac49412),
	.w5(32'h3a1b1610),
	.w6(32'hbb4cc966),
	.w7(32'hb9c6e3cd),
	.w8(32'h3a8ef26d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38abf6b1),
	.w1(32'h373a04c8),
	.w2(32'h3682cdc6),
	.w3(32'h380c2838),
	.w4(32'hb884ad4f),
	.w5(32'hb8457bcb),
	.w6(32'h381444d6),
	.w7(32'hb7f86b20),
	.w8(32'h37ac3d47),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919f422),
	.w1(32'h39781f64),
	.w2(32'h38df6497),
	.w3(32'h395a1f99),
	.w4(32'h3886dd12),
	.w5(32'hb8003235),
	.w6(32'h38c62924),
	.w7(32'hb9281c5c),
	.w8(32'hb8b53f7a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb727284f),
	.w1(32'h3630c6cb),
	.w2(32'h37175677),
	.w3(32'hb7537d06),
	.w4(32'h37b06943),
	.w5(32'h384d0181),
	.w6(32'h3824e432),
	.w7(32'h3819f54c),
	.w8(32'h37bb2b7e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65c3aaa),
	.w1(32'hb717b124),
	.w2(32'h36aa5bed),
	.w3(32'h37aa0895),
	.w4(32'h37e5a2a9),
	.w5(32'h3668630d),
	.w6(32'h381c6169),
	.w7(32'h38071623),
	.w8(32'h3704cafc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b90b1),
	.w1(32'h3a5e210f),
	.w2(32'hbafe0f87),
	.w3(32'h3a966090),
	.w4(32'h3ac1295d),
	.w5(32'hba4783fe),
	.w6(32'hb916621c),
	.w7(32'h391111e9),
	.w8(32'hba2e0edd),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a446e),
	.w1(32'hb9684d94),
	.w2(32'h3b5e1a88),
	.w3(32'h3a5ef5b7),
	.w4(32'hbae37f80),
	.w5(32'hbaff6aa1),
	.w6(32'hbb122421),
	.w7(32'h39c72d7a),
	.w8(32'hba4e4f99),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0c655),
	.w1(32'hbb42aeba),
	.w2(32'hb9f9500c),
	.w3(32'hbaaa3884),
	.w4(32'hbac1ac95),
	.w5(32'hb9ad202f),
	.w6(32'hbaebe1d4),
	.w7(32'h38843cfb),
	.w8(32'h3a7dde1f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4515d4),
	.w1(32'hbab2dd15),
	.w2(32'h3aa6e419),
	.w3(32'hba1977c2),
	.w4(32'hbae7a527),
	.w5(32'hba86670b),
	.w6(32'hbb25497f),
	.w7(32'hba0bc533),
	.w8(32'h3a07cdda),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dde2c0),
	.w1(32'h390324cf),
	.w2(32'h384949e6),
	.w3(32'h38d38e28),
	.w4(32'h391051ce),
	.w5(32'h38a536ae),
	.w6(32'h38307d58),
	.w7(32'h38ae600f),
	.w8(32'h3835fa4f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcf629),
	.w1(32'hb90dfc6b),
	.w2(32'h387b87e3),
	.w3(32'hb79bc253),
	.w4(32'hba0aca40),
	.w5(32'hb9b7cf69),
	.w6(32'h383b98d9),
	.w7(32'hb8668a20),
	.w8(32'hb9896755),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3847efca),
	.w1(32'h3832a51a),
	.w2(32'h383fd05a),
	.w3(32'h36bec02b),
	.w4(32'h37e10153),
	.w5(32'h3827a15e),
	.w6(32'hb6e1f13e),
	.w7(32'h381a4183),
	.w8(32'h384c1708),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37005bf7),
	.w1(32'hb775ea44),
	.w2(32'hb7e0468b),
	.w3(32'h3800039e),
	.w4(32'h371c8b3c),
	.w5(32'h3794f5a8),
	.w6(32'h38000ce9),
	.w7(32'h372035a2),
	.w8(32'hb64790b2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43af57),
	.w1(32'hbb42aa35),
	.w2(32'hbaa691b7),
	.w3(32'hbb3c9f0a),
	.w4(32'hbb5adb20),
	.w5(32'hbb40b5c0),
	.w6(32'hbae60f8a),
	.w7(32'hba3a3b6b),
	.w8(32'hbb1d3a7c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b5001a),
	.w1(32'hb800fa55),
	.w2(32'hb8c0156b),
	.w3(32'h3848dba1),
	.w4(32'hb7cb29ee),
	.w5(32'hb8e1084c),
	.w6(32'h38f3c428),
	.w7(32'h38148958),
	.w8(32'hb8df372a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a35276),
	.w1(32'h39203e94),
	.w2(32'hb78eea66),
	.w3(32'h38d9fee2),
	.w4(32'hb91308a0),
	.w5(32'hb8cab5e8),
	.w6(32'hb95b3c03),
	.w7(32'hb97fb48f),
	.w8(32'hb919504c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2a4bf),
	.w1(32'hbae7d380),
	.w2(32'hbaabed23),
	.w3(32'hbae002a2),
	.w4(32'hbabfe5f1),
	.w5(32'hba9c1c34),
	.w6(32'h3a0bff83),
	.w7(32'hb8e9b3d7),
	.w8(32'hb993a7b7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f5f93),
	.w1(32'h36a153f5),
	.w2(32'hb7bf9b5a),
	.w3(32'h385127d8),
	.w4(32'hb6d0a2ce),
	.w5(32'hb7b31c1f),
	.w6(32'h3863d98e),
	.w7(32'hb761f6d0),
	.w8(32'hb82a886e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394e60fa),
	.w1(32'h395cb055),
	.w2(32'hbaa969ff),
	.w3(32'h3a7b4ab6),
	.w4(32'h398f74cb),
	.w5(32'hbabee3d6),
	.w6(32'h3985ad95),
	.w7(32'hb9e7d4c3),
	.w8(32'hba99c81d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39baf71f),
	.w1(32'hb95a9bfc),
	.w2(32'hb9620fd7),
	.w3(32'h3a05bbf6),
	.w4(32'hb97bc3da),
	.w5(32'hb9f7e0b7),
	.w6(32'h39968c29),
	.w7(32'hb919c4f3),
	.w8(32'hb9ef0916),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1caefe),
	.w1(32'hbb8b3315),
	.w2(32'h3b0e378a),
	.w3(32'hbbd1c0cb),
	.w4(32'hbb82e9b1),
	.w5(32'hbb487811),
	.w6(32'hbbae057d),
	.w7(32'h3838f595),
	.w8(32'h3ab77cbe),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395aa830),
	.w1(32'h3802fba8),
	.w2(32'hb93c70e4),
	.w3(32'h387e2275),
	.w4(32'hb918c5eb),
	.w5(32'hb990de7a),
	.w6(32'h37dc0755),
	.w7(32'h3826d000),
	.w8(32'hb832f259),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13b6a4),
	.w1(32'hb8ea3a56),
	.w2(32'hbb2e5179),
	.w3(32'hbaa9472b),
	.w4(32'h3ae1dc9a),
	.w5(32'h3a01bf42),
	.w6(32'hbb121350),
	.w7(32'h398315b5),
	.w8(32'hbbb78523),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule