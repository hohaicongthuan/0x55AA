module layer_10_featuremap_363(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39104365),
	.w1(32'h39b58aa4),
	.w2(32'h3a41020c),
	.w3(32'h388bd0f4),
	.w4(32'h39bc87bf),
	.w5(32'hbaa7478c),
	.w6(32'h39845e49),
	.w7(32'h39f9722e),
	.w8(32'hbabcec4a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a5997),
	.w1(32'hba4db15a),
	.w2(32'hb8027580),
	.w3(32'hba40f396),
	.w4(32'hba8119e8),
	.w5(32'h39ae2d4a),
	.w6(32'hba6befd4),
	.w7(32'hba509587),
	.w8(32'hba16fed0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a075033),
	.w1(32'h39ed4f56),
	.w2(32'h3a56076b),
	.w3(32'hb8f8dd76),
	.w4(32'h379602a9),
	.w5(32'h38b5e432),
	.w6(32'hba727676),
	.w7(32'hb789f31f),
	.w8(32'hb8fcb1f0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abf77c),
	.w1(32'hb919f7ee),
	.w2(32'hb9996b70),
	.w3(32'h392e57bc),
	.w4(32'hb904e06d),
	.w5(32'hba950347),
	.w6(32'hba23dc07),
	.w7(32'hb9759387),
	.w8(32'hbac344ee),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c49ebc),
	.w1(32'hb9a0a193),
	.w2(32'h3a39807f),
	.w3(32'hbab200ff),
	.w4(32'h39e79a0a),
	.w5(32'h39e64fe0),
	.w6(32'hbaa895aa),
	.w7(32'hb897d148),
	.w8(32'h397d36c4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35b2c8),
	.w1(32'h3a0873c1),
	.w2(32'h3a567ab7),
	.w3(32'h39b7789b),
	.w4(32'h39d8d48c),
	.w5(32'hb8f16dd3),
	.w6(32'h39d3261d),
	.w7(32'h3a31f259),
	.w8(32'h3902c7ff),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f110e),
	.w1(32'hb9bfdbb0),
	.w2(32'h38b3971e),
	.w3(32'hb915bab3),
	.w4(32'h39793a33),
	.w5(32'h3908235a),
	.w6(32'hb723df28),
	.w7(32'h3903673a),
	.w8(32'hba432773),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28636f),
	.w1(32'hb8fbcdb1),
	.w2(32'hb95a3b0a),
	.w3(32'hba274441),
	.w4(32'hbab488e2),
	.w5(32'h3a684064),
	.w6(32'hbac1d9a7),
	.w7(32'hbad98e2c),
	.w8(32'h3a33bbea),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04b490),
	.w1(32'h3a5661ea),
	.w2(32'h3a3e0880),
	.w3(32'h3a8c9088),
	.w4(32'h3a70ab3d),
	.w5(32'h3a236028),
	.w6(32'h3a93a08f),
	.w7(32'h3a8b16e3),
	.w8(32'h39eb4734),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52449d),
	.w1(32'h39c1fe32),
	.w2(32'h3a502145),
	.w3(32'h395587fa),
	.w4(32'h39cd9bf6),
	.w5(32'h39f7c2ed),
	.w6(32'h3968aae1),
	.w7(32'h3a3fd0c7),
	.w8(32'h3a0c02a3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a766d55),
	.w1(32'h3a4ee08d),
	.w2(32'h3a54a1de),
	.w3(32'h39c4404b),
	.w4(32'h39bbdb8a),
	.w5(32'hba15e66f),
	.w6(32'h3a01942c),
	.w7(32'h3a0c0c15),
	.w8(32'hba1dde83),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38348155),
	.w1(32'h389d1f97),
	.w2(32'hb9c64c03),
	.w3(32'hba335fa8),
	.w4(32'hba185d0b),
	.w5(32'hbacd3fa4),
	.w6(32'hb9c20352),
	.w7(32'h3808a5cd),
	.w8(32'hbac8f2c1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada99a9),
	.w1(32'hbac09976),
	.w2(32'hbaa842e0),
	.w3(32'hbab2e81a),
	.w4(32'hba3be900),
	.w5(32'hb9f08ba5),
	.w6(32'hba0ce135),
	.w7(32'hb9d93255),
	.w8(32'hba08a78e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2a4f4),
	.w1(32'hb771cd7c),
	.w2(32'hb9eb4682),
	.w3(32'hbaa8a1c7),
	.w4(32'hb9fd72c7),
	.w5(32'h39aa789b),
	.w6(32'hba67cf54),
	.w7(32'hba502f89),
	.w8(32'h390b1db4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39984de0),
	.w1(32'h3908a46d),
	.w2(32'hb83c32a3),
	.w3(32'h3a0f16bb),
	.w4(32'h39bc5721),
	.w5(32'hb9cb78e9),
	.w6(32'h39b18e1c),
	.w7(32'h38b7b6d2),
	.w8(32'hba12e3cf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f7f90),
	.w1(32'hb9d5d547),
	.w2(32'h39b54a05),
	.w3(32'hb9e54299),
	.w4(32'h39dfa53b),
	.w5(32'h3904c046),
	.w6(32'h398ed8e3),
	.w7(32'h3a32064f),
	.w8(32'h3a0dfe48),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6da73),
	.w1(32'h3a0be393),
	.w2(32'h3a5db1c8),
	.w3(32'h39ace6b9),
	.w4(32'h3a310168),
	.w5(32'hba23ebc9),
	.w6(32'h3a2be69d),
	.w7(32'h3a291332),
	.w8(32'hb9f335e8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e1667),
	.w1(32'h37071a35),
	.w2(32'h3933fd05),
	.w3(32'h3884af72),
	.w4(32'h395b83dd),
	.w5(32'hba5cc44b),
	.w6(32'h38930ca5),
	.w7(32'h39997908),
	.w8(32'h39e5af9f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b85f07),
	.w1(32'hb7929486),
	.w2(32'h39c05f80),
	.w3(32'hb92b460e),
	.w4(32'h3a396f87),
	.w5(32'hba26af4e),
	.w6(32'h3a2e475a),
	.w7(32'h391c17df),
	.w8(32'hb9c993c5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8556d),
	.w1(32'hba4281f8),
	.w2(32'hba95352f),
	.w3(32'hba1f2d8b),
	.w4(32'hb98db6ef),
	.w5(32'h39f48342),
	.w6(32'hb99c9b20),
	.w7(32'hb9a82e49),
	.w8(32'hb8c9b236),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a716d64),
	.w1(32'hb9a61206),
	.w2(32'h3a0ffccf),
	.w3(32'hb9aecfc2),
	.w4(32'h3a213250),
	.w5(32'h3a8d0966),
	.w6(32'hb97d5ef8),
	.w7(32'h3a493e93),
	.w8(32'h3aa3d564),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf656a),
	.w1(32'h3aaa235a),
	.w2(32'h3ad265e6),
	.w3(32'h3a81cc2c),
	.w4(32'h3a85f3b1),
	.w5(32'hba43bbaf),
	.w6(32'h3a9e0fdb),
	.w7(32'h3ad6ed59),
	.w8(32'hba84235a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba071a8d),
	.w1(32'hb99398bc),
	.w2(32'hb9bed515),
	.w3(32'hb9c7515b),
	.w4(32'hba184ed2),
	.w5(32'hba709863),
	.w6(32'hba39d407),
	.w7(32'hb9f81a05),
	.w8(32'hbac2ed93),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d06a2),
	.w1(32'hba54d0cc),
	.w2(32'hba36a0e9),
	.w3(32'hbab704ee),
	.w4(32'hba242953),
	.w5(32'hba7ac7ff),
	.w6(32'hba9062b8),
	.w7(32'hba7fd099),
	.w8(32'hbaee0aa9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceb000),
	.w1(32'hbaa4fd7f),
	.w2(32'hba42c8e2),
	.w3(32'hba80d00a),
	.w4(32'hbaa10bbe),
	.w5(32'h3a86cf2d),
	.w6(32'hba34ac3b),
	.w7(32'hbad91b1d),
	.w8(32'h3aed4a22),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5aa46d),
	.w1(32'h39e09fbe),
	.w2(32'h396891b3),
	.w3(32'h3a92bd02),
	.w4(32'h3a6e2b16),
	.w5(32'hba2c4aa8),
	.w6(32'h3ac507f4),
	.w7(32'h3a725bf4),
	.w8(32'hb930a369),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7ed6c),
	.w1(32'h3929df97),
	.w2(32'hba0ac77e),
	.w3(32'hb84ffe1c),
	.w4(32'hba1a9618),
	.w5(32'h3aa2f421),
	.w6(32'hb8519e04),
	.w7(32'hba075550),
	.w8(32'h3a595330),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a576791),
	.w1(32'h3a2bdbc3),
	.w2(32'h3a936fec),
	.w3(32'h3993937b),
	.w4(32'h3a8a5b79),
	.w5(32'hbaf2f533),
	.w6(32'h3a58e8ab),
	.w7(32'h3ad2cea5),
	.w8(32'hba165cfc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e573c),
	.w1(32'hba98151f),
	.w2(32'hba224157),
	.w3(32'hbb0475f6),
	.w4(32'hba262b33),
	.w5(32'hba2d6368),
	.w6(32'hba55a5e6),
	.w7(32'hba2f8f27),
	.w8(32'hb953c8a5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4a1a8),
	.w1(32'hb947e42c),
	.w2(32'h38df63db),
	.w3(32'hba0cec7a),
	.w4(32'hb8d9dc1c),
	.w5(32'hb9e7acea),
	.w6(32'hb988bec0),
	.w7(32'h389d2a69),
	.w8(32'hbae491a9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72287c),
	.w1(32'hba9a1fdf),
	.w2(32'hbacabee7),
	.w3(32'hba7fd0b7),
	.w4(32'hba3b6f9a),
	.w5(32'hb9c6938b),
	.w6(32'hb9f86578),
	.w7(32'hbae7bf94),
	.w8(32'hba1e381d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6bae9),
	.w1(32'hb96e4d85),
	.w2(32'hb7354005),
	.w3(32'h38da8c62),
	.w4(32'hb93238ee),
	.w5(32'hb910ee65),
	.w6(32'hb8da1e59),
	.w7(32'h39f77fbe),
	.w8(32'hb68310db),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec1bd9),
	.w1(32'hba7dc7ea),
	.w2(32'hba4f6589),
	.w3(32'h39d694d7),
	.w4(32'h3986dcdc),
	.w5(32'hba737e30),
	.w6(32'hb9f2305e),
	.w7(32'hb971b4d3),
	.w8(32'hbaa220a2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aef67),
	.w1(32'hb9e1f775),
	.w2(32'h393a6f28),
	.w3(32'hb9b1e5fc),
	.w4(32'hba0cd74c),
	.w5(32'hba8082e1),
	.w6(32'hb97af164),
	.w7(32'hba06d613),
	.w8(32'hba9b0a88),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a683c),
	.w1(32'hba92c440),
	.w2(32'hba7a413d),
	.w3(32'hba01831d),
	.w4(32'hb9b3656b),
	.w5(32'h3a0b38de),
	.w6(32'hb9552319),
	.w7(32'hba894c35),
	.w8(32'hba5fd461),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7dc98),
	.w1(32'hba042cf2),
	.w2(32'h37c3600f),
	.w3(32'hb989d1ab),
	.w4(32'h3a05d517),
	.w5(32'hba364a5c),
	.w6(32'hba362394),
	.w7(32'hba34ace7),
	.w8(32'h3a64272b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4efcd),
	.w1(32'h39b86ff6),
	.w2(32'h396b1e43),
	.w3(32'hba6f525e),
	.w4(32'hba4b54b2),
	.w5(32'h3a29f6ec),
	.w6(32'h3b36a6a6),
	.w7(32'h39f63919),
	.w8(32'h3a26df59),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a332407),
	.w1(32'h3a18105a),
	.w2(32'h3a242c96),
	.w3(32'h39f36109),
	.w4(32'hb7b4453c),
	.w5(32'hba5a545b),
	.w6(32'h39f87550),
	.w7(32'hb97c8463),
	.w8(32'hbab88e41),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab69b46),
	.w1(32'hbab7221a),
	.w2(32'hba68a37e),
	.w3(32'hba09e1bd),
	.w4(32'hba28de27),
	.w5(32'h3a8ddefb),
	.w6(32'hba5b0ea1),
	.w7(32'hbaac87ae),
	.w8(32'h3a39c1ae),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ecfe4),
	.w1(32'h3a03d87f),
	.w2(32'h3a752f44),
	.w3(32'h3a737190),
	.w4(32'h3b0b164f),
	.w5(32'hba2e2756),
	.w6(32'h3a344909),
	.w7(32'h3b12f586),
	.w8(32'hba6ce303),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba567103),
	.w1(32'hb94fd7e5),
	.w2(32'hba22d94d),
	.w3(32'hba12fb02),
	.w4(32'hb9c75404),
	.w5(32'h3a7b2b1f),
	.w6(32'hba8886f8),
	.w7(32'hba0f3b53),
	.w8(32'h3abe0cf6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a580c63),
	.w1(32'h39705afc),
	.w2(32'h39f7bb7f),
	.w3(32'h39a8430b),
	.w4(32'h3a0da1ff),
	.w5(32'hba85c0b4),
	.w6(32'h3a2d4a91),
	.w7(32'h3aa59303),
	.w8(32'hba8733e3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab989eb),
	.w1(32'hbb00ee1c),
	.w2(32'hbafe7fe3),
	.w3(32'hbab2d596),
	.w4(32'hbabf3ea4),
	.w5(32'hba738c49),
	.w6(32'hbb1aa971),
	.w7(32'hbaef9489),
	.w8(32'hbb036aef),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99adff1),
	.w1(32'hba051c43),
	.w2(32'hb77c3326),
	.w3(32'hb9f5b66f),
	.w4(32'hba2ff87a),
	.w5(32'h3980df4b),
	.w6(32'hbacfa848),
	.w7(32'hbae05471),
	.w8(32'h38b3bcb9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997f137),
	.w1(32'hbaa1689f),
	.w2(32'hba52f571),
	.w3(32'hb9b96165),
	.w4(32'hba3db9ff),
	.w5(32'h3a8204bf),
	.w6(32'hba874d87),
	.w7(32'hb9581de8),
	.w8(32'h3aafc3c9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a628213),
	.w1(32'h391cb2c8),
	.w2(32'h3a0b1dfe),
	.w3(32'h3a71ca9d),
	.w4(32'h3a004318),
	.w5(32'hba2dbd84),
	.w6(32'h3a3dd664),
	.w7(32'h39e4d5f5),
	.w8(32'hba8b331b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba911246),
	.w1(32'hbaaa51ed),
	.w2(32'hba1783ce),
	.w3(32'hba65d3ef),
	.w4(32'hbab7b324),
	.w5(32'h3ac3975c),
	.w6(32'hbacac6f2),
	.w7(32'hba95faa2),
	.w8(32'h3ae50e59),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9b5d9),
	.w1(32'h3afbe542),
	.w2(32'h3ad940ee),
	.w3(32'h3af3de07),
	.w4(32'h3ad74cbe),
	.w5(32'hbade9daa),
	.w6(32'h3b0cd31b),
	.w7(32'h3b0afb2f),
	.w8(32'hbb0270ac),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e119),
	.w1(32'hbb133325),
	.w2(32'hbb126c7a),
	.w3(32'hbafddb80),
	.w4(32'hbab3912a),
	.w5(32'h3ae48b1c),
	.w6(32'hbab498d7),
	.w7(32'hbadf29eb),
	.w8(32'h3b0b7a1f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae47355),
	.w1(32'h3acc116f),
	.w2(32'h3b0217cc),
	.w3(32'h3a9b3ccc),
	.w4(32'h3acfd436),
	.w5(32'h39b58d89),
	.w6(32'h3aeec8ba),
	.w7(32'h3b10b633),
	.w8(32'hba7339dc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80a389),
	.w1(32'hba99605b),
	.w2(32'hba374e03),
	.w3(32'hb989959a),
	.w4(32'h3709e5bf),
	.w5(32'hb929ff86),
	.w6(32'hba9fb943),
	.w7(32'hba144eef),
	.w8(32'hb84dd007),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe6278),
	.w1(32'h3ab49446),
	.w2(32'h3a4c3391),
	.w3(32'h3a963183),
	.w4(32'h3a7536b6),
	.w5(32'hb934c6a6),
	.w6(32'hb9e2a0ec),
	.w7(32'hba0a5514),
	.w8(32'hba6be533),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb863294c),
	.w1(32'h393cfa8f),
	.w2(32'hb8b32327),
	.w3(32'hba0d77b2),
	.w4(32'hb9f1b4e7),
	.w5(32'hba89e38b),
	.w6(32'hba75b2b3),
	.w7(32'hba3f76dc),
	.w8(32'hba968832),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4754a),
	.w1(32'hba920d84),
	.w2(32'hba426d30),
	.w3(32'hba24cafb),
	.w4(32'h3964e36a),
	.w5(32'hba2febd7),
	.w6(32'hba5ffe91),
	.w7(32'h3a020501),
	.w8(32'hb9d635bc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cfc76),
	.w1(32'hb9c05152),
	.w2(32'hb9e4f663),
	.w3(32'hb981a19b),
	.w4(32'hb5d903c4),
	.w5(32'hba96c74e),
	.w6(32'h3905f50e),
	.w7(32'hb91ba085),
	.w8(32'hba898bfe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6997eb),
	.w1(32'hbaa35533),
	.w2(32'hba8e9466),
	.w3(32'hb9ef68dd),
	.w4(32'hba0f7ba0),
	.w5(32'hba409608),
	.w6(32'hba47b828),
	.w7(32'hba434274),
	.w8(32'hb8b485cc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d64744),
	.w1(32'hb9a7aabe),
	.w2(32'hba68d86c),
	.w3(32'hba168d65),
	.w4(32'hb9c4e1ac),
	.w5(32'hba289a54),
	.w6(32'hb929a5c1),
	.w7(32'hb9bffca0),
	.w8(32'hba8a763f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f229c),
	.w1(32'h372f649c),
	.w2(32'hba364198),
	.w3(32'hb9fe5e4d),
	.w4(32'hb946f332),
	.w5(32'h3afb5194),
	.w6(32'hb9356430),
	.w7(32'h394e4187),
	.w8(32'h3b0afde8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af292bd),
	.w1(32'h3abff0c6),
	.w2(32'h3acaa2b0),
	.w3(32'h3a99800f),
	.w4(32'h3ad9c0db),
	.w5(32'hb9bee24f),
	.w6(32'h3addb327),
	.w7(32'h3b0e8e0a),
	.w8(32'h3a6a0409),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7495f0),
	.w1(32'h3ab7db61),
	.w2(32'h3ab99f74),
	.w3(32'h3a3f9b24),
	.w4(32'h39e1c760),
	.w5(32'hb9b3a2b7),
	.w6(32'h3abe8671),
	.w7(32'h3a49ff51),
	.w8(32'hb9982a74),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fff48),
	.w1(32'hba0b8091),
	.w2(32'hba067be0),
	.w3(32'hb977027b),
	.w4(32'hb9abfdb2),
	.w5(32'h378f6124),
	.w6(32'hb98e8bbc),
	.w7(32'hba813a35),
	.w8(32'h3a890ed7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a9b41),
	.w1(32'h369b1faf),
	.w2(32'hb78849ec),
	.w3(32'hb99656f1),
	.w4(32'h39663728),
	.w5(32'hb97348f7),
	.w6(32'h3a49fcd1),
	.w7(32'h3a003937),
	.w8(32'hbaa2dbc8),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16df74),
	.w1(32'hba8a8f51),
	.w2(32'hb8b6e460),
	.w3(32'hb9c30a77),
	.w4(32'h3980b841),
	.w5(32'hba76bd94),
	.w6(32'hba9c05fd),
	.w7(32'hba848134),
	.w8(32'hba74ba05),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87cfd6),
	.w1(32'hba07fa78),
	.w2(32'hba1bcb2d),
	.w3(32'hba2f221b),
	.w4(32'hb97e6c11),
	.w5(32'hbaab32f2),
	.w6(32'hb985e0c3),
	.w7(32'hba0b6d08),
	.w8(32'hba1d3e43),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a35b74),
	.w1(32'hb98bf970),
	.w2(32'hb9ded009),
	.w3(32'hba02c055),
	.w4(32'hb8628369),
	.w5(32'hbab732d3),
	.w6(32'hb9235c39),
	.w7(32'hb9bde5c5),
	.w8(32'hbab986a1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba886c41),
	.w1(32'hbaabdf81),
	.w2(32'hba036740),
	.w3(32'hbaaec319),
	.w4(32'hba73a252),
	.w5(32'h39f5b8f2),
	.w6(32'hbaa2b928),
	.w7(32'hba66dce5),
	.w8(32'h39ce0f7f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3799e),
	.w1(32'h3a349ccd),
	.w2(32'h39e62966),
	.w3(32'h3a5a50b6),
	.w4(32'h39f3e602),
	.w5(32'hba35bd50),
	.w6(32'h3a4d990e),
	.w7(32'h389215fa),
	.w8(32'hb6dc67a6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9021abe),
	.w1(32'h39ad899e),
	.w2(32'hba8761e8),
	.w3(32'h3a1d22ae),
	.w4(32'hba240dd9),
	.w5(32'h39af7283),
	.w6(32'h3ab2c935),
	.w7(32'hb9335010),
	.w8(32'h3853320f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927ebc6),
	.w1(32'h39be0c40),
	.w2(32'hb99a15a2),
	.w3(32'hb84abaf2),
	.w4(32'hb8f657f8),
	.w5(32'h3a94db04),
	.w6(32'hb9acfe5f),
	.w7(32'hb8aa98f1),
	.w8(32'h3a016160),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a877297),
	.w1(32'h3a3b25ce),
	.w2(32'h39958383),
	.w3(32'h3a2d33f4),
	.w4(32'hb9d9cde9),
	.w5(32'hba02afdb),
	.w6(32'h39627f48),
	.w7(32'hb9e2e2b9),
	.w8(32'hb8935ca6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0860a7),
	.w1(32'hba7a9271),
	.w2(32'hba698226),
	.w3(32'hb9800782),
	.w4(32'hba48c2d7),
	.w5(32'hb985df94),
	.w6(32'hb8ad004b),
	.w7(32'hba519ea7),
	.w8(32'hb997048f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8805d0a),
	.w1(32'hba1cfba9),
	.w2(32'h38055753),
	.w3(32'hb9709fb4),
	.w4(32'hb945cacb),
	.w5(32'hb9c5f7d6),
	.w6(32'hb9a60bb6),
	.w7(32'hb9308af9),
	.w8(32'hb981c7a3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba560407),
	.w1(32'hb8dece78),
	.w2(32'hb92853f7),
	.w3(32'h37fd488b),
	.w4(32'h390d9905),
	.w5(32'hbb0a87c8),
	.w6(32'h3a776a3d),
	.w7(32'hb8cc66ca),
	.w8(32'hbadd8f7a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb7540),
	.w1(32'hba8590c1),
	.w2(32'hba151328),
	.w3(32'hbabbdde4),
	.w4(32'hbaa3b5ca),
	.w5(32'h39f0f94b),
	.w6(32'hba65d46c),
	.w7(32'hb9d56782),
	.w8(32'h3a0fa2fc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c2542),
	.w1(32'h3a20d79b),
	.w2(32'h39fd88bc),
	.w3(32'h3a3799cf),
	.w4(32'h397dda1a),
	.w5(32'hbb0729ed),
	.w6(32'h3a81cc6c),
	.w7(32'h39b0bd8a),
	.w8(32'hbb02a1f1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d3201),
	.w1(32'hbacbb24a),
	.w2(32'hbac4cf97),
	.w3(32'hbaf1fceb),
	.w4(32'hbac2a813),
	.w5(32'hba8af67b),
	.w6(32'hbab5cb0a),
	.w7(32'hbab64dd0),
	.w8(32'hbae44633),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7a82c),
	.w1(32'hba316c40),
	.w2(32'hb9bb8a7b),
	.w3(32'hba534d82),
	.w4(32'hb9d891f3),
	.w5(32'h386aee25),
	.w6(32'hbae27c67),
	.w7(32'hba779087),
	.w8(32'hba489e6f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21262b),
	.w1(32'hb96566e1),
	.w2(32'hba0bdd98),
	.w3(32'hb9ac8610),
	.w4(32'hba1a8606),
	.w5(32'hba174fc9),
	.w6(32'hba966c84),
	.w7(32'hba8478d3),
	.w8(32'hbaa1b1aa),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba471e35),
	.w1(32'hba34aeea),
	.w2(32'hba03747e),
	.w3(32'hb62ab8c4),
	.w4(32'h3924b032),
	.w5(32'hb953f069),
	.w6(32'hba873108),
	.w7(32'hb9f69066),
	.w8(32'hb992bbb5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c94b7a),
	.w1(32'hb8b11aca),
	.w2(32'hb97d56ce),
	.w3(32'h3a00aed0),
	.w4(32'h3a2010bc),
	.w5(32'hbaedc30a),
	.w6(32'h39e78de7),
	.w7(32'h395ef9cd),
	.w8(32'hbb1d89cb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04bbab),
	.w1(32'hbb0cc07c),
	.w2(32'hbabbde02),
	.w3(32'hbb1daa98),
	.w4(32'hbb2ba7b6),
	.w5(32'hba4764fb),
	.w6(32'hbb80dd13),
	.w7(32'hbb1ffcb0),
	.w8(32'hb9bf02fe),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f558a),
	.w1(32'hba40bc09),
	.w2(32'hba68e0e7),
	.w3(32'hba45a323),
	.w4(32'hb9706450),
	.w5(32'h3a4b7891),
	.w6(32'h391bd1e0),
	.w7(32'h36dba4f7),
	.w8(32'h38cf1143),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b0227),
	.w1(32'h395273c2),
	.w2(32'h390a376b),
	.w3(32'h3a1a4f95),
	.w4(32'h38449d05),
	.w5(32'hbb174cd3),
	.w6(32'hb7a3d75c),
	.w7(32'h38cdf2bd),
	.w8(32'hba9e9643),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3db1af),
	.w1(32'hb91dbe9c),
	.w2(32'hba2723ad),
	.w3(32'hba4a768e),
	.w4(32'hbabf5945),
	.w5(32'h39aa1c00),
	.w6(32'h398c2050),
	.w7(32'hb9f33a8c),
	.w8(32'h39b4aa19),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39529974),
	.w1(32'h3953503b),
	.w2(32'h39cbe34a),
	.w3(32'h3977620c),
	.w4(32'hb7a1198e),
	.w5(32'h38eb5f8f),
	.w6(32'h3980292c),
	.w7(32'h39b72363),
	.w8(32'hb921cd60),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad0780),
	.w1(32'hba470399),
	.w2(32'hba821c34),
	.w3(32'hba8437f8),
	.w4(32'hba8030fa),
	.w5(32'h3a6e449b),
	.w6(32'hba10b81d),
	.w7(32'hbabddb75),
	.w8(32'h39eb825f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d2bf58),
	.w1(32'hba5291ca),
	.w2(32'hb9103cdc),
	.w3(32'hba1ecc2f),
	.w4(32'hb9e8a104),
	.w5(32'hba212d41),
	.w6(32'hba7281a3),
	.w7(32'hb9b0d612),
	.w8(32'hba40de29),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961323f),
	.w1(32'hba3d225d),
	.w2(32'hb8fafc3e),
	.w3(32'hb9109fe8),
	.w4(32'h38061770),
	.w5(32'h3981860b),
	.w6(32'hb9cf299b),
	.w7(32'hb9d76fd2),
	.w8(32'h394a7a71),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37976b40),
	.w1(32'hb99b94bd),
	.w2(32'h393cb6ff),
	.w3(32'h39e1cca3),
	.w4(32'h3a24c9e2),
	.w5(32'hb98b8d61),
	.w6(32'h39a4f5aa),
	.w7(32'h3a036026),
	.w8(32'h3840a356),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f3da5),
	.w1(32'h39cd4663),
	.w2(32'hb97bc8dc),
	.w3(32'h39d3a242),
	.w4(32'h3a7a085c),
	.w5(32'hba71c0ec),
	.w6(32'hb9cc4cc4),
	.w7(32'h39abea8b),
	.w8(32'hbaba068e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04b32e),
	.w1(32'hba87dd40),
	.w2(32'hba6ee258),
	.w3(32'hba4f599c),
	.w4(32'hb949e13d),
	.w5(32'hbacd25a3),
	.w6(32'hba79b19d),
	.w7(32'hba5c4601),
	.w8(32'hba755bf7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba775951),
	.w1(32'hb9e86648),
	.w2(32'hba3b7978),
	.w3(32'h38915ee2),
	.w4(32'h39303d9b),
	.w5(32'hbae4b9f2),
	.w6(32'hb9ac17d1),
	.w7(32'h39792a1f),
	.w8(32'hbad67940),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86ec00),
	.w1(32'hba8dc0e6),
	.w2(32'hba28094d),
	.w3(32'hba80fe82),
	.w4(32'hba3c08d9),
	.w5(32'hb70b3250),
	.w6(32'hbab69d3c),
	.w7(32'hba5aa14a),
	.w8(32'h37fae8fb),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0b75d),
	.w1(32'h3a8b1c3b),
	.w2(32'h3acdb4b3),
	.w3(32'h39913724),
	.w4(32'h3a91b57a),
	.w5(32'h38ed9755),
	.w6(32'h38b4a0d0),
	.w7(32'h3a8238d5),
	.w8(32'hb9452c1f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39315f39),
	.w1(32'hb993537c),
	.w2(32'h39e30567),
	.w3(32'hb9c6bbd9),
	.w4(32'hb8f2aaa8),
	.w5(32'hba4da280),
	.w6(32'hba41e57d),
	.w7(32'hb60a56ef),
	.w8(32'hba74804f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934cb10),
	.w1(32'h38750bc8),
	.w2(32'hba1ec9fa),
	.w3(32'h3a804b44),
	.w4(32'hba10c4f7),
	.w5(32'hb988ba2c),
	.w6(32'hbab10715),
	.w7(32'hb946f98f),
	.w8(32'hba838edd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b10bc),
	.w1(32'hba92db0f),
	.w2(32'hba089604),
	.w3(32'hb88edc3c),
	.w4(32'h398be288),
	.w5(32'hb9259504),
	.w6(32'hba1d9427),
	.w7(32'hb833a584),
	.w8(32'hb8fc9bb6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828102a),
	.w1(32'hb9239131),
	.w2(32'hb9c80c56),
	.w3(32'h39e8d6a8),
	.w4(32'h39946200),
	.w5(32'h3b0c240a),
	.w6(32'hb9cb9bdb),
	.w7(32'hb9431dfe),
	.w8(32'h3b05517c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af45657),
	.w1(32'h3b72b577),
	.w2(32'h3b2049a2),
	.w3(32'h3b7a1b5b),
	.w4(32'h3af4c8d0),
	.w5(32'h3b8a6f3b),
	.w6(32'h3be40de4),
	.w7(32'h3b052d63),
	.w8(32'h3be11d32),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec35f9),
	.w1(32'hbbae459c),
	.w2(32'hbb18cf67),
	.w3(32'hba7640b8),
	.w4(32'hbba9f150),
	.w5(32'h3a9054c0),
	.w6(32'h3a3f4ec4),
	.w7(32'hbbd97562),
	.w8(32'h3aa42d4e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89e971),
	.w1(32'h3b0fe775),
	.w2(32'hbb61fd2a),
	.w3(32'h3b0c7b00),
	.w4(32'hbb274beb),
	.w5(32'hba47c8e3),
	.w6(32'hbb4d75bc),
	.w7(32'h385c86ae),
	.w8(32'hbc07e1a1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f2f70),
	.w1(32'h3aa63edf),
	.w2(32'h3b9deb8b),
	.w3(32'hb9e7c352),
	.w4(32'hbb252b3b),
	.w5(32'hba151f0d),
	.w6(32'hbbcc4716),
	.w7(32'h3932038b),
	.w8(32'h39b2efee),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e179fa),
	.w1(32'hbb64f17b),
	.w2(32'h3a1c8774),
	.w3(32'h3af76e3e),
	.w4(32'hbad4cf35),
	.w5(32'hbb2d03ea),
	.w6(32'h39a1883a),
	.w7(32'hbb33dfb3),
	.w8(32'h3a353816),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7755e7),
	.w1(32'h3b1e191f),
	.w2(32'hbaad60a1),
	.w3(32'hbbabeb35),
	.w4(32'hbbaa25c8),
	.w5(32'h3b820cad),
	.w6(32'hbb4b035e),
	.w7(32'hbb18b4d5),
	.w8(32'hbbd1c690),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56b5ee),
	.w1(32'h3b73f2b5),
	.w2(32'hbbaa9295),
	.w3(32'h3c24109f),
	.w4(32'h3b5fc471),
	.w5(32'hbba4c21a),
	.w6(32'h3c35739c),
	.w7(32'h3c2086f1),
	.w8(32'hbb8ba6ba),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070189),
	.w1(32'h3aa2dec3),
	.w2(32'h3a2e9810),
	.w3(32'hb77f20ec),
	.w4(32'h3b061299),
	.w5(32'h3b2b79f5),
	.w6(32'hbbaab787),
	.w7(32'h3a902b00),
	.w8(32'hbbcd4e67),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e6e53),
	.w1(32'hb9fe957b),
	.w2(32'h3b1f981b),
	.w3(32'hbbc86948),
	.w4(32'hba7a6d82),
	.w5(32'hba6e8129),
	.w6(32'h3bb10831),
	.w7(32'h3b894149),
	.w8(32'hbb11853a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b4e16),
	.w1(32'hbb8733cb),
	.w2(32'hbad44903),
	.w3(32'hbafca3d0),
	.w4(32'hbaf9f8f8),
	.w5(32'hbaa5a6fa),
	.w6(32'h3b38bcd0),
	.w7(32'hb8fad821),
	.w8(32'hbb280490),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1906a1),
	.w1(32'hbb19a61b),
	.w2(32'hbb16d00e),
	.w3(32'hba73f668),
	.w4(32'hbaf6da4e),
	.w5(32'hbadc2670),
	.w6(32'h3ac033d5),
	.w7(32'hbb0c6aa9),
	.w8(32'hba7db7b5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5936e8),
	.w1(32'h3aa38c83),
	.w2(32'h3abfc7ae),
	.w3(32'h39da0563),
	.w4(32'h3966f5cb),
	.w5(32'h3bd9854c),
	.w6(32'h3b87d410),
	.w7(32'h3b374059),
	.w8(32'hba08a88a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5b284),
	.w1(32'hbb322407),
	.w2(32'hba730717),
	.w3(32'h39e51343),
	.w4(32'hbafdcdc1),
	.w5(32'h3abad7f7),
	.w6(32'h3b0b9459),
	.w7(32'hbaa77925),
	.w8(32'h3ac6e5e5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f8917),
	.w1(32'h3b205604),
	.w2(32'h3b3ca183),
	.w3(32'hbab3a752),
	.w4(32'h3ad25f6f),
	.w5(32'hbb9a9ce6),
	.w6(32'h3b51ac61),
	.w7(32'h3bf1ad9e),
	.w8(32'hbb6ff2da),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d46ff),
	.w1(32'h3b102f49),
	.w2(32'h3b35649f),
	.w3(32'h3a2b1575),
	.w4(32'h3b220fc4),
	.w5(32'hbb144211),
	.w6(32'h3b64edf1),
	.w7(32'h3b0a556d),
	.w8(32'h3b171b86),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00354b),
	.w1(32'h3a5324be),
	.w2(32'h3b195a55),
	.w3(32'hbb0c9b42),
	.w4(32'hbb0e5d9a),
	.w5(32'h38838887),
	.w6(32'hba30b18e),
	.w7(32'hbb78e360),
	.w8(32'h3bf0f163),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41268d),
	.w1(32'h3b119664),
	.w2(32'hbacbe453),
	.w3(32'hbbfe9c6b),
	.w4(32'h3c0fd72b),
	.w5(32'h3a875281),
	.w6(32'h3c36a7be),
	.w7(32'hbb6497f2),
	.w8(32'hbacedbd7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a599c94),
	.w1(32'h3c1864ef),
	.w2(32'hba6be0ae),
	.w3(32'hb9823d6c),
	.w4(32'hbbb2338a),
	.w5(32'hb9f830ad),
	.w6(32'h3ac0df3e),
	.w7(32'h3b6a70b7),
	.w8(32'hba0c015d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55ab61),
	.w1(32'h3a42345e),
	.w2(32'h3a97f743),
	.w3(32'hba3354d7),
	.w4(32'h3b9456d5),
	.w5(32'h38ed92ae),
	.w6(32'h3a15ff61),
	.w7(32'h3b0baec5),
	.w8(32'hbb21764e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fa321),
	.w1(32'hbbde639a),
	.w2(32'h3b3d11ce),
	.w3(32'h3b3fccd5),
	.w4(32'hbb6fe9fe),
	.w5(32'h3a20b5ef),
	.w6(32'hbaf4f986),
	.w7(32'h3ba2a07e),
	.w8(32'h3adccd9d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4afa8f),
	.w1(32'h391c0882),
	.w2(32'h39ba8532),
	.w3(32'hba01eef3),
	.w4(32'hbb4e0d95),
	.w5(32'h3b9ab268),
	.w6(32'h3b2bb855),
	.w7(32'hbb3374d4),
	.w8(32'h3c0e878a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ffa44),
	.w1(32'h3bd791c6),
	.w2(32'h3baabbee),
	.w3(32'h3bbbcd94),
	.w4(32'h3ba75658),
	.w5(32'hbb0dc9d7),
	.w6(32'h3a62e874),
	.w7(32'h3b8e318e),
	.w8(32'hbb059b5a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4609e4),
	.w1(32'h3b784360),
	.w2(32'h3bdda1fb),
	.w3(32'h3992b2a1),
	.w4(32'h3a1a5146),
	.w5(32'hb92f72e1),
	.w6(32'hba5ad968),
	.w7(32'h3c0adcae),
	.w8(32'hba94381e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a561e),
	.w1(32'hbb1581e4),
	.w2(32'h3b2c4994),
	.w3(32'hbaa1bc66),
	.w4(32'h3aadd562),
	.w5(32'hba6ae5d5),
	.w6(32'hbbf63269),
	.w7(32'hbaa95da7),
	.w8(32'hbbbb0e5a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a59f4c),
	.w1(32'h3ae1611f),
	.w2(32'hbb82a3cc),
	.w3(32'hb91d2b9f),
	.w4(32'hbb47ce13),
	.w5(32'hba551920),
	.w6(32'hbb80e3f6),
	.w7(32'hbabae820),
	.w8(32'h3ab15de6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54983a),
	.w1(32'hbabe7475),
	.w2(32'h3ae78bbc),
	.w3(32'h39a3269c),
	.w4(32'h3afe266c),
	.w5(32'hbb6e4a69),
	.w6(32'h3acaf914),
	.w7(32'hbb9188f1),
	.w8(32'h3ac3bcdd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb218e94),
	.w1(32'hba70a27c),
	.w2(32'h39937ebb),
	.w3(32'hb9a1832c),
	.w4(32'hbbb1245d),
	.w5(32'h3c0af389),
	.w6(32'h3b7cdb4e),
	.w7(32'hbb3661fb),
	.w8(32'hbae389d6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a395dba),
	.w1(32'h3ad5918c),
	.w2(32'h3c082994),
	.w3(32'h3b2d8397),
	.w4(32'h3b303688),
	.w5(32'hbaa1fa71),
	.w6(32'h3a064c0f),
	.w7(32'h3b9dbc84),
	.w8(32'hba8cc35a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443e9f),
	.w1(32'hbb9d73af),
	.w2(32'hbb8a60a7),
	.w3(32'hba258e86),
	.w4(32'hbb052ebb),
	.w5(32'hb9d593c7),
	.w6(32'h3ba07ea6),
	.w7(32'hbab45cdf),
	.w8(32'hba1eb38d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a9409),
	.w1(32'hbb2515e9),
	.w2(32'h3aa3a3d7),
	.w3(32'hba7853e8),
	.w4(32'h3ab22ad5),
	.w5(32'hbbafb716),
	.w6(32'hbbebb034),
	.w7(32'h3b02ba32),
	.w8(32'hbbc112af),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9c416),
	.w1(32'hbb9ad663),
	.w2(32'hbb0a0c81),
	.w3(32'hbb272a31),
	.w4(32'hba4ed2e6),
	.w5(32'h3b256351),
	.w6(32'hbba15cac),
	.w7(32'hbb2b87ce),
	.w8(32'h3bd09882),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef8b51),
	.w1(32'h3b1b4e15),
	.w2(32'h3b9955a3),
	.w3(32'h3bdb60b8),
	.w4(32'h3c10001b),
	.w5(32'hbbba18f6),
	.w6(32'h3c7f57f2),
	.w7(32'h3c25eeef),
	.w8(32'hbb47bf8f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2051c7),
	.w1(32'h3b793015),
	.w2(32'h3a77a9b5),
	.w3(32'hbb4c696d),
	.w4(32'hbbf27da9),
	.w5(32'h3b39860b),
	.w6(32'hbaa58075),
	.w7(32'h3a7c7de7),
	.w8(32'h3a77602c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896d936),
	.w1(32'h39d6855d),
	.w2(32'hb9c0f272),
	.w3(32'hbacdee8c),
	.w4(32'hbb35d636),
	.w5(32'h3b8f2a7b),
	.w6(32'h3b8f2727),
	.w7(32'hbaae4c9b),
	.w8(32'hbaad18c5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955422a),
	.w1(32'hbc168b4f),
	.w2(32'hbb0184a3),
	.w3(32'hbb1e4f32),
	.w4(32'hbb8292eb),
	.w5(32'hbb0be007),
	.w6(32'hbbb6385a),
	.w7(32'hbb5b20d7),
	.w8(32'hbb38b659),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ed71a),
	.w1(32'h39f72fc2),
	.w2(32'h387d22c8),
	.w3(32'h39bb7d9c),
	.w4(32'hbac177db),
	.w5(32'hbb9e76d8),
	.w6(32'h3bc397cc),
	.w7(32'h3988db35),
	.w8(32'hbb853abe),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4469db),
	.w1(32'hbbb03766),
	.w2(32'hbb8a0a60),
	.w3(32'hba1d7e9f),
	.w4(32'hbb36a37d),
	.w5(32'hbbe5ab41),
	.w6(32'h3b17b7df),
	.w7(32'hbb1eec92),
	.w8(32'hbc030f1c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39278e),
	.w1(32'hbb97acb7),
	.w2(32'hbb957c53),
	.w3(32'hbc08b16a),
	.w4(32'hbb4c478c),
	.w5(32'hbb9bc385),
	.w6(32'hbbbc00ec),
	.w7(32'hbab53d85),
	.w8(32'hbbb0ccdf),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88cfc6),
	.w1(32'hbb02d8ca),
	.w2(32'hba8d1747),
	.w3(32'hbb577f24),
	.w4(32'hba57b2ec),
	.w5(32'hba72afd2),
	.w6(32'hbb2c1732),
	.w7(32'h370eb4a5),
	.w8(32'hbac7c137),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b3928),
	.w1(32'h39fb5d78),
	.w2(32'hba15534e),
	.w3(32'h37af7c8c),
	.w4(32'hbac0dbf2),
	.w5(32'h398402ac),
	.w6(32'h3bb4d175),
	.w7(32'hba384621),
	.w8(32'hb9b7c40b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48507e),
	.w1(32'hba8ed08e),
	.w2(32'h3a0529cb),
	.w3(32'h3a329b72),
	.w4(32'hbb052ddc),
	.w5(32'hbae67625),
	.w6(32'h3bf7b90f),
	.w7(32'hbb159a97),
	.w8(32'hbb68bd70),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadcaa9),
	.w1(32'hb97a7c33),
	.w2(32'hba53adfc),
	.w3(32'hbba034cc),
	.w4(32'h39df4e0a),
	.w5(32'h3ac96781),
	.w6(32'hbad5e060),
	.w7(32'hbb92fb94),
	.w8(32'h3b2e7659),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0e35d),
	.w1(32'h3c16335a),
	.w2(32'h3b2b1969),
	.w3(32'h3ba5eb1c),
	.w4(32'h3bec0514),
	.w5(32'hba0c5e70),
	.w6(32'h3c68f466),
	.w7(32'h3b9b4598),
	.w8(32'hb8d1cf60),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a282d8e),
	.w1(32'hba5bdaf7),
	.w2(32'h3a224e0d),
	.w3(32'hbba792b6),
	.w4(32'h3b688b50),
	.w5(32'h3adab092),
	.w6(32'hba14e19e),
	.w7(32'h3b664c76),
	.w8(32'hba8e8039),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90de9e),
	.w1(32'hbb38d3b6),
	.w2(32'hbab73799),
	.w3(32'h3b2b9557),
	.w4(32'hba91eba5),
	.w5(32'hbb196cf0),
	.w6(32'h3b967988),
	.w7(32'h3b15dc35),
	.w8(32'h3aedc824),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5ccaa),
	.w1(32'hbabb6b74),
	.w2(32'h3b008f92),
	.w3(32'h3b198672),
	.w4(32'hbb8b9701),
	.w5(32'hbb91656b),
	.w6(32'h3aab53a0),
	.w7(32'h3b0c1143),
	.w8(32'hbb661d72),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed3054),
	.w1(32'hbbd3a462),
	.w2(32'hbb0a738b),
	.w3(32'h3aa2cf23),
	.w4(32'hbaa07e2d),
	.w5(32'hbb0679ad),
	.w6(32'h3bb4e47c),
	.w7(32'h3a90c311),
	.w8(32'hbb0e85a9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05178c),
	.w1(32'hba460322),
	.w2(32'hbae4a396),
	.w3(32'hbb6b7784),
	.w4(32'hbac23d92),
	.w5(32'h3ae3f8f0),
	.w6(32'hbafc4068),
	.w7(32'hb9acf996),
	.w8(32'hbb071ae6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910e73),
	.w1(32'h3a5e0932),
	.w2(32'h3a563bdb),
	.w3(32'hbb86072d),
	.w4(32'hbbe7f680),
	.w5(32'hb9d3351f),
	.w6(32'h396d0703),
	.w7(32'hbb2aff65),
	.w8(32'hbb7460ac),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35987095),
	.w1(32'hbbc95981),
	.w2(32'h3b29b4fa),
	.w3(32'h38cc956b),
	.w4(32'hbb89b8ba),
	.w5(32'hba9a911d),
	.w6(32'hb98ead02),
	.w7(32'h3994d3f8),
	.w8(32'h3b122bdb),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17cc45),
	.w1(32'h3a3e3d41),
	.w2(32'hba45b370),
	.w3(32'hb9b40f51),
	.w4(32'hbb2ed943),
	.w5(32'h38d8c4f0),
	.w6(32'hbb2b3ffb),
	.w7(32'h3aead7d9),
	.w8(32'hbaa7a51b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85acfc),
	.w1(32'hbad4a385),
	.w2(32'hbb017470),
	.w3(32'hba66bcb2),
	.w4(32'h3a8b1ef4),
	.w5(32'h394c7fa8),
	.w6(32'h39546645),
	.w7(32'hba6f522e),
	.w8(32'h3b409d99),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28128a),
	.w1(32'h3b574bec),
	.w2(32'h3b68e7bf),
	.w3(32'h3b4c7e13),
	.w4(32'h3ae70c77),
	.w5(32'h3b988af9),
	.w6(32'h3c0a160d),
	.w7(32'hbb48bb0e),
	.w8(32'h3b9e74d3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23321d),
	.w1(32'hbb38ff17),
	.w2(32'hbab9ac0e),
	.w3(32'h396b7e81),
	.w4(32'hbb994598),
	.w5(32'hbb20f155),
	.w6(32'h3a144efd),
	.w7(32'hbb8aed6f),
	.w8(32'hba955893),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bf337),
	.w1(32'h3c187107),
	.w2(32'h3911bb42),
	.w3(32'hba5e80cb),
	.w4(32'h394629f0),
	.w5(32'h3b03536f),
	.w6(32'hbb078a7a),
	.w7(32'h3b16ffa6),
	.w8(32'hba25bc68),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe2f5c),
	.w1(32'hbb67da5b),
	.w2(32'h391e6cc4),
	.w3(32'hba8b1baf),
	.w4(32'hbb1c9d48),
	.w5(32'h3b948b89),
	.w6(32'hb9db3585),
	.w7(32'h3b47effd),
	.w8(32'hbb839abf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65a2cb),
	.w1(32'hbb6752a5),
	.w2(32'hbb281edc),
	.w3(32'hbb86d120),
	.w4(32'hbbb39e74),
	.w5(32'hbb6620e2),
	.w6(32'hbb7e75ce),
	.w7(32'hbb2a76da),
	.w8(32'hbb4a7c1d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4512f1),
	.w1(32'h3a540051),
	.w2(32'h3a7cb36c),
	.w3(32'hbad38931),
	.w4(32'hbab5998b),
	.w5(32'h3b3726a0),
	.w6(32'hb90db952),
	.w7(32'h3a17d146),
	.w8(32'hbad332f5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf31ad),
	.w1(32'hbaccd701),
	.w2(32'hb94d1a52),
	.w3(32'hbb80970e),
	.w4(32'h3b1b8490),
	.w5(32'hbb3167bf),
	.w6(32'hbb870ae8),
	.w7(32'h3a00af98),
	.w8(32'hbb84a6a2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098597),
	.w1(32'hbb53d69f),
	.w2(32'h3b3ca5a8),
	.w3(32'hbb1de51e),
	.w4(32'h3b28b196),
	.w5(32'h3b0b64cc),
	.w6(32'hbb6e7801),
	.w7(32'h3b58a21e),
	.w8(32'h3c26dea9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b5632),
	.w1(32'hbaa25005),
	.w2(32'h3a697af9),
	.w3(32'h3c2da815),
	.w4(32'hbb59c547),
	.w5(32'hbb8ffcfb),
	.w6(32'h3ba268dc),
	.w7(32'hbbd9719a),
	.w8(32'hbba33d48),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee7d90),
	.w1(32'hbbd1b440),
	.w2(32'hbb578e88),
	.w3(32'hbba4a48b),
	.w4(32'hbaf5c381),
	.w5(32'h3b76cd10),
	.w6(32'h3ad7f8d2),
	.w7(32'hbb12c78c),
	.w8(32'hbb36bbe7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2233b4),
	.w1(32'h3c4085cf),
	.w2(32'h3c00fff3),
	.w3(32'hbbddcdf2),
	.w4(32'h3ae00f15),
	.w5(32'hba1c3878),
	.w6(32'hb9fe87c7),
	.w7(32'h3c25188b),
	.w8(32'h3b238518),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2919c2),
	.w1(32'hbae29c7b),
	.w2(32'hba0a01e5),
	.w3(32'hb8e02760),
	.w4(32'h3bac6af2),
	.w5(32'h3b1247c0),
	.w6(32'hba60c689),
	.w7(32'h3b37c175),
	.w8(32'hb882f4a0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb055832),
	.w1(32'h3ab5d8f3),
	.w2(32'hb9cd3bd7),
	.w3(32'h3a478156),
	.w4(32'h3aad33f7),
	.w5(32'hbb6763b1),
	.w6(32'hbae4adb5),
	.w7(32'h3b11c044),
	.w8(32'h3bef9964),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ea9f8),
	.w1(32'h3b7d37dd),
	.w2(32'h3992d54f),
	.w3(32'h3c252ec4),
	.w4(32'hb99b6410),
	.w5(32'h3b1b8538),
	.w6(32'h3b222854),
	.w7(32'hba71eac9),
	.w8(32'hba4d8981),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1b034),
	.w1(32'hbb39483e),
	.w2(32'hbb18d087),
	.w3(32'h3b569053),
	.w4(32'hbb903634),
	.w5(32'hbb05e058),
	.w6(32'hbc103a6e),
	.w7(32'h3b816788),
	.w8(32'hbb9b9888),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7d5f8),
	.w1(32'hba860f54),
	.w2(32'h3ad6acea),
	.w3(32'hbb4cc6a7),
	.w4(32'hbb2a166b),
	.w5(32'hb9baa91f),
	.w6(32'h3b69c04a),
	.w7(32'h3a65341e),
	.w8(32'hb98e175c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e0d6a),
	.w1(32'h3a386ec2),
	.w2(32'h3a6e8995),
	.w3(32'h3b08ff8a),
	.w4(32'h3a9ab675),
	.w5(32'hbb79a858),
	.w6(32'h3b3e02e8),
	.w7(32'h3ae3dec2),
	.w8(32'hbb4af0c3),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb419915),
	.w1(32'hbb52e523),
	.w2(32'hbc12f0e6),
	.w3(32'h3a51537a),
	.w4(32'hbb589240),
	.w5(32'h3a35bad4),
	.w6(32'h3a94f2e6),
	.w7(32'hbb84d3cc),
	.w8(32'h3ab6742d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab11af1),
	.w1(32'h38436680),
	.w2(32'h3a77900e),
	.w3(32'h3a025012),
	.w4(32'h3b96dfb6),
	.w5(32'hba20961f),
	.w6(32'h3b81cb0b),
	.w7(32'h3a807208),
	.w8(32'hb9f0c5ce),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82c659),
	.w1(32'hbbb83e9d),
	.w2(32'hbb0e5ca7),
	.w3(32'hba31308f),
	.w4(32'hba3848ef),
	.w5(32'h3b859fd6),
	.w6(32'h3b568ddf),
	.w7(32'hb93628d3),
	.w8(32'h3acaf4c4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3a1f7),
	.w1(32'h3bfbf798),
	.w2(32'h3b8fafc1),
	.w3(32'h3c1d8e93),
	.w4(32'h3b686e5a),
	.w5(32'hbac84351),
	.w6(32'h3c1053bc),
	.w7(32'h3b16283c),
	.w8(32'h3b97af55),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89988a),
	.w1(32'h3bbc1668),
	.w2(32'h3be5c1d9),
	.w3(32'h3c40d882),
	.w4(32'h3bdaab24),
	.w5(32'h3b28d8e7),
	.w6(32'h3d181f04),
	.w7(32'h3b87c279),
	.w8(32'h3b1acc86),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec86b),
	.w1(32'h3b6810fe),
	.w2(32'hbb08ba5c),
	.w3(32'h3ae1c6a8),
	.w4(32'h3a7a5e1d),
	.w5(32'hbb96d736),
	.w6(32'h3b29f8f5),
	.w7(32'h3b29ec03),
	.w8(32'hba8f6bc1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc4bf9),
	.w1(32'hbc045ee3),
	.w2(32'hbb84d8b5),
	.w3(32'hbc075420),
	.w4(32'hbbd5984d),
	.w5(32'h3ad05755),
	.w6(32'hbb87a4b8),
	.w7(32'hbb5af36f),
	.w8(32'h3b15a181),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac6345),
	.w1(32'hbbcfadeb),
	.w2(32'hbb1b21ca),
	.w3(32'hbc150e0e),
	.w4(32'hbc0a66f2),
	.w5(32'h3b62a23d),
	.w6(32'hbabfe534),
	.w7(32'h3b0b6cb5),
	.w8(32'h3bf2452d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba130d9),
	.w1(32'h3bd67efb),
	.w2(32'h3bae74c0),
	.w3(32'h3b8ad9af),
	.w4(32'h3bbf5da1),
	.w5(32'hbab392f1),
	.w6(32'h3c176401),
	.w7(32'h3b59b44d),
	.w8(32'h3b517ae2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06a0ff),
	.w1(32'h3c00f370),
	.w2(32'hb9bc1c4d),
	.w3(32'h3b3b1b8b),
	.w4(32'h3bb86a8f),
	.w5(32'hbb0d3a61),
	.w6(32'h3bc4eccc),
	.w7(32'hbb041169),
	.w8(32'hbb0db09f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ccc51),
	.w1(32'hbb831c51),
	.w2(32'hbb8baab9),
	.w3(32'hbae59507),
	.w4(32'hbae5d943),
	.w5(32'h3adecfa9),
	.w6(32'h39718dbb),
	.w7(32'hbb170490),
	.w8(32'h3b5bd8ef),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0bc17),
	.w1(32'hbb7627ca),
	.w2(32'hbad845ed),
	.w3(32'hbc02d207),
	.w4(32'hba860d78),
	.w5(32'hbb97c0bf),
	.w6(32'hbbec5303),
	.w7(32'hbb020fd7),
	.w8(32'hbb923fd8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab76986),
	.w1(32'hbaa50454),
	.w2(32'h35496ac4),
	.w3(32'hbb899e40),
	.w4(32'hb8f73569),
	.w5(32'h3b89cdaf),
	.w6(32'h3ae7af73),
	.w7(32'hba3cbd96),
	.w8(32'h3b6041b8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e75fc),
	.w1(32'hba0c51cf),
	.w2(32'h3bd6725d),
	.w3(32'h3baad547),
	.w4(32'h3bed4e56),
	.w5(32'h3b9ade6a),
	.w6(32'hba1b239f),
	.w7(32'h3b48cb0b),
	.w8(32'h3b8e4589),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44ea78),
	.w1(32'hbafb8ade),
	.w2(32'h3c08845e),
	.w3(32'hbb31588d),
	.w4(32'h3bf6ba2c),
	.w5(32'hbb3178b1),
	.w6(32'hbbae3df6),
	.w7(32'h3c209db4),
	.w8(32'hbbf9a343),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87c698),
	.w1(32'hbbb7e299),
	.w2(32'h3998cbf2),
	.w3(32'hba8c352b),
	.w4(32'hbbb5b1c9),
	.w5(32'hbb42241c),
	.w6(32'h3a2a21c2),
	.w7(32'hbb97f70a),
	.w8(32'hbb086adb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88cfab),
	.w1(32'hbb009d44),
	.w2(32'hbbb83127),
	.w3(32'hbbbbb88c),
	.w4(32'h3a0404e3),
	.w5(32'h397bc6c5),
	.w6(32'h3a29017b),
	.w7(32'hbb886b75),
	.w8(32'hb9b6cdde),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b23b8),
	.w1(32'h3b0abb17),
	.w2(32'h3ab918c7),
	.w3(32'h37fc7f1b),
	.w4(32'h3bbf726a),
	.w5(32'hba0ffa7d),
	.w6(32'h3b98451e),
	.w7(32'h3b9b3740),
	.w8(32'hbb139203),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9e14e),
	.w1(32'h3b073292),
	.w2(32'h3c6b5853),
	.w3(32'h3b1dbbf8),
	.w4(32'h3c1bb649),
	.w5(32'hbb1c8656),
	.w6(32'h3c369f09),
	.w7(32'h3c6735e7),
	.w8(32'hbb8907be),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb969a72),
	.w1(32'hbb6da2cc),
	.w2(32'hbaf87f34),
	.w3(32'hbac8823d),
	.w4(32'hba086077),
	.w5(32'hbb0494d5),
	.w6(32'hba30090c),
	.w7(32'hbb1b1343),
	.w8(32'hbaeb9b10),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb946e85),
	.w1(32'hbb5dcb79),
	.w2(32'hbb3dde23),
	.w3(32'hbacee42f),
	.w4(32'hbb1a31d2),
	.w5(32'h398db8b4),
	.w6(32'h3b82c57e),
	.w7(32'h3b0c5b33),
	.w8(32'hba9f02a8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b0aca),
	.w1(32'hbb65ab0f),
	.w2(32'hbb01d72a),
	.w3(32'hbab6878e),
	.w4(32'hbb92e3cc),
	.w5(32'hba37cbe2),
	.w6(32'h3b667bf2),
	.w7(32'h3b08f701),
	.w8(32'h3b199812),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b47fe),
	.w1(32'hbbf8c4dd),
	.w2(32'hbbbfe510),
	.w3(32'hbb576bb5),
	.w4(32'hbbe8228d),
	.w5(32'h3b0b9db0),
	.w6(32'h3bd583f0),
	.w7(32'h38fb7962),
	.w8(32'hbb1ff8ba),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab02f21),
	.w1(32'h3b2754ce),
	.w2(32'h369c81c7),
	.w3(32'h398b72c1),
	.w4(32'hbb5a788b),
	.w5(32'hbae43169),
	.w6(32'hbbc3e627),
	.w7(32'hbb8741b3),
	.w8(32'h3a8260ea),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d2e73),
	.w1(32'hbabdc327),
	.w2(32'hbacf429f),
	.w3(32'hbb09d5c0),
	.w4(32'h3ad11fe6),
	.w5(32'hba84f996),
	.w6(32'hbb2a44cd),
	.w7(32'h3ad20839),
	.w8(32'hbb9a7f2d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf24cd),
	.w1(32'hbbf742ca),
	.w2(32'h3ad44ef9),
	.w3(32'hbb203199),
	.w4(32'hbba9a1b8),
	.w5(32'h3a85df39),
	.w6(32'hbb89b1b5),
	.w7(32'hbb1f2bde),
	.w8(32'hbbb4be1a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc20dcf),
	.w1(32'hbc005990),
	.w2(32'hbab457b0),
	.w3(32'h3af5a1b0),
	.w4(32'hbaa42353),
	.w5(32'hbb0d451e),
	.w6(32'hbabf4d5d),
	.w7(32'hbbcca3bb),
	.w8(32'hbb79409e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb988c82),
	.w1(32'hbb3bbb0f),
	.w2(32'hbab0112c),
	.w3(32'hbabcf9a8),
	.w4(32'hbb47cede),
	.w5(32'h3a9c1193),
	.w6(32'hbb6e7230),
	.w7(32'hbb3c8452),
	.w8(32'h3c6bd625),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c816b44),
	.w1(32'h3c45972e),
	.w2(32'h3b40620f),
	.w3(32'h3c3ed84f),
	.w4(32'h3c02d81c),
	.w5(32'hbb328115),
	.w6(32'h3cec5a3d),
	.w7(32'h3b9b994f),
	.w8(32'hbbe49a33),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ea1f8),
	.w1(32'hbbd39c87),
	.w2(32'hbb5a7c93),
	.w3(32'hbc213d97),
	.w4(32'hba993362),
	.w5(32'hbb076d1f),
	.w6(32'hbb26c83b),
	.w7(32'hba371d5c),
	.w8(32'hbabf20ac),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dc260),
	.w1(32'h3b041661),
	.w2(32'h3c014384),
	.w3(32'h3bf7a427),
	.w4(32'h3b9c7c98),
	.w5(32'h3baf72cb),
	.w6(32'h3c6adf84),
	.w7(32'h3b42d67d),
	.w8(32'h3bb73848),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1e9d2),
	.w1(32'h3ba857fb),
	.w2(32'h3b4f2298),
	.w3(32'h3beefbb7),
	.w4(32'h3a907bfe),
	.w5(32'hb9a1904b),
	.w6(32'h3aaba510),
	.w7(32'h3b5817c6),
	.w8(32'h3960e369),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b6b40),
	.w1(32'hba64b74e),
	.w2(32'hbb0b0d4d),
	.w3(32'h3b4b159c),
	.w4(32'hbb418999),
	.w5(32'hbaccf081),
	.w6(32'hbad6324c),
	.w7(32'h3ab9c207),
	.w8(32'h3b374b77),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad89873),
	.w1(32'h3b282d32),
	.w2(32'h3b607253),
	.w3(32'h3a048a52),
	.w4(32'h3b8f510f),
	.w5(32'h39f6eddd),
	.w6(32'h3b622917),
	.w7(32'hba433920),
	.w8(32'h3bd745aa),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6add0b),
	.w1(32'h3ab41392),
	.w2(32'h3bf07762),
	.w3(32'h3c2dba73),
	.w4(32'h3c0b51e9),
	.w5(32'hbb3397f7),
	.w6(32'h3c421951),
	.w7(32'h3c64702e),
	.w8(32'hbb7de8c3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce386),
	.w1(32'h3b309f04),
	.w2(32'h3b70e4ca),
	.w3(32'h38456e98),
	.w4(32'hb9867e2a),
	.w5(32'hbb0ed123),
	.w6(32'h3b9396b6),
	.w7(32'h3a1c7a62),
	.w8(32'h3b4dae1b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7390e),
	.w1(32'h3c074f15),
	.w2(32'h3b9d90fb),
	.w3(32'h39a1f37e),
	.w4(32'h3be5ef22),
	.w5(32'h3a1a01fe),
	.w6(32'h3bf14aff),
	.w7(32'h3af5e5cc),
	.w8(32'h3b13dac1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08529c),
	.w1(32'hbb260bea),
	.w2(32'h39043514),
	.w3(32'h3b544985),
	.w4(32'hbaa0d6ca),
	.w5(32'hbb5c6475),
	.w6(32'h3ba61e51),
	.w7(32'hbbfe3931),
	.w8(32'hbaa9875c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93cdbd),
	.w1(32'hbbb4e43c),
	.w2(32'hbaef4981),
	.w3(32'hbb771e7a),
	.w4(32'hba17e707),
	.w5(32'hbad314f6),
	.w6(32'h3aa5c59c),
	.w7(32'hbb53eb08),
	.w8(32'hb9be3aff),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb770d34),
	.w1(32'hbb732383),
	.w2(32'hbbe0ce93),
	.w3(32'hba8c55c8),
	.w4(32'hbb8b27a5),
	.w5(32'hbba52a68),
	.w6(32'h3a45c4ee),
	.w7(32'hbad3b7ab),
	.w8(32'hbb3097cd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92d0b0),
	.w1(32'hbb8a45c2),
	.w2(32'hbb047012),
	.w3(32'hbb56ef66),
	.w4(32'hbb6d767e),
	.w5(32'hbb48ed4a),
	.w6(32'h3b8f6c20),
	.w7(32'hbabdc2b3),
	.w8(32'hb98a5c4c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bceacb9),
	.w1(32'h3bcb3425),
	.w2(32'hbaec3162),
	.w3(32'h3a451415),
	.w4(32'h3c0729f8),
	.w5(32'hbb10c4f0),
	.w6(32'h3ace16f5),
	.w7(32'hbb0cfb55),
	.w8(32'h3b049854),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31cbf1),
	.w1(32'h3acf57c5),
	.w2(32'h3a6ecd24),
	.w3(32'h39947f07),
	.w4(32'h3a934e09),
	.w5(32'hba0d857b),
	.w6(32'hb920f8b4),
	.w7(32'hbae1dd4e),
	.w8(32'hba72f490),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39488dd4),
	.w1(32'hbb7a1586),
	.w2(32'hbb517157),
	.w3(32'h3bb87dd0),
	.w4(32'h3a6698ca),
	.w5(32'h3bd78c6c),
	.w6(32'hba855aa9),
	.w7(32'hbb47c4d0),
	.w8(32'h3bc30380),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2da918),
	.w1(32'h3b84af39),
	.w2(32'h3c02514d),
	.w3(32'h3b64fb55),
	.w4(32'h3ba564ec),
	.w5(32'h3b02b947),
	.w6(32'h3c8c9a9b),
	.w7(32'h3bd0a9ab),
	.w8(32'h3b899fd6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3f2f8),
	.w1(32'h3af5cacf),
	.w2(32'h39187872),
	.w3(32'h3ba71725),
	.w4(32'h3bc4c392),
	.w5(32'h3ab3f80a),
	.w6(32'h3b0f063b),
	.w7(32'hb875c71b),
	.w8(32'hb8518393),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c18af),
	.w1(32'hbb4a7a9e),
	.w2(32'hba6f8c0b),
	.w3(32'hbb09e59d),
	.w4(32'hbb8979d7),
	.w5(32'hba29cadd),
	.w6(32'h3ba1155f),
	.w7(32'hba62f8c8),
	.w8(32'hbbbb4a7a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb57528),
	.w1(32'hbb905202),
	.w2(32'h3bd04c86),
	.w3(32'h3b6186e5),
	.w4(32'h39c3d33f),
	.w5(32'h3aea3ad8),
	.w6(32'hba6492dd),
	.w7(32'h3c571b8b),
	.w8(32'hbad41722),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9b1f9),
	.w1(32'hba1bcad6),
	.w2(32'h3a9283dd),
	.w3(32'hb9a9bf07),
	.w4(32'hbaecd22b),
	.w5(32'hbb347025),
	.w6(32'hbadf8d2f),
	.w7(32'hbb410b00),
	.w8(32'hbb61f039),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba33b9d),
	.w1(32'hbb656cca),
	.w2(32'hbade7e99),
	.w3(32'hba57011e),
	.w4(32'hbb538218),
	.w5(32'hbac34641),
	.w6(32'h3bc1108c),
	.w7(32'hb9d257ba),
	.w8(32'hbb626cfe),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a8ac3),
	.w1(32'hbbae3010),
	.w2(32'hbb42eb96),
	.w3(32'hbba0e60a),
	.w4(32'hbb2ac95a),
	.w5(32'h3a094e28),
	.w6(32'hbc165338),
	.w7(32'hbb8100e5),
	.w8(32'h3ab4c329),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2bd1e),
	.w1(32'hb9c91479),
	.w2(32'hba994153),
	.w3(32'hb7b7af86),
	.w4(32'h39096ee2),
	.w5(32'h3bc3834b),
	.w6(32'h3b525a54),
	.w7(32'h3b2a4f27),
	.w8(32'h3bdc96c8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fea3b),
	.w1(32'hba9f39fa),
	.w2(32'h396ea98d),
	.w3(32'hb8ec30ae),
	.w4(32'h3bb23a45),
	.w5(32'hba31f189),
	.w6(32'h3aa5d667),
	.w7(32'h3b232651),
	.w8(32'h3c2261a1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8826db),
	.w1(32'hba8e61ce),
	.w2(32'hbb0b942b),
	.w3(32'hbb0ffc44),
	.w4(32'h3955ba5b),
	.w5(32'hbb832cab),
	.w6(32'h3ac610c6),
	.w7(32'hb92f1733),
	.w8(32'hba5b7bf6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85557e),
	.w1(32'hbab75661),
	.w2(32'hbb2928db),
	.w3(32'hbb3ef58a),
	.w4(32'hbb00e5ca),
	.w5(32'hba93e8fa),
	.w6(32'h3bc127de),
	.w7(32'h3b29741f),
	.w8(32'h3a6a80ab),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3df89f),
	.w1(32'hba2183f3),
	.w2(32'hba8de6ef),
	.w3(32'hb95692e8),
	.w4(32'hba756394),
	.w5(32'hbb50bb76),
	.w6(32'h3b2b9100),
	.w7(32'h3b3acc8d),
	.w8(32'hbc1bf269),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1434ab),
	.w1(32'hb897b51f),
	.w2(32'h38d399d0),
	.w3(32'hbb92ebce),
	.w4(32'hbb871b27),
	.w5(32'hbb8b5378),
	.w6(32'h3b48bbad),
	.w7(32'h3757d1c3),
	.w8(32'h3b33b42d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826757),
	.w1(32'h3b158c72),
	.w2(32'hbbc525a7),
	.w3(32'hbb2af424),
	.w4(32'hbb56ac61),
	.w5(32'h39d2f5b2),
	.w6(32'h3bbf43b3),
	.w7(32'hba74c83c),
	.w8(32'hbb2041aa),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2c85c),
	.w1(32'hbb29d954),
	.w2(32'hbb8fd110),
	.w3(32'hbbafa51c),
	.w4(32'hb88df03d),
	.w5(32'hbf3bf51e),
	.w6(32'hbbad1eae),
	.w7(32'hbb08b7f4),
	.w8(32'hbea7c35a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbee21ac9),
	.w1(32'hbf852c73),
	.w2(32'hbe660805),
	.w3(32'hbf1622a2),
	.w4(32'hbeffd459),
	.w5(32'h3e02c44c),
	.w6(32'hbd8e8784),
	.w7(32'hbeeda331),
	.w8(32'hbf1b3cbf),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3ae7a2),
	.w1(32'hbf8dfdf8),
	.w2(32'hbeb9e80e),
	.w3(32'hbddd8016),
	.w4(32'hbee2d8e3),
	.w5(32'hbee90ae1),
	.w6(32'h3d50d9a1),
	.w7(32'hbf7b3064),
	.w8(32'hbf35f334),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec673cf),
	.w1(32'h3dd36cd0),
	.w2(32'hbe93c7d3),
	.w3(32'hbebc97f1),
	.w4(32'h3e29430f),
	.w5(32'hbe5d214f),
	.w6(32'hbf846f3b),
	.w7(32'hbf563d91),
	.w8(32'hbf693f7b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf976069),
	.w1(32'hbe9eea89),
	.w2(32'hbf0386db),
	.w3(32'hbf763bd4),
	.w4(32'hbf0995c4),
	.w5(32'hbe11f1c3),
	.w6(32'hbeb8fb75),
	.w7(32'hbf04b07f),
	.w8(32'hbd5411d1),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbef538d6),
	.w1(32'hbf49842d),
	.w2(32'hbf2d675e),
	.w3(32'hbf12ae64),
	.w4(32'hbdf5fc44),
	.w5(32'hbdebdbd3),
	.w6(32'hbec7deb8),
	.w7(32'hbea610a5),
	.w8(32'hbeb9fbf5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe910457),
	.w1(32'hbf23b2d9),
	.w2(32'hbe94480b),
	.w3(32'h3e9c23d1),
	.w4(32'hbeb4e699),
	.w5(32'h3e0f2952),
	.w6(32'hbecdf57d),
	.w7(32'hbf4dbe1e),
	.w8(32'hbeb8fd4e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe817602),
	.w1(32'hbe8d6a7d),
	.w2(32'hbed28162),
	.w3(32'hbf080abb),
	.w4(32'hbecde37b),
	.w5(32'hbe8ef7f0),
	.w6(32'hbf491c6e),
	.w7(32'hbf22e938),
	.w8(32'hbe41ad74),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbea8619e),
	.w1(32'hbed83836),
	.w2(32'hbea8fc2f),
	.w3(32'h3e9e40a5),
	.w4(32'hbec093e1),
	.w5(32'hbf07bb38),
	.w6(32'hbf423b8a),
	.w7(32'hbd6da239),
	.w8(32'hbe9784b1),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbde14c80),
	.w1(32'hbe174b7f),
	.w2(32'hbf625523),
	.w3(32'hbf7db69d),
	.w4(32'hbf8179ed),
	.w5(32'hbf42d47c),
	.w6(32'hbe112c40),
	.w7(32'hbde7b9fb),
	.w8(32'hbebfbc1d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf3399f9),
	.w1(32'hbeada4d3),
	.w2(32'hbf8735cd),
	.w3(32'hbf6bfe3e),
	.w4(32'hbf54d0e3),
	.w5(32'hbf08040d),
	.w6(32'hbf1a7c2b),
	.w7(32'hbca4aab0),
	.w8(32'hbf3e0421),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbea8b21d),
	.w1(32'hbf2a693d),
	.w2(32'hbed15b7a),
	.w3(32'h3e80edc9),
	.w4(32'hbeb520e5),
	.w5(32'hbe8e86d7),
	.w6(32'h3e286cea),
	.w7(32'hbd44808c),
	.w8(32'hbe956955),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec26601),
	.w1(32'hbe542392),
	.w2(32'h3e15cc51),
	.w3(32'hbeba8689),
	.w4(32'hbeaba183),
	.w5(32'h3e76b6bf),
	.w6(32'hbef663e4),
	.w7(32'hbea851f8),
	.w8(32'hbe5bd484),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbee801ad),
	.w1(32'hbee046cd),
	.w2(32'hbf3f49db),
	.w3(32'h3cddabf1),
	.w4(32'hbf0e8694),
	.w5(32'hbf3b001d),
	.w6(32'h3d6b3e56),
	.w7(32'hbe78e109),
	.w8(32'hbf271fa1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf5eb4e0),
	.w1(32'hbe8e3784),
	.w2(32'hbf70bf32),
	.w3(32'hbe9df45d),
	.w4(32'h3f7bf131),
	.w5(32'hbf649f9f),
	.w6(32'hbe4679e5),
	.w7(32'hbd15352b),
	.w8(32'hbf052091),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f5a86c8),
	.w1(32'h3f5ad17f),
	.w2(32'h3f36eae4),
	.w3(32'h3f11a2fa),
	.w4(32'h3f17a629),
	.w5(32'h3f502fab),
	.w6(32'h3f81d0ba),
	.w7(32'h3f80b25c),
	.w8(32'h3f74962e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f22895b),
	.w1(32'h3f0592fb),
	.w2(32'h3f480598),
	.w3(32'h3f380b6b),
	.w4(32'h3f15563e),
	.w5(32'h3f83dea5),
	.w6(32'h3f03460b),
	.w7(32'h3f892e51),
	.w8(32'h3f6a01ec),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f88feef),
	.w1(32'h3f309727),
	.w2(32'h3f21a47e),
	.w3(32'h3f526a70),
	.w4(32'h3f847b5b),
	.w5(32'h3f6f660a),
	.w6(32'h3f386bb6),
	.w7(32'h3f311314),
	.w8(32'h3f8009cc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3f0f51),
	.w1(32'h3f719dd9),
	.w2(32'h3f82ea7c),
	.w3(32'h3f91ade3),
	.w4(32'h3f490a6d),
	.w5(32'h3f8be176),
	.w6(32'h3f9e3095),
	.w7(32'h3f392cf9),
	.w8(32'h3f84fb33),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ee63078),
	.w1(32'h3f6f8738),
	.w2(32'h3f160562),
	.w3(32'h3f134169),
	.w4(32'h3f793567),
	.w5(32'h3f5272a7),
	.w6(32'h3f4b2812),
	.w7(32'h3f6c58a8),
	.w8(32'h3f96df5c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f35d897),
	.w1(32'h3f31909a),
	.w2(32'h3f3bbaeb),
	.w3(32'h3f078a70),
	.w4(32'h3f5798f7),
	.w5(32'h3f72cae7),
	.w6(32'h3f442ae6),
	.w7(32'h3f996f91),
	.w8(32'h3f478719),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f37fb99),
	.w1(32'h3f55fc73),
	.w2(32'h3f1f70a3),
	.w3(32'h3f82a411),
	.w4(32'h3f363d55),
	.w5(32'h3f97c4df),
	.w6(32'h3f42d8c5),
	.w7(32'h3f3473e8),
	.w8(32'h3f767634),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f16f01b),
	.w1(32'h3f47bcd1),
	.w2(32'h3f12af28),
	.w3(32'h3f28fbf0),
	.w4(32'h3fadfbcd),
	.w5(32'h3f17922d),
	.w6(32'h3f433ae8),
	.w7(32'h3f45f645),
	.w8(32'h3f7bf3b0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f7da491),
	.w1(32'h3f6673db),
	.w2(32'h3f82d42f),
	.w3(32'h3f385d32),
	.w4(32'h3f3d5850),
	.w5(32'h3f23bb30),
	.w6(32'h3f004135),
	.w7(32'h3f1b424c),
	.w8(32'h3f6d7b32),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f55181f),
	.w1(32'h3f9057be),
	.w2(32'h3f65ad14),
	.w3(32'h3f3be3ef),
	.w4(32'h3f592154),
	.w5(32'h3f293520),
	.w6(32'h3f697c40),
	.w7(32'h3f1ca01a),
	.w8(32'h3f855209),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f81e917),
	.w1(32'h3f5ba2eb),
	.w2(32'h3f514461),
	.w3(32'h3f7dd24e),
	.w4(32'h3f0dc073),
	.w5(32'h3f438215),
	.w6(32'h3f3a593e),
	.w7(32'h3f314ab2),
	.w8(32'h3f4f1cf7),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f80c909),
	.w1(32'h3f464391),
	.w2(32'h3f623c02),
	.w3(32'h3f33fc1b),
	.w4(32'h3f2822ce),
	.w5(32'h3f1fa006),
	.w6(32'h3f5a8c8d),
	.w7(32'h3f0ff336),
	.w8(32'h3f38cba8),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f50f83c),
	.w1(32'h3f1b6f6e),
	.w2(32'h3f8b1bd1),
	.w3(32'h3f261cd5),
	.w4(32'h3f52ae78),
	.w5(32'h3f1d49c2),
	.w6(32'h3f383092),
	.w7(32'h3f543ecf),
	.w8(32'h3f5a27c0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f4ab69f),
	.w1(32'h3f2e094f),
	.w2(32'h3e863285),
	.w3(32'h3f63205d),
	.w4(32'h3f41ef61),
	.w5(32'h3f355682),
	.w6(32'h3f81a71b),
	.w7(32'h3f1f7940),
	.w8(32'h3f6c8c6a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f8a5f35),
	.w1(32'hbd86ce73),
	.w2(32'hbe9a688f),
	.w3(32'h3f4012dc),
	.w4(32'hbe0ef667),
	.w5(32'h3eaa4f03),
	.w6(32'hbd25f9c0),
	.w7(32'hbd9a113b),
	.w8(32'hbe3ec42a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe177970),
	.w1(32'hbdc1b234),
	.w2(32'hbecff725),
	.w3(32'hbe1084a8),
	.w4(32'hbee0cc4a),
	.w5(32'hbe50001c),
	.w6(32'hbe9edf20),
	.w7(32'h3d372b93),
	.w8(32'hbd9df27b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule