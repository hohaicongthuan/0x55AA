module layer_10_featuremap_505(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a96b6a),
	.w1(32'hb88737b0),
	.w2(32'hb915a5c5),
	.w3(32'hb894f4af),
	.w4(32'hb984ed0e),
	.w5(32'hb91b8242),
	.w6(32'hb9a3f8fd),
	.w7(32'hb961503e),
	.w8(32'hba0b23a1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c37ad),
	.w1(32'h3a70a076),
	.w2(32'h3ac1a25d),
	.w3(32'h3af2d51d),
	.w4(32'hba2277d0),
	.w5(32'h390a34f9),
	.w6(32'h3a4aa76a),
	.w7(32'hba9e34d8),
	.w8(32'h391094c3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982b819),
	.w1(32'h39754f52),
	.w2(32'hb9b6bd0d),
	.w3(32'h37dcc4fe),
	.w4(32'h3a4248f2),
	.w5(32'h391c0d03),
	.w6(32'hb98946f8),
	.w7(32'h3945e65e),
	.w8(32'hba52415a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946e2e6),
	.w1(32'hb8bde0b3),
	.w2(32'hba39b968),
	.w3(32'h390fad8c),
	.w4(32'h39ace1cc),
	.w5(32'hbb01a7f2),
	.w6(32'h39c16b7f),
	.w7(32'h3a249b38),
	.w8(32'h39c44490),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37872ab6),
	.w1(32'h396f3f92),
	.w2(32'hb996820f),
	.w3(32'h39ad7200),
	.w4(32'h3816924b),
	.w5(32'h39c3a8b0),
	.w6(32'hb91dfeac),
	.w7(32'h3856c6f1),
	.w8(32'h390cc2d0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc6998),
	.w1(32'h39e68389),
	.w2(32'h392a4e71),
	.w3(32'hb9701349),
	.w4(32'h3a3c1e6a),
	.w5(32'h3aa28540),
	.w6(32'hb8dfe8a5),
	.w7(32'h3a29d9e6),
	.w8(32'h39e7f93a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39ffa2),
	.w1(32'h3b43d98b),
	.w2(32'h3b90eda2),
	.w3(32'h3900e463),
	.w4(32'h3b2779b2),
	.w5(32'h3b4bf54c),
	.w6(32'hb915958b),
	.w7(32'h3b4d74ed),
	.w8(32'h3ba0a7ee),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83277c),
	.w1(32'h3b54ae31),
	.w2(32'h3aae88ff),
	.w3(32'h3abc167b),
	.w4(32'h3af54e1e),
	.w5(32'hb929f544),
	.w6(32'h3b81d0de),
	.w7(32'h3b0d5753),
	.w8(32'hba456cb4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3ecc5),
	.w1(32'h38d74b1f),
	.w2(32'hb942b3d5),
	.w3(32'h39abb435),
	.w4(32'hba5e94d9),
	.w5(32'hbadaeb78),
	.w6(32'h3a04c375),
	.w7(32'hba4e92cc),
	.w8(32'hb9a0b82e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc35916),
	.w1(32'h3bacc74f),
	.w2(32'h3c128199),
	.w3(32'h39708d53),
	.w4(32'hbac0867f),
	.w5(32'h3a259a15),
	.w6(32'hb9c72416),
	.w7(32'hbb06fc78),
	.w8(32'h3adf3271),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94dac49),
	.w1(32'h395357b7),
	.w2(32'h3953427f),
	.w3(32'h3819a920),
	.w4(32'h391c21a0),
	.w5(32'h3a46f377),
	.w6(32'hb94df7ce),
	.w7(32'h37e085c7),
	.w8(32'h3a725dd9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165707),
	.w1(32'hbb3703b8),
	.w2(32'h39f1ce97),
	.w3(32'hbb39b74b),
	.w4(32'hbb2b8804),
	.w5(32'h3abca46e),
	.w6(32'hbac7603d),
	.w7(32'hbad971a5),
	.w8(32'h3b5b84c2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a3739),
	.w1(32'h3b2077e4),
	.w2(32'h3bd65141),
	.w3(32'hbb3eb651),
	.w4(32'hbb4be3e9),
	.w5(32'hba0d802f),
	.w6(32'hbb4a65e3),
	.w7(32'hbae9f029),
	.w8(32'h3adeb9dd),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab953af),
	.w1(32'h3b139963),
	.w2(32'h3ac5d8cf),
	.w3(32'h3a876fb2),
	.w4(32'h3b1a97bb),
	.w5(32'h3ac1f4f7),
	.w6(32'h39f13247),
	.w7(32'h3a3b5d73),
	.w8(32'h3a9baf9e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b522cc7),
	.w1(32'h3a23e828),
	.w2(32'h3b0da2cb),
	.w3(32'h3b23cc11),
	.w4(32'hbae18a9e),
	.w5(32'h39dd033a),
	.w6(32'h3b30b322),
	.w7(32'hbaf8ec11),
	.w8(32'hb9f7a2ed),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2360e),
	.w1(32'h3ba5deec),
	.w2(32'h3be6a932),
	.w3(32'h3abf0436),
	.w4(32'hba6af172),
	.w5(32'h3a0dfbc2),
	.w6(32'hb9818dea),
	.w7(32'hbabef700),
	.w8(32'h3a330569),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c367d),
	.w1(32'h38f1b041),
	.w2(32'h39898e27),
	.w3(32'hb80d86a7),
	.w4(32'h39879757),
	.w5(32'hb8b05f41),
	.w6(32'hb963e2a2),
	.w7(32'h39f03991),
	.w8(32'hb805fc1c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baab910),
	.w1(32'h3b916d64),
	.w2(32'h3bbe57df),
	.w3(32'hba81c1f5),
	.w4(32'hb9e63539),
	.w5(32'h3afad480),
	.w6(32'h3b60a693),
	.w7(32'h3acbe7df),
	.w8(32'h3b568f00),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e792a),
	.w1(32'h3b116c61),
	.w2(32'h3b7483bd),
	.w3(32'hbaa239c9),
	.w4(32'hba571720),
	.w5(32'h3a346b88),
	.w6(32'h37eb6ef5),
	.w7(32'hb8dcd4b1),
	.w8(32'h3aadee09),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88e8faa),
	.w1(32'hb99e81e0),
	.w2(32'hb947ff6b),
	.w3(32'hb995bce8),
	.w4(32'hb906fd9c),
	.w5(32'hba0bc929),
	.w6(32'hb94b3c69),
	.w7(32'hb946170e),
	.w8(32'hb9ecbeb4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d9f49),
	.w1(32'h392094df),
	.w2(32'h39231551),
	.w3(32'h39860030),
	.w4(32'hba0f8d5a),
	.w5(32'hb9793861),
	.w6(32'hb97d3a71),
	.w7(32'hb9ab030e),
	.w8(32'hb9301e82),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d6f0d),
	.w1(32'hbb3b52e3),
	.w2(32'hba1caebb),
	.w3(32'hba81eff8),
	.w4(32'hbb51b081),
	.w5(32'hb9919dd1),
	.w6(32'h3864eb30),
	.w7(32'hbb39ab28),
	.w8(32'hb99fe76a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6377e2),
	.w1(32'h3bc5b6ab),
	.w2(32'h3c26db10),
	.w3(32'h3bb05f5f),
	.w4(32'hbb8bacf9),
	.w5(32'h3ac3fc36),
	.w6(32'h3be0c6a1),
	.w7(32'hbb2ab024),
	.w8(32'h3bf3570b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a613a),
	.w1(32'h3b92321c),
	.w2(32'h3bcd88c3),
	.w3(32'h3b34d926),
	.w4(32'hbb043fde),
	.w5(32'h390994f6),
	.w6(32'h3ac042e8),
	.w7(32'hbad85a0e),
	.w8(32'h3a986fbd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf15fc9),
	.w1(32'h3af57b8b),
	.w2(32'h3b8901fa),
	.w3(32'h3b62e229),
	.w4(32'hbaddcbd5),
	.w5(32'h39d9b4cd),
	.w6(32'h3b8dca73),
	.w7(32'hbb336167),
	.w8(32'hb9efefe6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922a08e),
	.w1(32'h38b6a45d),
	.w2(32'h3a25845b),
	.w3(32'h398c4cbb),
	.w4(32'h39b3e268),
	.w5(32'h3abcdce0),
	.w6(32'h39d20473),
	.w7(32'hb9025e8d),
	.w8(32'h3966cc86),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b8554),
	.w1(32'hb855fe39),
	.w2(32'hb8a7a4d8),
	.w3(32'h3a9bbec9),
	.w4(32'hb9ce021e),
	.w5(32'hba196d41),
	.w6(32'h3993f943),
	.w7(32'h39a09e47),
	.w8(32'h395294a3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba690ca4),
	.w1(32'hbaf0fb6f),
	.w2(32'h3b097e8c),
	.w3(32'h399008a4),
	.w4(32'hb9e2eceb),
	.w5(32'hb9fb841b),
	.w6(32'h3a2111da),
	.w7(32'h3a3dd3a8),
	.w8(32'hba345490),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad42f00),
	.w1(32'hbb1588cb),
	.w2(32'hbb1a5e40),
	.w3(32'hba958236),
	.w4(32'hbb1a2535),
	.w5(32'hbb1032bc),
	.w6(32'h3a2d0d55),
	.w7(32'hbac67917),
	.w8(32'hbb259fff),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b484273),
	.w1(32'h3a986ec1),
	.w2(32'h3ba84f34),
	.w3(32'h3ac632c3),
	.w4(32'hba52c730),
	.w5(32'h3b0101cd),
	.w6(32'h39701da1),
	.w7(32'hbb0521c5),
	.w8(32'h3a2c5db7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ad0e0),
	.w1(32'h39449b1d),
	.w2(32'h3a2307cf),
	.w3(32'hb9f6e82a),
	.w4(32'h39b75901),
	.w5(32'h376a41d5),
	.w6(32'hb8a37b9c),
	.w7(32'h3989b6b8),
	.w8(32'h38776b9a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962bdc7),
	.w1(32'hb9b11618),
	.w2(32'hb9a60998),
	.w3(32'h397d81f4),
	.w4(32'h391db92f),
	.w5(32'hb99fa576),
	.w6(32'h398f3638),
	.w7(32'h396e07b1),
	.w8(32'hb9b550af),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b825f2c),
	.w1(32'h3b1a2489),
	.w2(32'h3b8390b8),
	.w3(32'h3aa9760a),
	.w4(32'h3932b3d3),
	.w5(32'h3a9f4c3e),
	.w6(32'h3a6265b4),
	.w7(32'h3a02b61a),
	.w8(32'h3b2511d8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6f6d8),
	.w1(32'h39a470f4),
	.w2(32'h3a46e13d),
	.w3(32'h3ac8a3e7),
	.w4(32'hb8a3988b),
	.w5(32'hba9d3c64),
	.w6(32'h3a443a06),
	.w7(32'hb99a380b),
	.w8(32'hb9a49439),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb5290),
	.w1(32'hb8f56a28),
	.w2(32'hb94a1403),
	.w3(32'hb8c5ad8a),
	.w4(32'hb958a17c),
	.w5(32'hb97134f3),
	.w6(32'h39726656),
	.w7(32'h3a1a7a96),
	.w8(32'hb9483cf6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a446eaf),
	.w1(32'h3ac820fd),
	.w2(32'h3b0446a1),
	.w3(32'hba5469c9),
	.w4(32'hb88cf481),
	.w5(32'h3a0440a5),
	.w6(32'h3a6d08d0),
	.w7(32'h3a8d4dae),
	.w8(32'h3af9d2ba),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac1dcf),
	.w1(32'hbaa4ff2d),
	.w2(32'h3bbdeae9),
	.w3(32'h39e206a2),
	.w4(32'hbbc5eb61),
	.w5(32'hbaca0997),
	.w6(32'hbb32024e),
	.w7(32'hbc1aa746),
	.w8(32'h395618af),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba56d2f),
	.w1(32'hbb98252c),
	.w2(32'h3b3244dc),
	.w3(32'h3b861963),
	.w4(32'hbbf12871),
	.w5(32'hbaeae6f1),
	.w6(32'h3b7e43c8),
	.w7(32'hbc051b3b),
	.w8(32'hba85a000),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31d952),
	.w1(32'hbb65e0e0),
	.w2(32'h3b1ab4d8),
	.w3(32'h3bbae50d),
	.w4(32'hbb2ffb54),
	.w5(32'h3a9954cd),
	.w6(32'h3bdca236),
	.w7(32'hba66b8ca),
	.w8(32'h3aeb4034),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098d6e),
	.w1(32'h3a931424),
	.w2(32'h3a36ee2f),
	.w3(32'h3b015cf3),
	.w4(32'h3aa23b23),
	.w5(32'hb9012235),
	.w6(32'h3a6801f1),
	.w7(32'h38c5e309),
	.w8(32'h38918017),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38059da1),
	.w1(32'h36b08578),
	.w2(32'hb7cfbcf9),
	.w3(32'h3a0d6ba7),
	.w4(32'h391a43c0),
	.w5(32'h3977e014),
	.w6(32'h3889f325),
	.w7(32'h39831b3c),
	.w8(32'h39ac8236),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39403b15),
	.w1(32'hba1e383c),
	.w2(32'hb9159ab1),
	.w3(32'h39c434df),
	.w4(32'hba18c299),
	.w5(32'hb9ead75b),
	.w6(32'hb984140d),
	.w7(32'hb98bf062),
	.w8(32'hb9d2b828),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac571cf),
	.w1(32'hbb6d5d63),
	.w2(32'hbadcf15b),
	.w3(32'hba77e4b2),
	.w4(32'hbb7074cd),
	.w5(32'hbaecdbef),
	.w6(32'hb9bd46e4),
	.w7(32'hbb51ef0b),
	.w8(32'hb9ba675a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3f69),
	.w1(32'h3bc74ae0),
	.w2(32'h3c1d880d),
	.w3(32'h3a81d7ef),
	.w4(32'h3903cf06),
	.w5(32'h3b5ecbdc),
	.w6(32'h39909431),
	.w7(32'hb902fece),
	.w8(32'h3b492cbe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd08df),
	.w1(32'h3b4c8020),
	.w2(32'h3bc61041),
	.w3(32'h3b819d5c),
	.w4(32'hbac4f2fe),
	.w5(32'h3a2ced34),
	.w6(32'h3af9888b),
	.w7(32'hbb38dcac),
	.w8(32'h3a940778),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1867c6),
	.w1(32'h3ba3c064),
	.w2(32'h3bd3d085),
	.w3(32'h3b1d9ed4),
	.w4(32'hbb3b9e12),
	.w5(32'hb9feb74b),
	.w6(32'h3b0ec4b1),
	.w7(32'hbb1cbe58),
	.w8(32'h39ed5c45),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc467d8),
	.w1(32'h3b2ee439),
	.w2(32'h3bb78d45),
	.w3(32'h3b07865c),
	.w4(32'hbad886cd),
	.w5(32'hb91c69cd),
	.w6(32'h3abdf186),
	.w7(32'hbad42cd8),
	.w8(32'h3a5039be),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7115a7),
	.w1(32'h3b83d87f),
	.w2(32'h3c021428),
	.w3(32'hbb86a548),
	.w4(32'hbaf70684),
	.w5(32'h3aa7ca01),
	.w6(32'hba80bc8d),
	.w7(32'hba3ddb4d),
	.w8(32'h3b322536),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b5d6e),
	.w1(32'h398e420a),
	.w2(32'h39987256),
	.w3(32'hba90b40f),
	.w4(32'hb8c72503),
	.w5(32'hb947aad0),
	.w6(32'hba673d48),
	.w7(32'h38f1d615),
	.w8(32'h39f4999b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e1407),
	.w1(32'h3a11750c),
	.w2(32'h3a061d15),
	.w3(32'hb99db924),
	.w4(32'h3897efd3),
	.w5(32'hb980e3fa),
	.w6(32'h398cc15d),
	.w7(32'h3a0c6cb1),
	.w8(32'h3a0849b6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e36207),
	.w1(32'h39a7faf3),
	.w2(32'hb9c2d97e),
	.w3(32'hb948bc21),
	.w4(32'h39d54165),
	.w5(32'hb997f9ae),
	.w6(32'h39ace0e9),
	.w7(32'h3a356e38),
	.w8(32'hb7f2c087),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43d24),
	.w1(32'h3b2b5b31),
	.w2(32'h3b63d52d),
	.w3(32'h3a84bb29),
	.w4(32'hba81cd85),
	.w5(32'hb8421b67),
	.w6(32'hb96a876e),
	.w7(32'hba90da4e),
	.w8(32'h3aa23943),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae35ffa),
	.w1(32'h3a8c76d3),
	.w2(32'h3a52cae1),
	.w3(32'h395a2493),
	.w4(32'hb97ec684),
	.w5(32'h38f8097c),
	.w6(32'hb9051aec),
	.w7(32'hb9e26f61),
	.w8(32'h399b355e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb38ae8),
	.w1(32'h3ba6d213),
	.w2(32'h3bef2ffd),
	.w3(32'h39b5fca8),
	.w4(32'h39974e4b),
	.w5(32'h3aecd48e),
	.w6(32'h3b602872),
	.w7(32'h3b15d4f5),
	.w8(32'h3b96799f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1299dc),
	.w1(32'hba23e575),
	.w2(32'h3891578f),
	.w3(32'hb909b120),
	.w4(32'hb92fd3fc),
	.w5(32'hb967dea4),
	.w6(32'h3a8e4ab3),
	.w7(32'h3a031a02),
	.w8(32'h3965f876),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954a91d),
	.w1(32'h398b076a),
	.w2(32'h39cdf02c),
	.w3(32'hb9b21468),
	.w4(32'h390a57fb),
	.w5(32'h3986697c),
	.w6(32'hb9a4c8a4),
	.w7(32'hb960eb8c),
	.w8(32'hb915de94),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ef4bb),
	.w1(32'h389b5e3e),
	.w2(32'h38923133),
	.w3(32'hb9cd78d1),
	.w4(32'hb8e64378),
	.w5(32'h395f9acf),
	.w6(32'hb92f174d),
	.w7(32'hb8065a45),
	.w8(32'h3849a9dc),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939f4b3),
	.w1(32'hb99eb46a),
	.w2(32'h390866dd),
	.w3(32'hb89b0280),
	.w4(32'hb989a6ab),
	.w5(32'h3a1346b7),
	.w6(32'h392c30c1),
	.w7(32'hb95960ec),
	.w8(32'h3a0c4449),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12ad65),
	.w1(32'hbb138d33),
	.w2(32'hbb003a7f),
	.w3(32'hb999920f),
	.w4(32'hbb12cc1e),
	.w5(32'hbad623b9),
	.w6(32'hb8b86e5b),
	.w7(32'hbb1d10a7),
	.w8(32'hbb1f6918),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba461948),
	.w1(32'hb6e4af91),
	.w2(32'hb940fd7a),
	.w3(32'hba8ee118),
	.w4(32'hba4416ee),
	.w5(32'hb99ca155),
	.w6(32'hba89bd52),
	.w7(32'hb9c00ce9),
	.w8(32'h391eeed2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2cf21),
	.w1(32'h3aa04d60),
	.w2(32'h3b0669f0),
	.w3(32'hba8e8b5a),
	.w4(32'hba85b498),
	.w5(32'h39303c3c),
	.w6(32'hba1e0e0f),
	.w7(32'h39a6a22c),
	.w8(32'h3a95a540),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75c3c1),
	.w1(32'h3aa164a7),
	.w2(32'h3b10d7a5),
	.w3(32'h3a24ea6d),
	.w4(32'h38c6871a),
	.w5(32'h39fda723),
	.w6(32'h3abaf1ee),
	.w7(32'h397a18ab),
	.w8(32'h3aa89e2a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb166b),
	.w1(32'hb941cd2b),
	.w2(32'hba25a847),
	.w3(32'h390044db),
	.w4(32'hba0f0740),
	.w5(32'hba447385),
	.w6(32'hb8587541),
	.w7(32'hb8fe7e87),
	.w8(32'hb7a7cbe1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33831a),
	.w1(32'h3997acb9),
	.w2(32'hb9632ed7),
	.w3(32'h3a16e18f),
	.w4(32'hb6b81ac6),
	.w5(32'h37c92ab9),
	.w6(32'h39e625b2),
	.w7(32'hb6d129c4),
	.w8(32'hb7e6896f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981f519),
	.w1(32'h3aac7320),
	.w2(32'h3a46588d),
	.w3(32'h39f116ad),
	.w4(32'h3a6bd5a8),
	.w5(32'hb7d3eadc),
	.w6(32'hb81244aa),
	.w7(32'h3a6e9fbe),
	.w8(32'h3a5d3d6e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c8932),
	.w1(32'h399eab56),
	.w2(32'h39f91ece),
	.w3(32'h39a2d5d0),
	.w4(32'h3909d491),
	.w5(32'h37a03a6a),
	.w6(32'h3a4b0be9),
	.w7(32'h39bb0e44),
	.w8(32'hb9290aa2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b5b56),
	.w1(32'h3bb0e5ed),
	.w2(32'h3bd99a6e),
	.w3(32'h3a369e64),
	.w4(32'h3a9e9bd7),
	.w5(32'h39216b1f),
	.w6(32'h3b0fd120),
	.w7(32'h39c3b680),
	.w8(32'h3ad16ddc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07faac),
	.w1(32'h3b9e46f4),
	.w2(32'h3bcdaf02),
	.w3(32'hb9a940ee),
	.w4(32'hbb4bd124),
	.w5(32'h39c8afc0),
	.w6(32'h3ba2eed9),
	.w7(32'h3b1800e7),
	.w8(32'h3ba2254f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be13c82),
	.w1(32'h3ae6a50a),
	.w2(32'h3b94ec1e),
	.w3(32'h3ae7859c),
	.w4(32'hbb4f9dbf),
	.w5(32'h3aa20b35),
	.w6(32'h3b987a4e),
	.w7(32'h39fcafb3),
	.w8(32'h3b405202),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ccffd),
	.w1(32'h3a6b7e9e),
	.w2(32'h3c496b44),
	.w3(32'h3bdafdf0),
	.w4(32'hbc071919),
	.w5(32'hbbe30fef),
	.w6(32'h3bf4a5de),
	.w7(32'hbc67b2ac),
	.w8(32'hbb82d3de),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b252f89),
	.w1(32'h3b696c9c),
	.w2(32'hb98da7e7),
	.w3(32'hbb97d4f5),
	.w4(32'hbb585199),
	.w5(32'h3bcc5c02),
	.w6(32'h3bc49530),
	.w7(32'h3b08798d),
	.w8(32'h3c06ca3c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad78e88),
	.w1(32'h3b08331d),
	.w2(32'h3a8b90eb),
	.w3(32'h3b63f992),
	.w4(32'h3ba8902f),
	.w5(32'h3c961cb0),
	.w6(32'h3bb7e0d7),
	.w7(32'h3ac20ef3),
	.w8(32'hbac8c6f5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac48c48),
	.w1(32'h3a8d73ff),
	.w2(32'hba267b98),
	.w3(32'h3aed678c),
	.w4(32'hbb8dfd59),
	.w5(32'hbbe83a7c),
	.w6(32'hbbf51b69),
	.w7(32'hbba13cc7),
	.w8(32'hbb9a9767),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00c66e),
	.w1(32'h3bae6765),
	.w2(32'h3c7ad366),
	.w3(32'hbbc04111),
	.w4(32'h3ba55bbb),
	.w5(32'h3cf94ac4),
	.w6(32'hbb6533e4),
	.w7(32'h3c80c16c),
	.w8(32'h3d04ead5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9801f1),
	.w1(32'hbb25cdd3),
	.w2(32'hbb926fff),
	.w3(32'h3ca7ae7a),
	.w4(32'hbc5b53ad),
	.w5(32'hbcb18774),
	.w6(32'h3cab5166),
	.w7(32'hbc645891),
	.w8(32'hbbc76ab4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50338b),
	.w1(32'hbcc3a1be),
	.w2(32'hbc9855af),
	.w3(32'hbc5e0ac6),
	.w4(32'hbba52caa),
	.w5(32'h3cc721e1),
	.w6(32'hba9eb8b6),
	.w7(32'h3bb2b68d),
	.w8(32'h3c967654),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc481f67),
	.w1(32'h3b4f176a),
	.w2(32'h3b6b27c4),
	.w3(32'h3b25b4ed),
	.w4(32'h3b99427e),
	.w5(32'hbc15223c),
	.w6(32'hbb9208ff),
	.w7(32'hbba124db),
	.w8(32'hba2410df),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0b17),
	.w1(32'hbb2add3b),
	.w2(32'h3bb447b9),
	.w3(32'h3a944a15),
	.w4(32'hbc64de8a),
	.w5(32'hbb320e52),
	.w6(32'h3a90a65d),
	.w7(32'hbbfeabed),
	.w8(32'hbb6b4333),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd398f),
	.w1(32'h3b0628b0),
	.w2(32'h3c63c9d6),
	.w3(32'hbb5d50f6),
	.w4(32'hbb59251b),
	.w5(32'h3c60cb1e),
	.w6(32'hbbb292b0),
	.w7(32'hbadf21f9),
	.w8(32'h3b876ff1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80c348),
	.w1(32'h3abd9458),
	.w2(32'h3c08c62d),
	.w3(32'h3bd4ad70),
	.w4(32'hba69817e),
	.w5(32'h3b3c73e9),
	.w6(32'hbc083435),
	.w7(32'hba21f633),
	.w8(32'h3bddbbce),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae13819),
	.w1(32'h3c8bb824),
	.w2(32'h3c69066a),
	.w3(32'h3bac1a34),
	.w4(32'h3ab8f87c),
	.w5(32'hbab3a67d),
	.w6(32'h3b2e51ec),
	.w7(32'hbb0f3209),
	.w8(32'hbb2a2492),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61a7cf),
	.w1(32'hbb5340d0),
	.w2(32'hb94673a1),
	.w3(32'h3b398591),
	.w4(32'hbb2ff960),
	.w5(32'h3bc8b60d),
	.w6(32'hbb28d8ba),
	.w7(32'hbbb447e5),
	.w8(32'h3ab6d5fc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb032457),
	.w1(32'hbbc9d220),
	.w2(32'hbc98f23d),
	.w3(32'h3b903b87),
	.w4(32'hbc3239e3),
	.w5(32'hbcfb9810),
	.w6(32'hbae22b5b),
	.w7(32'hbc822e39),
	.w8(32'hbc8b9333),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca57509),
	.w1(32'h3c37bf2e),
	.w2(32'hba32ed85),
	.w3(32'hbc45f6c9),
	.w4(32'h3b3d8245),
	.w5(32'h3c4887b3),
	.w6(32'hbb82f0bb),
	.w7(32'h3b7f2916),
	.w8(32'h3ad0460d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbc2c3),
	.w1(32'h3b0b954d),
	.w2(32'h3bca9667),
	.w3(32'h3b3999fb),
	.w4(32'hbb5b0784),
	.w5(32'h3a8d6230),
	.w6(32'hbb444aad),
	.w7(32'hbc217adc),
	.w8(32'hbb9b31c7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed9033),
	.w1(32'hbabbc828),
	.w2(32'h3b918688),
	.w3(32'hbb1b2844),
	.w4(32'h3b965062),
	.w5(32'h3c31d0ed),
	.w6(32'hbc38181d),
	.w7(32'h3bffdb89),
	.w8(32'h3bd50594),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e6128),
	.w1(32'hbb92b570),
	.w2(32'h398bd542),
	.w3(32'h3c274ed3),
	.w4(32'hbc147c40),
	.w5(32'hbb28b37e),
	.w6(32'hba1db6a9),
	.w7(32'hbb257386),
	.w8(32'hbbc55cd7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7b6c0),
	.w1(32'h3b7cf582),
	.w2(32'hbb254dea),
	.w3(32'hbb6470b6),
	.w4(32'h3b20820d),
	.w5(32'h3b939a0c),
	.w6(32'hbbbcc9c7),
	.w7(32'h3afb622a),
	.w8(32'hbc94910b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5355b6),
	.w1(32'h3a269614),
	.w2(32'h3a5d28bd),
	.w3(32'hbc0282cf),
	.w4(32'h39b9191a),
	.w5(32'hbb36a9ff),
	.w6(32'hbbbddf77),
	.w7(32'hba0a6701),
	.w8(32'h3bd731cc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcd1da),
	.w1(32'hbaa8fa13),
	.w2(32'h3ba6121a),
	.w3(32'h3b2d93ca),
	.w4(32'hba5be30d),
	.w5(32'h3c1c7dcd),
	.w6(32'h3b913a15),
	.w7(32'h3bb3a662),
	.w8(32'h3bc765f5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadad09),
	.w1(32'hbbe4a75e),
	.w2(32'hbbbc82db),
	.w3(32'h3b5f02c0),
	.w4(32'hbb896496),
	.w5(32'hbbf768ba),
	.w6(32'hbb715a4b),
	.w7(32'hbc0bd237),
	.w8(32'hbc34e823),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a307380),
	.w1(32'h3b78c56e),
	.w2(32'h3bf66177),
	.w3(32'h3ae41d95),
	.w4(32'hbb26926a),
	.w5(32'h3bb09ac2),
	.w6(32'h3bcb19ea),
	.w7(32'h3982240e),
	.w8(32'hba9a7e77),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab0c61),
	.w1(32'h3c26b6b0),
	.w2(32'h3c49ee36),
	.w3(32'h3c1e78db),
	.w4(32'h3bed1a9e),
	.w5(32'h3c4a95e9),
	.w6(32'h3be6e562),
	.w7(32'h3bf18dc3),
	.w8(32'h3c41d29e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e65ab),
	.w1(32'h3c41e833),
	.w2(32'h3ceef028),
	.w3(32'h3c3263a9),
	.w4(32'h3c8852eb),
	.w5(32'h3d1be843),
	.w6(32'h3c2f4279),
	.w7(32'h3c48d831),
	.w8(32'h3cbdee6c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a32ab),
	.w1(32'h3abc6528),
	.w2(32'h3bcf1cf8),
	.w3(32'h3c9b5caf),
	.w4(32'h3baffd46),
	.w5(32'h3be16fc8),
	.w6(32'h3c4ca445),
	.w7(32'h3b7c6f02),
	.w8(32'hbb64b70b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44a901),
	.w1(32'h3bc6d5a3),
	.w2(32'hbb50f94f),
	.w3(32'h3bf1b7b4),
	.w4(32'h3b33db41),
	.w5(32'h38159ff0),
	.w6(32'h3b522483),
	.w7(32'h3a1827a4),
	.w8(32'hbbc2ee07),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e661d),
	.w1(32'hbc0b68cb),
	.w2(32'hbbcb729c),
	.w3(32'hbb07f8ca),
	.w4(32'hbbd44a20),
	.w5(32'h3b231014),
	.w6(32'h3b960579),
	.w7(32'hbbf4c8ba),
	.w8(32'hbb78061d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ae2a77),
	.w1(32'h3c86240f),
	.w2(32'h3c5d483b),
	.w3(32'hbbd46b0a),
	.w4(32'h3922f0bd),
	.w5(32'h393cc272),
	.w6(32'h3bc53262),
	.w7(32'hbb5ace25),
	.w8(32'hbb46ed77),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d4031),
	.w1(32'h39e6cc8e),
	.w2(32'h3afb1156),
	.w3(32'h39b29e22),
	.w4(32'h3a948f8b),
	.w5(32'hba2495ef),
	.w6(32'hba760c29),
	.w7(32'hb91d5745),
	.w8(32'hbaeb1fda),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f9e8f),
	.w1(32'h3ae012f6),
	.w2(32'h3bb192cc),
	.w3(32'hbb11ce57),
	.w4(32'hb94e0dc1),
	.w5(32'h3bc7829d),
	.w6(32'h3b4f8d45),
	.w7(32'h3b3552e1),
	.w8(32'h3bb27fae),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0166c5),
	.w1(32'h3b53628e),
	.w2(32'h3c0db73f),
	.w3(32'h3c3a45bd),
	.w4(32'hbc1c633b),
	.w5(32'h3c5aeb03),
	.w6(32'h3c4a84ab),
	.w7(32'hbbf20de2),
	.w8(32'h3c06327b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75cc96),
	.w1(32'h3c21cc3b),
	.w2(32'h3c6d9280),
	.w3(32'h3b58e252),
	.w4(32'h3bb88994),
	.w5(32'h3c1759cd),
	.w6(32'h3b2145ac),
	.w7(32'hbaf60f71),
	.w8(32'h3b1eed99),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dffad),
	.w1(32'hbad7e637),
	.w2(32'h3c011849),
	.w3(32'h3c45f81e),
	.w4(32'h3c58e8fe),
	.w5(32'h3cae1d82),
	.w6(32'h3c3f0c34),
	.w7(32'hbbcdd512),
	.w8(32'h39b0dace),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4a3dd),
	.w1(32'hbcd46b36),
	.w2(32'hbb28916a),
	.w3(32'h3b18527a),
	.w4(32'hbc0e0c53),
	.w5(32'h3c6c5033),
	.w6(32'hbb0babf4),
	.w7(32'h39605dc9),
	.w8(32'h3b9c7e02),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef728e),
	.w1(32'h3c1b7c69),
	.w2(32'h3baf9f6e),
	.w3(32'hbb296576),
	.w4(32'h3ae1a3f4),
	.w5(32'h3ba8b22a),
	.w6(32'hbcd6d71e),
	.w7(32'hbc00d53b),
	.w8(32'h3b06de0f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c04a8),
	.w1(32'h39bc4bb4),
	.w2(32'h3b6821f6),
	.w3(32'h3b30f632),
	.w4(32'hbab2fcff),
	.w5(32'h3b82ee24),
	.w6(32'hbac7acdc),
	.w7(32'hbba59ebe),
	.w8(32'hbb8ed33e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9837f73),
	.w1(32'h3b790245),
	.w2(32'hbb9642ea),
	.w3(32'h3b093bb5),
	.w4(32'h3b61a464),
	.w5(32'h3aa21dd6),
	.w6(32'hbbaf872c),
	.w7(32'h3bccd029),
	.w8(32'h3b9d071b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a322606),
	.w1(32'h3c04b190),
	.w2(32'h3bc5d14e),
	.w3(32'h3bf8aed4),
	.w4(32'h3b91ab81),
	.w5(32'hb92b01fe),
	.w6(32'hbab5524e),
	.w7(32'hbbaf6620),
	.w8(32'hbbe7b731),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb62cc5),
	.w1(32'h3af961ad),
	.w2(32'hba4d7058),
	.w3(32'hbb2c7255),
	.w4(32'hbb77820a),
	.w5(32'h3b26c98a),
	.w6(32'h3b20e5ba),
	.w7(32'hbb54f006),
	.w8(32'hbbb7c8fd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc672c6),
	.w1(32'h3ae83bd8),
	.w2(32'h3c42d32a),
	.w3(32'h3b2df11b),
	.w4(32'h3b4a3c2a),
	.w5(32'h3c8d413b),
	.w6(32'h393bec4c),
	.w7(32'hbabacb02),
	.w8(32'h3c0c9423),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6575c1),
	.w1(32'hbc137b59),
	.w2(32'hba120625),
	.w3(32'h3c064118),
	.w4(32'h3b6463b6),
	.w5(32'h3c61a9b9),
	.w6(32'h3c239a13),
	.w7(32'h3b218b11),
	.w8(32'hbb6952eb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe3258),
	.w1(32'hb8f15fc0),
	.w2(32'h3b621655),
	.w3(32'h3b32b5ca),
	.w4(32'hbb2d54af),
	.w5(32'h3b1b7708),
	.w6(32'hba536564),
	.w7(32'h3b30cd7a),
	.w8(32'h39468630),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe1106),
	.w1(32'h3c248623),
	.w2(32'hbbd770c3),
	.w3(32'hbb9787da),
	.w4(32'hbbead5ff),
	.w5(32'hbc98a142),
	.w6(32'hbb1772af),
	.w7(32'hbc0d276a),
	.w8(32'hbc1f8a36),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73ca8f),
	.w1(32'hbcb22382),
	.w2(32'hbd295833),
	.w3(32'hbbe96b9f),
	.w4(32'hbcc858b2),
	.w5(32'h3c756db3),
	.w6(32'h3c0159a4),
	.w7(32'h3bc051a7),
	.w8(32'h3d4f55e6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43745f),
	.w1(32'hbbadf2d2),
	.w2(32'hbb083d2c),
	.w3(32'h3bf327f5),
	.w4(32'hbbbacb4e),
	.w5(32'h3b5a195b),
	.w6(32'h3c518265),
	.w7(32'hbc445791),
	.w8(32'hbb9be927),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987427),
	.w1(32'h3bf2cf52),
	.w2(32'h3aeea568),
	.w3(32'h3bf41600),
	.w4(32'h3b9ee0a2),
	.w5(32'hbb9da051),
	.w6(32'h3ad804fa),
	.w7(32'hba988b41),
	.w8(32'hbac901d1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0617ba),
	.w1(32'hba19b167),
	.w2(32'hbc7098b9),
	.w3(32'hbadfa3ba),
	.w4(32'h3c0ac582),
	.w5(32'hbbd5bada),
	.w6(32'hba8b60ce),
	.w7(32'hbba26d38),
	.w8(32'hbb92a129),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe536e1),
	.w1(32'h3c62a480),
	.w2(32'h3cefe53d),
	.w3(32'h3c2abf9d),
	.w4(32'h3ca7b9f8),
	.w5(32'h3d181125),
	.w6(32'h3c3fe90e),
	.w7(32'h3c974417),
	.w8(32'h3cb5fa6a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0d1fd),
	.w1(32'hb9536aa1),
	.w2(32'hbba51110),
	.w3(32'h3cb870f8),
	.w4(32'hbbf2d06b),
	.w5(32'h3a8776bf),
	.w6(32'h3c0f727e),
	.w7(32'hbc1dd7fe),
	.w8(32'hbc6a6365),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f3c2f),
	.w1(32'h3c153a0d),
	.w2(32'hbca11f00),
	.w3(32'hbbdcf321),
	.w4(32'h3bab39e5),
	.w5(32'hbc970a54),
	.w6(32'hbb587cd3),
	.w7(32'hbc2fdee4),
	.w8(32'hbca38f3f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb86ad5),
	.w1(32'h3afc74ea),
	.w2(32'hba1fac66),
	.w3(32'h3b227e62),
	.w4(32'h3b128cdc),
	.w5(32'hbab4b040),
	.w6(32'h3bbda2fd),
	.w7(32'h3bd577dd),
	.w8(32'h3bbd2ebd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86a362),
	.w1(32'h3a69a0e1),
	.w2(32'h3b9c4f61),
	.w3(32'h3bc8dcb3),
	.w4(32'hbb47594e),
	.w5(32'hbb2aaeb3),
	.w6(32'h3aa7a4d7),
	.w7(32'h3b3b360e),
	.w8(32'h3a5ae80a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc9d0e),
	.w1(32'h3b27197b),
	.w2(32'hbaf10f6b),
	.w3(32'hba5d2d42),
	.w4(32'h39a20d88),
	.w5(32'hbbb94419),
	.w6(32'h38adc875),
	.w7(32'hbc2982ce),
	.w8(32'hbbf97afd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc823c06),
	.w1(32'h3b86264c),
	.w2(32'h3ad5972a),
	.w3(32'hbc0a3e95),
	.w4(32'h3bf12b8d),
	.w5(32'h3a9f9734),
	.w6(32'h3bd4145f),
	.w7(32'hbacbbf81),
	.w8(32'h3b77733e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7a729),
	.w1(32'h399cfa7a),
	.w2(32'h3b7ad06b),
	.w3(32'hbb8f9418),
	.w4(32'h3c093b75),
	.w5(32'h3cf55353),
	.w6(32'h3becd984),
	.w7(32'h3c34af02),
	.w8(32'h3c4cd67e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac97b8c),
	.w1(32'hbc747502),
	.w2(32'hbc2318fa),
	.w3(32'h3c1760fb),
	.w4(32'hbc874330),
	.w5(32'h3d181d02),
	.w6(32'h3b49af2b),
	.w7(32'hbaafaa7a),
	.w8(32'h3cd5fba3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba700488),
	.w1(32'hbaa55bac),
	.w2(32'hbad9c56c),
	.w3(32'h3c01a4b8),
	.w4(32'h3bd48f11),
	.w5(32'h3ba4bc34),
	.w6(32'h3b84316c),
	.w7(32'hbaad5dde),
	.w8(32'hbb49b85f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9ceb6),
	.w1(32'h3bdea352),
	.w2(32'h3a429e8b),
	.w3(32'hbbe72a8e),
	.w4(32'hbbbb7b92),
	.w5(32'hbbb99f67),
	.w6(32'hbb76a42b),
	.w7(32'hbc26c59c),
	.w8(32'hbc02907d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5af62),
	.w1(32'hbafe6b0a),
	.w2(32'h3b916611),
	.w3(32'hbc1fb320),
	.w4(32'hba5ea601),
	.w5(32'h3b2d39d8),
	.w6(32'hbb21040d),
	.w7(32'h3b72db88),
	.w8(32'h3bde0ca3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38267a),
	.w1(32'hbbc07d33),
	.w2(32'hbc149fcb),
	.w3(32'h3b65815e),
	.w4(32'hbaecb453),
	.w5(32'h3b8d1ff7),
	.w6(32'h3b53eb0c),
	.w7(32'h3bcf2b99),
	.w8(32'h3c31db84),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc310835),
	.w1(32'h3bac9670),
	.w2(32'h3ba48558),
	.w3(32'hba91da28),
	.w4(32'h3b79d560),
	.w5(32'h3d03e2a3),
	.w6(32'h3ab3e2ec),
	.w7(32'h3c6c6f85),
	.w8(32'h3cf08273),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941292),
	.w1(32'h3c4531a7),
	.w2(32'h3c109abe),
	.w3(32'h3c3a5ffe),
	.w4(32'h3b46aa1a),
	.w5(32'h3ca5a475),
	.w6(32'h3c2d8c87),
	.w7(32'h3b98bc43),
	.w8(32'h3c11a8fc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54ac7e),
	.w1(32'h3b4176fb),
	.w2(32'h3bd59a79),
	.w3(32'h3c038f94),
	.w4(32'h3aa31ecf),
	.w5(32'hbb3c2123),
	.w6(32'h3b517808),
	.w7(32'hb9c64e45),
	.w8(32'hb9c5b858),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07835f),
	.w1(32'hba7cf0e8),
	.w2(32'h3b9ab37b),
	.w3(32'h3b2eb2a3),
	.w4(32'h3c03724e),
	.w5(32'h3bb2ed94),
	.w6(32'h3bbe00ca),
	.w7(32'h3c0c8560),
	.w8(32'h3c105bbd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7eb97),
	.w1(32'h3b0cd301),
	.w2(32'hbbbd55f7),
	.w3(32'h3a8a7b38),
	.w4(32'hbc283434),
	.w5(32'hbbb36070),
	.w6(32'h3bc64d4e),
	.w7(32'hba782da4),
	.w8(32'h3b7e32d2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c2010),
	.w1(32'h3c29777e),
	.w2(32'h3cb719d2),
	.w3(32'hbbc894f8),
	.w4(32'h3bf91a40),
	.w5(32'h3d078603),
	.w6(32'h3badc612),
	.w7(32'h3c75de9a),
	.w8(32'h3ccab7a6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72c9ee),
	.w1(32'h3b484aa6),
	.w2(32'h3c34ad7d),
	.w3(32'h3c8fdbfe),
	.w4(32'hbbfba088),
	.w5(32'h3d000f45),
	.w6(32'h3cdf42f4),
	.w7(32'h3bdac2b3),
	.w8(32'h3caad2f1),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce6481f),
	.w1(32'h3be53d3a),
	.w2(32'h3be7274a),
	.w3(32'h3c832087),
	.w4(32'h3c463f29),
	.w5(32'h3cbb3073),
	.w6(32'hbc7377ea),
	.w7(32'h3bc5ee3e),
	.w8(32'h3be1f4a6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5c505),
	.w1(32'hbbd41e45),
	.w2(32'h3b05cfd2),
	.w3(32'h3ac860bf),
	.w4(32'hbc3e24b6),
	.w5(32'hba8bcb95),
	.w6(32'h3b7e01bc),
	.w7(32'hbcbf448f),
	.w8(32'hbc80deaa),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31ecf1),
	.w1(32'hba9beca0),
	.w2(32'hb8cef7c5),
	.w3(32'hbb39e51f),
	.w4(32'h3a8b6862),
	.w5(32'h3b28426b),
	.w6(32'hbc01d22f),
	.w7(32'hb9e8c0d2),
	.w8(32'h3bfbcd02),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb078a86),
	.w1(32'h3aefcf50),
	.w2(32'hbbc3302e),
	.w3(32'h3c00aaa2),
	.w4(32'hbb7f6675),
	.w5(32'h3c3d00ba),
	.w6(32'h3b403427),
	.w7(32'h3bceff11),
	.w8(32'h3c8a2b75),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc961ca),
	.w1(32'hbc4c45cf),
	.w2(32'h3a40d32d),
	.w3(32'h3c73ae8f),
	.w4(32'hbc64b56c),
	.w5(32'hbc831f1f),
	.w6(32'h3bef03de),
	.w7(32'hbba018e2),
	.w8(32'hbb5de8a6),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b459a66),
	.w1(32'h3b62ff6a),
	.w2(32'hbb1c2c9e),
	.w3(32'hbc285eb1),
	.w4(32'h3c162545),
	.w5(32'hba20ba22),
	.w6(32'hbc045779),
	.w7(32'hbadf4bd9),
	.w8(32'hbb3c73e2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0148bd),
	.w1(32'hbb4d4ee5),
	.w2(32'hbbef5bbb),
	.w3(32'h3bfd4d46),
	.w4(32'hbaedd671),
	.w5(32'h3a5da325),
	.w6(32'h3c42e5da),
	.w7(32'hba63fc51),
	.w8(32'h3bc7bb1e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d108d),
	.w1(32'hbb152741),
	.w2(32'h3b3a661b),
	.w3(32'h3b5e5668),
	.w4(32'hbc4cb2d2),
	.w5(32'hbc180bd6),
	.w6(32'h3c1ee809),
	.w7(32'hba95fcb9),
	.w8(32'h3b3cb1c6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c097d3e),
	.w1(32'hbc16c8ab),
	.w2(32'hbbbcc95e),
	.w3(32'h3adb172e),
	.w4(32'hbb8e6684),
	.w5(32'hbb38f2ff),
	.w6(32'h3bd970a2),
	.w7(32'h394fbef6),
	.w8(32'hbb043216),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37a4a9),
	.w1(32'h3b046a8e),
	.w2(32'h3aee535d),
	.w3(32'h39856701),
	.w4(32'hbb8cac1a),
	.w5(32'h3be2fa36),
	.w6(32'h3aed593c),
	.w7(32'hbb855582),
	.w8(32'h3c08ff08),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e23a2),
	.w1(32'h3b0b5d66),
	.w2(32'h3c076744),
	.w3(32'h3aea3e47),
	.w4(32'hbac6df81),
	.w5(32'hbae7bcfa),
	.w6(32'hbaa903f4),
	.w7(32'h39a506d8),
	.w8(32'h3ba1141a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f17123),
	.w1(32'hbb0110ad),
	.w2(32'hbbe7c061),
	.w3(32'hbaec4f36),
	.w4(32'h3ba9ffbd),
	.w5(32'h3bcd2a82),
	.w6(32'h3b884987),
	.w7(32'h3bce06c6),
	.w8(32'h3c0ecfb2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0af53),
	.w1(32'h3ba01510),
	.w2(32'h3bbed6f3),
	.w3(32'h3a0e48f2),
	.w4(32'h3b8c578a),
	.w5(32'h3b9a9e86),
	.w6(32'hbb0a41ef),
	.w7(32'hbb91ca87),
	.w8(32'h3b8f0012),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92c42a),
	.w1(32'h3a3c2ba6),
	.w2(32'hbb113e45),
	.w3(32'h3af26de7),
	.w4(32'hba9fecf1),
	.w5(32'h390d0053),
	.w6(32'h3c22d561),
	.w7(32'hba912288),
	.w8(32'h3a32d574),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af939cb),
	.w1(32'hbc095ef6),
	.w2(32'hbbeb7681),
	.w3(32'hb58335f9),
	.w4(32'hbbfd2e72),
	.w5(32'hba25f4ca),
	.w6(32'h3b62ff03),
	.w7(32'hbb0a5a6d),
	.w8(32'h3b91ec02),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fdbf8),
	.w1(32'h3bd90c68),
	.w2(32'h3ba77e79),
	.w3(32'h3b1c485f),
	.w4(32'h3bedb805),
	.w5(32'h3bf31918),
	.w6(32'h3c0bac52),
	.w7(32'hbbd4b0fd),
	.w8(32'hbbe85470),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74ee07),
	.w1(32'h39b29a93),
	.w2(32'hba9e659e),
	.w3(32'h3b0d8f40),
	.w4(32'h3bcad3e1),
	.w5(32'hbb8c1569),
	.w6(32'hba74c3f4),
	.w7(32'h3b027c62),
	.w8(32'hbb57b342),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9bd2b),
	.w1(32'h3c552276),
	.w2(32'h3c0b0468),
	.w3(32'hbb32804b),
	.w4(32'h3c1ab485),
	.w5(32'h3af91597),
	.w6(32'hbb92bcda),
	.w7(32'h39c043a5),
	.w8(32'hbb88a678),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25f5b7),
	.w1(32'hbaeabd36),
	.w2(32'h3af4c3cf),
	.w3(32'hbb108965),
	.w4(32'h3b0b0942),
	.w5(32'h3b640bb8),
	.w6(32'h3b8600d0),
	.w7(32'hbbba0e07),
	.w8(32'hbbf4dc24),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79b524),
	.w1(32'h3a173a45),
	.w2(32'hb8ca1d71),
	.w3(32'hba74987f),
	.w4(32'hbb0a74d9),
	.w5(32'hbba9ed47),
	.w6(32'hbb090349),
	.w7(32'h3a14a32a),
	.w8(32'hba4394df),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8ebeb),
	.w1(32'hbbe91836),
	.w2(32'hbae4ed93),
	.w3(32'hbc3b55a7),
	.w4(32'hbb0cf8ce),
	.w5(32'h3b3697af),
	.w6(32'hbb03bdde),
	.w7(32'h3a311806),
	.w8(32'h3abd1c9a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c98ad),
	.w1(32'h3aa7283d),
	.w2(32'hb8b85278),
	.w3(32'h3b77fe94),
	.w4(32'hbb624bc0),
	.w5(32'hbb2d28b1),
	.w6(32'hbb2b847d),
	.w7(32'hb9df61eb),
	.w8(32'h3b1199c6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba914701),
	.w1(32'h3cb4cdbe),
	.w2(32'hbc08ac6a),
	.w3(32'hbb5d9b44),
	.w4(32'h3c588b9b),
	.w5(32'hbc5ddac8),
	.w6(32'h3b699d39),
	.w7(32'hba7b98eb),
	.w8(32'hbc0c67a9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9010e7),
	.w1(32'h3b70db24),
	.w2(32'h3c14d6f6),
	.w3(32'h3c0f03c7),
	.w4(32'hb9664124),
	.w5(32'h3b1d6ffa),
	.w6(32'h3c9f6dbf),
	.w7(32'h3bda0025),
	.w8(32'h3b839d37),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b548833),
	.w1(32'hb9a22a35),
	.w2(32'hbaddcf43),
	.w3(32'hbb3d32a6),
	.w4(32'h37f06dd2),
	.w5(32'h3a423d44),
	.w6(32'hbb038039),
	.w7(32'hbb90c475),
	.w8(32'hbbf1f115),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96c689),
	.w1(32'hbc4e918b),
	.w2(32'hbcdaae58),
	.w3(32'hb9f1b11b),
	.w4(32'hbd210e5a),
	.w5(32'hbd837b65),
	.w6(32'h3ba06edf),
	.w7(32'hbcb964a0),
	.w8(32'hbcec3d26),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcceb0b8),
	.w1(32'hbb1af168),
	.w2(32'h3b8894cb),
	.w3(32'hbd31a1e0),
	.w4(32'hbb83b512),
	.w5(32'h3c8c4b99),
	.w6(32'hbcbd0d35),
	.w7(32'h39feaab9),
	.w8(32'h3c77f4d5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b802d17),
	.w1(32'hbced2dd9),
	.w2(32'hbcd9adb9),
	.w3(32'h3c0aa5bb),
	.w4(32'hbc9749e8),
	.w5(32'hbba54496),
	.w6(32'h3ad33da0),
	.w7(32'hbbab627c),
	.w8(32'hbaec05b6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc420c15),
	.w1(32'hbb25c7d9),
	.w2(32'hbc4f49fd),
	.w3(32'h3bad4f05),
	.w4(32'hba6d6338),
	.w5(32'hbbe33783),
	.w6(32'h3b71cd7e),
	.w7(32'h3bc98652),
	.w8(32'h3aa4ea7f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f9dfa),
	.w1(32'h3acf9366),
	.w2(32'hbb0f7ba4),
	.w3(32'hbbe84fe5),
	.w4(32'h3ac8b860),
	.w5(32'hbb620dff),
	.w6(32'hbbc1cf78),
	.w7(32'hbc1d29d6),
	.w8(32'hbc0fae4c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d02145),
	.w1(32'h3ac03747),
	.w2(32'h3b995156),
	.w3(32'h3bb50775),
	.w4(32'h39ed3b3a),
	.w5(32'hb9a3716a),
	.w6(32'h3bd26de5),
	.w7(32'h3b16beab),
	.w8(32'hbb3e1888),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94810a),
	.w1(32'h3ae63733),
	.w2(32'h3d1739a0),
	.w3(32'h3b638676),
	.w4(32'h3adec429),
	.w5(32'hbb2b1525),
	.w6(32'hbb36eb59),
	.w7(32'hbc8cedac),
	.w8(32'hbccb82a8),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb44d),
	.w1(32'hbba68925),
	.w2(32'hbc069479),
	.w3(32'hbc20e892),
	.w4(32'h3bf8423a),
	.w5(32'hbbcec03b),
	.w6(32'hba09cd35),
	.w7(32'hba1cc95b),
	.w8(32'hbc546263),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4de125),
	.w1(32'h3a7ed69a),
	.w2(32'h3b00d372),
	.w3(32'h3bbd5113),
	.w4(32'hbb5b3003),
	.w5(32'h3c6d5996),
	.w6(32'h38b55ceb),
	.w7(32'h3ac5a33f),
	.w8(32'h3c809d03),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2ab93),
	.w1(32'h3b868810),
	.w2(32'h3c21229d),
	.w3(32'h3c426648),
	.w4(32'h3a162137),
	.w5(32'hbbe6554b),
	.w6(32'h3c1d2216),
	.w7(32'h3b942a2a),
	.w8(32'hba880769),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfadc2a),
	.w1(32'h3be1215a),
	.w2(32'h3bd13f65),
	.w3(32'h3b61a00d),
	.w4(32'hba604049),
	.w5(32'h3c216188),
	.w6(32'h3b0cb7c0),
	.w7(32'h3b93834a),
	.w8(32'h3bef058a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20702d),
	.w1(32'hba6d0cd9),
	.w2(32'hbaecb13b),
	.w3(32'h3a8053a2),
	.w4(32'hbbcaa9b0),
	.w5(32'h3b931dff),
	.w6(32'hba6a8921),
	.w7(32'hbb860bb5),
	.w8(32'hbaeb7adc),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cc41e),
	.w1(32'h3c1534b1),
	.w2(32'h3c06e392),
	.w3(32'h3ade7c6f),
	.w4(32'h3ba6f4eb),
	.w5(32'h3c860e0e),
	.w6(32'h3b914eb6),
	.w7(32'h3b4dba04),
	.w8(32'h3c4313d3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85ba0c),
	.w1(32'h3c18224d),
	.w2(32'h3b9d1781),
	.w3(32'h3b0921be),
	.w4(32'h3b3d06a0),
	.w5(32'h3b333e5d),
	.w6(32'h3b63f234),
	.w7(32'h3b72df0f),
	.w8(32'hbb83ee4e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb9ebd),
	.w1(32'hbb89ec28),
	.w2(32'h3b61e7b0),
	.w3(32'h3b990443),
	.w4(32'h391686dc),
	.w5(32'h3c2a3e5e),
	.w6(32'h3abb602c),
	.w7(32'h3c2fd03e),
	.w8(32'h3c6e64d3),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2395ed),
	.w1(32'h3b21b592),
	.w2(32'hbc95fe31),
	.w3(32'hb9d0a774),
	.w4(32'h39e6f4dc),
	.w5(32'hbcead77d),
	.w6(32'hbbe8772a),
	.w7(32'hbc92f1bf),
	.w8(32'hbcb7ae63),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d7150),
	.w1(32'h3b946ff0),
	.w2(32'h3ba30d4d),
	.w3(32'hbb31e287),
	.w4(32'h38aa1dab),
	.w5(32'h3aaf68a1),
	.w6(32'h3b900555),
	.w7(32'hbb38dba9),
	.w8(32'h3b00353d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30ba3a),
	.w1(32'hba9e5824),
	.w2(32'hbac43c12),
	.w3(32'h3a839f29),
	.w4(32'hbbc51259),
	.w5(32'hbae8e58a),
	.w6(32'hbb9b0e64),
	.w7(32'hbaff6ed0),
	.w8(32'h3ba213f6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fdf220),
	.w1(32'h3bf67341),
	.w2(32'h3bebd7f6),
	.w3(32'hbb982493),
	.w4(32'hbbf9d456),
	.w5(32'hbbf23049),
	.w6(32'h3b3370a1),
	.w7(32'hbc59339a),
	.w8(32'hbc8fb42c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef0621),
	.w1(32'hbc176b01),
	.w2(32'hbc6bd279),
	.w3(32'hbbb9336b),
	.w4(32'hbca01d0c),
	.w5(32'hbcd71ba6),
	.w6(32'hbc095ca4),
	.w7(32'hbbf94443),
	.w8(32'hbc4fb2b6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6eadcb),
	.w1(32'h3b365830),
	.w2(32'h39a973de),
	.w3(32'hbc5c95bc),
	.w4(32'hbbbd41e0),
	.w5(32'hbbb17420),
	.w6(32'hbc48b3b0),
	.w7(32'h3bc7d570),
	.w8(32'h3bc54602),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52adba),
	.w1(32'hbcdff5e9),
	.w2(32'hbc8ebac5),
	.w3(32'h3b93e4b6),
	.w4(32'hbc74caee),
	.w5(32'h3c2da7da),
	.w6(32'h3b218b5b),
	.w7(32'h3ac544f0),
	.w8(32'h3c887204),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd97866),
	.w1(32'hb9db852f),
	.w2(32'h3b4cb398),
	.w3(32'h3c1e8c41),
	.w4(32'hba422a0a),
	.w5(32'h3b975c13),
	.w6(32'hbbe8b893),
	.w7(32'hbbfcc23b),
	.w8(32'hbb85d5e8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67e7ea),
	.w1(32'hbbccb125),
	.w2(32'h3a01d309),
	.w3(32'h3acd3e57),
	.w4(32'hbbf0b659),
	.w5(32'h3a293ceb),
	.w6(32'hbba4f564),
	.w7(32'hbaf5561e),
	.w8(32'hbb9db483),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f3333),
	.w1(32'hbb6346e0),
	.w2(32'h3b89d045),
	.w3(32'h3a1611bf),
	.w4(32'h3b2f3687),
	.w5(32'h3b7a4082),
	.w6(32'hb984040f),
	.w7(32'h3af28ff9),
	.w8(32'h3bea4bd8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d99cf),
	.w1(32'h3ae5f5d5),
	.w2(32'h3bc2a81a),
	.w3(32'hba0b5ae3),
	.w4(32'h3ab8ec99),
	.w5(32'h3c0ce349),
	.w6(32'hb9ca9d05),
	.w7(32'h3c095bd5),
	.w8(32'h3c3e3876),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04a1a5),
	.w1(32'h3b5ffd2a),
	.w2(32'h3b6c377c),
	.w3(32'h3b78e653),
	.w4(32'h3c0becfe),
	.w5(32'h3b00ad1b),
	.w6(32'h3b888fbc),
	.w7(32'hbb7305b5),
	.w8(32'hbc1d8df4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49f066),
	.w1(32'hbba749b0),
	.w2(32'hbc67d6de),
	.w3(32'hbb8a1866),
	.w4(32'hba5bb6fb),
	.w5(32'hbc1a8436),
	.w6(32'hb9efa4a1),
	.w7(32'hbc1169f5),
	.w8(32'hbbf5abb6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86d51e),
	.w1(32'h3ad54e39),
	.w2(32'h3b74a3a2),
	.w3(32'hbacc84ca),
	.w4(32'h3c06b148),
	.w5(32'h3c2fa96b),
	.w6(32'h3c5741f0),
	.w7(32'h3b15f430),
	.w8(32'h3b96e700),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049516),
	.w1(32'h3b2d9730),
	.w2(32'h3bac70fb),
	.w3(32'hbb4f2920),
	.w4(32'hbb09479c),
	.w5(32'hbbbcf62a),
	.w6(32'hbbb77163),
	.w7(32'hbbea9bf6),
	.w8(32'hbb8bb338),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb64175),
	.w1(32'h3b8484a2),
	.w2(32'h3c385c50),
	.w3(32'hbae9a2e9),
	.w4(32'hba996f29),
	.w5(32'h3b7a4c2f),
	.w6(32'h3b21ae67),
	.w7(32'hbb06e3e6),
	.w8(32'hbaa04e93),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ccef8),
	.w1(32'hb8de1ab7),
	.w2(32'h3a41a6c0),
	.w3(32'h3a4ff362),
	.w4(32'hba9f15ac),
	.w5(32'hb9cdb324),
	.w6(32'hbbdaff04),
	.w7(32'hbba3fd36),
	.w8(32'hbb98d91f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2ade0),
	.w1(32'hbc08a6c3),
	.w2(32'hbba42a2f),
	.w3(32'h3b9baa0d),
	.w4(32'h3b0965a4),
	.w5(32'h3c48d138),
	.w6(32'h3b646965),
	.w7(32'hba5df972),
	.w8(32'hbb662872),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc174ac0),
	.w1(32'hbb90a144),
	.w2(32'hbc18f9a5),
	.w3(32'hbbc852fb),
	.w4(32'hbb2204f3),
	.w5(32'h3b645f01),
	.w6(32'hbc85fe0b),
	.w7(32'h3a0a9dd5),
	.w8(32'h399d17a8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf24bc),
	.w1(32'hbb7e5fa2),
	.w2(32'hbb7716a8),
	.w3(32'h3b41b02e),
	.w4(32'hbbb04f3e),
	.w5(32'h3ad85e3b),
	.w6(32'hbb1fff68),
	.w7(32'h3b588877),
	.w8(32'h3b833d59),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af47e93),
	.w1(32'h3b2c705b),
	.w2(32'h3bbb1db6),
	.w3(32'h3aff16cd),
	.w4(32'hbaffe1ab),
	.w5(32'h3af06459),
	.w6(32'hb905d3c4),
	.w7(32'hbab88028),
	.w8(32'h3b2ed30b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5d13c),
	.w1(32'h398db730),
	.w2(32'h3a50997e),
	.w3(32'h3a371cea),
	.w4(32'hb9cddf8c),
	.w5(32'h38f47c39),
	.w6(32'h38ee3242),
	.w7(32'hb8967e92),
	.w8(32'h39532d1d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a96912),
	.w1(32'hb82bf001),
	.w2(32'hb89fec60),
	.w3(32'hb838b907),
	.w4(32'hb60c97ae),
	.w5(32'hb805f20a),
	.w6(32'hb8374b56),
	.w7(32'hb6e0646f),
	.w8(32'hb826e31d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93acd8),
	.w1(32'h3a876940),
	.w2(32'h399fb8bb),
	.w3(32'h3a2f7949),
	.w4(32'h38af6b4d),
	.w5(32'hb9da850d),
	.w6(32'h396510a2),
	.w7(32'hb99a054d),
	.w8(32'hb93a00d1),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9212ada),
	.w1(32'hb8b3d7c7),
	.w2(32'hb9272e7c),
	.w3(32'hb8839a1c),
	.w4(32'h3708da39),
	.w5(32'hb88de84f),
	.w6(32'hb8ddabb7),
	.w7(32'hb6b6e29f),
	.w8(32'hb8d92f67),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb691ec),
	.w1(32'h3b937e7f),
	.w2(32'h3bd353b6),
	.w3(32'h3a935257),
	.w4(32'hb939b508),
	.w5(32'h3b1e968f),
	.w6(32'h3a51867b),
	.w7(32'hb95e341d),
	.w8(32'h3b2b8cd2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfab4ca),
	.w1(32'h3ae3bcd8),
	.w2(32'h3b21be70),
	.w3(32'h3bcdf0a4),
	.w4(32'hb9ca672a),
	.w5(32'h39cec2c4),
	.w6(32'h3bae8160),
	.w7(32'hba320ecc),
	.w8(32'hb94f762b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e1443),
	.w1(32'h3ae11fb5),
	.w2(32'h3b6ad96b),
	.w3(32'h3b250b79),
	.w4(32'hba377bcc),
	.w5(32'h3a9eadd8),
	.w6(32'h3ac21ec9),
	.w7(32'hbaa7a411),
	.w8(32'h3aaa8528),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00c57a),
	.w1(32'hbaae014a),
	.w2(32'hba03d212),
	.w3(32'hb9ab88bd),
	.w4(32'hba86d763),
	.w5(32'hb9bac0a5),
	.w6(32'h39e3e920),
	.w7(32'hba0ace51),
	.w8(32'hb9ca9236),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf34d9),
	.w1(32'h3b186919),
	.w2(32'h3b933244),
	.w3(32'h3b489bfc),
	.w4(32'hba4f60cf),
	.w5(32'h3a56c587),
	.w6(32'h3ac08d58),
	.w7(32'hbb13816d),
	.w8(32'h39709889),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2129ac),
	.w1(32'h3ab9ecb9),
	.w2(32'h3b3ee2c8),
	.w3(32'h3a60ec65),
	.w4(32'hba1c9eb2),
	.w5(32'h39a71fc4),
	.w6(32'h3a21a506),
	.w7(32'hba6a7ad4),
	.w8(32'h3a324da8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a22f1),
	.w1(32'h3b000c5c),
	.w2(32'h3ba53bf7),
	.w3(32'hba543f4b),
	.w4(32'hbb383a31),
	.w5(32'hb8c76dac),
	.w6(32'hbacd6de2),
	.w7(32'hbb02686b),
	.w8(32'h3a8f79da),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fd9fb),
	.w1(32'hb6347151),
	.w2(32'hb829d252),
	.w3(32'hb7dda080),
	.w4(32'h369260ec),
	.w5(32'hb80a23f3),
	.w6(32'hb7e6397b),
	.w7(32'hb70a7064),
	.w8(32'hb7ffaf83),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81034b1),
	.w1(32'hb7c3fb88),
	.w2(32'h3793742c),
	.w3(32'h38093675),
	.w4(32'hb73c7f8c),
	.w5(32'h388cc563),
	.w6(32'h388d01c9),
	.w7(32'hb587b27f),
	.w8(32'h38115efc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac8300),
	.w1(32'h3ae8fcfb),
	.w2(32'h3b56119d),
	.w3(32'h390e83fa),
	.w4(32'hbafbde0b),
	.w5(32'h39c7f97a),
	.w6(32'h3b41433c),
	.w7(32'h3a1af170),
	.w8(32'h3b0fb9b1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf48c27),
	.w1(32'h3ba60774),
	.w2(32'h3be4ae6a),
	.w3(32'h3b2efb9e),
	.w4(32'hba8ccfb8),
	.w5(32'h3b34702c),
	.w6(32'h3b86ca3d),
	.w7(32'h3abadb5f),
	.w8(32'h3b9354b6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0f968),
	.w1(32'h3b59e643),
	.w2(32'h3b9e3e0b),
	.w3(32'h3b1dafd1),
	.w4(32'hba3fa8a2),
	.w5(32'h39815f08),
	.w6(32'h3b083f9b),
	.w7(32'hba92546b),
	.w8(32'h39d452b3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a803b3),
	.w1(32'h3b00b902),
	.w2(32'h3b1af993),
	.w3(32'hb9a9b402),
	.w4(32'h3a1034dc),
	.w5(32'h39e5b170),
	.w6(32'hba971a2c),
	.w7(32'hb9a2f578),
	.w8(32'h3b17a406),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e075bb),
	.w1(32'h39017913),
	.w2(32'h383036d6),
	.w3(32'hb80b0a2b),
	.w4(32'h38896dd3),
	.w5(32'h3914ac72),
	.w6(32'h378697ce),
	.w7(32'h39307d51),
	.w8(32'h391608c3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a003cd8),
	.w1(32'h3a1d3717),
	.w2(32'h39e45ff9),
	.w3(32'h389aed42),
	.w4(32'h387b288b),
	.w5(32'h393969e9),
	.w6(32'h3905be6c),
	.w7(32'h3990935d),
	.w8(32'h39a91374),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bca76),
	.w1(32'hbaa31763),
	.w2(32'h3b5e0cde),
	.w3(32'hbaaff98c),
	.w4(32'hba82808d),
	.w5(32'h3b86baab),
	.w6(32'hb9288dba),
	.w7(32'hba0dffa8),
	.w8(32'h3b8ddd48),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b634821),
	.w1(32'h3b24b364),
	.w2(32'h3b571df4),
	.w3(32'hbacae873),
	.w4(32'hba99bbf7),
	.w5(32'h3a5b8c89),
	.w6(32'h3921c231),
	.w7(32'h3a516e3d),
	.w8(32'h3b4a7b38),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c314c),
	.w1(32'h3b1e3f44),
	.w2(32'h3b44c81a),
	.w3(32'h3a291a67),
	.w4(32'hb99842a8),
	.w5(32'h3a52732c),
	.w6(32'h39f6bdda),
	.w7(32'h3a216ff8),
	.w8(32'h3aeea206),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdf9b2),
	.w1(32'hbad2ab7f),
	.w2(32'h3a00690f),
	.w3(32'h3aebbbd1),
	.w4(32'hbaed166a),
	.w5(32'hb999d1e3),
	.w6(32'h3b0673a4),
	.w7(32'hbb138a1b),
	.w8(32'hb87d347a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba53baa),
	.w1(32'h3b0cfce5),
	.w2(32'h3b7c3c5b),
	.w3(32'h3b5da4f0),
	.w4(32'hb9a5dfc3),
	.w5(32'h3a00e526),
	.w6(32'h3b35823a),
	.w7(32'hbaab7ad4),
	.w8(32'h388fa384),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb812de22),
	.w1(32'hb7dec0f1),
	.w2(32'hb80facde),
	.w3(32'hb7b0b1fd),
	.w4(32'hb7211a63),
	.w5(32'hb7894aa4),
	.w6(32'hb7c40458),
	.w7(32'hb75d1c13),
	.w8(32'hb7b796c6),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a79095),
	.w1(32'hb8640819),
	.w2(32'hb89268eb),
	.w3(32'hb889ff5a),
	.w4(32'hb828d02f),
	.w5(32'hb859ae60),
	.w6(32'hb87a7093),
	.w7(32'hb819f7a2),
	.w8(32'hb8562aca),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a580cc),
	.w1(32'h376a316f),
	.w2(32'h3807aae4),
	.w3(32'hba76a0cf),
	.w4(32'hb99cacbf),
	.w5(32'hb80694c2),
	.w6(32'hb8333cd6),
	.w7(32'h3a4e2053),
	.w8(32'h3a0bd7a4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a653a8),
	.w1(32'hb84e988d),
	.w2(32'hb8909816),
	.w3(32'hb868f9e4),
	.w4(32'hb79b3b30),
	.w5(32'hb7e84ae5),
	.w6(32'hb84dbc89),
	.w7(32'hb7c66e21),
	.w8(32'hb807fc27),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fd050a),
	.w1(32'h3a3eb1f3),
	.w2(32'h3a898592),
	.w3(32'hba63a947),
	.w4(32'h39a6a756),
	.w5(32'h3a4340d5),
	.w6(32'h3843987d),
	.w7(32'h3a805efe),
	.w8(32'h3a8b8574),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6ce72),
	.w1(32'h3b2b08ef),
	.w2(32'h3b8b3eb8),
	.w3(32'h3ad71824),
	.w4(32'hba88edf8),
	.w5(32'h3a78ef12),
	.w6(32'h3b2a8b4c),
	.w7(32'h3a156cbe),
	.w8(32'h3b3ae07d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62279f),
	.w1(32'h3ab20bae),
	.w2(32'h3b0e0151),
	.w3(32'h3b18aa07),
	.w4(32'hba124ebc),
	.w5(32'h3a3f4e10),
	.w6(32'h3a9306fa),
	.w7(32'hba561862),
	.w8(32'h3a76b038),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85270af),
	.w1(32'hb82e1d9b),
	.w2(32'hb82cd8f7),
	.w3(32'hb84a434f),
	.w4(32'hb7fe13cc),
	.w5(32'hb8297c88),
	.w6(32'hb7fec863),
	.w7(32'hb8036376),
	.w8(32'hb83e6691),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d890d),
	.w1(32'h3a25e011),
	.w2(32'h3ba9e810),
	.w3(32'hbabd0344),
	.w4(32'hbb5c42e1),
	.w5(32'h3a902111),
	.w6(32'hbac484ee),
	.w7(32'hbaf758a2),
	.w8(32'h3b4a8882),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b319aae),
	.w1(32'h3b16ad82),
	.w2(32'h3b3badad),
	.w3(32'h39ca5623),
	.w4(32'h3a11e7c9),
	.w5(32'h3aa14463),
	.w6(32'h388f06fd),
	.w7(32'h3a8fd08a),
	.w8(32'h3b0c7019),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f21afe),
	.w1(32'h36bbd71b),
	.w2(32'hb8a3f80c),
	.w3(32'h37ec97df),
	.w4(32'h389eeba6),
	.w5(32'hb68b960e),
	.w6(32'h380d73c5),
	.w7(32'h389f2702),
	.w8(32'h378d9bcb),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd495b),
	.w1(32'h3a363d96),
	.w2(32'h3b109434),
	.w3(32'hba90d096),
	.w4(32'hba32ffdf),
	.w5(32'h3a8b086c),
	.w6(32'hba488b5b),
	.w7(32'hb9b24e65),
	.w8(32'h3ac7496e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884f1ce),
	.w1(32'hb88c7c8b),
	.w2(32'hb8a35dbf),
	.w3(32'h370b2e32),
	.w4(32'hb7f4f86f),
	.w5(32'hb80a61c1),
	.w6(32'hb8509c0d),
	.w7(32'hb8cd5268),
	.w8(32'hb8c741fb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dee431),
	.w1(32'h391ba843),
	.w2(32'h39dc9125),
	.w3(32'hb7c9172d),
	.w4(32'hb872fc7c),
	.w5(32'hb88dbdfb),
	.w6(32'h3957fef8),
	.w7(32'h3903b02c),
	.w8(32'h39a462bf),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fc513c),
	.w1(32'hb712d0b3),
	.w2(32'hb80739e0),
	.w3(32'hb76dd7c2),
	.w4(32'h3736d09c),
	.w5(32'hb78e3d15),
	.w6(32'hb77dd264),
	.w7(32'hb65e3290),
	.w8(32'hb7cc0217),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88438d9),
	.w1(32'hb826ec2d),
	.w2(32'hb84c4ad4),
	.w3(32'hb841e5fa),
	.w4(32'hb7eadcd2),
	.w5(32'hb7f8b84b),
	.w6(32'hb8273da7),
	.w7(32'hb7e58b31),
	.w8(32'hb7fa6f63),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c2e3b),
	.w1(32'hba840cae),
	.w2(32'hb92d7271),
	.w3(32'h3a10af8a),
	.w4(32'hba86268e),
	.w5(32'hb921e959),
	.w6(32'h3a9db9fc),
	.w7(32'hba3cebd2),
	.w8(32'h37d5908f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfe193),
	.w1(32'h3bd6212f),
	.w2(32'h3c0e059f),
	.w3(32'h3b2e6370),
	.w4(32'h3adb73f8),
	.w5(32'h3b2b480a),
	.w6(32'h3a58f7ea),
	.w7(32'h39ab8ee4),
	.w8(32'h3b48a12b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4efe00),
	.w1(32'h3b0c359d),
	.w2(32'h3b79cb01),
	.w3(32'h3a1ed18f),
	.w4(32'hb87b9f9c),
	.w5(32'h3a85e428),
	.w6(32'h3a4b3fac),
	.w7(32'h3a0f3f15),
	.w8(32'h3af86115),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b391537),
	.w1(32'h3b579c73),
	.w2(32'h3b94bc02),
	.w3(32'h388a9c5f),
	.w4(32'hb9801385),
	.w5(32'h3a055f3b),
	.w6(32'h396d2d96),
	.w7(32'hba165939),
	.w8(32'h3a899252),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb938acbd),
	.w1(32'hb9506dba),
	.w2(32'hb8f1c3b3),
	.w3(32'hb91f1c77),
	.w4(32'hb948aed5),
	.w5(32'hb9185204),
	.w6(32'hb7812058),
	.w7(32'hb8eb511f),
	.w8(32'hb8929903),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ac1bf),
	.w1(32'h39934632),
	.w2(32'h38c1312c),
	.w3(32'h3826c415),
	.w4(32'hb588ca2f),
	.w5(32'hb8ccb7ea),
	.w6(32'h37236d70),
	.w7(32'h38b6cbd0),
	.w8(32'hb79ada4f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a8b217),
	.w1(32'hb60c8bcc),
	.w2(32'hb7b3b1f4),
	.w3(32'h36aaa6ad),
	.w4(32'h37b31cd9),
	.w5(32'h3640efe2),
	.w6(32'hb683cef8),
	.w7(32'h375fd7af),
	.w8(32'hb6c75114),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb880ac4e),
	.w1(32'hb82138d0),
	.w2(32'hb6857db8),
	.w3(32'hb82c25ba),
	.w4(32'hb7ca3c21),
	.w5(32'hb80efd37),
	.w6(32'hb7dc1bd0),
	.w7(32'h36ce08d4),
	.w8(32'h37985d25),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8a50b),
	.w1(32'h3b49d8c1),
	.w2(32'h3b6c1e59),
	.w3(32'h3b3a9a80),
	.w4(32'h39daf148),
	.w5(32'h3aae2e10),
	.w6(32'h3ac1a37b),
	.w7(32'h393ca7a1),
	.w8(32'h3affc347),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abb21c),
	.w1(32'hb8a0e2d1),
	.w2(32'hb8b7a79e),
	.w3(32'hb84c595f),
	.w4(32'hb7fce0b0),
	.w5(32'hb8458e7f),
	.w6(32'hb886c7de),
	.w7(32'hb806b7e5),
	.w8(32'hb8b3b911),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e8c9c7),
	.w1(32'hba87ee28),
	.w2(32'h3a00902f),
	.w3(32'hb7b7fd18),
	.w4(32'hb9ca00d2),
	.w5(32'h3a053208),
	.w6(32'h3a8f7545),
	.w7(32'h394b7811),
	.w8(32'h3a263b67),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d38d6),
	.w1(32'hb8b52935),
	.w2(32'h39047613),
	.w3(32'h39df3555),
	.w4(32'hb9b03fdf),
	.w5(32'hb9e906a9),
	.w6(32'h39a8c578),
	.w7(32'hb9488fd8),
	.w8(32'hba30b11d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ed0d50),
	.w1(32'hb7bfc8b0),
	.w2(32'hb7b179ed),
	.w3(32'hb78cfe22),
	.w4(32'hb7717dee),
	.w5(32'hb59c101d),
	.w6(32'hb7d29533),
	.w7(32'hb797f617),
	.w8(32'hb72e047f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d81a5),
	.w1(32'h3a5b244c),
	.w2(32'h3a829b96),
	.w3(32'hb9b5194e),
	.w4(32'hba06fbbc),
	.w5(32'hb9d644b8),
	.w6(32'hb9812e7e),
	.w7(32'hb9536f80),
	.w8(32'h383d7aa2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3822b39d),
	.w1(32'h386659ba),
	.w2(32'h38820b3a),
	.w3(32'hb8b3f765),
	.w4(32'hb87c2f8e),
	.w5(32'hb78958cf),
	.w6(32'hb8936d6c),
	.w7(32'h3873840e),
	.w8(32'h38d28466),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b13de),
	.w1(32'h3b8c6ca7),
	.w2(32'h3babadb9),
	.w3(32'h3afba9cd),
	.w4(32'h39550b93),
	.w5(32'hb9ed1a7d),
	.w6(32'h3ae0e3c8),
	.w7(32'hb98e5e05),
	.w8(32'hb81a1fce),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61449f2),
	.w1(32'h3863872f),
	.w2(32'h381bfd27),
	.w3(32'hb7d75abe),
	.w4(32'h37d3ee78),
	.w5(32'h3609fba8),
	.w6(32'h37f5e23a),
	.w7(32'h389b5ed0),
	.w8(32'h35834902),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9808b9),
	.w1(32'hbb3cf8fe),
	.w2(32'hbb2343cf),
	.w3(32'h394cc947),
	.w4(32'hbb4c926d),
	.w5(32'hbb498112),
	.w6(32'h3ba664f3),
	.w7(32'h3a8c4329),
	.w8(32'hba257824),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule