module layer_10_featuremap_182(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8cb1c),
	.w1(32'h395c7b58),
	.w2(32'hb96be165),
	.w3(32'hb96f63d3),
	.w4(32'h3a6d769a),
	.w5(32'h39b3e380),
	.w6(32'h37bbf971),
	.w7(32'h37964402),
	.w8(32'h3a321769),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9100bc),
	.w1(32'h39c73945),
	.w2(32'h39404d57),
	.w3(32'h3a9f3dc9),
	.w4(32'h39036135),
	.w5(32'hb9d18040),
	.w6(32'h3a7b101d),
	.w7(32'h3a215df7),
	.w8(32'hb9993032),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe9cfb),
	.w1(32'hba8db216),
	.w2(32'hba76804e),
	.w3(32'hba184cfa),
	.w4(32'hba9af774),
	.w5(32'hba85113d),
	.w6(32'hba37841a),
	.w7(32'hba2eca96),
	.w8(32'hba3a9cb0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba571750),
	.w1(32'hba61a129),
	.w2(32'hba769a34),
	.w3(32'hba818055),
	.w4(32'hba06d4a8),
	.w5(32'hb9dc202b),
	.w6(32'hb9b4b7f5),
	.w7(32'hb8e5f1c8),
	.w8(32'hb8bf6810),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c41ae),
	.w1(32'h3a3d4218),
	.w2(32'h3a001df9),
	.w3(32'hb9abc0b6),
	.w4(32'h3a3f72b7),
	.w5(32'h39b7c97b),
	.w6(32'h3a2e0da0),
	.w7(32'h39e53275),
	.w8(32'h3a0bb6d0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a333eba),
	.w1(32'hba0e96f7),
	.w2(32'hba2daba9),
	.w3(32'h38888c81),
	.w4(32'hb92750c7),
	.w5(32'hb9e4945d),
	.w6(32'hb97c503f),
	.w7(32'hba0b3099),
	.w8(32'hb9d46e9a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39821846),
	.w1(32'h3a35778d),
	.w2(32'h3849f179),
	.w3(32'h39d7996c),
	.w4(32'h3999d77e),
	.w5(32'hb9af15f1),
	.w6(32'h3a25d3f6),
	.w7(32'h39ab9f26),
	.w8(32'hb9603a0a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa223bc),
	.w1(32'h3a12d856),
	.w2(32'hb9eec19a),
	.w3(32'hbaae7613),
	.w4(32'hba017354),
	.w5(32'hb9a8cdf3),
	.w6(32'hba77b085),
	.w7(32'hb9be5239),
	.w8(32'h3968b66b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75a321),
	.w1(32'hb97971a1),
	.w2(32'hb9f8f737),
	.w3(32'hba396077),
	.w4(32'hb8f66e82),
	.w5(32'hb963c8b8),
	.w6(32'hba5fa186),
	.w7(32'hba1d7a8a),
	.w8(32'hb901096f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb605e),
	.w1(32'hba7ee01f),
	.w2(32'hbab36592),
	.w3(32'hbb17440f),
	.w4(32'hbab9261d),
	.w5(32'hbafb0b8c),
	.w6(32'hba614392),
	.w7(32'hbb04075c),
	.w8(32'hbb1979e1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39196785),
	.w1(32'hba357883),
	.w2(32'hba8bc024),
	.w3(32'hb941943a),
	.w4(32'hba0deb35),
	.w5(32'hb9d5f95d),
	.w6(32'hba34f86c),
	.w7(32'hba3b6d29),
	.w8(32'hba37633b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15838a),
	.w1(32'h3affc59e),
	.w2(32'h3afd379c),
	.w3(32'h395a38b1),
	.w4(32'h3aab7757),
	.w5(32'h3b0c665b),
	.w6(32'h394f0d11),
	.w7(32'h3a1b4ead),
	.w8(32'h3ac4cb69),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafabdfd),
	.w1(32'hbaff9ad1),
	.w2(32'hbab9c2ec),
	.w3(32'hbabd9de1),
	.w4(32'hbafe562d),
	.w5(32'hba8b2ed9),
	.w6(32'hbaa1586d),
	.w7(32'hbb03bdbc),
	.w8(32'hba4b69fb),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e60e23),
	.w1(32'hba5b1e3f),
	.w2(32'hba8a346d),
	.w3(32'h3a31f227),
	.w4(32'hba5e191a),
	.w5(32'hba7f450d),
	.w6(32'h3a23b2ea),
	.w7(32'hba839d69),
	.w8(32'hba673b1b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d98658),
	.w1(32'h3a1c46e4),
	.w2(32'hba0094dc),
	.w3(32'hb99d1563),
	.w4(32'h39926e35),
	.w5(32'hb980eff0),
	.w6(32'hba4d67c1),
	.w7(32'hb9f2b71c),
	.w8(32'hb9a96efb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3755bcc9),
	.w1(32'hbaf7a6f7),
	.w2(32'hbb1524da),
	.w3(32'hba60b02e),
	.w4(32'hbb04f3b7),
	.w5(32'hbb23976e),
	.w6(32'hba711735),
	.w7(32'hbadc09bd),
	.w8(32'hbb02e78d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891ba27),
	.w1(32'hba360085),
	.w2(32'hba585c5a),
	.w3(32'hb986b8cf),
	.w4(32'hb9e066f6),
	.w5(32'hb9d2648d),
	.w6(32'hba45e0e2),
	.w7(32'hba523b6d),
	.w8(32'hba60a448),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcae77),
	.w1(32'hbb2f7d56),
	.w2(32'hbb494a2b),
	.w3(32'hbb13076c),
	.w4(32'hbb0200ab),
	.w5(32'hbaa8c0f6),
	.w6(32'hb9ec880a),
	.w7(32'hba8c090a),
	.w8(32'hbabd6767),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb157340),
	.w1(32'hbb56f4cc),
	.w2(32'hbb3aa228),
	.w3(32'hbb2e50c9),
	.w4(32'hbb508709),
	.w5(32'hbb0310ab),
	.w6(32'hbae48899),
	.w7(32'hbb20dd8b),
	.w8(32'hbad4ba93),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7c924),
	.w1(32'hb953410b),
	.w2(32'hba1ba8f4),
	.w3(32'hba09df92),
	.w4(32'hb926091f),
	.w5(32'hb9e15793),
	.w6(32'hb9324b92),
	.w7(32'hba0ad982),
	.w8(32'hb992c036),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97183d9),
	.w1(32'h38daa85d),
	.w2(32'hb99e05f0),
	.w3(32'hb889fddf),
	.w4(32'h39d8d103),
	.w5(32'hb735d542),
	.w6(32'h39b7ed53),
	.w7(32'h37aac963),
	.w8(32'h39a987fe),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d319a),
	.w1(32'hbb04b203),
	.w2(32'hbaea97a2),
	.w3(32'h393cfa25),
	.w4(32'hbab9fe1f),
	.w5(32'hba8fdb81),
	.w6(32'hbadea676),
	.w7(32'hbaa05393),
	.w8(32'hbabe61aa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0af7f),
	.w1(32'hb9e37a14),
	.w2(32'hbb983a53),
	.w3(32'h39965095),
	.w4(32'hb8032209),
	.w5(32'hbacd4c2b),
	.w6(32'h37b2d5ab),
	.w7(32'hba865c27),
	.w8(32'hba9aabbc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002272),
	.w1(32'hba2d40c0),
	.w2(32'hba61db4b),
	.w3(32'hbab27add),
	.w4(32'hba122dcc),
	.w5(32'hbaa61871),
	.w6(32'hba363a6e),
	.w7(32'hba8212cc),
	.w8(32'hbac13f5a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4c841),
	.w1(32'hba1a8ab9),
	.w2(32'hba753b33),
	.w3(32'hb837a910),
	.w4(32'hb93f7dd7),
	.w5(32'hba8742ea),
	.w6(32'hba0bf78b),
	.w7(32'hb9eaa0ee),
	.w8(32'hba65604c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba443579),
	.w1(32'hb990f144),
	.w2(32'hb9e2940c),
	.w3(32'hb981d85e),
	.w4(32'hb8995e10),
	.w5(32'h3955568b),
	.w6(32'hb978a23f),
	.w7(32'hb8d402d4),
	.w8(32'hb8507c50),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f0811),
	.w1(32'hb8c91335),
	.w2(32'hb9d7ad1a),
	.w3(32'hb8a3785f),
	.w4(32'h36c892ea),
	.w5(32'hb9693012),
	.w6(32'h371c0f35),
	.w7(32'hb977f4ad),
	.w8(32'hb61bd501),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e243c3),
	.w1(32'h398a2437),
	.w2(32'h38a95362),
	.w3(32'h3a214a2e),
	.w4(32'hb97d419b),
	.w5(32'h38acc2b9),
	.w6(32'h38a18fb3),
	.w7(32'hba107b9d),
	.w8(32'h397ae5e7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9214dd0),
	.w1(32'h3a2f409e),
	.w2(32'hba5e9b01),
	.w3(32'h3926637b),
	.w4(32'h3aa4170e),
	.w5(32'hb9ace65d),
	.w6(32'h399b7992),
	.w7(32'hb8d3e842),
	.w8(32'h39ce5aca),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40af18),
	.w1(32'hbaac1e2e),
	.w2(32'hba809c12),
	.w3(32'hbb1a1a70),
	.w4(32'hba806e23),
	.w5(32'hba3785a7),
	.w6(32'hbaead43e),
	.w7(32'hbacf6f9c),
	.w8(32'hba9d4d13),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8942f8),
	.w1(32'hb73a9cfa),
	.w2(32'hb984beed),
	.w3(32'hba65012e),
	.w4(32'h39011a66),
	.w5(32'hb8aa79f1),
	.w6(32'h392d062c),
	.w7(32'hb8bdf4d6),
	.w8(32'h383ce3e3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953868a),
	.w1(32'h3973f21f),
	.w2(32'h38f6f307),
	.w3(32'hb81a4e6a),
	.w4(32'h39e0f417),
	.w5(32'h39a155ba),
	.w6(32'h39cfb922),
	.w7(32'h39eac6db),
	.w8(32'h39f604f6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81c19cc),
	.w1(32'h39a81568),
	.w2(32'hba325f14),
	.w3(32'hb70de417),
	.w4(32'h38d75c15),
	.w5(32'hba3eeda9),
	.w6(32'hb85e0af2),
	.w7(32'hb9df1393),
	.w8(32'hba854629),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa88530),
	.w1(32'hba1d72c8),
	.w2(32'hb8fb6712),
	.w3(32'hba510dfe),
	.w4(32'hba0a103c),
	.w5(32'hb96ae3f8),
	.w6(32'hba765a71),
	.w7(32'hba00be2e),
	.w8(32'h389d709b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382c3656),
	.w1(32'h381f8dd9),
	.w2(32'h384520ee),
	.w3(32'hb9dbb4b6),
	.w4(32'hb954ccff),
	.w5(32'hb8c073d2),
	.w6(32'hb91fb877),
	.w7(32'h38aad81c),
	.w8(32'h385ec3d1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96786f1),
	.w1(32'h3903fabc),
	.w2(32'hb9cefd4b),
	.w3(32'hb9c3e688),
	.w4(32'h3923af87),
	.w5(32'hb8d9917a),
	.w6(32'h38aba871),
	.w7(32'h391a51e2),
	.w8(32'h388bf51b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19f05b),
	.w1(32'h38ed8b83),
	.w2(32'hba8ebd49),
	.w3(32'hba9f1156),
	.w4(32'hba413337),
	.w5(32'hba791ce6),
	.w6(32'hbae917f7),
	.w7(32'hbaa6ade3),
	.w8(32'hba26f78a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e474c1),
	.w1(32'h3b072c53),
	.w2(32'h399f6667),
	.w3(32'h3ad0c2a1),
	.w4(32'h3b34e61b),
	.w5(32'h3ac3ee50),
	.w6(32'hb95106f1),
	.w7(32'h3ad2f0cf),
	.w8(32'h3889aa83),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ad7c9),
	.w1(32'h3b7b6944),
	.w2(32'h3b8dfc48),
	.w3(32'h3b0920a4),
	.w4(32'h3b92aee2),
	.w5(32'h3b81ae7b),
	.w6(32'h3ad976ff),
	.w7(32'h3b2f25f0),
	.w8(32'h3b19811a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34a3b1),
	.w1(32'hb89ec2f5),
	.w2(32'hba3160e1),
	.w3(32'h3a58723f),
	.w4(32'hb91a6bec),
	.w5(32'hbaadf01e),
	.w6(32'h3a476331),
	.w7(32'h39fb31b3),
	.w8(32'hba7c83fd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dc6b8),
	.w1(32'hba2fb1ec),
	.w2(32'hba1565fe),
	.w3(32'hba8203e8),
	.w4(32'hb9e6473b),
	.w5(32'hba191b21),
	.w6(32'hba6f18ac),
	.w7(32'hba148793),
	.w8(32'hb9a95f0a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba860614),
	.w1(32'hba10c7a4),
	.w2(32'hb9830f60),
	.w3(32'hba6107d3),
	.w4(32'hba65008e),
	.w5(32'hb9d2127d),
	.w6(32'hba09289c),
	.w7(32'hb9dfb64b),
	.w8(32'hb9e72094),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27a8be),
	.w1(32'h39a0e352),
	.w2(32'h39d2dfc0),
	.w3(32'hba282e52),
	.w4(32'h3a1a0ea0),
	.w5(32'h3a33d643),
	.w6(32'h399f6958),
	.w7(32'h399079c7),
	.w8(32'h3a4e9838),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf03a1b),
	.w1(32'hbaa910ee),
	.w2(32'hbb186b4e),
	.w3(32'hba0963a5),
	.w4(32'hba55ec7e),
	.w5(32'hbb07bc2b),
	.w6(32'h3a9a5440),
	.w7(32'hb8bfe33c),
	.w8(32'hba7a70d9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad554b4),
	.w1(32'hba5d6cf4),
	.w2(32'hb9a6acc1),
	.w3(32'hba69fee1),
	.w4(32'hb9fc543e),
	.w5(32'hba103032),
	.w6(32'hba2de177),
	.w7(32'hba2185db),
	.w8(32'hba7a139e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91b511),
	.w1(32'hba8bdd7f),
	.w2(32'hbaa07c9b),
	.w3(32'hb9a0d04f),
	.w4(32'hba2382a6),
	.w5(32'hbaa53201),
	.w6(32'hba80bfdf),
	.w7(32'hba9b67ec),
	.w8(32'hbaea5ca2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33c309),
	.w1(32'h3890ff2d),
	.w2(32'h39f38ad9),
	.w3(32'hbaffdce7),
	.w4(32'hb88acd75),
	.w5(32'hb813aaf2),
	.w6(32'hba7dd650),
	.w7(32'hb83c4e95),
	.w8(32'hb99bb669),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafaad65),
	.w1(32'hbb7b2783),
	.w2(32'hbbb039a9),
	.w3(32'hbb2ed708),
	.w4(32'hbb6b1cd7),
	.w5(32'hbb56bb9b),
	.w6(32'hbb2fac7c),
	.w7(32'hbb812f44),
	.w8(32'hbb25a4d5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab6273),
	.w1(32'h39d4d132),
	.w2(32'hb9569676),
	.w3(32'hba22ccc2),
	.w4(32'h3a2ab94e),
	.w5(32'h3872d3a3),
	.w6(32'h3a14a542),
	.w7(32'h39f5635b),
	.w8(32'h39994cdd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36be925c),
	.w1(32'h39e1ff0c),
	.w2(32'h3992701d),
	.w3(32'h3a0b0236),
	.w4(32'h39fa32f0),
	.w5(32'h38e15401),
	.w6(32'h3a084a90),
	.w7(32'h3988a32b),
	.w8(32'h39acc770),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01b18e),
	.w1(32'h3aa24cd4),
	.w2(32'h3a1ed9df),
	.w3(32'h3a80c755),
	.w4(32'h3a8d5f03),
	.w5(32'h3a1cb47e),
	.w6(32'h3adc5438),
	.w7(32'h3a9477cb),
	.w8(32'h3a2d268d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6f73a),
	.w1(32'h3a1b7ef3),
	.w2(32'hba5b49b6),
	.w3(32'h3988cebb),
	.w4(32'hba37e169),
	.w5(32'hba8c59d0),
	.w6(32'hb9216510),
	.w7(32'hba25d7e7),
	.w8(32'hba840564),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388111b2),
	.w1(32'hbab6f450),
	.w2(32'hbafe1ebb),
	.w3(32'h3a5a339b),
	.w4(32'hba972441),
	.w5(32'hbaf350de),
	.w6(32'hba8a5eca),
	.w7(32'hbab81bc3),
	.w8(32'hbacc4675),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aac6d1),
	.w1(32'h3a2ac436),
	.w2(32'hbb21c9d7),
	.w3(32'hba5396fc),
	.w4(32'hba27f625),
	.w5(32'hbb3888ef),
	.w6(32'h3a68d5e3),
	.w7(32'h39cbb696),
	.w8(32'hbb046a91),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37a0bd),
	.w1(32'hb948b51d),
	.w2(32'hb9d97aeb),
	.w3(32'hb814282a),
	.w4(32'hb93acd61),
	.w5(32'hb96667be),
	.w6(32'h376ce014),
	.w7(32'hb9857b4d),
	.w8(32'hb9abe90b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc585e),
	.w1(32'hba1c78f6),
	.w2(32'hba981bb2),
	.w3(32'hb9835a91),
	.w4(32'hba2a94e4),
	.w5(32'hba6e32be),
	.w6(32'hba333593),
	.w7(32'hba547630),
	.w8(32'hba7fcb0e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa650bd),
	.w1(32'hba503988),
	.w2(32'hba42b1b3),
	.w3(32'hba638045),
	.w4(32'hba4d43f4),
	.w5(32'hba375859),
	.w6(32'hb9e29dec),
	.w7(32'hba3dd057),
	.w8(32'hba3c4d32),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e8112),
	.w1(32'h3935eb5e),
	.w2(32'hb980770d),
	.w3(32'hba4984ca),
	.w4(32'h38c5b302),
	.w5(32'hb993375b),
	.w6(32'hb90b34b8),
	.w7(32'hb9f7f865),
	.w8(32'hb8f2ed5f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3869c668),
	.w1(32'h39d2b50d),
	.w2(32'h3a311cb2),
	.w3(32'hb9ea4e4f),
	.w4(32'h38455063),
	.w5(32'h390629f0),
	.w6(32'hb8c912bb),
	.w7(32'h393ee7a4),
	.w8(32'h38e3d4a7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d389fe),
	.w1(32'h394455b2),
	.w2(32'hb88b0632),
	.w3(32'hba10e21b),
	.w4(32'h394ca32b),
	.w5(32'h386aba55),
	.w6(32'hb9026c18),
	.w7(32'hb957dba5),
	.w8(32'h39123e5b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae975b9),
	.w1(32'hbb2ae555),
	.w2(32'hbaba194b),
	.w3(32'hbb0d88c6),
	.w4(32'hbb48a0eb),
	.w5(32'hbaf24bb6),
	.w6(32'hbb296d6d),
	.w7(32'hbb0074f9),
	.w8(32'hbaccade4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a3cac),
	.w1(32'hba1e8ee2),
	.w2(32'hba5f9be0),
	.w3(32'hba8218de),
	.w4(32'hb9918a7d),
	.w5(32'hba41cb18),
	.w6(32'h388f7451),
	.w7(32'hb9741d86),
	.w8(32'hb8d210b3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a8bcf),
	.w1(32'h399fd303),
	.w2(32'hba17ef65),
	.w3(32'h37fa9560),
	.w4(32'h39b083f4),
	.w5(32'hb9357603),
	.w6(32'h38166ca2),
	.w7(32'hb96587fc),
	.w8(32'hba0dcaa1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c12b4),
	.w1(32'h39fab138),
	.w2(32'h38f194a8),
	.w3(32'h3902d1bc),
	.w4(32'h39efa29f),
	.w5(32'h38ea10dc),
	.w6(32'h3a690341),
	.w7(32'h39d840cd),
	.w8(32'h39c56efc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbea15),
	.w1(32'hb94fcacb),
	.w2(32'hba1b3467),
	.w3(32'h39b79996),
	.w4(32'hb96ac209),
	.w5(32'hba369ae9),
	.w6(32'h382bb2a6),
	.w7(32'hb9902316),
	.w8(32'hba15c89b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee0a69),
	.w1(32'hb8c6f722),
	.w2(32'hb9c1a3da),
	.w3(32'hba094f40),
	.w4(32'h3774017a),
	.w5(32'hb91ffe51),
	.w6(32'hb72eb66f),
	.w7(32'hb9cdd1ec),
	.w8(32'hb919f8bb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab28bb8),
	.w1(32'hbab3ec05),
	.w2(32'hbac64d68),
	.w3(32'h3828a510),
	.w4(32'hbb042519),
	.w5(32'hbb1c3257),
	.w6(32'hba8ac1f5),
	.w7(32'hbac26278),
	.w8(32'hbb1e22a1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad73848),
	.w1(32'hba90fd95),
	.w2(32'hbb0711b0),
	.w3(32'hbac1ffcb),
	.w4(32'hba677adc),
	.w5(32'hbb0baf52),
	.w6(32'hbabe4dd2),
	.w7(32'hbac79045),
	.w8(32'hbadb107e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb7a64),
	.w1(32'h3a4b6ded),
	.w2(32'hba214741),
	.w3(32'h3a6beb76),
	.w4(32'h3a8c6a3d),
	.w5(32'hb9fc18ce),
	.w6(32'h370728ce),
	.w7(32'h391414ef),
	.w8(32'hba15576f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0428f2),
	.w1(32'h3a022260),
	.w2(32'hba363b49),
	.w3(32'hbab93a96),
	.w4(32'h3a22e831),
	.w5(32'hb9f04a66),
	.w6(32'hb9d83bf8),
	.w7(32'hb7da3769),
	.w8(32'hba82dceb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a194a),
	.w1(32'hb8a68eb5),
	.w2(32'hb91233d5),
	.w3(32'h39597e1b),
	.w4(32'hb9885df0),
	.w5(32'hb9c37b80),
	.w6(32'h385313b0),
	.w7(32'hb8bf5c56),
	.w8(32'hb9bd6e95),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2063e),
	.w1(32'hb983f198),
	.w2(32'hb9cea25e),
	.w3(32'hb9e184dd),
	.w4(32'hb750757a),
	.w5(32'hb9855a59),
	.w6(32'hb8f9fe18),
	.w7(32'hb9ad277a),
	.w8(32'hb92ea7f2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2aa89),
	.w1(32'hb98ad136),
	.w2(32'hb9b41777),
	.w3(32'hb96b25d3),
	.w4(32'hb84071a0),
	.w5(32'hb957d3ca),
	.w6(32'hb9199c32),
	.w7(32'hb996d2c2),
	.w8(32'hb810065b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51735b),
	.w1(32'hba117412),
	.w2(32'hba5c335b),
	.w3(32'hba685dce),
	.w4(32'hb9a227de),
	.w5(32'hb8cc4668),
	.w6(32'hb9f7d057),
	.w7(32'hba14037e),
	.w8(32'hb885b0d0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb705caec),
	.w1(32'hb9d1f07b),
	.w2(32'hb92a2a38),
	.w3(32'h39eaff5a),
	.w4(32'hba3d743f),
	.w5(32'hba2fd660),
	.w6(32'hb96706a0),
	.w7(32'hb9bd6360),
	.w8(32'hba004f3d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8953353),
	.w1(32'hb8443c49),
	.w2(32'hba55dbc0),
	.w3(32'hb9e79253),
	.w4(32'hba26eb0c),
	.w5(32'hb9fda50f),
	.w6(32'hb9fba0fc),
	.w7(32'hb8869aea),
	.w8(32'hba883de1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd29b),
	.w1(32'hba9beac7),
	.w2(32'hbb0a07e1),
	.w3(32'hbab3f615),
	.w4(32'hba97e092),
	.w5(32'hbad41f42),
	.w6(32'hba9db7d4),
	.w7(32'hba54587d),
	.w8(32'hb98dee23),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c5fc),
	.w1(32'hbb1d40a6),
	.w2(32'hbb0e0839),
	.w3(32'hbb3c6a54),
	.w4(32'hbb2dfaa3),
	.w5(32'hbab9988b),
	.w6(32'hbb3223d0),
	.w7(32'hbb16e43f),
	.w8(32'hbaa8037f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3a471),
	.w1(32'hba4e16d7),
	.w2(32'hbad6e03c),
	.w3(32'hba1011f2),
	.w4(32'hba7b4c37),
	.w5(32'hbad264b8),
	.w6(32'hb9e01f3f),
	.w7(32'hbac06c8d),
	.w8(32'hbb045c84),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b3c899),
	.w1(32'h38f7f275),
	.w2(32'hba9215d9),
	.w3(32'hba21b0e9),
	.w4(32'hb985853c),
	.w5(32'hbac24df6),
	.w6(32'h3939ca2b),
	.w7(32'hba0ae512),
	.w8(32'hba589a5e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba175540),
	.w1(32'hba7199db),
	.w2(32'hba2d58f1),
	.w3(32'hb9f84411),
	.w4(32'hba4fc41d),
	.w5(32'hba4d9d30),
	.w6(32'hbb0394e3),
	.w7(32'hbacfa801),
	.w8(32'hba7a1359),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca791f),
	.w1(32'hba686087),
	.w2(32'hba691403),
	.w3(32'hbad8804e),
	.w4(32'hbaa936c9),
	.w5(32'hba56a320),
	.w6(32'hba29b6dc),
	.w7(32'hba486da3),
	.w8(32'hba66990e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c34ea3),
	.w1(32'hb9da3e3f),
	.w2(32'hba3ffe16),
	.w3(32'hba023249),
	.w4(32'hb9dfe69f),
	.w5(32'hba2f270e),
	.w6(32'hb9e3bab4),
	.w7(32'hba36d50a),
	.w8(32'hba04673a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34465e),
	.w1(32'hb9742e3d),
	.w2(32'hb8a5307d),
	.w3(32'hb9c354f7),
	.w4(32'hb9c1dd6c),
	.w5(32'hb99fab51),
	.w6(32'hb993f87b),
	.w7(32'hb953da9c),
	.w8(32'hba084aa1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11506e),
	.w1(32'hb9385a53),
	.w2(32'hb8eb12b4),
	.w3(32'hba19e776),
	.w4(32'hb9c5a594),
	.w5(32'hb85e2d3f),
	.w6(32'hb95938e2),
	.w7(32'h391d838f),
	.w8(32'hb9d53cdf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ca629),
	.w1(32'hba60a630),
	.w2(32'hba33b672),
	.w3(32'hb9b8f9fe),
	.w4(32'hba2d96db),
	.w5(32'hba3255c1),
	.w6(32'hba531fc5),
	.w7(32'hba4d8e86),
	.w8(32'hba683873),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba193ad5),
	.w1(32'h3ad5549a),
	.w2(32'h3a819f77),
	.w3(32'h3a424e7c),
	.w4(32'h3b000050),
	.w5(32'h3a055d1c),
	.w6(32'h3a945b1b),
	.w7(32'h3a43d0e3),
	.w8(32'hb9a8056b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9765890),
	.w1(32'hb98e11ca),
	.w2(32'h385ff973),
	.w3(32'h38183a72),
	.w4(32'h3949eb92),
	.w5(32'h3a10eb07),
	.w6(32'hb9702685),
	.w7(32'hb7a73eb5),
	.w8(32'h3a1fa555),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a752f19),
	.w1(32'hb9c0d2a9),
	.w2(32'hbaad0ad1),
	.w3(32'h3ab1162b),
	.w4(32'hba151313),
	.w5(32'hbae2ed87),
	.w6(32'h3aa1cb78),
	.w7(32'hb8ed9b72),
	.w8(32'hbad7cdb8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5497f0),
	.w1(32'hba17d322),
	.w2(32'hbad755af),
	.w3(32'hba98c3fb),
	.w4(32'hba50d26f),
	.w5(32'hbaaaee3e),
	.w6(32'hb9fcc5fd),
	.w7(32'hba2c3391),
	.w8(32'hb9be1f87),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83f8d22),
	.w1(32'h3a63fae1),
	.w2(32'hb9ece980),
	.w3(32'h3a225396),
	.w4(32'h3ac9f041),
	.w5(32'h38eecce1),
	.w6(32'h39a88194),
	.w7(32'h3a330bf9),
	.w8(32'h39412c85),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399188f8),
	.w1(32'h398db01e),
	.w2(32'hb9de2fa9),
	.w3(32'hb9ea8bca),
	.w4(32'hb94129ac),
	.w5(32'hba276bf1),
	.w6(32'hb9ac1385),
	.w7(32'hba24b6fe),
	.w8(32'hba92dc47),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae290f3),
	.w1(32'h3a0acc44),
	.w2(32'hba3abd22),
	.w3(32'h3abb92f0),
	.w4(32'h39825df8),
	.w5(32'hba890870),
	.w6(32'h3a7cc4d6),
	.w7(32'h391ea64f),
	.w8(32'hbaab3df8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65ba7e),
	.w1(32'hb8a01ce1),
	.w2(32'hbb30efb1),
	.w3(32'h3a67e1e5),
	.w4(32'hb9835f6b),
	.w5(32'hbb61149d),
	.w6(32'h39cdc314),
	.w7(32'hba5b54eb),
	.w8(32'hbb4137a6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb4524),
	.w1(32'h39699e97),
	.w2(32'hbae0a9a3),
	.w3(32'h3b0875f3),
	.w4(32'hb7856f06),
	.w5(32'hbb2151d8),
	.w6(32'h3b036dd2),
	.w7(32'h39e80c39),
	.w8(32'hbb187f24),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba810222),
	.w1(32'hb986288a),
	.w2(32'hba8cef23),
	.w3(32'hb9a5c0bd),
	.w4(32'hb906c3b4),
	.w5(32'hba6cda17),
	.w6(32'hb80b7ac1),
	.w7(32'hb84d1fa1),
	.w8(32'hbad2af69),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977c40c),
	.w1(32'hb9ee8752),
	.w2(32'hba3e9889),
	.w3(32'h3a21362b),
	.w4(32'hb971320a),
	.w5(32'hba1b7121),
	.w6(32'h37271c42),
	.w7(32'hb9ed12c2),
	.w8(32'h3a1dd4c8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd2677),
	.w1(32'hb8997532),
	.w2(32'hbb584f68),
	.w3(32'h3a072f69),
	.w4(32'hb816cb26),
	.w5(32'hbb0e0af4),
	.w6(32'h3a312e45),
	.w7(32'hba9a9766),
	.w8(32'hba566ab7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc513),
	.w1(32'h3b2ce2df),
	.w2(32'h3a2a0f74),
	.w3(32'h3b6152d9),
	.w4(32'h3ae5fefb),
	.w5(32'h3903e70a),
	.w6(32'h3af0b720),
	.w7(32'h3a8cb934),
	.w8(32'h375ea206),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbb8e3),
	.w1(32'hba8fe454),
	.w2(32'hbb212a48),
	.w3(32'hbb00f937),
	.w4(32'hbad1c5b3),
	.w5(32'hbb16d19d),
	.w6(32'hba884faa),
	.w7(32'hb9cce3f8),
	.w8(32'hbaa22c4b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a715f3a),
	.w1(32'h3bf473f0),
	.w2(32'h3b59293b),
	.w3(32'h3bb2a334),
	.w4(32'h3c02b79b),
	.w5(32'h3baf1741),
	.w6(32'h3b5c0123),
	.w7(32'h3b1337a8),
	.w8(32'h3b4c527d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffe2ac),
	.w1(32'hbab62553),
	.w2(32'hbab14396),
	.w3(32'hbaa89c8f),
	.w4(32'hbad0917f),
	.w5(32'hba9dd6f6),
	.w6(32'hb98aac8c),
	.w7(32'hba61310c),
	.w8(32'hbb06310c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37f1ad),
	.w1(32'h3b5b085d),
	.w2(32'hba994719),
	.w3(32'h3b2ebee7),
	.w4(32'h3b60fa5d),
	.w5(32'hb9fa60d1),
	.w6(32'h3ae36ee2),
	.w7(32'h3aa3eff7),
	.w8(32'hb8d3169e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b3ca9),
	.w1(32'h3a1f2e86),
	.w2(32'hba3d5b6d),
	.w3(32'h3ab92731),
	.w4(32'h3a8240e1),
	.w5(32'hba037de4),
	.w6(32'h3a2c7b8d),
	.w7(32'h39ee3320),
	.w8(32'h3a9b73cc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba932ae9),
	.w1(32'h3a1d127d),
	.w2(32'hbaa18a4e),
	.w3(32'hbade0336),
	.w4(32'hb8559a4c),
	.w5(32'hb9c38ecc),
	.w6(32'hba282a30),
	.w7(32'hb9e6e6d1),
	.w8(32'h3a4831ac),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71827c),
	.w1(32'hb8bca26f),
	.w2(32'h381b0530),
	.w3(32'hb8403f43),
	.w4(32'h38c9cb75),
	.w5(32'h39376ec2),
	.w6(32'hb99dd087),
	.w7(32'h393c0e7c),
	.w8(32'h3971c9c4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a5e9e6),
	.w1(32'hba70cc9b),
	.w2(32'hba8118b4),
	.w3(32'hb7feae68),
	.w4(32'hba845282),
	.w5(32'hba7a0544),
	.w6(32'hba652649),
	.w7(32'hba5be391),
	.w8(32'hba7d9aa7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d98f5),
	.w1(32'hb90e5caa),
	.w2(32'hba23900b),
	.w3(32'hba5a2793),
	.w4(32'h39f470a7),
	.w5(32'h372a0702),
	.w6(32'h39a9a83e),
	.w7(32'h38d6f379),
	.w8(32'h38f664a7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3f025),
	.w1(32'hbaa7eb70),
	.w2(32'hbb0ba33a),
	.w3(32'hba514cb6),
	.w4(32'hba25f2c8),
	.w5(32'hbac6877f),
	.w6(32'h39d89f2a),
	.w7(32'hba8d50d1),
	.w8(32'hba3e2155),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03cbb1),
	.w1(32'hb949a005),
	.w2(32'hba40de49),
	.w3(32'h3a03e1a4),
	.w4(32'h37eb4337),
	.w5(32'hba87793d),
	.w6(32'h3a0ea6e3),
	.w7(32'h38b5c4a8),
	.w8(32'hba97ea95),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14792a),
	.w1(32'h3a4bae8c),
	.w2(32'hb954c63c),
	.w3(32'h3a64a5ab),
	.w4(32'h3a50d274),
	.w5(32'h3a3a4220),
	.w6(32'h3a23c22e),
	.w7(32'h3a21973c),
	.w8(32'h3a02539b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9485246),
	.w1(32'h3aca6764),
	.w2(32'h3a8fc172),
	.w3(32'h3a0eb986),
	.w4(32'h3ac79c16),
	.w5(32'h3a518b9f),
	.w6(32'h3a3267aa),
	.w7(32'h3a646b7c),
	.w8(32'h3a25b28f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bca4b),
	.w1(32'h39d767a1),
	.w2(32'h39d38373),
	.w3(32'h3a13d0e1),
	.w4(32'h381e29e5),
	.w5(32'h399de861),
	.w6(32'hba8c0cb3),
	.w7(32'hba212f49),
	.w8(32'hb8407442),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cfaaf),
	.w1(32'hba43fe7a),
	.w2(32'hba8e0ffe),
	.w3(32'hba9f84cf),
	.w4(32'hbacb49c8),
	.w5(32'hbae1c2fb),
	.w6(32'hba8866e6),
	.w7(32'hba931588),
	.w8(32'hbb075f2d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba662a3b),
	.w1(32'h38b7c509),
	.w2(32'hb9e568bd),
	.w3(32'hba284ec9),
	.w4(32'h39b9b899),
	.w5(32'hb9cc158f),
	.w6(32'h39052612),
	.w7(32'hb8e7278a),
	.w8(32'hba06c945),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ee084),
	.w1(32'h3910d638),
	.w2(32'hb9a512a6),
	.w3(32'h374b10ac),
	.w4(32'h3a13c982),
	.w5(32'hb6e66a23),
	.w6(32'h3a069b22),
	.w7(32'hb7f598d0),
	.w8(32'h39ffa621),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87b4b4e),
	.w1(32'hb9a9195d),
	.w2(32'hb9f80a5d),
	.w3(32'h39b16af7),
	.w4(32'hb8bd460d),
	.w5(32'hb9a4470f),
	.w6(32'hb8eea0b9),
	.w7(32'hb9b5eee0),
	.w8(32'hb918f161),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9847ea3),
	.w1(32'hb918ad26),
	.w2(32'hb9fa71a7),
	.w3(32'h37d47028),
	.w4(32'h3940d187),
	.w5(32'hb98652d7),
	.w6(32'h38d95ed1),
	.w7(32'hb9629a98),
	.w8(32'hb85ee1fa),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98da178),
	.w1(32'hba2bc52e),
	.w2(32'hb9aaadd4),
	.w3(32'hb83466a4),
	.w4(32'h37d1c75a),
	.w5(32'h390d9e8b),
	.w6(32'hb9d67291),
	.w7(32'hb9910114),
	.w8(32'h373c310c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16cae5),
	.w1(32'hba1474c7),
	.w2(32'hb9df85ac),
	.w3(32'h399bbcf3),
	.w4(32'hba1cd049),
	.w5(32'hb9e73878),
	.w6(32'hba90960f),
	.w7(32'hba9554b0),
	.w8(32'hba6cc8e5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b9d20),
	.w1(32'hba29d271),
	.w2(32'hba4c4358),
	.w3(32'hba0c29b2),
	.w4(32'hba07f4b1),
	.w5(32'hba322579),
	.w6(32'hba81ecda),
	.w7(32'hba7bfc2d),
	.w8(32'hba347fcf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad9435),
	.w1(32'hba7b2e2d),
	.w2(32'hbadf4cd7),
	.w3(32'hba97f03f),
	.w4(32'hba85d189),
	.w5(32'hbab1078f),
	.w6(32'hba8f9f34),
	.w7(32'hbadc8fe8),
	.w8(32'hbabd4bde),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba961dd2),
	.w1(32'h3a033d55),
	.w2(32'hb94a1948),
	.w3(32'hba0beacf),
	.w4(32'h3a366ea7),
	.w5(32'h3851215d),
	.w6(32'h3924f9a7),
	.w7(32'h396c5b13),
	.w8(32'hb8d92800),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0234e),
	.w1(32'hb8224674),
	.w2(32'h39855800),
	.w3(32'h38b786e6),
	.w4(32'h398d14ad),
	.w5(32'h3a340e47),
	.w6(32'h37a5a231),
	.w7(32'h380f42fa),
	.w8(32'hb99a4303),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39438ae8),
	.w1(32'hbad04836),
	.w2(32'hbadb97d4),
	.w3(32'h3a0b3413),
	.w4(32'hbaa40ba5),
	.w5(32'hbacb7b7c),
	.w6(32'hbaab4623),
	.w7(32'hbad70fd2),
	.w8(32'hbacfc445),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7503e),
	.w1(32'hb9a26dc3),
	.w2(32'hba344445),
	.w3(32'hba9d82ef),
	.w4(32'h38dd9065),
	.w5(32'hb984a146),
	.w6(32'hb84bafea),
	.w7(32'hb9c07cd7),
	.w8(32'h370e6140),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c512c),
	.w1(32'hb9213dc1),
	.w2(32'hba4759e5),
	.w3(32'hb8af2b57),
	.w4(32'hb97af478),
	.w5(32'hb9fb21f3),
	.w6(32'h39cdbe15),
	.w7(32'hb6d9ad82),
	.w8(32'hb98c03ec),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8a2b7),
	.w1(32'hb727419d),
	.w2(32'hb987144b),
	.w3(32'hba3cc15f),
	.w4(32'hb9dc264d),
	.w5(32'hba3bf620),
	.w6(32'hb9f78f4b),
	.w7(32'hb9bed872),
	.w8(32'hba329657),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372e8afb),
	.w1(32'hbacdb2b4),
	.w2(32'hbb667db8),
	.w3(32'hba08274b),
	.w4(32'hbab1ed4a),
	.w5(32'hbb64b8f0),
	.w6(32'h3a2cada3),
	.w7(32'hba04cb59),
	.w8(32'hbb36ab71),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f3c6f8),
	.w1(32'h382f82ad),
	.w2(32'hb879e31c),
	.w3(32'h37bb05ef),
	.w4(32'hb7fee27c),
	.w5(32'hb8217f39),
	.w6(32'hb8272ce7),
	.w7(32'hb723ce1b),
	.w8(32'hb7cc1091),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e05bd4),
	.w1(32'hb908a4ef),
	.w2(32'hb9a676f7),
	.w3(32'hb9c34612),
	.w4(32'hb92b7a1f),
	.w5(32'hb94cdbe4),
	.w6(32'hb9dbca69),
	.w7(32'hb96cc240),
	.w8(32'hb9054cf5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389610d8),
	.w1(32'h3992c05f),
	.w2(32'hb9d673ef),
	.w3(32'h395745f7),
	.w4(32'h39582270),
	.w5(32'hba0a57cc),
	.w6(32'h391456c1),
	.w7(32'h38b52e9c),
	.w8(32'hba38edb0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710634d),
	.w1(32'hb939bee7),
	.w2(32'hba406d3b),
	.w3(32'h38b4fc44),
	.w4(32'hb8bc5040),
	.w5(32'hb9f13c68),
	.w6(32'h39386c58),
	.w7(32'hb61da15e),
	.w8(32'hb9c5cb6c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a169a3d),
	.w1(32'h3979c3b8),
	.w2(32'hbaa7c4a3),
	.w3(32'h3a40ce11),
	.w4(32'h39a6459e),
	.w5(32'hbaba094d),
	.w6(32'h3a4156c5),
	.w7(32'h3989c336),
	.w8(32'hba9571f6),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90485b2),
	.w1(32'h3828e098),
	.w2(32'hbae92a26),
	.w3(32'hba30225b),
	.w4(32'hba2624f3),
	.w5(32'hba60f4a4),
	.w6(32'hb941c33d),
	.w7(32'hb9e10668),
	.w8(32'hb9fe2bce),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391dba0d),
	.w1(32'h37eac26e),
	.w2(32'hba0161cb),
	.w3(32'h3a386a8b),
	.w4(32'hb8672bce),
	.w5(32'hba17f5f7),
	.w6(32'h39c206e3),
	.w7(32'hb86f2a3c),
	.w8(32'hba893a42),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79b865),
	.w1(32'h3a52085d),
	.w2(32'h398d0c5d),
	.w3(32'h3b078c59),
	.w4(32'h3aecab79),
	.w5(32'h397bb55a),
	.w6(32'h3ad26c51),
	.w7(32'h3a073d2c),
	.w8(32'hba2bbc09),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb0b8),
	.w1(32'h3ad15505),
	.w2(32'hba25f501),
	.w3(32'h3ab95652),
	.w4(32'h3a843182),
	.w5(32'hba1ea44c),
	.w6(32'h3a556cbc),
	.w7(32'h3a6230af),
	.w8(32'hba18f9e2),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c3c9b),
	.w1(32'h39bf8d62),
	.w2(32'hb8155450),
	.w3(32'h39b7ab89),
	.w4(32'h39824044),
	.w5(32'hb99dfc05),
	.w6(32'h392df34b),
	.w7(32'h3921e878),
	.w8(32'hba0f210f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fc0ab),
	.w1(32'hb75ebbf0),
	.w2(32'hba8eb10a),
	.w3(32'hb9da1d69),
	.w4(32'hb942f60e),
	.w5(32'hba8f99ce),
	.w6(32'h39d6b581),
	.w7(32'hb996a97b),
	.w8(32'hbaacd436),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d6959),
	.w1(32'hb834a927),
	.w2(32'hb916a4b3),
	.w3(32'hb8ceb9f0),
	.w4(32'hb6ec2cc8),
	.w5(32'hb90fc38a),
	.w6(32'hb8c48cc7),
	.w7(32'hb8697040),
	.w8(32'hb90cb980),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4c8a5),
	.w1(32'h3a8c5cd3),
	.w2(32'h3912d13e),
	.w3(32'h3b007f1e),
	.w4(32'h3a68f632),
	.w5(32'h38c86eeb),
	.w6(32'h3a944932),
	.w7(32'hb8c6b586),
	.w8(32'hbaac524e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ebb10),
	.w1(32'h3a8b6688),
	.w2(32'hba858017),
	.w3(32'h3b22c33e),
	.w4(32'h3a574002),
	.w5(32'hbab9d09f),
	.w6(32'h3b19a43f),
	.w7(32'h3a7cb40f),
	.w8(32'hbaa7eefe),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4ccc085),
	.w1(32'h370727e0),
	.w2(32'h3677f809),
	.w3(32'h3726d304),
	.w4(32'h3717776c),
	.w5(32'h36bc0a6b),
	.w6(32'h37db7207),
	.w7(32'h37fbc4ea),
	.w8(32'h37d71d7c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371b8e75),
	.w1(32'h35150e58),
	.w2(32'h360664b8),
	.w3(32'h37a925a7),
	.w4(32'h379673c5),
	.w5(32'h37437494),
	.w6(32'h37f0fb9d),
	.w7(32'h37e3e03e),
	.w8(32'h373eac34),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c157e6),
	.w1(32'h38f985ab),
	.w2(32'h38d32bfa),
	.w3(32'hb8bba6f1),
	.w4(32'hb721bf02),
	.w5(32'h3924c8bd),
	.w6(32'hb8ef5b0e),
	.w7(32'hb7e0fe3b),
	.w8(32'h397055ca),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa4705),
	.w1(32'h3a7c9b76),
	.w2(32'hb9b7ed03),
	.w3(32'h3b2943a8),
	.w4(32'h3a9423e3),
	.w5(32'hba8017fa),
	.w6(32'h3b0425c5),
	.w7(32'h3a8312cc),
	.w8(32'hba8a58da),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fe82e),
	.w1(32'hbb074a0f),
	.w2(32'hbab5e7b4),
	.w3(32'hbb200b6b),
	.w4(32'hbb025749),
	.w5(32'hbaacfc9f),
	.w6(32'hbb14eebb),
	.w7(32'hbb03c10e),
	.w8(32'hba729401),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb726d44c),
	.w1(32'h36f97c62),
	.w2(32'h3757e929),
	.w3(32'hb737a400),
	.w4(32'hb69edc28),
	.w5(32'h375a5b85),
	.w6(32'hb79f2175),
	.w7(32'hb747c3a8),
	.w8(32'h3766d113),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba575187),
	.w1(32'hba5b5135),
	.w2(32'hbabb1b90),
	.w3(32'hba77eb01),
	.w4(32'hba7b890b),
	.w5(32'hbab5d26e),
	.w6(32'hba0539c0),
	.w7(32'hba93be3c),
	.w8(32'hbabfa6fa),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d80d6),
	.w1(32'hba7326ea),
	.w2(32'hbb06a4ae),
	.w3(32'h37c28b10),
	.w4(32'hba3a0f85),
	.w5(32'hbb069f16),
	.w6(32'h3a3a007d),
	.w7(32'hba18ffe6),
	.w8(32'hbb0146cc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02658c),
	.w1(32'hbaaa7f60),
	.w2(32'hbb1ff686),
	.w3(32'hbb4ce073),
	.w4(32'hbadbe68b),
	.w5(32'hba8287df),
	.w6(32'hbafe9112),
	.w7(32'hbb199fd8),
	.w8(32'hbaaeaf04),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55cf4a),
	.w1(32'hb9a73013),
	.w2(32'hba1acb1f),
	.w3(32'hb98ec610),
	.w4(32'hb9305a39),
	.w5(32'hb9c49e7c),
	.w6(32'hb95ae621),
	.w7(32'hb99d332d),
	.w8(32'hb9882aea),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48eae4),
	.w1(32'h3b0d61a8),
	.w2(32'h398087f1),
	.w3(32'h3b4093d3),
	.w4(32'h3ac45686),
	.w5(32'hb99a7d38),
	.w6(32'h3af78d4d),
	.w7(32'h3aa71e9a),
	.w8(32'h38553eee),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39549efe),
	.w1(32'h3a89b6cf),
	.w2(32'h391a575f),
	.w3(32'h3a450a02),
	.w4(32'h3ae24d03),
	.w5(32'h3a970a86),
	.w6(32'h3aa9bb2c),
	.w7(32'h3adf465f),
	.w8(32'h3a92e634),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2109),
	.w1(32'hb9a99274),
	.w2(32'h3aae96f4),
	.w3(32'hbb01a671),
	.w4(32'hb886f650),
	.w5(32'h3aa3ae1d),
	.w6(32'hbb0816fd),
	.w7(32'hba1c8581),
	.w8(32'h399da86b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba90c33),
	.w1(32'h3b376974),
	.w2(32'h39a1c2b5),
	.w3(32'h3bbcf02a),
	.w4(32'h3b3bed28),
	.w5(32'hba11837b),
	.w6(32'h3b8a3e31),
	.w7(32'h3b2be3be),
	.w8(32'hbaa59682),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a32ea8),
	.w1(32'h3a885c9d),
	.w2(32'h3aaf2623),
	.w3(32'h399c7c2a),
	.w4(32'h3a8c182f),
	.w5(32'h3aa7f69b),
	.w6(32'h38d6f1b0),
	.w7(32'h3a2d3a35),
	.w8(32'h3a6ae1e0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d73e78),
	.w1(32'h3836ac64),
	.w2(32'hb8c9b6cf),
	.w3(32'hb734f84b),
	.w4(32'hb71acb50),
	.w5(32'hb83559d1),
	.w6(32'h379b9173),
	.w7(32'h380981f2),
	.w8(32'hb891e826),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb762b281),
	.w1(32'hb80cfba5),
	.w2(32'hb768c8b8),
	.w3(32'hb6e82e35),
	.w4(32'h385f76b9),
	.w5(32'h389b7303),
	.w6(32'hb6e6fb89),
	.w7(32'h380a1775),
	.w8(32'h387616a8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba122967),
	.w1(32'hb993a158),
	.w2(32'hba9d81e5),
	.w3(32'hb9c3a9bc),
	.w4(32'hba17b580),
	.w5(32'hbaade0e5),
	.w6(32'hb86cb745),
	.w7(32'hba17722b),
	.w8(32'hba4099e7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c78b79),
	.w1(32'h389b301f),
	.w2(32'h38827fe7),
	.w3(32'h37612205),
	.w4(32'h38c4f114),
	.w5(32'h3865b447),
	.w6(32'h3846cc79),
	.w7(32'h38e9c345),
	.w8(32'h389259f5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba134073),
	.w1(32'hb7eb797a),
	.w2(32'h38abeb3b),
	.w3(32'hb9b1aba0),
	.w4(32'h37a7af10),
	.w5(32'h38a26f6b),
	.w6(32'hb93e552a),
	.w7(32'h381504f1),
	.w8(32'h387aafa2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8846c75),
	.w1(32'h38cfa903),
	.w2(32'h37bc1008),
	.w3(32'h38514de6),
	.w4(32'h39719de8),
	.w5(32'h38fe86a6),
	.w6(32'hb903dd4a),
	.w7(32'h37f23433),
	.w8(32'h3855152a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e37c58),
	.w1(32'h3a97508d),
	.w2(32'h3ae9862e),
	.w3(32'h39f7ca7e),
	.w4(32'h3ad5a82a),
	.w5(32'h3b081063),
	.w6(32'h39ae5620),
	.w7(32'h3ab9eb74),
	.w8(32'h3af91ddc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c975e0),
	.w1(32'h387de7cf),
	.w2(32'h391f5106),
	.w3(32'hb7f1732e),
	.w4(32'h392b5b4e),
	.w5(32'h39501e53),
	.w6(32'h37e85107),
	.w7(32'h39583b8b),
	.w8(32'h39708c73),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab7059),
	.w1(32'h392ea64f),
	.w2(32'hb9133fd4),
	.w3(32'h39721a93),
	.w4(32'h38a9b4f2),
	.w5(32'hb908d20e),
	.w6(32'h390a7431),
	.w7(32'h39227c28),
	.w8(32'h36430538),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977b65f),
	.w1(32'h39bac048),
	.w2(32'hba95b7e8),
	.w3(32'h3a06bb18),
	.w4(32'h39f99019),
	.w5(32'hba8da355),
	.w6(32'h3a87b92b),
	.w7(32'h39f2a68c),
	.w8(32'hba89e735),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba999757),
	.w1(32'hba566858),
	.w2(32'hbab3ab11),
	.w3(32'hbab6abde),
	.w4(32'hbaaf4b0a),
	.w5(32'hbb03c37f),
	.w6(32'hbabe9fc1),
	.w7(32'hba9b251a),
	.w8(32'hbb008c37),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22fa68),
	.w1(32'h3a874be2),
	.w2(32'h3a1260ad),
	.w3(32'h39b9c941),
	.w4(32'h3a650b85),
	.w5(32'h39e2be24),
	.w6(32'h39a7ba4f),
	.w7(32'h3a304365),
	.w8(32'h39b260fd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba666877),
	.w1(32'hba320023),
	.w2(32'hbad75693),
	.w3(32'hba20ffb4),
	.w4(32'hba0257b8),
	.w5(32'hbaa9ca12),
	.w6(32'h394b85b6),
	.w7(32'hb8da0d2c),
	.w8(32'hbaa5d25a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b4e1b),
	.w1(32'hb8270fb4),
	.w2(32'hb9fc7a47),
	.w3(32'h390546b5),
	.w4(32'hb8a520e4),
	.w5(32'hb9fc5e8d),
	.w6(32'h397b79c5),
	.w7(32'hb8ae45e6),
	.w8(32'hb9e65569),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0b6a8),
	.w1(32'hbaff9081),
	.w2(32'hba58bb68),
	.w3(32'h3a1c013f),
	.w4(32'hbaddfae9),
	.w5(32'hbac84c60),
	.w6(32'h3a477922),
	.w7(32'hba817afd),
	.w8(32'hbad8038d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e99f2e),
	.w1(32'hb91643a3),
	.w2(32'hba594be0),
	.w3(32'hba03ce42),
	.w4(32'h37041405),
	.w5(32'hba237533),
	.w6(32'hba183086),
	.w7(32'hb8b330c5),
	.w8(32'hb9fa95b1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05d9de),
	.w1(32'hb9ef466a),
	.w2(32'hbae7369f),
	.w3(32'hb9940af7),
	.w4(32'hb9c946b6),
	.w5(32'hbae075bb),
	.w6(32'h382a3b17),
	.w7(32'hb9c9f8ff),
	.w8(32'hbace6ede),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365cf31f),
	.w1(32'h3937beea),
	.w2(32'h39546bba),
	.w3(32'h391be578),
	.w4(32'h3a1671f0),
	.w5(32'h39a42cec),
	.w6(32'h39980d88),
	.w7(32'h3a2db48d),
	.w8(32'h39df5085),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacb50c),
	.w1(32'h39f99bab),
	.w2(32'hbac910c7),
	.w3(32'h3a7db38c),
	.w4(32'h39005b98),
	.w5(32'hbb0f222d),
	.w6(32'h3a79bbb0),
	.w7(32'hb83e856c),
	.w8(32'hbb1641b0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fc6ae7),
	.w1(32'h36d2539e),
	.w2(32'h36b541dd),
	.w3(32'h37dc1035),
	.w4(32'h3648299c),
	.w5(32'hb6978d81),
	.w6(32'h3809cff7),
	.w7(32'h373c558a),
	.w8(32'h372abe72),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2ee51),
	.w1(32'hba3d9107),
	.w2(32'hb9fc0789),
	.w3(32'hb9f299dc),
	.w4(32'hba4ab223),
	.w5(32'hb96db2d1),
	.w6(32'hb9f012e1),
	.w7(32'hb9eae220),
	.w8(32'hb756833d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380b79b4),
	.w1(32'h386be802),
	.w2(32'h37b99ff1),
	.w3(32'h3904a92d),
	.w4(32'h3929c0bd),
	.w5(32'h393195cf),
	.w6(32'hb661300f),
	.w7(32'h38cbf045),
	.w8(32'h3903e1d6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba877653),
	.w1(32'hba5cda87),
	.w2(32'hba97c9ee),
	.w3(32'hba324716),
	.w4(32'hba4e2745),
	.w5(32'hba894d9f),
	.w6(32'hba2b2880),
	.w7(32'hba841423),
	.w8(32'hba9d03d0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b6408e),
	.w1(32'hb4944b4b),
	.w2(32'h358bd821),
	.w3(32'h3690d001),
	.w4(32'hb43b6a33),
	.w5(32'h35a8c38c),
	.w6(32'h36a5d756),
	.w7(32'h3544940e),
	.w8(32'hb60edc65),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901a29b),
	.w1(32'h37f84918),
	.w2(32'hb7b74212),
	.w3(32'h37f664d2),
	.w4(32'h38ce0cb6),
	.w5(32'hb82e4916),
	.w6(32'h38a650c5),
	.w7(32'h385cf008),
	.w8(32'h37576322),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a0be1),
	.w1(32'h3a1974d1),
	.w2(32'h3a66c4ed),
	.w3(32'hb8345b36),
	.w4(32'h39ffd1ba),
	.w5(32'h3a4ca3f5),
	.w6(32'hb9867c05),
	.w7(32'h39667822),
	.w8(32'h3a0c247c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a744f02),
	.w1(32'h3b00999d),
	.w2(32'h3a6c378c),
	.w3(32'h3aad607e),
	.w4(32'h3adc8751),
	.w5(32'h3a5e7d8c),
	.w6(32'h3a1c9f11),
	.w7(32'hb84e76e8),
	.w8(32'h390b950b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ce41e),
	.w1(32'h3944c43d),
	.w2(32'hb8f14346),
	.w3(32'hb81474b0),
	.w4(32'hb82472c7),
	.w5(32'hb7c944b0),
	.w6(32'hb939890d),
	.w7(32'hb8aa0d5f),
	.w8(32'h3781cc50),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3869edff),
	.w1(32'hb89911ce),
	.w2(32'hb931c51e),
	.w3(32'h388aa234),
	.w4(32'hb7e0a403),
	.w5(32'hb9145051),
	.w6(32'h38fdb2dd),
	.w7(32'h3884a9ab),
	.w8(32'hb88c8622),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcb3de),
	.w1(32'hbc0743ea),
	.w2(32'hbb518c32),
	.w3(32'hbc034f75),
	.w4(32'hbbe9ac01),
	.w5(32'hbb6d65d8),
	.w6(32'hbbd3250d),
	.w7(32'hbbc2afcc),
	.w8(32'hbb0ca19e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04afdd),
	.w1(32'hb97ed5da),
	.w2(32'hbaf7e71b),
	.w3(32'h3ac4cb25),
	.w4(32'h3629e940),
	.w5(32'hbb925810),
	.w6(32'h3ab3849b),
	.w7(32'hba83b629),
	.w8(32'hbba5ef2d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947bdb9),
	.w1(32'h398ee7e8),
	.w2(32'h38bd6ec5),
	.w3(32'h3935be89),
	.w4(32'h396a5483),
	.w5(32'h38fac914),
	.w6(32'h39884e1c),
	.w7(32'h39b585d9),
	.w8(32'h398040a6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ab3d7b),
	.w1(32'h375f0e13),
	.w2(32'h369e0ac8),
	.w3(32'h36e1872c),
	.w4(32'h37839c39),
	.w5(32'h376bddaf),
	.w6(32'h37e0be70),
	.w7(32'h369fb478),
	.w8(32'h381ac316),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b358b),
	.w1(32'h392621cf),
	.w2(32'hb8fb5987),
	.w3(32'h39247a70),
	.w4(32'h39624f33),
	.w5(32'hb91e592a),
	.w6(32'h397c65b3),
	.w7(32'h36131dbe),
	.w8(32'hb92234ee),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38579bb0),
	.w1(32'h372b12ce),
	.w2(32'hb67ce80d),
	.w3(32'h37fd0d9e),
	.w4(32'hb724f8ce),
	.w5(32'hb7d78e74),
	.w6(32'h38141793),
	.w7(32'h36a024e1),
	.w8(32'hb5d6f8b2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a392803),
	.w1(32'h3a5ffd99),
	.w2(32'hb9488e4c),
	.w3(32'h3a305fde),
	.w4(32'h39fecf4d),
	.w5(32'hb99715e6),
	.w6(32'h3a1e50e7),
	.w7(32'h39602dc3),
	.w8(32'hb95b0b42),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dce0f),
	.w1(32'h3a9acdd9),
	.w2(32'hbaa7a01a),
	.w3(32'h3b4e3ea5),
	.w4(32'h3ab64b12),
	.w5(32'hba4855fe),
	.w6(32'h3b2cdcfc),
	.w7(32'h3acd76ec),
	.w8(32'hba1140fb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4154c),
	.w1(32'hbb2f66a0),
	.w2(32'hbae615af),
	.w3(32'hba9bddb0),
	.w4(32'hbb036b57),
	.w5(32'hbae52804),
	.w6(32'hba9a0719),
	.w7(32'hbaaf6b86),
	.w8(32'hbaae00de),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9961456),
	.w1(32'hb9409056),
	.w2(32'h3916a2dc),
	.w3(32'hb980495d),
	.w4(32'h365ab10a),
	.w5(32'h398d9bae),
	.w6(32'hb94671dd),
	.w7(32'h383a0c98),
	.w8(32'h397b5baf),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ebe67),
	.w1(32'hbaff477d),
	.w2(32'hbb0dc320),
	.w3(32'hbb25be0e),
	.w4(32'hbb0ed297),
	.w5(32'hbaa1cde2),
	.w6(32'hbadbdcc0),
	.w7(32'hbae68177),
	.w8(32'hba312b74),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ebf82),
	.w1(32'h38fb82e2),
	.w2(32'h38c85cf5),
	.w3(32'hb98b43ff),
	.w4(32'h372a800a),
	.w5(32'h3a002832),
	.w6(32'hb9e4caaf),
	.w7(32'hb9b63a02),
	.w8(32'h39021f39),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36daca03),
	.w1(32'h369918c7),
	.w2(32'h378a20b8),
	.w3(32'h36969bf7),
	.w4(32'h35e1ae43),
	.w5(32'h3752eefa),
	.w6(32'h374bb666),
	.w7(32'h373030a4),
	.w8(32'h379cbc05),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398062cf),
	.w1(32'h3991c3ce),
	.w2(32'hb6a184d5),
	.w3(32'h37ea7039),
	.w4(32'hb8cdb7f9),
	.w5(32'hb941b392),
	.w6(32'hb89c365c),
	.w7(32'hb86fac10),
	.w8(32'h359c0cf4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f200c2),
	.w1(32'hb76578c2),
	.w2(32'h36a3a2c8),
	.w3(32'h379f3ac6),
	.w4(32'hb766f81e),
	.w5(32'hb754e243),
	.w6(32'h3810ce71),
	.w7(32'h370373a7),
	.w8(32'h36d6e641),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d6b51),
	.w1(32'hb960f3df),
	.w2(32'hba005b9f),
	.w3(32'hb9e3624c),
	.w4(32'hb91ae0c0),
	.w5(32'hb9ca46a0),
	.w6(32'hba1d7771),
	.w7(32'hb9cdc83f),
	.w8(32'hb9f369ed),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b270e93),
	.w1(32'h3a967c95),
	.w2(32'hba7090fd),
	.w3(32'h3b1a0cbe),
	.w4(32'h3aced126),
	.w5(32'hbac32d5c),
	.w6(32'h3ae85a98),
	.w7(32'h3ae00598),
	.w8(32'hba83de40),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9416067),
	.w1(32'hb9931346),
	.w2(32'hba8f689f),
	.w3(32'hb62e25d3),
	.w4(32'hb913f132),
	.w5(32'hba8159f1),
	.w6(32'hb8926ff5),
	.w7(32'hb9dd62fb),
	.w8(32'hbac4f1d9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad2d1d),
	.w1(32'h3a761a72),
	.w2(32'h3a97fc0f),
	.w3(32'h39d151f5),
	.w4(32'h3a6415f5),
	.w5(32'h3a9d0e7f),
	.w6(32'h3936f3e4),
	.w7(32'h39c4ebf7),
	.w8(32'h3a46a366),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a3a6c),
	.w1(32'hba300c7b),
	.w2(32'hba5ffedb),
	.w3(32'hb819e77c),
	.w4(32'hba55617d),
	.w5(32'hba06f753),
	.w6(32'h3985f6d7),
	.w7(32'hba14c7ca),
	.w8(32'hba46025f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8374b9),
	.w1(32'hba0e1c80),
	.w2(32'hbaa77b75),
	.w3(32'hba210fb1),
	.w4(32'hb9ed2968),
	.w5(32'hbaa76803),
	.w6(32'h398075e6),
	.w7(32'hb9f295ed),
	.w8(32'hba6c8f4b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fde8c),
	.w1(32'hbaa85661),
	.w2(32'h3a353a62),
	.w3(32'hbb4ab8a9),
	.w4(32'hbacd9782),
	.w5(32'h3a000d57),
	.w6(32'hbb717838),
	.w7(32'hbb0d3ff4),
	.w8(32'hb716c265),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3823445e),
	.w1(32'h3780a8e0),
	.w2(32'hb7845f6f),
	.w3(32'h37fb45de),
	.w4(32'h37d6518b),
	.w5(32'h369463b2),
	.w6(32'h380a6c3d),
	.w7(32'h37e7ad13),
	.w8(32'h3763e7a5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b3d105),
	.w1(32'h37dfc214),
	.w2(32'h37477f26),
	.w3(32'hb600da82),
	.w4(32'h365348ee),
	.w5(32'h37d384ed),
	.w6(32'h36175dfb),
	.w7(32'hb52775c8),
	.w8(32'h38050eb5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9395e86),
	.w1(32'h39d4fbc0),
	.w2(32'hb9290666),
	.w3(32'h388824a2),
	.w4(32'h393656aa),
	.w5(32'hb83ef203),
	.w6(32'hb9baaa90),
	.w7(32'hb9659202),
	.w8(32'hb96b7fb6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23a0ff),
	.w1(32'hba0c5f81),
	.w2(32'hba856c19),
	.w3(32'hba850e06),
	.w4(32'hba8991b6),
	.w5(32'hbab52945),
	.w6(32'hba61d226),
	.w7(32'hba5a3252),
	.w8(32'hba89caa4),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dc4e1),
	.w1(32'hba2a3c41),
	.w2(32'hba9c8b38),
	.w3(32'hba137a5f),
	.w4(32'hba2ffae0),
	.w5(32'hbad7cfc6),
	.w6(32'hba006b83),
	.w7(32'hba884e0c),
	.w8(32'hbb08ccea),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a487993),
	.w1(32'h3a0b6147),
	.w2(32'h39cac91c),
	.w3(32'hb90a32de),
	.w4(32'hb776ee71),
	.w5(32'h38a78eb1),
	.w6(32'h37ed86b3),
	.w7(32'h393310d9),
	.w8(32'h39cddee2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383eb7d7),
	.w1(32'hb675c39f),
	.w2(32'hb8375d55),
	.w3(32'h3887d8a5),
	.w4(32'h36876cd9),
	.w5(32'hb893a226),
	.w6(32'h3884f215),
	.w7(32'h3872f58b),
	.w8(32'hb7f92e32),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4c8f6),
	.w1(32'h3697b46f),
	.w2(32'h37851c28),
	.w3(32'hb898bef8),
	.w4(32'hb6eb22e0),
	.w5(32'h37c40071),
	.w6(32'hb8bbb549),
	.w7(32'h36a1cf85),
	.w8(32'h389075da),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f24029),
	.w1(32'h3a14dc74),
	.w2(32'hb92dc23e),
	.w3(32'hba26fd5a),
	.w4(32'hb8c78566),
	.w5(32'h397c1a51),
	.w6(32'hba2e4da8),
	.w7(32'h37cf03f5),
	.w8(32'h3a834370),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cf098),
	.w1(32'hbb390d5b),
	.w2(32'hbadafe9d),
	.w3(32'hbb259850),
	.w4(32'hbb116a5d),
	.w5(32'hbaa32419),
	.w6(32'hbb009060),
	.w7(32'hbae353d2),
	.w8(32'hb967cefe),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e777b7),
	.w1(32'hb85fc2cf),
	.w2(32'hbaeab7fb),
	.w3(32'h3936e884),
	.w4(32'hba6f9e2e),
	.w5(32'hba9714fc),
	.w6(32'h3a0ef3cf),
	.w7(32'hb97add65),
	.w8(32'hbaa3031a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fdcb0),
	.w1(32'h3aac4dba),
	.w2(32'hb89042ae),
	.w3(32'h3ad11a0d),
	.w4(32'h3aab71ec),
	.w5(32'h3933be99),
	.w6(32'h3a80988f),
	.w7(32'h3aa214bd),
	.w8(32'hb800b7db),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bad8e),
	.w1(32'hba441536),
	.w2(32'h3a080333),
	.w3(32'hbae19da4),
	.w4(32'hb9d75305),
	.w5(32'h3a55851e),
	.w6(32'hbafb33b4),
	.w7(32'hba90f341),
	.w8(32'h390a38bb),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379ddcaf),
	.w1(32'h374703cc),
	.w2(32'h373f8812),
	.w3(32'h370436d6),
	.w4(32'h3619d5ec),
	.w5(32'h368611f3),
	.w6(32'h37472da7),
	.w7(32'h3723e78b),
	.w8(32'h37214288),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e77e6a),
	.w1(32'hb6b076e3),
	.w2(32'h37547332),
	.w3(32'hb7056c19),
	.w4(32'hb6873727),
	.w5(32'h377d4215),
	.w6(32'hb61e2f75),
	.w7(32'hb2a5a32b),
	.w8(32'h378682ec),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3764289a),
	.w1(32'h38a505ec),
	.w2(32'h388ffe03),
	.w3(32'h384a9546),
	.w4(32'h37791a55),
	.w5(32'h35a20394),
	.w6(32'h38724508),
	.w7(32'h382fe8f2),
	.w8(32'h383766e3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367e59de),
	.w1(32'h36e1f00b),
	.w2(32'h37207f46),
	.w3(32'hb69aa369),
	.w4(32'h35aebe91),
	.w5(32'h3729878b),
	.w6(32'h37897c4f),
	.w7(32'h37856a9d),
	.w8(32'h37cd244f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85ce1f6),
	.w1(32'h39c69f37),
	.w2(32'h389b976b),
	.w3(32'hb6a3b2df),
	.w4(32'h39938c40),
	.w5(32'h3965dd11),
	.w6(32'hb89865b4),
	.w7(32'h38d1e3ac),
	.w8(32'h391334c1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba221b52),
	.w1(32'hb99f26d6),
	.w2(32'hba29645f),
	.w3(32'hba8208c6),
	.w4(32'hba718492),
	.w5(32'hba894838),
	.w6(32'hba6fa5f7),
	.w7(32'hba89e01a),
	.w8(32'hbad20924),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f08c3c),
	.w1(32'hba0a32ac),
	.w2(32'hba4fead8),
	.w3(32'hba1d9a05),
	.w4(32'hba0d3400),
	.w5(32'hba666a30),
	.w6(32'hba12df5e),
	.w7(32'hba52b89c),
	.w8(32'hbaa7f340),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64be65f),
	.w1(32'h37be3908),
	.w2(32'h37e81bba),
	.w3(32'hb6bd6127),
	.w4(32'h37e6611c),
	.w5(32'h380b4103),
	.w6(32'hb74e9529),
	.w7(32'h37ed7def),
	.w8(32'h3802c0f1),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bc37d),
	.w1(32'h367f37e0),
	.w2(32'hbb0a2931),
	.w3(32'hbad7a0cb),
	.w4(32'hba9dce03),
	.w5(32'hba3b9525),
	.w6(32'hba4f7694),
	.w7(32'hba4de1d6),
	.w8(32'hb931d748),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7df947b),
	.w1(32'hba05719b),
	.w2(32'hba5056b9),
	.w3(32'hb8e85f36),
	.w4(32'hb9dca1a5),
	.w5(32'hba47e963),
	.w6(32'hb7928cf6),
	.w7(32'hb95b6719),
	.w8(32'hba0f04d8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb824e0b2),
	.w1(32'hb895e3e5),
	.w2(32'h37814ca1),
	.w3(32'hb7ca676a),
	.w4(32'hb88207c9),
	.w5(32'h36ba9729),
	.w6(32'h3804a766),
	.w7(32'hb80c1f10),
	.w8(32'h373964c7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f99b3b),
	.w1(32'hb8116528),
	.w2(32'hb9d04f57),
	.w3(32'hba1acdb6),
	.w4(32'hb91ef25e),
	.w5(32'hb98ebcd6),
	.w6(32'hb9d6454f),
	.w7(32'hb910dd0a),
	.w8(32'hb9014b26),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b4c19),
	.w1(32'h38ebd8a6),
	.w2(32'h387ea15f),
	.w3(32'h39462f58),
	.w4(32'h38d05181),
	.w5(32'h38615e66),
	.w6(32'h390eb12e),
	.w7(32'h38019547),
	.w8(32'h3784914d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38438382),
	.w1(32'h393ebcc6),
	.w2(32'h37a48156),
	.w3(32'h360d5f48),
	.w4(32'h3965d931),
	.w5(32'h389a8ef9),
	.w6(32'h389ff791),
	.w7(32'h3947ad86),
	.w8(32'h394e73ea),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379214d9),
	.w1(32'h3700eb9d),
	.w2(32'h3716deff),
	.w3(32'h35de33a9),
	.w4(32'hb6cbff53),
	.w5(32'h3722f29d),
	.w6(32'h36d15e6c),
	.w7(32'h366dd5fb),
	.w8(32'h365099ba),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384241fb),
	.w1(32'h380edc7d),
	.w2(32'h37669bbb),
	.w3(32'h379fabc7),
	.w4(32'hb6245c5a),
	.w5(32'hb70e12d7),
	.w6(32'h3768dbb0),
	.w7(32'h36cb230b),
	.w8(32'hb623ad85),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37defc15),
	.w1(32'h3a364900),
	.w2(32'h3a2fbb28),
	.w3(32'h378ed470),
	.w4(32'h39c91fcf),
	.w5(32'h3a04e482),
	.w6(32'hba092e65),
	.w7(32'hb8d92165),
	.w8(32'hb7fdd97b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388114c7),
	.w1(32'hb9985d52),
	.w2(32'hba9953d5),
	.w3(32'hb99366ce),
	.w4(32'hba07487b),
	.w5(32'hbacbf7ae),
	.w6(32'hb901eebf),
	.w7(32'hba5c5fe0),
	.w8(32'hbafa629e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bea588),
	.w1(32'hb9d69fe8),
	.w2(32'hbaa5f6cb),
	.w3(32'hb98b11fb),
	.w4(32'hb9f014b0),
	.w5(32'hbab42684),
	.w6(32'hb9998d23),
	.w7(32'hba30a80d),
	.w8(32'hbaa385aa),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f5718),
	.w1(32'hbb31932f),
	.w2(32'hbb0d016f),
	.w3(32'hbb47f66f),
	.w4(32'hbb36eac3),
	.w5(32'hbb02bed5),
	.w6(32'hbb08ec97),
	.w7(32'hbb157d19),
	.w8(32'hbadd6e05),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38abacb6),
	.w1(32'h384bb292),
	.w2(32'hb6cdff45),
	.w3(32'h384fdeb8),
	.w4(32'h38870c06),
	.w5(32'h33331f16),
	.w6(32'h38590bb4),
	.w7(32'h38ad7bc7),
	.w8(32'h37d42fb0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38058ce9),
	.w1(32'hb5a48227),
	.w2(32'hb8231ec2),
	.w3(32'h37d3049d),
	.w4(32'hb6a42a7c),
	.w5(32'hb8681ee9),
	.w6(32'h37883614),
	.w7(32'hb71df3d7),
	.w8(32'hb8590af8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb824f96b),
	.w1(32'h3827f3c7),
	.w2(32'h37bde49e),
	.w3(32'hb77cfe20),
	.w4(32'h382207ce),
	.w5(32'h381d1007),
	.w6(32'hb78b91df),
	.w7(32'h37a89aa2),
	.w8(32'h383b75d2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb684726d),
	.w1(32'h3729f6f7),
	.w2(32'h35a65721),
	.w3(32'h37a50c26),
	.w4(32'h37910285),
	.w5(32'h37a2b072),
	.w6(32'h37bcefe3),
	.w7(32'h373f22f5),
	.w8(32'h37644a15),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3971a7),
	.w1(32'hb9085557),
	.w2(32'hbaec75a7),
	.w3(32'h3a535b10),
	.w4(32'hb98262f6),
	.w5(32'hbb04eb37),
	.w6(32'h3a76cda3),
	.w7(32'h374f464a),
	.w8(32'hbae6b6e8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a87506),
	.w1(32'h36d4de09),
	.w2(32'hb857c9a8),
	.w3(32'hb91bddd7),
	.w4(32'h3800345f),
	.w5(32'hb8da948e),
	.w6(32'hb8c18297),
	.w7(32'hb8ae01a7),
	.w8(32'hb9545b67),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eaaba2),
	.w1(32'h39ebafb3),
	.w2(32'h3950e1c9),
	.w3(32'h3a005ba9),
	.w4(32'h39d5743c),
	.w5(32'h398c82c1),
	.w6(32'h3a0ec1d0),
	.w7(32'h39e5029a),
	.w8(32'h391b052c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39629763),
	.w1(32'h39dccb68),
	.w2(32'h39c65ccd),
	.w3(32'h39be3a78),
	.w4(32'h39d67dc2),
	.w5(32'h39f928fa),
	.w6(32'h3952d8d0),
	.w7(32'h3981d8f6),
	.w8(32'h39a07ca9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3824e593),
	.w1(32'h37b859e4),
	.w2(32'h37d42351),
	.w3(32'h38677c10),
	.w4(32'h36d21d4c),
	.w5(32'h3828851a),
	.w6(32'h37b8e92b),
	.w7(32'hb7f8b153),
	.w8(32'h381f6ede),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba004784),
	.w1(32'hba626e41),
	.w2(32'hb99f7219),
	.w3(32'hba23e031),
	.w4(32'hba4be35b),
	.w5(32'hb9f57129),
	.w6(32'hba0ac150),
	.w7(32'hba22f916),
	.w8(32'hba0fa1a7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3850cbb4),
	.w1(32'h3891984c),
	.w2(32'h3793bf34),
	.w3(32'h38665326),
	.w4(32'h3885a210),
	.w5(32'h381fbfb7),
	.w6(32'h38513b7f),
	.w7(32'h38991b17),
	.w8(32'h3883d6c0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d69a7a),
	.w1(32'hbaae97a0),
	.w2(32'hbb1d6ffe),
	.w3(32'hb9058ca7),
	.w4(32'hba79f8f5),
	.w5(32'hbb1da7b4),
	.w6(32'hb886a79b),
	.w7(32'hba95acee),
	.w8(32'hbb076101),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a53d0),
	.w1(32'h37bc6603),
	.w2(32'h375a915f),
	.w3(32'h387ffd28),
	.w4(32'hb4b1db24),
	.w5(32'hb844cc79),
	.w6(32'hb680931c),
	.w7(32'hb8671fd3),
	.w8(32'hb8a4f808),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acea54d),
	.w1(32'h3ad8dcd7),
	.w2(32'h3ad4a387),
	.w3(32'h3af214ab),
	.w4(32'h3af8ad2d),
	.w5(32'h39d7431e),
	.w6(32'h39a03faf),
	.w7(32'h3aa9531a),
	.w8(32'hb91303f2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule