module layer_10_featuremap_331(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a6b46),
	.w1(32'hba6b6776),
	.w2(32'hba1f446f),
	.w3(32'hbacf9f3c),
	.w4(32'hb98d2e7d),
	.w5(32'h3b00912b),
	.w6(32'hbb216598),
	.w7(32'hba57bd0f),
	.w8(32'h3a5f8c18),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5431c),
	.w1(32'hb9a5d564),
	.w2(32'h398e8001),
	.w3(32'h3ac66a8a),
	.w4(32'h3a1d854e),
	.w5(32'hba57ae34),
	.w6(32'h39425b0f),
	.w7(32'hba6082f6),
	.w8(32'hbae9e1d8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82b37a),
	.w1(32'h3a504ec6),
	.w2(32'h3a7f76fa),
	.w3(32'h39b21ed7),
	.w4(32'h3a55aded),
	.w5(32'hb93e68d6),
	.w6(32'hb7a3d6a9),
	.w7(32'h3a04d511),
	.w8(32'h39fbd052),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b9057),
	.w1(32'hb91ed7ec),
	.w2(32'hb84225e8),
	.w3(32'h37a7f0cb),
	.w4(32'hba859d08),
	.w5(32'hb9587b6d),
	.w6(32'h3a9fdbce),
	.w7(32'hba129071),
	.w8(32'h3a592adb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcae8e),
	.w1(32'hb90f17b7),
	.w2(32'h3b15ce3f),
	.w3(32'hbb1328bb),
	.w4(32'hba384f99),
	.w5(32'hb6f295ba),
	.w6(32'hb9af00d3),
	.w7(32'h3b0cec6a),
	.w8(32'h39501832),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb970ef0d),
	.w1(32'hba39dafa),
	.w2(32'hba271665),
	.w3(32'hba703f03),
	.w4(32'hba8b065f),
	.w5(32'h39c1aed7),
	.w6(32'h399e6904),
	.w7(32'hba5d72c3),
	.w8(32'hba6d47c1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba595fa8),
	.w1(32'hb989a3ac),
	.w2(32'h3a20dbc4),
	.w3(32'hba68359f),
	.w4(32'hb9615bd7),
	.w5(32'hbb05cadb),
	.w6(32'hb95f6f5c),
	.w7(32'hba116532),
	.w8(32'hbafa6ff5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb033f32),
	.w1(32'hbb2bfe1f),
	.w2(32'hbb048007),
	.w3(32'hbb0bb658),
	.w4(32'hba5963e9),
	.w5(32'hba30aa82),
	.w6(32'hbafd3776),
	.w7(32'hbaed680e),
	.w8(32'hbaa176e3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcb4b5),
	.w1(32'hba2235ef),
	.w2(32'hb81aceae),
	.w3(32'hba892a09),
	.w4(32'h3971827e),
	.w5(32'h3a0667b4),
	.w6(32'hbaa26182),
	.w7(32'hba205902),
	.w8(32'h3a3b9377),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96543d2),
	.w1(32'hba2feb01),
	.w2(32'hbb3f28e5),
	.w3(32'hba03de1b),
	.w4(32'hbab375e8),
	.w5(32'hbb35f992),
	.w6(32'hb955496c),
	.w7(32'hba304163),
	.w8(32'hbad12967),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a9a5c),
	.w1(32'h3a03d972),
	.w2(32'h3a98d7b1),
	.w3(32'h396dcdb4),
	.w4(32'h3a0563e9),
	.w5(32'h3ad21c83),
	.w6(32'h3a95d529),
	.w7(32'hba18bfe7),
	.w8(32'h3a40283d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5f4ae),
	.w1(32'h3a799258),
	.w2(32'hba6c88e9),
	.w3(32'h3aa8311f),
	.w4(32'h3b28f363),
	.w5(32'h39b6ee5a),
	.w6(32'h392ee5ed),
	.w7(32'h3a75558b),
	.w8(32'h3a6b3506),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a6b14),
	.w1(32'h3ada94ca),
	.w2(32'hba7d250c),
	.w3(32'h38495b94),
	.w4(32'h3a32fd39),
	.w5(32'hbb1a513d),
	.w6(32'hb9b95a46),
	.w7(32'h3a3718c8),
	.w8(32'hbac14768),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba998f9a),
	.w1(32'hbae3ea42),
	.w2(32'hba40aad1),
	.w3(32'hba40e34b),
	.w4(32'hba09107c),
	.w5(32'hb6f1c688),
	.w6(32'hb9f6cd69),
	.w7(32'h3aa739bb),
	.w8(32'h3a4af352),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a835b1f),
	.w1(32'hb7f70476),
	.w2(32'hba6e7fa4),
	.w3(32'h3a4d897e),
	.w4(32'h3a9a34eb),
	.w5(32'h3a03ffe1),
	.w6(32'h3a0ed048),
	.w7(32'hb94784f7),
	.w8(32'hb93ac48e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9480e02),
	.w1(32'hba7e000d),
	.w2(32'hbb29f3b5),
	.w3(32'h3893f9f5),
	.w4(32'hba8d643f),
	.w5(32'hbb580929),
	.w6(32'h3a1e2b6c),
	.w7(32'hba0ad023),
	.w8(32'hbb5dc721),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a3d16),
	.w1(32'hbb324295),
	.w2(32'hbb220a7e),
	.w3(32'hba2cf542),
	.w4(32'hba990288),
	.w5(32'hbad18937),
	.w6(32'hba518537),
	.w7(32'hbb3f1328),
	.w8(32'hba5bac00),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a12247),
	.w1(32'h389fb0c5),
	.w2(32'hbb159839),
	.w3(32'hbb03ee51),
	.w4(32'hbaf06155),
	.w5(32'hba8cdf2c),
	.w6(32'hbafff778),
	.w7(32'hba36bcaa),
	.w8(32'h3a603133),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940b158),
	.w1(32'hba0ac054),
	.w2(32'hbae44bc3),
	.w3(32'hbb16b47d),
	.w4(32'hba345ad0),
	.w5(32'hba9b6666),
	.w6(32'h3a4af512),
	.w7(32'h3b100607),
	.w8(32'hbaaa6a4a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7b646),
	.w1(32'h38566f6a),
	.w2(32'hb8ae9bfc),
	.w3(32'hba429e40),
	.w4(32'hb7d5cf46),
	.w5(32'h3adafd94),
	.w6(32'hbad607ba),
	.w7(32'hba0363ea),
	.w8(32'h3a0a91aa),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1871e5),
	.w1(32'h3a742c05),
	.w2(32'h3a8009fd),
	.w3(32'h3aa53967),
	.w4(32'h39d02aa2),
	.w5(32'h399e6f49),
	.w6(32'h3adb8592),
	.w7(32'h3a95b6a7),
	.w8(32'h3944cfb2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb80ad),
	.w1(32'hb899142e),
	.w2(32'hb9bfb48f),
	.w3(32'hb95e81f9),
	.w4(32'h391e8e03),
	.w5(32'hb9bbaef3),
	.w6(32'hb9ee0a4a),
	.w7(32'hb9a08221),
	.w8(32'hba44d4c3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38683180),
	.w1(32'hba8549df),
	.w2(32'hbb81b36b),
	.w3(32'hbb4ed678),
	.w4(32'hbb89bdd6),
	.w5(32'hbb679002),
	.w6(32'hbb9f8e42),
	.w7(32'hbb875ff6),
	.w8(32'hbaf19df4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2588da),
	.w1(32'hba94b500),
	.w2(32'hbb02055f),
	.w3(32'hba0ab0d5),
	.w4(32'hbac1b0a0),
	.w5(32'hbb05e70e),
	.w6(32'hbab98e31),
	.w7(32'hb9754f52),
	.w8(32'h3a081153),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb14a0),
	.w1(32'h3ad06e42),
	.w2(32'h39a25fa8),
	.w3(32'hbad0abb9),
	.w4(32'hb98239ec),
	.w5(32'hbb195480),
	.w6(32'h3a8c6f40),
	.w7(32'h3af4bff2),
	.w8(32'hbb1a766d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c285d),
	.w1(32'h39148b61),
	.w2(32'h386efe73),
	.w3(32'h388d2bd7),
	.w4(32'h39c71529),
	.w5(32'hbabbfd31),
	.w6(32'h3a7a188d),
	.w7(32'hba431745),
	.w8(32'hbad6c4a1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac93163),
	.w1(32'hbb3a422c),
	.w2(32'hbaea8c26),
	.w3(32'hbae27308),
	.w4(32'hbad3426d),
	.w5(32'hbacd9569),
	.w6(32'hbae862c8),
	.w7(32'hbafdc353),
	.w8(32'hbb05ac80),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4e62f),
	.w1(32'hbae3ea56),
	.w2(32'hbacec295),
	.w3(32'hbb2d09dc),
	.w4(32'hba8e7915),
	.w5(32'hba23e548),
	.w6(32'hbb32b316),
	.w7(32'hbad91e38),
	.w8(32'hba11e588),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba213174),
	.w1(32'hba41bb84),
	.w2(32'hbafdf127),
	.w3(32'h39f48d06),
	.w4(32'hbb0727cc),
	.w5(32'hbb32d3d1),
	.w6(32'hb986f0bd),
	.w7(32'hba5b6f14),
	.w8(32'hbb1fccc7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95510c),
	.w1(32'hbb0a1dbb),
	.w2(32'hbb5a46c7),
	.w3(32'hbaea79ca),
	.w4(32'hba6e12bb),
	.w5(32'hbb084029),
	.w6(32'hbb0f0b7b),
	.w7(32'h39336abc),
	.w8(32'hb8bb6689),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a874a59),
	.w1(32'h3aafe860),
	.w2(32'h3a770858),
	.w3(32'h399d43f1),
	.w4(32'hb7f67c92),
	.w5(32'h3b12e35c),
	.w6(32'h3b2a6ecf),
	.w7(32'h39a95ae1),
	.w8(32'h3a70575a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e7208),
	.w1(32'h389110dc),
	.w2(32'hb9c1b250),
	.w3(32'h3b6ca38e),
	.w4(32'h3af5b8e3),
	.w5(32'hb9fd3dbc),
	.w6(32'h39aed926),
	.w7(32'hbaad1f5d),
	.w8(32'h3ada581e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51884e),
	.w1(32'hb9ae5681),
	.w2(32'hb877009c),
	.w3(32'hb9d32a52),
	.w4(32'hb9c5802c),
	.w5(32'hbb62e12c),
	.w6(32'hba43d64c),
	.w7(32'hb9665b62),
	.w8(32'hbb3b4338),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2def1),
	.w1(32'h3844c0b7),
	.w2(32'hba9c62d1),
	.w3(32'hbadfc09b),
	.w4(32'hbb33b8f8),
	.w5(32'hba818196),
	.w6(32'hbaa312e1),
	.w7(32'hbabb0ac6),
	.w8(32'h3a3fc2ed),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7032ef),
	.w1(32'h3a1197b7),
	.w2(32'h3a6eee33),
	.w3(32'hbad72fef),
	.w4(32'hbaba84ff),
	.w5(32'hba84599a),
	.w6(32'h3a29e16e),
	.w7(32'hb822ab97),
	.w8(32'hba704171),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c66d47),
	.w1(32'h3a31e8e1),
	.w2(32'h3a3801c0),
	.w3(32'hbb1bd9cb),
	.w4(32'hbaa7264a),
	.w5(32'hb7ae01df),
	.w6(32'hba82dc97),
	.w7(32'h3995037f),
	.w8(32'hbab6d863),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7a697),
	.w1(32'h3a6b7729),
	.w2(32'h3aa82ec6),
	.w3(32'h3ae29f7c),
	.w4(32'h3a7d7c63),
	.w5(32'hb8a9c4aa),
	.w6(32'hbab6721b),
	.w7(32'hb96267ad),
	.w8(32'h3a82e370),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b196644),
	.w1(32'h3b095eff),
	.w2(32'h3ab9bcde),
	.w3(32'h38f40a83),
	.w4(32'h3af71fa1),
	.w5(32'h3975bd7d),
	.w6(32'h3aa04ba1),
	.w7(32'hb9dab4d4),
	.w8(32'hbb57076c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa80e2d),
	.w1(32'h3b2fd46e),
	.w2(32'hba0d9620),
	.w3(32'h3b30c8a5),
	.w4(32'h3b0098be),
	.w5(32'hbb592f5f),
	.w6(32'h3aa0b40f),
	.w7(32'h3a34d709),
	.w8(32'hbb05d0a7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac21832),
	.w1(32'hbb048ddd),
	.w2(32'hbb0483cb),
	.w3(32'hbad8761c),
	.w4(32'hbb0b7d92),
	.w5(32'hba8ee01d),
	.w6(32'hb90eacb4),
	.w7(32'hb9c61177),
	.w8(32'hba6408d9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba686d0f),
	.w1(32'hbabf82c4),
	.w2(32'hba88bfe4),
	.w3(32'h3a28d86c),
	.w4(32'h3a320593),
	.w5(32'hba84ead7),
	.w6(32'hba2700a1),
	.w7(32'hb9ac849c),
	.w8(32'hbacdef04),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaae40e),
	.w1(32'hba64661b),
	.w2(32'hb90fb262),
	.w3(32'h3987165d),
	.w4(32'hb9499728),
	.w5(32'h3aa5e057),
	.w6(32'h3ac4f3e2),
	.w7(32'hba35068f),
	.w8(32'h3b138d5c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88746a),
	.w1(32'h3b0d597f),
	.w2(32'h3b2a2b72),
	.w3(32'h3b123c5d),
	.w4(32'h3b7e2d4c),
	.w5(32'hbb415411),
	.w6(32'h3b67ddd5),
	.w7(32'h3bb4b54f),
	.w8(32'hbaf605ef),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1f5d),
	.w1(32'hbbac44af),
	.w2(32'hbb8ad707),
	.w3(32'hbb42f029),
	.w4(32'hbacd28fa),
	.w5(32'hbbb5363c),
	.w6(32'h3ab9bc66),
	.w7(32'hba518822),
	.w8(32'hbb94b32c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961b347),
	.w1(32'h386fa865),
	.w2(32'hbb2d0c1a),
	.w3(32'hbaff17ef),
	.w4(32'hbb2671fd),
	.w5(32'hbb77f252),
	.w6(32'hbb19d921),
	.w7(32'hbaf73c30),
	.w8(32'hbb89941d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61bd81),
	.w1(32'hbadb51d3),
	.w2(32'hbb9df0ec),
	.w3(32'h38ed7322),
	.w4(32'hbae2caf0),
	.w5(32'hbb406822),
	.w6(32'h3a0221a3),
	.w7(32'hbaec739e),
	.w8(32'hbb4414ac),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3416d8fe),
	.w1(32'hb891f6b8),
	.w2(32'hbb1d70d1),
	.w3(32'h3a106647),
	.w4(32'h3a0dcc5d),
	.w5(32'h3a92d2c9),
	.w6(32'h3a777d58),
	.w7(32'h3a3bd300),
	.w8(32'h3a6c69b1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5777e),
	.w1(32'hbaac1586),
	.w2(32'hbae109b0),
	.w3(32'hbb0069cd),
	.w4(32'hb94cb18e),
	.w5(32'h396b6aaa),
	.w6(32'hbb5dbfb8),
	.w7(32'hba9f3807),
	.w8(32'h39d9122e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac788ac),
	.w1(32'h3a6e420e),
	.w2(32'h39fe189a),
	.w3(32'h393f824c),
	.w4(32'h3a716b77),
	.w5(32'h3a6479fa),
	.w6(32'hb99ccc8b),
	.w7(32'h39a97160),
	.w8(32'h3a1c2bc6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39249119),
	.w1(32'h38debb42),
	.w2(32'h3a732d1f),
	.w3(32'h39859392),
	.w4(32'h3a415c13),
	.w5(32'hba2f9008),
	.w6(32'hb79311a4),
	.w7(32'h39555ceb),
	.w8(32'h3a4cdcd5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64d5e1),
	.w1(32'h3aa9235f),
	.w2(32'h3afdb0fb),
	.w3(32'h3938ba01),
	.w4(32'hba826ad3),
	.w5(32'hbaaaad46),
	.w6(32'h3af25516),
	.w7(32'h3ae665be),
	.w8(32'hb9c937fc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08d826),
	.w1(32'h392a0d68),
	.w2(32'hba16fb52),
	.w3(32'hba85cda9),
	.w4(32'hba881b66),
	.w5(32'hbac0e609),
	.w6(32'h3adb81e6),
	.w7(32'h3a0b24a1),
	.w8(32'hbad49177),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc1566),
	.w1(32'hbaa20c2f),
	.w2(32'hbab52b38),
	.w3(32'h39dedb5d),
	.w4(32'h393367c6),
	.w5(32'hbadfd46c),
	.w6(32'h3a54cae1),
	.w7(32'hba0c77fb),
	.w8(32'hba9e8558),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27e115),
	.w1(32'hbadc588c),
	.w2(32'hba7d1a5f),
	.w3(32'hbb63a058),
	.w4(32'hba8c2324),
	.w5(32'h3a88bc2d),
	.w6(32'hbb674e31),
	.w7(32'hb9a9d62f),
	.w8(32'h3a82e871),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a761782),
	.w1(32'h3a846994),
	.w2(32'hb8aed55a),
	.w3(32'h3aa905a3),
	.w4(32'h3b0f65fc),
	.w5(32'hbb0f2cc4),
	.w6(32'h3a6eebeb),
	.w7(32'h3a116cf2),
	.w8(32'h3923a8ab),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71dd17),
	.w1(32'h3a073e01),
	.w2(32'h39701001),
	.w3(32'hbb4792e8),
	.w4(32'hbb3ddb94),
	.w5(32'hbaa8929f),
	.w6(32'hb93c936a),
	.w7(32'hbaa7dfca),
	.w8(32'hba738c3c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1c2e9),
	.w1(32'hba10b7dd),
	.w2(32'hba4a75a5),
	.w3(32'hba009d6f),
	.w4(32'h39557fb7),
	.w5(32'hba3d5684),
	.w6(32'hba91cdaf),
	.w7(32'hba0097cf),
	.w8(32'hb938f2c4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074221),
	.w1(32'hba99429a),
	.w2(32'hb8fa4927),
	.w3(32'hba02d3c4),
	.w4(32'hba186c5b),
	.w5(32'h3a0a4e44),
	.w6(32'h39e02096),
	.w7(32'hb8a8e774),
	.w8(32'hb9cebcd8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce67b5),
	.w1(32'h395a4711),
	.w2(32'h3a8439c1),
	.w3(32'h3969adae),
	.w4(32'h3a622c03),
	.w5(32'h3affb0ec),
	.w6(32'h391ec167),
	.w7(32'h38a56927),
	.w8(32'h3b00e35d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9be4ff),
	.w1(32'h3aa5dfd3),
	.w2(32'hb870292a),
	.w3(32'h3a852065),
	.w4(32'h3adddda6),
	.w5(32'h3912ab33),
	.w6(32'h3b338b87),
	.w7(32'h3a560aae),
	.w8(32'hb8a983fa),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad3675),
	.w1(32'h3a1ac525),
	.w2(32'hb9342d4f),
	.w3(32'h3acf7a79),
	.w4(32'h396666cb),
	.w5(32'hb9dc6226),
	.w6(32'h3ac5b6c8),
	.w7(32'h392934a0),
	.w8(32'hbaa3b699),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c88bf),
	.w1(32'h3aca6cce),
	.w2(32'h39289ac0),
	.w3(32'h3b37ebad),
	.w4(32'h3a73d50f),
	.w5(32'hb9711b58),
	.w6(32'h3b58ec02),
	.w7(32'hb94bfa03),
	.w8(32'h3b0c16c6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b115bf3),
	.w1(32'h3a9bf5bf),
	.w2(32'h3b024ede),
	.w3(32'hbb1289e5),
	.w4(32'hbad3d96f),
	.w5(32'hbaf56837),
	.w6(32'h3b4ac764),
	.w7(32'h3b04d5af),
	.w8(32'hbaadc1a6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952b102),
	.w1(32'hba8ff509),
	.w2(32'hba852dc5),
	.w3(32'hbad31e6c),
	.w4(32'hbae53c5e),
	.w5(32'hb9b8488d),
	.w6(32'hbb0e7774),
	.w7(32'hbb179513),
	.w8(32'hb820421e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38273e4b),
	.w1(32'hba83248d),
	.w2(32'hba8210e1),
	.w3(32'hbabaf15d),
	.w4(32'hba7f33d1),
	.w5(32'h3ae892f6),
	.w6(32'hb98822bc),
	.w7(32'hba9f4d42),
	.w8(32'h3a8f992b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9329829),
	.w1(32'hba0505d7),
	.w2(32'hba151a3e),
	.w3(32'h3a97f9f1),
	.w4(32'h3ae4b484),
	.w5(32'hb9a2ee4d),
	.w6(32'h3aeeb90b),
	.w7(32'h3813399e),
	.w8(32'hb9c503f2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac70a1b),
	.w1(32'hbaa910b2),
	.w2(32'hba8abfe1),
	.w3(32'hbada3647),
	.w4(32'hba55d096),
	.w5(32'hbae5a146),
	.w6(32'h394c9fe6),
	.w7(32'hba7ab3f0),
	.w8(32'hbad1b0b8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d7d33),
	.w1(32'hba80617b),
	.w2(32'hbad60af7),
	.w3(32'hbae4b9d3),
	.w4(32'h3a31ed10),
	.w5(32'hbadc0a4b),
	.w6(32'hbaa7733e),
	.w7(32'hba7a54f1),
	.w8(32'hbadd8213),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389eb220),
	.w1(32'h3a1cff14),
	.w2(32'hba27b962),
	.w3(32'h39a6d899),
	.w4(32'h3a8d3551),
	.w5(32'hbb4e1945),
	.w6(32'hba97f8f0),
	.w7(32'h39b99132),
	.w8(32'hbb2f0568),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91109f),
	.w1(32'hba7302f1),
	.w2(32'hbb1c0cb8),
	.w3(32'hbade64d1),
	.w4(32'h38cade7b),
	.w5(32'hba8e47c1),
	.w6(32'h3925fcf3),
	.w7(32'h3a09058a),
	.w8(32'hba5b38a3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa15058),
	.w1(32'h3a053521),
	.w2(32'h3aad8a57),
	.w3(32'h3a833112),
	.w4(32'h3ab0235a),
	.w5(32'hb84fa671),
	.w6(32'hba31f2b5),
	.w7(32'h39abe4ec),
	.w8(32'h37d6a4a0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5219ab),
	.w1(32'hba0089ea),
	.w2(32'h3a8364a0),
	.w3(32'h36e5efbd),
	.w4(32'h385fe6c8),
	.w5(32'h3a3d2af8),
	.w6(32'hba16d1c9),
	.w7(32'hb7d99745),
	.w8(32'h3a1898da),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9f493),
	.w1(32'h3b3351ff),
	.w2(32'h3af2b275),
	.w3(32'h3b256a77),
	.w4(32'h3aa19116),
	.w5(32'h39611058),
	.w6(32'h392ae640),
	.w7(32'hbaa218af),
	.w8(32'h3a6ce02f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01bf3f),
	.w1(32'h3967fe99),
	.w2(32'h3a7614e5),
	.w3(32'h3a757961),
	.w4(32'h3b163ddc),
	.w5(32'h3adca303),
	.w6(32'hb8ab09ef),
	.w7(32'h3b0d6532),
	.w8(32'h3abd31ba),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3957b69b),
	.w1(32'h38b748bc),
	.w2(32'h39c9358a),
	.w3(32'h39e488df),
	.w4(32'h3a2961fe),
	.w5(32'h3a126a18),
	.w6(32'h3ac0ce8c),
	.w7(32'h3a4c7f4b),
	.w8(32'h3ad817ed),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad54278),
	.w1(32'h3b01a048),
	.w2(32'h3aa078d7),
	.w3(32'hb9e56f1c),
	.w4(32'h3a0779f0),
	.w5(32'hba8f64ae),
	.w6(32'h39ed5951),
	.w7(32'h3ae49b00),
	.w8(32'hba442c5e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6659e0),
	.w1(32'hbaa976d2),
	.w2(32'hbabb343e),
	.w3(32'hbb0c4c1f),
	.w4(32'hbb11564d),
	.w5(32'hbb742ee4),
	.w6(32'hbb24076b),
	.w7(32'hbb1a60ef),
	.w8(32'hbb6a741f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57f2ee),
	.w1(32'hbaa23c87),
	.w2(32'hbac4c91f),
	.w3(32'hbb4a360c),
	.w4(32'hbb605aae),
	.w5(32'hbabf8dd7),
	.w6(32'hbab42475),
	.w7(32'hbaa831e8),
	.w8(32'h3a541eb7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c7fd8),
	.w1(32'h3ac864ce),
	.w2(32'hba6da2f4),
	.w3(32'h3a8a1bd5),
	.w4(32'hb9c378af),
	.w5(32'h3955f1eb),
	.w6(32'h3aeefae2),
	.w7(32'h3a34a1e5),
	.w8(32'hb7a2d7cd),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba843f45),
	.w1(32'hb96f359c),
	.w2(32'hba998506),
	.w3(32'hba85498a),
	.w4(32'hba715f46),
	.w5(32'h3b6707c1),
	.w6(32'hba0171f7),
	.w7(32'hbb16da5a),
	.w8(32'h3b9d9c17),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b785),
	.w1(32'h3b5b6043),
	.w2(32'h3b05f27a),
	.w3(32'h3ba90ccb),
	.w4(32'h3bbaa82a),
	.w5(32'hba098fc9),
	.w6(32'h3b901da8),
	.w7(32'h3bb0f9a9),
	.w8(32'h399f3ede),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb975c377),
	.w1(32'h3a314bc3),
	.w2(32'hb995651e),
	.w3(32'hb9e7f344),
	.w4(32'hb8a95297),
	.w5(32'hbaaff8b4),
	.w6(32'h3991da43),
	.w7(32'h3ae74dbe),
	.w8(32'hbab4b4ba),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f64c5),
	.w1(32'h3ae83c22),
	.w2(32'h3ae81024),
	.w3(32'h38aac9d0),
	.w4(32'h35edb871),
	.w5(32'h3a4ea67b),
	.w6(32'hb86772ed),
	.w7(32'h3a43cada),
	.w8(32'h3b10f4a8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2dfc1),
	.w1(32'hba46bc58),
	.w2(32'h39aaaf66),
	.w3(32'h390ff358),
	.w4(32'hb9c61f41),
	.w5(32'hb9829db3),
	.w6(32'h3aa3a31b),
	.w7(32'h3ace8c20),
	.w8(32'hb9c264cf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af70061),
	.w1(32'h3b273f56),
	.w2(32'h3b295779),
	.w3(32'hba531643),
	.w4(32'hb8a1af13),
	.w5(32'hb9e6d315),
	.w6(32'h387609ba),
	.w7(32'h3a944f30),
	.w8(32'hbab36283),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07d929),
	.w1(32'h3aa64aa5),
	.w2(32'hb9ca4f4c),
	.w3(32'h3ae748e4),
	.w4(32'h3a8337cf),
	.w5(32'hbb165951),
	.w6(32'h3b7eb836),
	.w7(32'h3a506b15),
	.w8(32'hbb39781f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac475bc),
	.w1(32'h39d555d9),
	.w2(32'h399612b9),
	.w3(32'hba1d07bc),
	.w4(32'hba892f9d),
	.w5(32'hba1c9d55),
	.w6(32'hbb1501aa),
	.w7(32'hbafef1a2),
	.w8(32'h39a25c53),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a547965),
	.w1(32'h3a9c2f15),
	.w2(32'h3a18b1f1),
	.w3(32'hba19365e),
	.w4(32'hba5c4540),
	.w5(32'hba00465e),
	.w6(32'h38fa916f),
	.w7(32'h39d6ceb0),
	.w8(32'hba8b1189),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd562c),
	.w1(32'hbab8d2da),
	.w2(32'hbac44257),
	.w3(32'hba89c464),
	.w4(32'hbab5619c),
	.w5(32'hb9e083f8),
	.w6(32'hbadc2371),
	.w7(32'hbae9a7b4),
	.w8(32'h3ac39968),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921ad8b),
	.w1(32'hba3ea001),
	.w2(32'hbab27e7a),
	.w3(32'hbaaeaba3),
	.w4(32'hbaf59e1b),
	.w5(32'h3937fb51),
	.w6(32'hbaee3c1d),
	.w7(32'hba83fe9f),
	.w8(32'h3a19b0f1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb7fd5),
	.w1(32'h3a801bfe),
	.w2(32'hba247c5f),
	.w3(32'h3a613668),
	.w4(32'h38bfcb88),
	.w5(32'hbafcd3ec),
	.w6(32'hb91d0972),
	.w7(32'hb9dce62b),
	.w8(32'hbabc2513),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a866e9d),
	.w1(32'h3aa8eabb),
	.w2(32'h3b8723fc),
	.w3(32'hba9a8633),
	.w4(32'hba4adf1d),
	.w5(32'h3a4fb02c),
	.w6(32'hbad3a848),
	.w7(32'h3a4665aa),
	.w8(32'hbab6e04e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1b027),
	.w1(32'hba31b17b),
	.w2(32'h39b1a729),
	.w3(32'h3914ab2e),
	.w4(32'h3a2831ef),
	.w5(32'hb8d46e1c),
	.w6(32'hbadc964d),
	.w7(32'h38cec2cc),
	.w8(32'h38e91220),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78af27),
	.w1(32'hbacdc751),
	.w2(32'hbb8241d0),
	.w3(32'hb91585f6),
	.w4(32'hbac06d7b),
	.w5(32'hba4223ef),
	.w6(32'h3a4b103e),
	.w7(32'hb960e094),
	.w8(32'h3ac901e0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1959cb),
	.w1(32'hb9422627),
	.w2(32'h39ac9ca7),
	.w3(32'hb97b453d),
	.w4(32'hb97cc722),
	.w5(32'hbaa71305),
	.w6(32'hbafcb46e),
	.w7(32'hbaa22587),
	.w8(32'hb8c5746f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac28de5),
	.w1(32'hb95517f1),
	.w2(32'h3aa2801e),
	.w3(32'hb9be5ce5),
	.w4(32'h39974662),
	.w5(32'h39d8ca77),
	.w6(32'h3af63f42),
	.w7(32'h3b03c0ec),
	.w8(32'h3b23f0f1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc6d6f),
	.w1(32'h3aafc238),
	.w2(32'hb8779909),
	.w3(32'h3aba71e9),
	.w4(32'hba8694e3),
	.w5(32'h3a110890),
	.w6(32'h3b2cdf61),
	.w7(32'h39df3826),
	.w8(32'h3abd138b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21a5e3),
	.w1(32'hba8e1436),
	.w2(32'hbadb4d27),
	.w3(32'hba66d23a),
	.w4(32'h394ca4ae),
	.w5(32'h3b4cab62),
	.w6(32'hbaaa2d0f),
	.w7(32'h3984e175),
	.w8(32'h3a83f9f1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a606cc2),
	.w1(32'h3a4e5609),
	.w2(32'h3b32ca6e),
	.w3(32'h3af873f0),
	.w4(32'h3b1c6cad),
	.w5(32'hbb30f1a2),
	.w6(32'hba234a15),
	.w7(32'h3abd33bf),
	.w8(32'hbbe83ed7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf56f9),
	.w1(32'h3bf786f4),
	.w2(32'h3bbb30b3),
	.w3(32'h3c114227),
	.w4(32'h3b69dba3),
	.w5(32'hbb892fb5),
	.w6(32'h3c5458a1),
	.w7(32'h3bccd0b6),
	.w8(32'hbb360be9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ef021),
	.w1(32'h3b1d35ba),
	.w2(32'h3c1b0331),
	.w3(32'hb60e7c2f),
	.w4(32'h3b86c8c9),
	.w5(32'hbc8993dd),
	.w6(32'hbbcf5be7),
	.w7(32'h3ae01d4a),
	.w8(32'hbc5f29a3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88bc1a),
	.w1(32'hbbc5bc8d),
	.w2(32'hbbffe738),
	.w3(32'hbc1bb5aa),
	.w4(32'hbbb25196),
	.w5(32'h3b9fe431),
	.w6(32'hbb8fc436),
	.w7(32'h3b1d860b),
	.w8(32'h3c4ef28b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2ebc7),
	.w1(32'h3c45ca69),
	.w2(32'hba5ad0f2),
	.w3(32'h3ca953b0),
	.w4(32'h3b6deb98),
	.w5(32'hbaf86380),
	.w6(32'h3cb97069),
	.w7(32'hb9a2e905),
	.w8(32'hbb7c7855),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cae494),
	.w1(32'hbad258e5),
	.w2(32'h3b5245c0),
	.w3(32'hbb011315),
	.w4(32'hbaef6192),
	.w5(32'hbbb69bc2),
	.w6(32'h39947ddf),
	.w7(32'hb9dcae40),
	.w8(32'h3a9d3ba9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba237541),
	.w1(32'hbb42a306),
	.w2(32'hbb2a5ed0),
	.w3(32'hbbef1a96),
	.w4(32'h39b3ceff),
	.w5(32'hbb22f5a1),
	.w6(32'hbb334881),
	.w7(32'hbc0cefcf),
	.w8(32'hbb60dafc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb21627),
	.w1(32'hb9a85a39),
	.w2(32'h3b457765),
	.w3(32'hbb224874),
	.w4(32'h3ae06073),
	.w5(32'hbbd3c7c4),
	.w6(32'hbb72c6da),
	.w7(32'h3bd1a58d),
	.w8(32'hbbbb1732),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3ccd4),
	.w1(32'hbad6b1da),
	.w2(32'h3c0595b0),
	.w3(32'hbb75c55c),
	.w4(32'hbbca40a8),
	.w5(32'h3ad3ab89),
	.w6(32'h3b95b600),
	.w7(32'h3ba31baf),
	.w8(32'h3ba8dffa),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddc2e6),
	.w1(32'h3ccfe55f),
	.w2(32'hba2c0581),
	.w3(32'h3c9d80b3),
	.w4(32'hba7a5583),
	.w5(32'h3b17e155),
	.w6(32'h3c9e8da6),
	.w7(32'hbbc41343),
	.w8(32'h38b6a2f4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae22a12),
	.w1(32'h3ba689b6),
	.w2(32'hbb5811fe),
	.w3(32'h3be8c123),
	.w4(32'hbb256fc8),
	.w5(32'h3a92f596),
	.w6(32'h3bc38ad7),
	.w7(32'h3ac8a638),
	.w8(32'h3b588b9e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13d145),
	.w1(32'hbaeae84a),
	.w2(32'hbb7dff07),
	.w3(32'hbb1cf405),
	.w4(32'hbabad9ad),
	.w5(32'hbbcea9c9),
	.w6(32'hba1cef6e),
	.w7(32'hbb156d6d),
	.w8(32'h392d775b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaee2e),
	.w1(32'hb996d673),
	.w2(32'hb9d481c2),
	.w3(32'hbba69ae6),
	.w4(32'hbb519c0f),
	.w5(32'hbbdf0f75),
	.w6(32'hbb2ab14a),
	.w7(32'h38f4e845),
	.w8(32'hbc412a80),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc192315),
	.w1(32'hbc366bb4),
	.w2(32'hb86a4de2),
	.w3(32'hbc180674),
	.w4(32'h3b3c211d),
	.w5(32'hbb3c3cdb),
	.w6(32'hbae1d301),
	.w7(32'hbbbe1a6d),
	.w8(32'hbb54c6d5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f407c),
	.w1(32'hbba4d602),
	.w2(32'h3b32a02f),
	.w3(32'hbb898ff3),
	.w4(32'h3b58ff0b),
	.w5(32'hbc0223c2),
	.w6(32'hbb8ab432),
	.w7(32'h3bb551ad),
	.w8(32'hba3aa360),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944acc3),
	.w1(32'hbb37417b),
	.w2(32'hbb16056b),
	.w3(32'hbbce2e46),
	.w4(32'hbb8e62bc),
	.w5(32'h3b0edd7b),
	.w6(32'h3a62e08f),
	.w7(32'hba6dec37),
	.w8(32'h3b3093e8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb972f91),
	.w1(32'h3be6fae9),
	.w2(32'h3bf1c1f0),
	.w3(32'hbbd54726),
	.w4(32'h3ac6a2be),
	.w5(32'hbbbdfc78),
	.w6(32'h3b23f5bc),
	.w7(32'h3b1bd4d7),
	.w8(32'hbc1dd5eb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1657a7),
	.w1(32'hbc0a515e),
	.w2(32'h3b1f09eb),
	.w3(32'hbc38dff6),
	.w4(32'h3b2c6342),
	.w5(32'h3ac320f1),
	.w6(32'hbbce3276),
	.w7(32'h38ab01b4),
	.w8(32'h3b27d27d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20a803),
	.w1(32'hbabb1b50),
	.w2(32'h3b3213b1),
	.w3(32'hbb670524),
	.w4(32'h3b4f7f4e),
	.w5(32'hbb9c6337),
	.w6(32'hbb107d64),
	.w7(32'h3a85f251),
	.w8(32'hbbc72124),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1e826),
	.w1(32'hbbe87714),
	.w2(32'hbbb2661c),
	.w3(32'hbb6f6403),
	.w4(32'h3afb6bb8),
	.w5(32'hbacca640),
	.w6(32'hbbc05380),
	.w7(32'hbb566b95),
	.w8(32'hbb9ed649),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba904313),
	.w1(32'h3c2e7924),
	.w2(32'h3b409a05),
	.w3(32'h3c0283d6),
	.w4(32'h3afb0aed),
	.w5(32'hbaa57188),
	.w6(32'h3c89aeef),
	.w7(32'hba25170b),
	.w8(32'hbaea29c7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb495475),
	.w1(32'hb9de4321),
	.w2(32'hbb877652),
	.w3(32'h3a8a8a17),
	.w4(32'hbc2afd5b),
	.w5(32'hbc039eac),
	.w6(32'h3b631289),
	.w7(32'hbb801ad4),
	.w8(32'hbbebaf54),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfed013),
	.w1(32'hbc0e38bf),
	.w2(32'h3b06bad9),
	.w3(32'hbb4a8044),
	.w4(32'hba6d19ea),
	.w5(32'hbbb13d31),
	.w6(32'hbb00338b),
	.w7(32'hbbe85ece),
	.w8(32'hbba3d6c0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0131b9),
	.w1(32'hbbdfa5c6),
	.w2(32'hbb5516d5),
	.w3(32'hbbdd77cb),
	.w4(32'hbba1af27),
	.w5(32'hbb1d888a),
	.w6(32'hbb3c0900),
	.w7(32'hbbc04a97),
	.w8(32'hbc133e51),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1734b1),
	.w1(32'h3b8ec271),
	.w2(32'h39c0ad0c),
	.w3(32'hbaee6855),
	.w4(32'hbb20b5a0),
	.w5(32'hbc2f5714),
	.w6(32'hbb4068b6),
	.w7(32'h39d4e61d),
	.w8(32'hbbc156a6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd89e77),
	.w1(32'hbbcd6059),
	.w2(32'hba972d6b),
	.w3(32'hbae373f9),
	.w4(32'hba1ada5f),
	.w5(32'hbb0daf7d),
	.w6(32'hbb8f9981),
	.w7(32'h3b70dc67),
	.w8(32'hbba02bcd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea774e),
	.w1(32'hbaaffe19),
	.w2(32'h38514629),
	.w3(32'hbb5359e6),
	.w4(32'hbba87978),
	.w5(32'hbb89d7dc),
	.w6(32'hbb7ef92e),
	.w7(32'hbba658dd),
	.w8(32'hbb82d3cd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12ca72),
	.w1(32'h3b78dc9c),
	.w2(32'hbb82178e),
	.w3(32'hbb91b9c0),
	.w4(32'hbba4d4bb),
	.w5(32'hbb7f5cc1),
	.w6(32'h3bce6a20),
	.w7(32'hbb4e3746),
	.w8(32'hb9bc2b3c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e94eb),
	.w1(32'h3b1daa8d),
	.w2(32'hba545c34),
	.w3(32'hbb8a94cb),
	.w4(32'hbab385fb),
	.w5(32'h3ba97b34),
	.w6(32'hbb1a762e),
	.w7(32'hba44ef86),
	.w8(32'h3be01fea),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd458d4),
	.w1(32'hbb247c7c),
	.w2(32'hbb5d228f),
	.w3(32'hba8da422),
	.w4(32'hbb9c4c08),
	.w5(32'hbac81723),
	.w6(32'hbb51e3aa),
	.w7(32'hbba556a5),
	.w8(32'hbb0319e6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0cf1b),
	.w1(32'hbb1c15e4),
	.w2(32'h3a4d8d3f),
	.w3(32'hbbbdd71f),
	.w4(32'h3ac3a140),
	.w5(32'h3b449bcd),
	.w6(32'hbba20ebd),
	.w7(32'h3ab5862d),
	.w8(32'h3a59abc3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda37a4),
	.w1(32'h3b1bc40f),
	.w2(32'hba4894e6),
	.w3(32'h39cc99cf),
	.w4(32'h3aa27613),
	.w5(32'h3c1e9e3f),
	.w6(32'hbb2e9676),
	.w7(32'hbab6bd09),
	.w8(32'h3bc115f3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c099382),
	.w1(32'hbc417939),
	.w2(32'h3bd8e7b6),
	.w3(32'hbc380a95),
	.w4(32'hbc137d15),
	.w5(32'hbaf48e60),
	.w6(32'hbc4406e9),
	.w7(32'hbc259734),
	.w8(32'hbb9ad579),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8b600),
	.w1(32'h3af06f52),
	.w2(32'h3a26a66c),
	.w3(32'hbb247398),
	.w4(32'hb9e3fc97),
	.w5(32'hbc519631),
	.w6(32'hb9bc68a9),
	.w7(32'h3a2e3223),
	.w8(32'hbc1bca5a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3a1c8),
	.w1(32'hbc48a8b4),
	.w2(32'hbbcf78d9),
	.w3(32'hbbda6c3d),
	.w4(32'hb96c59f9),
	.w5(32'hb9f0553e),
	.w6(32'hbac175d0),
	.w7(32'h3a7d2858),
	.w8(32'h3ac25c7b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924f347),
	.w1(32'h3b45279e),
	.w2(32'hbab09526),
	.w3(32'h38e2a33e),
	.w4(32'hb9454aec),
	.w5(32'hbb639dbf),
	.w6(32'h3aadf72a),
	.w7(32'hbab28894),
	.w8(32'hbb4ff439),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9683f3),
	.w1(32'hb98c9637),
	.w2(32'hbac4820e),
	.w3(32'hbb7176d0),
	.w4(32'h3a1b2dc9),
	.w5(32'hbb525158),
	.w6(32'hbb44f500),
	.w7(32'hbb4af3ba),
	.w8(32'hbb81fb66),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a72cf),
	.w1(32'hbbde16ee),
	.w2(32'h3b448de1),
	.w3(32'hbbe11a8a),
	.w4(32'h3b4e35a0),
	.w5(32'h39639654),
	.w6(32'hbbf36feb),
	.w7(32'h3bc469e5),
	.w8(32'h3a20ab5b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa323),
	.w1(32'hbb56ee28),
	.w2(32'h3b8245d6),
	.w3(32'hbb49795d),
	.w4(32'h3ba59bb6),
	.w5(32'hbb060499),
	.w6(32'hbb96c744),
	.w7(32'h3b7cecff),
	.w8(32'h39d7470e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a083ea0),
	.w1(32'h3b80f5f1),
	.w2(32'h38f80ca0),
	.w3(32'h3a62fdc4),
	.w4(32'h3b03a4eb),
	.w5(32'hbb8cafd5),
	.w6(32'h3ae4cd90),
	.w7(32'hb9871f2d),
	.w8(32'hbae731df),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53b695),
	.w1(32'h3c0555ad),
	.w2(32'h3b217e08),
	.w3(32'h3be75f38),
	.w4(32'h3a43ca56),
	.w5(32'hbc2c9c86),
	.w6(32'h3c42b78e),
	.w7(32'h3ae999c2),
	.w8(32'hbc2fa907),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3acd1),
	.w1(32'hbadf9ea1),
	.w2(32'hba254cb2),
	.w3(32'hbb4236e5),
	.w4(32'hbc3a8e87),
	.w5(32'hbae6b81e),
	.w6(32'hba84b5fc),
	.w7(32'hba85a658),
	.w8(32'hbb8eee4a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a758f),
	.w1(32'hba39385e),
	.w2(32'h3c1bf93b),
	.w3(32'h3a0d4898),
	.w4(32'h3a4523e6),
	.w5(32'h3bbe8011),
	.w6(32'hba4b6a93),
	.w7(32'h3c1af686),
	.w8(32'h3c4e994a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb783c0),
	.w1(32'h3cb0b7a8),
	.w2(32'h3c3105d2),
	.w3(32'h3cad4618),
	.w4(32'h3bc393d2),
	.w5(32'hbb891212),
	.w6(32'h3c9afebe),
	.w7(32'h3c0ed01e),
	.w8(32'h3a475e97),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941a027),
	.w1(32'hbb4a2a99),
	.w2(32'hbb106659),
	.w3(32'hbba9406d),
	.w4(32'hbba507d2),
	.w5(32'hbb8ef9f5),
	.w6(32'hbb8a7b9e),
	.w7(32'hbaa9bbec),
	.w8(32'hbbfbdf37),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc02979),
	.w1(32'h3c0035f8),
	.w2(32'h3b571889),
	.w3(32'h3bc3948a),
	.w4(32'h3af3d726),
	.w5(32'h389d6c42),
	.w6(32'h3be1ee80),
	.w7(32'h3c0f872a),
	.w8(32'hba7d94e5),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380dd268),
	.w1(32'h3b257e63),
	.w2(32'h3b7a6849),
	.w3(32'hbb6bac68),
	.w4(32'h3b51d3e2),
	.w5(32'h3826bec7),
	.w6(32'hbba3e900),
	.w7(32'h3b1af4a5),
	.w8(32'h3a33f0a0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a5ab5),
	.w1(32'hb9a987d6),
	.w2(32'h3b79a21b),
	.w3(32'hba119edf),
	.w4(32'h3ada71dc),
	.w5(32'hbbdaa3dd),
	.w6(32'h3b6c7403),
	.w7(32'h3a49dc8f),
	.w8(32'hbb73aa3e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84830d),
	.w1(32'hba4a0f79),
	.w2(32'hbbb84e05),
	.w3(32'h3a9d063c),
	.w4(32'h3b352235),
	.w5(32'hbbc66451),
	.w6(32'hbb826612),
	.w7(32'h3b1bd38b),
	.w8(32'hbbda088e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad853bd),
	.w1(32'hbc426092),
	.w2(32'h3945da40),
	.w3(32'hbc2cb5da),
	.w4(32'h3c01ce1e),
	.w5(32'h3af4bd15),
	.w6(32'hbba9ca6a),
	.w7(32'hbb667755),
	.w8(32'hb97240de),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf0bb7),
	.w1(32'h3c45313e),
	.w2(32'hbb591ef3),
	.w3(32'h3bb129bb),
	.w4(32'h3b0ef363),
	.w5(32'hba23a6cb),
	.w6(32'h3c2d772b),
	.w7(32'h3b68b4e6),
	.w8(32'hbb82bd76),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad05188),
	.w1(32'hbac37398),
	.w2(32'hba83af83),
	.w3(32'hbb4c5279),
	.w4(32'h3a1e4945),
	.w5(32'hbc0b6c56),
	.w6(32'hbb89e048),
	.w7(32'hba165895),
	.w8(32'hbb9fa09a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d7f77),
	.w1(32'hbb0fe52b),
	.w2(32'hbb931dd4),
	.w3(32'h3bb40779),
	.w4(32'hbbc6fc4a),
	.w5(32'h3c20ac2f),
	.w6(32'h3b8ae527),
	.w7(32'hbb58d473),
	.w8(32'h3c6a5fd4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f3915),
	.w1(32'h3b9201b5),
	.w2(32'h3baea996),
	.w3(32'h3ab384ec),
	.w4(32'h3b87049a),
	.w5(32'hbb750442),
	.w6(32'h39ae1b3e),
	.w7(32'h3be76024),
	.w8(32'h3c6d8064),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902231f),
	.w1(32'hbb6aecb8),
	.w2(32'hbba80ede),
	.w3(32'hbbc44d12),
	.w4(32'h3b619974),
	.w5(32'hbb764ce7),
	.w6(32'hbb4902b0),
	.w7(32'h3b391336),
	.w8(32'h39d448c5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3755921a),
	.w1(32'h39612271),
	.w2(32'h3b95b1d8),
	.w3(32'hbb8ec1df),
	.w4(32'h3ae1a9fc),
	.w5(32'hbba1aeae),
	.w6(32'hbb457deb),
	.w7(32'h3ba62d47),
	.w8(32'hbb20b82c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf4b76),
	.w1(32'h3b9f83f6),
	.w2(32'hbbbe8c4a),
	.w3(32'h3b31be84),
	.w4(32'hbc0f973a),
	.w5(32'h3b5d6b88),
	.w6(32'h3b83185b),
	.w7(32'hbbdbe984),
	.w8(32'h3b5e1557),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5da733),
	.w1(32'hbb441cb4),
	.w2(32'hba4918c3),
	.w3(32'hbb078848),
	.w4(32'h3b48db72),
	.w5(32'h3af19a86),
	.w6(32'hbab96595),
	.w7(32'h3a8f756b),
	.w8(32'h3c0d6e82),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2427f4),
	.w1(32'h3c331013),
	.w2(32'h3bbfbece),
	.w3(32'hbb3f9d68),
	.w4(32'hbb22c514),
	.w5(32'hbc18f2fc),
	.w6(32'h3bc6e21d),
	.w7(32'h3c1f496b),
	.w8(32'hbc0f4c12),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd74921),
	.w1(32'hbc60f3e4),
	.w2(32'h3b883035),
	.w3(32'hbc47405c),
	.w4(32'h3ab15757),
	.w5(32'hbba707d5),
	.w6(32'hbbf8d97a),
	.w7(32'h3afbf79a),
	.w8(32'h3c5b59c7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b394e16),
	.w1(32'hbbbb1127),
	.w2(32'hba2cbdd9),
	.w3(32'h3be2b1d3),
	.w4(32'h3c32f9ef),
	.w5(32'h3b8742ee),
	.w6(32'h3bc824fe),
	.w7(32'h3b5e1da6),
	.w8(32'h3c41f68a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a2b41),
	.w1(32'h3ca26ecd),
	.w2(32'h3c47aa3d),
	.w3(32'hbb6d4a96),
	.w4(32'hbb502c1f),
	.w5(32'hbb0e7ca6),
	.w6(32'h3be1de52),
	.w7(32'hbb9cffaa),
	.w8(32'hbb67fd3d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc560bd4),
	.w1(32'hbc3589c1),
	.w2(32'hbc202c65),
	.w3(32'hbbc51793),
	.w4(32'hbb9d09ef),
	.w5(32'hb9753731),
	.w6(32'hbc3204fc),
	.w7(32'hbb8755e1),
	.w8(32'hbb4aa8b9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23b902),
	.w1(32'hbaac6523),
	.w2(32'h3b4c8ab4),
	.w3(32'h3ae03186),
	.w4(32'h3b50bf85),
	.w5(32'h3998644b),
	.w6(32'h3bed591a),
	.w7(32'h3b71bdac),
	.w8(32'h3c85a53c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5242bd),
	.w1(32'h3c11d76c),
	.w2(32'h3b1b1ab2),
	.w3(32'h3b0e3b63),
	.w4(32'hbb1f146d),
	.w5(32'h3a97fde0),
	.w6(32'h3c662fd1),
	.w7(32'hba4eb85b),
	.w8(32'hba1f00b5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f7f4a),
	.w1(32'h3a138054),
	.w2(32'hbbaf44fd),
	.w3(32'hb93698da),
	.w4(32'h3b901d2c),
	.w5(32'hbc49a493),
	.w6(32'h3b93ece0),
	.w7(32'h3b547697),
	.w8(32'hbb471e0b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ceff2),
	.w1(32'hbc33d955),
	.w2(32'hbc1f209e),
	.w3(32'hb80ee204),
	.w4(32'hba856ae4),
	.w5(32'hbc02ad62),
	.w6(32'h3a9de5f7),
	.w7(32'h3af3a611),
	.w8(32'hbc0c2ac3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc6a3),
	.w1(32'h3ad8a888),
	.w2(32'h3b0655d1),
	.w3(32'h3a10e7ed),
	.w4(32'hba895cf6),
	.w5(32'hbbf6ef3a),
	.w6(32'hba183999),
	.w7(32'hba93beda),
	.w8(32'hbbbcc001),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1b670),
	.w1(32'hbb216161),
	.w2(32'hbbbdd6b1),
	.w3(32'h3b06609e),
	.w4(32'h3b3a2b10),
	.w5(32'h3b622d4b),
	.w6(32'h3a99d1e6),
	.w7(32'h395f1047),
	.w8(32'hbba8c080),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca5330),
	.w1(32'hbbbcadc2),
	.w2(32'h3b085e23),
	.w3(32'hbbe1c57c),
	.w4(32'hb85d1081),
	.w5(32'hbba18ab9),
	.w6(32'hbb908585),
	.w7(32'hb83d13a2),
	.w8(32'hbb04c365),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8542a7),
	.w1(32'h3ab86432),
	.w2(32'hb9e0ed5d),
	.w3(32'h3b858bce),
	.w4(32'hbb5695dd),
	.w5(32'hbc0a358d),
	.w6(32'hbc155f5b),
	.w7(32'hba5d51d3),
	.w8(32'hbc05be35),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da699),
	.w1(32'h3aece69a),
	.w2(32'h3aebc2d7),
	.w3(32'hbb461293),
	.w4(32'hb95ce54a),
	.w5(32'hbba55372),
	.w6(32'hbb4c4db0),
	.w7(32'h3aa93d57),
	.w8(32'hbb65fed8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae998),
	.w1(32'hbb19ca91),
	.w2(32'hbb8d82ed),
	.w3(32'hbbd6db85),
	.w4(32'hbb74074d),
	.w5(32'hbbbf28b8),
	.w6(32'hbac86e68),
	.w7(32'h3bb074d0),
	.w8(32'hba738b0e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d3ea8),
	.w1(32'h3bec7979),
	.w2(32'hbc0b61a7),
	.w3(32'h3b1bc3cc),
	.w4(32'hbbb04dec),
	.w5(32'h3c0b3ffe),
	.w6(32'h3bd67168),
	.w7(32'hbc0f3a48),
	.w8(32'h3bf201be),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6bf02),
	.w1(32'h3bb2aadc),
	.w2(32'h3b7cbd77),
	.w3(32'h399126d8),
	.w4(32'h3ac233ba),
	.w5(32'h3adb7c13),
	.w6(32'h3a1e2711),
	.w7(32'h3b24a334),
	.w8(32'h3b7c575d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b5269),
	.w1(32'hbb37b99e),
	.w2(32'hbaf77e2b),
	.w3(32'hbbe6bd6e),
	.w4(32'hb97292ac),
	.w5(32'h38538ecc),
	.w6(32'hbc2aeb9e),
	.w7(32'hbb4a98ae),
	.w8(32'hba0835e8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba587b02),
	.w1(32'h3b882a1b),
	.w2(32'h3992bea6),
	.w3(32'h3bac6f31),
	.w4(32'hbb68c35c),
	.w5(32'hbbe8b7fb),
	.w6(32'h3b68eebe),
	.w7(32'hbb69b50c),
	.w8(32'hbbea5851),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb264d92),
	.w1(32'hbb0fd88e),
	.w2(32'h3b2f7103),
	.w3(32'hbb217203),
	.w4(32'h3b5a8ccb),
	.w5(32'hba94ea18),
	.w6(32'hbb8468e2),
	.w7(32'h3ba52aeb),
	.w8(32'h3acf9740),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba642456),
	.w1(32'hb9a73a21),
	.w2(32'h3b751a9d),
	.w3(32'hba2292da),
	.w4(32'h3b648e13),
	.w5(32'hbb9d2f50),
	.w6(32'hb94f8c75),
	.w7(32'h3c01ed3e),
	.w8(32'hbbcfc75c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea735a),
	.w1(32'hbaeb96f2),
	.w2(32'hbaa8b752),
	.w3(32'hbb9b0814),
	.w4(32'hbb24bd0b),
	.w5(32'hbc06cefe),
	.w6(32'hbb7627fd),
	.w7(32'hbb1cb85f),
	.w8(32'hbc30a1af),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51dc04),
	.w1(32'h3b9e0c7e),
	.w2(32'h3a7fecdf),
	.w3(32'h3c3117b1),
	.w4(32'h3b9c9638),
	.w5(32'hba6efec8),
	.w6(32'h3cc946f8),
	.w7(32'h3bc711d4),
	.w8(32'hbb869dd7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb783762),
	.w1(32'h3b6d75ea),
	.w2(32'h3b42eee2),
	.w3(32'hba83702c),
	.w4(32'hbb5b90fe),
	.w5(32'hbbd0affe),
	.w6(32'hbb940649),
	.w7(32'hbba9c1f6),
	.w8(32'h3b16f27d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b2df9),
	.w1(32'h3b30f5ab),
	.w2(32'h3c0985e5),
	.w3(32'h3c643dac),
	.w4(32'h3bb9b35b),
	.w5(32'hbc43f046),
	.w6(32'h3c723390),
	.w7(32'h3c605bc8),
	.w8(32'hbc1c891c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cea91),
	.w1(32'hbbacb528),
	.w2(32'hb9b5d916),
	.w3(32'hb7a30049),
	.w4(32'hbb940a2e),
	.w5(32'hbb90872e),
	.w6(32'hbb5fe39e),
	.w7(32'h39b98086),
	.w8(32'hbbd75548),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5203ba),
	.w1(32'hbc726b52),
	.w2(32'hbab4a85b),
	.w3(32'hbc47efd7),
	.w4(32'hb9d52199),
	.w5(32'h3c0aca67),
	.w6(32'hbc13cac2),
	.w7(32'hbbba9424),
	.w8(32'h3cfc8cf5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c006fcd),
	.w1(32'h3d431a38),
	.w2(32'h3c8701d6),
	.w3(32'h3c8f1ca8),
	.w4(32'h3bf30289),
	.w5(32'h3c4d85b6),
	.w6(32'h3d1599bb),
	.w7(32'h3c128a38),
	.w8(32'h3c590ef8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ae5a4),
	.w1(32'h3c8d7216),
	.w2(32'h3bd9c284),
	.w3(32'h3c2d2379),
	.w4(32'h3a16a9c4),
	.w5(32'h3a67e17d),
	.w6(32'h398f62f2),
	.w7(32'hbb991714),
	.w8(32'hbb3af05a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6b96b),
	.w1(32'h3bccbc53),
	.w2(32'h3ba1d233),
	.w3(32'h3c5531b0),
	.w4(32'h3c1f8ebd),
	.w5(32'hbbb92991),
	.w6(32'h3cae4f6b),
	.w7(32'h3b8138f2),
	.w8(32'hbbaf53a5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19f722),
	.w1(32'hb9bb8291),
	.w2(32'h3b51ad5c),
	.w3(32'hbb8bf23c),
	.w4(32'h3a6e4ac5),
	.w5(32'h381df828),
	.w6(32'hbb55eb22),
	.w7(32'h39c614f2),
	.w8(32'hbc06c543),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0fc36),
	.w1(32'h3b4bb5eb),
	.w2(32'h3b9a0ca4),
	.w3(32'h3b2c62cd),
	.w4(32'h3b98824a),
	.w5(32'hbb4613ec),
	.w6(32'hbb15a356),
	.w7(32'h3c0a93b2),
	.w8(32'h3b294aa5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f71bd),
	.w1(32'hbbc30728),
	.w2(32'hbb192eb9),
	.w3(32'hbb552683),
	.w4(32'hba791219),
	.w5(32'hbb327528),
	.w6(32'hbb21479c),
	.w7(32'hbad45f4c),
	.w8(32'hbaebd952),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c4a1),
	.w1(32'hbb3ff2b9),
	.w2(32'h3a912d62),
	.w3(32'hbb46595b),
	.w4(32'h3a288e17),
	.w5(32'hbc27eb4b),
	.w6(32'hbc06b5df),
	.w7(32'h3b300cf0),
	.w8(32'hba427663),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b9617),
	.w1(32'hbb59134c),
	.w2(32'hbb8047ba),
	.w3(32'hbbc33d25),
	.w4(32'hbba19251),
	.w5(32'hbb7a0eb9),
	.w6(32'hbba8901c),
	.w7(32'hbbddc11e),
	.w8(32'h3b8beab8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25e35),
	.w1(32'h3c553991),
	.w2(32'h3c06dfbc),
	.w3(32'h3c6d5fdc),
	.w4(32'h3b98563e),
	.w5(32'hbaac6fda),
	.w6(32'h39edec47),
	.w7(32'h3c2b3522),
	.w8(32'h394d93a6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0039b4),
	.w1(32'h3bbc400d),
	.w2(32'h3ba1b94a),
	.w3(32'hbbd0750c),
	.w4(32'h3b358324),
	.w5(32'hbbafadfa),
	.w6(32'h3c291313),
	.w7(32'h3a422916),
	.w8(32'hbb6025bd),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fbfb2),
	.w1(32'hbb9bd062),
	.w2(32'hbab0bb14),
	.w3(32'h3a57abe8),
	.w4(32'hbbe8b69a),
	.w5(32'hbb622e61),
	.w6(32'h3b0fc8fd),
	.w7(32'h39bd9af9),
	.w8(32'hbbb1ffd6),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7937a),
	.w1(32'hbc0ae44f),
	.w2(32'hbac61030),
	.w3(32'hbbc462f2),
	.w4(32'hbbd51aeb),
	.w5(32'hba283bd1),
	.w6(32'hbc109799),
	.w7(32'hbadeeb4b),
	.w8(32'hbb7b1748),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc74539),
	.w1(32'h3af8016c),
	.w2(32'h3b09ab8a),
	.w3(32'h3b1ab21f),
	.w4(32'h3b3402af),
	.w5(32'hbb4f2060),
	.w6(32'h3b84c8eb),
	.w7(32'h3c1187c4),
	.w8(32'hbc2783da),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad01a),
	.w1(32'hbca106e1),
	.w2(32'h39987df2),
	.w3(32'hbc87fc21),
	.w4(32'h3ab4a492),
	.w5(32'h3b700440),
	.w6(32'hbaf8577f),
	.w7(32'hbaff851e),
	.w8(32'h38921979),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d6ed),
	.w1(32'hbc08f462),
	.w2(32'hbba7ee8b),
	.w3(32'hbba155bb),
	.w4(32'hb8a8d3f4),
	.w5(32'hbbf16342),
	.w6(32'hbca5e7e4),
	.w7(32'hbb86cb88),
	.w8(32'hbaa8c303),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7621ef),
	.w1(32'hbb7b161a),
	.w2(32'hbb11629f),
	.w3(32'hbb303cfa),
	.w4(32'hbb5179bf),
	.w5(32'hbae58d8b),
	.w6(32'hbba567c8),
	.w7(32'h3a152711),
	.w8(32'hbb98b70d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb067acf),
	.w1(32'h3b24a032),
	.w2(32'hb9f516a9),
	.w3(32'h3b8d8a35),
	.w4(32'h3babc030),
	.w5(32'hbae70075),
	.w6(32'h3b9e5128),
	.w7(32'h3a83850a),
	.w8(32'hbb4d8a07),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2667b2),
	.w1(32'h3b6d8dde),
	.w2(32'hb95b70c0),
	.w3(32'hba79ea04),
	.w4(32'hbad7f1a4),
	.w5(32'h39084610),
	.w6(32'h3ad35e3b),
	.w7(32'h3b8268b8),
	.w8(32'hbb004d9d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcadb94),
	.w1(32'hbbea51d8),
	.w2(32'h39587ce5),
	.w3(32'hbb8db2a2),
	.w4(32'h3b6d7b63),
	.w5(32'hbadc7c19),
	.w6(32'hbbaef5ba),
	.w7(32'h3b96020e),
	.w8(32'hbb138d73),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba373984),
	.w1(32'hb907455f),
	.w2(32'hbb0702d5),
	.w3(32'h3a46f13a),
	.w4(32'hbb6e10cf),
	.w5(32'hbb95fdd9),
	.w6(32'hbae7373e),
	.w7(32'h3aa16bdb),
	.w8(32'hbb914810),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6265c),
	.w1(32'h3b94109b),
	.w2(32'h3bd447d1),
	.w3(32'h3b0572c2),
	.w4(32'h3b5ed880),
	.w5(32'hbb1e5454),
	.w6(32'h3bbc0c6f),
	.w7(32'h3bfff38f),
	.w8(32'h3c6e2ac0),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6befb1),
	.w1(32'h3c47902c),
	.w2(32'h3adb7a24),
	.w3(32'h3c5f55db),
	.w4(32'hb700904c),
	.w5(32'h3a758f23),
	.w6(32'h3ca43859),
	.w7(32'h3bdca0b8),
	.w8(32'hba95546e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a4001),
	.w1(32'h3c0f6070),
	.w2(32'h3bc164d2),
	.w3(32'h3b7ad1a3),
	.w4(32'h3b15ab8f),
	.w5(32'hbc202d91),
	.w6(32'h3c0c8c7c),
	.w7(32'h3b310c5f),
	.w8(32'hbc263724),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae312c3),
	.w1(32'hbba7f211),
	.w2(32'hba9199ca),
	.w3(32'hbbf16c56),
	.w4(32'hbbb28385),
	.w5(32'h3aae4e98),
	.w6(32'hbc539a5e),
	.w7(32'hbb3ab3a4),
	.w8(32'h3acd50ca),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba739023),
	.w1(32'hbb86fe62),
	.w2(32'hbb4a1b32),
	.w3(32'hbb42e20f),
	.w4(32'h3a8cd6cf),
	.w5(32'h3ad8b464),
	.w6(32'hbb9d4f2b),
	.w7(32'h3b22dca8),
	.w8(32'h3b6dde55),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be20983),
	.w1(32'h3a8280bd),
	.w2(32'h3abbc587),
	.w3(32'h3aba0bab),
	.w4(32'h3b363a35),
	.w5(32'hbbd9ee87),
	.w6(32'hba9471b5),
	.w7(32'h3baff572),
	.w8(32'hbbf1251e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96910f),
	.w1(32'hbb19acc1),
	.w2(32'h3a152526),
	.w3(32'hbb530666),
	.w4(32'h3bd5945d),
	.w5(32'hbbe0a468),
	.w6(32'hbae94466),
	.w7(32'h3be4d05e),
	.w8(32'hbbe3fc0c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95c876),
	.w1(32'hbb175f86),
	.w2(32'h3a9747cc),
	.w3(32'h3bc8b540),
	.w4(32'h396d8485),
	.w5(32'h3b1ca029),
	.w6(32'h3c7a7ddf),
	.w7(32'h3a47ba31),
	.w8(32'h3aa444f8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6d3f9),
	.w1(32'h3af87f6e),
	.w2(32'hbb9e813f),
	.w3(32'h3a7e8d26),
	.w4(32'h350ff542),
	.w5(32'hbb592c5e),
	.w6(32'hb9fe7c58),
	.w7(32'hbb554c95),
	.w8(32'hbb8d6d85),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395971ac),
	.w1(32'hbb84b474),
	.w2(32'hbba50e4c),
	.w3(32'h3a04db83),
	.w4(32'hbb9511ba),
	.w5(32'hbb8fdd41),
	.w6(32'h3b5a66f0),
	.w7(32'hbb9397ea),
	.w8(32'h3af7c804),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6538bc),
	.w1(32'h3b9f7ff4),
	.w2(32'h3b2f922f),
	.w3(32'h3b5ba89f),
	.w4(32'h3ad0447e),
	.w5(32'h3b899ffe),
	.w6(32'h3be3a32c),
	.w7(32'h3b89cfc7),
	.w8(32'h3a97ca11),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada5c2d),
	.w1(32'hbbfeb521),
	.w2(32'h3bfd8278),
	.w3(32'hbb8aa53b),
	.w4(32'h37a98473),
	.w5(32'hbb44213d),
	.w6(32'h3b0e3090),
	.w7(32'hbad0c379),
	.w8(32'hbacc6141),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93ec49),
	.w1(32'hbbb4ba6c),
	.w2(32'hba880af4),
	.w3(32'hbb4b1d96),
	.w4(32'h397d4219),
	.w5(32'hba66d782),
	.w6(32'h3a8d226e),
	.w7(32'h3b2c6a15),
	.w8(32'hba80d986),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe74e7),
	.w1(32'hbabc267e),
	.w2(32'h3a78a5a1),
	.w3(32'hbb33a502),
	.w4(32'h39138068),
	.w5(32'hba8e9b46),
	.w6(32'hbb3a851b),
	.w7(32'h389a0284),
	.w8(32'h3a195adf),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18fd6b),
	.w1(32'hba8da003),
	.w2(32'h3b091312),
	.w3(32'hba9d81ab),
	.w4(32'hbb26c060),
	.w5(32'h3bce478d),
	.w6(32'hbc04c3ac),
	.w7(32'h3a3ecdc9),
	.w8(32'h3bea5ae8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a28ea),
	.w1(32'h39160ed4),
	.w2(32'hbb7b5ed1),
	.w3(32'h39ed984f),
	.w4(32'h3b698b74),
	.w5(32'hba98f185),
	.w6(32'h3a8d1bab),
	.w7(32'hbaf2001d),
	.w8(32'h3b03289d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fdf25),
	.w1(32'hbb9d16e8),
	.w2(32'h3ae9ecb8),
	.w3(32'hbc0bc490),
	.w4(32'h396281c1),
	.w5(32'h3b976a60),
	.w6(32'hba99f574),
	.w7(32'h3afdbbad),
	.w8(32'h3c99739f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce797a),
	.w1(32'h3c20ecef),
	.w2(32'h3c2ce140),
	.w3(32'hbbe523df),
	.w4(32'h374ce415),
	.w5(32'h3c1b3027),
	.w6(32'h3a6f0cbd),
	.w7(32'hba8dcd48),
	.w8(32'h3c087d46),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aaddf),
	.w1(32'h3c59c592),
	.w2(32'hbba66cfa),
	.w3(32'h3c34815b),
	.w4(32'hbb3ab22c),
	.w5(32'hbb841251),
	.w6(32'h3c8a21ab),
	.w7(32'hbc0e18c8),
	.w8(32'hbb9e2793),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d75c0),
	.w1(32'hbbc1938f),
	.w2(32'hbb379a41),
	.w3(32'hbbd01581),
	.w4(32'hbb82b4a3),
	.w5(32'hbc0c8cb2),
	.w6(32'hbbf66263),
	.w7(32'hbb1d57ca),
	.w8(32'hbc038472),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9a6b6),
	.w1(32'h3bc8a3de),
	.w2(32'h3b3f2a53),
	.w3(32'hbbb4fe6b),
	.w4(32'hbc0b2ec0),
	.w5(32'hbb9c6ef1),
	.w6(32'hbba9e3ac),
	.w7(32'hbb18f9b8),
	.w8(32'hbc4a1f96),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e8635),
	.w1(32'hbb3ae1ce),
	.w2(32'hbab52105),
	.w3(32'hba9df5e5),
	.w4(32'hbb33bce2),
	.w5(32'h3cdc1938),
	.w6(32'hbc201926),
	.w7(32'hbb0dbf3a),
	.w8(32'h3d59d2f3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf099ed),
	.w1(32'h3c612de9),
	.w2(32'hbbcae9d9),
	.w3(32'h3cfa990f),
	.w4(32'hbb0aff72),
	.w5(32'h3b90f170),
	.w6(32'h3c2f7e46),
	.w7(32'hbbcdfb26),
	.w8(32'h3badfe26),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2077f),
	.w1(32'h3c026f33),
	.w2(32'h3bc765a9),
	.w3(32'h3be4b157),
	.w4(32'h3b4ac84f),
	.w5(32'hbb583ec8),
	.w6(32'h3c0c9630),
	.w7(32'h3b9b1e70),
	.w8(32'hbbd149fc),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841d93),
	.w1(32'hbbc546a1),
	.w2(32'hbbe905cc),
	.w3(32'hbb3707ea),
	.w4(32'hbb259f56),
	.w5(32'hbc251208),
	.w6(32'hbb180393),
	.w7(32'h3a780736),
	.w8(32'hbc0fc6a0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdca3f1),
	.w1(32'hbb800b42),
	.w2(32'hbb288cbe),
	.w3(32'hbbab8c98),
	.w4(32'hbb21bc42),
	.w5(32'hbb27b04c),
	.w6(32'hbaf0478d),
	.w7(32'hb90e69ab),
	.w8(32'hbbac8408),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2506f5),
	.w1(32'hbc00cd3d),
	.w2(32'hbb9b8399),
	.w3(32'h3aba0d59),
	.w4(32'hbad0de37),
	.w5(32'h3a1eb5fd),
	.w6(32'hbb266e3e),
	.w7(32'hb9f29e3f),
	.w8(32'hba85ea3e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3542a8),
	.w1(32'hbb0c502c),
	.w2(32'h3a38f516),
	.w3(32'hbb472f5c),
	.w4(32'hb973c7b8),
	.w5(32'hbc1a6d1f),
	.w6(32'hbb0abafa),
	.w7(32'hba4c27c9),
	.w8(32'hbbc2b7d1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3493),
	.w1(32'hbc2df1e2),
	.w2(32'hbc1f1630),
	.w3(32'hbc0912c5),
	.w4(32'hbc17aa56),
	.w5(32'hbbc57f90),
	.w6(32'hbbfe7e12),
	.w7(32'hbc09e5d2),
	.w8(32'hbb9ffe01),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0055cb),
	.w1(32'hbb6727a6),
	.w2(32'hbb5644b7),
	.w3(32'h3b304ce5),
	.w4(32'h3b590e30),
	.w5(32'hbab79431),
	.w6(32'h3b7d9d44),
	.w7(32'h3b123a81),
	.w8(32'hbb60c1b1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3717fd),
	.w1(32'h3706264b),
	.w2(32'h3a0973fb),
	.w3(32'hb9f018de),
	.w4(32'hbb234428),
	.w5(32'hbb27862a),
	.w6(32'hbb4cd2fe),
	.w7(32'hbac8bef2),
	.w8(32'hbb6bc340),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb79520),
	.w1(32'hbb386669),
	.w2(32'hbb0392a6),
	.w3(32'hba00a843),
	.w4(32'h392d12df),
	.w5(32'h3b73c9a9),
	.w6(32'hb96c5706),
	.w7(32'hb83d0c91),
	.w8(32'h3b6faca4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3fe4b),
	.w1(32'h3b9f0469),
	.w2(32'h3bbc31a2),
	.w3(32'h3b93c3c1),
	.w4(32'h3b9ec725),
	.w5(32'h39b37694),
	.w6(32'h3c27bb40),
	.w7(32'h3c30ef72),
	.w8(32'h3a82dd9e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f7e66),
	.w1(32'h3b356384),
	.w2(32'h3b1a633b),
	.w3(32'h3aba4eb8),
	.w4(32'h38bfc10f),
	.w5(32'h3c1fecff),
	.w6(32'h3b9629e1),
	.w7(32'h3acd0ec8),
	.w8(32'h3bf2bec0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09587d),
	.w1(32'h3c712eef),
	.w2(32'h3bc9c2b8),
	.w3(32'h3c6e6776),
	.w4(32'h3c02de83),
	.w5(32'hbbe4cbfa),
	.w6(32'h3c4cd86f),
	.w7(32'h3bdf4733),
	.w8(32'hbc0f28dd),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d3ab8),
	.w1(32'hb7f26c14),
	.w2(32'hbb2d61bf),
	.w3(32'hbb606d7a),
	.w4(32'h3aa185c4),
	.w5(32'h3af29045),
	.w6(32'h3b347974),
	.w7(32'h3b6509f9),
	.w8(32'h3acc7230),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50a049),
	.w1(32'hba48fc68),
	.w2(32'hb9f410ac),
	.w3(32'h3b044b22),
	.w4(32'hbb19636f),
	.w5(32'h3981406d),
	.w6(32'h3ab3faf9),
	.w7(32'hbb51b967),
	.w8(32'hb98b0c00),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a2095),
	.w1(32'hb8dde1e8),
	.w2(32'h3ae5d534),
	.w3(32'hba638e2d),
	.w4(32'h3ad60b08),
	.w5(32'hba2fe084),
	.w6(32'hbbc14ed2),
	.w7(32'hbb271c44),
	.w8(32'h399dd1a2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2acd78),
	.w1(32'h3b888336),
	.w2(32'hbad1880a),
	.w3(32'h3b77d176),
	.w4(32'h3aacf60f),
	.w5(32'h3ad352f8),
	.w6(32'h3a57fb87),
	.w7(32'h3b3ee939),
	.w8(32'h3a5a76b0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a985d37),
	.w1(32'h3b6b4639),
	.w2(32'h3b88283f),
	.w3(32'hbaedd713),
	.w4(32'hbb304110),
	.w5(32'hbbb6e81f),
	.w6(32'h3b2e22da),
	.w7(32'h3a293242),
	.w8(32'hbbded18a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7ce8b),
	.w1(32'hbb2c4242),
	.w2(32'hbb64ba4d),
	.w3(32'h3b8bda68),
	.w4(32'hbb2eecca),
	.w5(32'h3bda97b2),
	.w6(32'h3b0fca4f),
	.w7(32'hbb985d4a),
	.w8(32'h3b9efd25),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddd713),
	.w1(32'h3b599632),
	.w2(32'h3a0a0136),
	.w3(32'h3b89d5ec),
	.w4(32'h3ac53914),
	.w5(32'hbb8afe38),
	.w6(32'hba9a5dcb),
	.w7(32'hba90ddd8),
	.w8(32'hbb68dece),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33e1a8),
	.w1(32'hbb8d1478),
	.w2(32'hbb28d558),
	.w3(32'hbba0b734),
	.w4(32'hbb21503a),
	.w5(32'hbab825d3),
	.w6(32'hbbb8cb58),
	.w7(32'h3a1e6468),
	.w8(32'hbb3d81a4),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8eccd),
	.w1(32'hbbd7ae78),
	.w2(32'hbbe6b535),
	.w3(32'hba8806a1),
	.w4(32'hbb98c815),
	.w5(32'h3bcea874),
	.w6(32'hbb8d1c5a),
	.w7(32'hbb99f425),
	.w8(32'h3c4edb27),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49b414),
	.w1(32'h3c5a93b1),
	.w2(32'h3c3de47a),
	.w3(32'h3c2996a3),
	.w4(32'h3b8ee378),
	.w5(32'hbb8ca422),
	.w6(32'h3c921491),
	.w7(32'h3c46168a),
	.w8(32'hbaaf0e21),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcd23a),
	.w1(32'hbb8ef49c),
	.w2(32'hba80bb8e),
	.w3(32'hba91b3d7),
	.w4(32'hba8ef77d),
	.w5(32'h3b41bdee),
	.w6(32'hba83f01e),
	.w7(32'hbb0e7239),
	.w8(32'h3b304a88),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e0219),
	.w1(32'hbb4d7216),
	.w2(32'hbb89219e),
	.w3(32'hbbe7d616),
	.w4(32'hbb26a524),
	.w5(32'hbc050785),
	.w6(32'hb9e05a3d),
	.w7(32'hbb982d57),
	.w8(32'hbbd640e4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7cdf),
	.w1(32'hba18abaa),
	.w2(32'hbb1356ad),
	.w3(32'hbba9c24b),
	.w4(32'h3a76e2e8),
	.w5(32'h3b39161b),
	.w6(32'hbb6917f4),
	.w7(32'h39ddc918),
	.w8(32'h3b24ccbc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f85f1),
	.w1(32'hba48ea09),
	.w2(32'hbb365f27),
	.w3(32'hbba446ec),
	.w4(32'h398974d0),
	.w5(32'hbc05ec23),
	.w6(32'h3ab71071),
	.w7(32'h3a765f0b),
	.w8(32'hbc37c311),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd433f9),
	.w1(32'hba4a17b9),
	.w2(32'hba6e20b7),
	.w3(32'hbab65f26),
	.w4(32'hbb00ad1c),
	.w5(32'hbb222521),
	.w6(32'hbb24da18),
	.w7(32'h3b16a346),
	.w8(32'hbbb32c12),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc1e27),
	.w1(32'hbbad438f),
	.w2(32'hbbd85df8),
	.w3(32'hbb39bfa1),
	.w4(32'hbba79b8d),
	.w5(32'h3b9d2fc9),
	.w6(32'hbbc6120b),
	.w7(32'hbb9ab415),
	.w8(32'h3c09f1bb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19c21f),
	.w1(32'h3c02d54f),
	.w2(32'hbaae9ebf),
	.w3(32'hba79f281),
	.w4(32'hbb2fb308),
	.w5(32'h3a6ce503),
	.w6(32'h3c0e15dd),
	.w7(32'h3ba1d85e),
	.w8(32'h3a8448ca),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad72eb0),
	.w1(32'h3b9e8152),
	.w2(32'hbb0d377c),
	.w3(32'h3b4efdcf),
	.w4(32'hbb10e5ad),
	.w5(32'h3b7ab4c9),
	.w6(32'h3b8f9858),
	.w7(32'hbb185df6),
	.w8(32'h3b104f64),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule