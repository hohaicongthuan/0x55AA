module layer_10_featuremap_408(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8595830),
	.w1(32'h37064301),
	.w2(32'h375be1c9),
	.w3(32'hb8341b49),
	.w4(32'h37d261d7),
	.w5(32'h38286487),
	.w6(32'hb83f138c),
	.w7(32'h37e28a43),
	.w8(32'h37b44346),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba466be),
	.w1(32'h3acf93d5),
	.w2(32'h3ab770ad),
	.w3(32'h3b68388b),
	.w4(32'hba19a0ad),
	.w5(32'hba23c9b9),
	.w6(32'h3b4ad718),
	.w7(32'hb9e54942),
	.w8(32'hb90687ca),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fd24e1),
	.w1(32'hb6d79943),
	.w2(32'hb766c18f),
	.w3(32'hb7db929d),
	.w4(32'hb67621bd),
	.w5(32'hb74480d1),
	.w6(32'hb7f80d60),
	.w7(32'hb731c996),
	.w8(32'hb7895d66),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95afcd3),
	.w1(32'hb98448e3),
	.w2(32'hba5a4bdb),
	.w3(32'h389758e2),
	.w4(32'h37b981e9),
	.w5(32'hb9c74003),
	.w6(32'h38efa54e),
	.w7(32'h394a8dd5),
	.w8(32'hba1934dc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9702416),
	.w1(32'hb8ad2d72),
	.w2(32'hb8e2af29),
	.w3(32'hb93b6bc2),
	.w4(32'hb862a411),
	.w5(32'hb8c4524a),
	.w6(32'hb9367421),
	.w7(32'hb89d0e67),
	.w8(32'hb9042974),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b4ab7),
	.w1(32'hb799d0b1),
	.w2(32'hb7045904),
	.w3(32'hb88f4a8d),
	.w4(32'hb79e4a9a),
	.w5(32'hb787bbf7),
	.w6(32'hb8885cc4),
	.w7(32'hb74128e8),
	.w8(32'hb7fe3ac1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba722050),
	.w1(32'h3afb5b37),
	.w2(32'h3b7af87e),
	.w3(32'h393f1e4d),
	.w4(32'h3b4aebad),
	.w5(32'h3b8eb749),
	.w6(32'hba9258bc),
	.w7(32'h3b1c7c6a),
	.w8(32'h3b59e822),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa412a),
	.w1(32'h3bd8cd7f),
	.w2(32'h3b65e078),
	.w3(32'h3bd4542f),
	.w4(32'h3bfea42a),
	.w5(32'h3bcc9505),
	.w6(32'h3bac7396),
	.w7(32'h3af58a1d),
	.w8(32'h3b2685b0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b791c),
	.w1(32'hba4293a0),
	.w2(32'hb9f87832),
	.w3(32'hb8f82273),
	.w4(32'hba3bbb55),
	.w5(32'hb95cdf13),
	.w6(32'h39442174),
	.w7(32'hb88ee5b2),
	.w8(32'h3a3d2955),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c08e8),
	.w1(32'h3a64409a),
	.w2(32'h3ae4158b),
	.w3(32'h3c0b5560),
	.w4(32'h39c98e25),
	.w5(32'hba9123d3),
	.w6(32'h3c09314f),
	.w7(32'h39e56469),
	.w8(32'h3a6919c4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39623a7e),
	.w1(32'hb966c2be),
	.w2(32'hb7792987),
	.w3(32'h382cc5a1),
	.w4(32'hb9520b9d),
	.w5(32'hb8684f2a),
	.w6(32'h38f421b7),
	.w7(32'hb8ac6344),
	.w8(32'h39034c56),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab760dc),
	.w1(32'hbb2a55e8),
	.w2(32'h3a735276),
	.w3(32'h39f45291),
	.w4(32'hba47a3ac),
	.w5(32'h3b34e922),
	.w6(32'h38c340fc),
	.w7(32'hb96ddc2b),
	.w8(32'h3b894eb3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0cf7c),
	.w1(32'h3a6d4821),
	.w2(32'h3b3deddb),
	.w3(32'h3bade2d1),
	.w4(32'h3b09e918),
	.w5(32'h3afc10c8),
	.w6(32'h3bb0dc35),
	.w7(32'h3b20620f),
	.w8(32'h3b678c4e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38cfb2),
	.w1(32'h3b268197),
	.w2(32'h3b3b8518),
	.w3(32'h3abfa54b),
	.w4(32'h3b14dd03),
	.w5(32'h3b22fb8b),
	.w6(32'h3aee433d),
	.w7(32'h3ab00d8f),
	.w8(32'h3b1912ae),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b985f5c),
	.w1(32'h36c89727),
	.w2(32'hba323bf0),
	.w3(32'h3b5112c0),
	.w4(32'hbb435835),
	.w5(32'hbb3bae02),
	.w6(32'h3b8b3e1c),
	.w7(32'hbaa994ed),
	.w8(32'hbabf291b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c108187),
	.w1(32'h3ad03950),
	.w2(32'h3b251c4b),
	.w3(32'h3c0532ac),
	.w4(32'h3b08a7fb),
	.w5(32'hb97a9ea3),
	.w6(32'h3bf4e440),
	.w7(32'h3b3b8d9a),
	.w8(32'h3acd3f88),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3969560e),
	.w1(32'hb959e450),
	.w2(32'hb994e903),
	.w3(32'h39564844),
	.w4(32'hb9a0df30),
	.w5(32'hb99cd42b),
	.w6(32'hb85838aa),
	.w7(32'hb9d7bc4b),
	.w8(32'hba242a5a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf69b26),
	.w1(32'h3b654954),
	.w2(32'h3ba099b7),
	.w3(32'h3bcfe428),
	.w4(32'h3b1c3aae),
	.w5(32'h3bac3d77),
	.w6(32'h3bcd7f93),
	.w7(32'h3a586c8c),
	.w8(32'h3b35f514),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c1150),
	.w1(32'h3b06f475),
	.w2(32'h3b850603),
	.w3(32'h3b0e009c),
	.w4(32'h3aab75c0),
	.w5(32'h3b382584),
	.w6(32'h3b1e8670),
	.w7(32'h3a897e98),
	.w8(32'h3b067b5f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb877dc25),
	.w1(32'hb8267f23),
	.w2(32'hb889f1bc),
	.w3(32'hb8f62bf7),
	.w4(32'hb8c6b8b5),
	.w5(32'hb8db61d3),
	.w6(32'hb8aea9db),
	.w7(32'h36a77c52),
	.w8(32'hb518a23a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb930ffc2),
	.w1(32'hb519b8c9),
	.w2(32'hb78c9382),
	.w3(32'hb9206b29),
	.w4(32'hb391d9e9),
	.w5(32'hb827a30e),
	.w6(32'hb930dadc),
	.w7(32'hb7d31f7e),
	.w8(32'hb8dc2a65),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd1bfd),
	.w1(32'hba7358d1),
	.w2(32'h3a75ae55),
	.w3(32'hb697ec78),
	.w4(32'hbad8cc1b),
	.w5(32'h39710228),
	.w6(32'h38ca0499),
	.w7(32'hba9cf576),
	.w8(32'h3a3859d1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c768438),
	.w1(32'h3aeecd40),
	.w2(32'h3b887218),
	.w3(32'h3c669a37),
	.w4(32'h3b01fee9),
	.w5(32'h3b054eb3),
	.w6(32'h3c376193),
	.w7(32'h3aff5370),
	.w8(32'h3b908c3c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1312b0),
	.w1(32'hba02dc02),
	.w2(32'hb8ea2f2c),
	.w3(32'h3befc5e5),
	.w4(32'hbb07e352),
	.w5(32'hbb06f7fc),
	.w6(32'h3c143ecf),
	.w7(32'hba2e062a),
	.w8(32'hb80e9251),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c426ba0),
	.w1(32'hb8957d8c),
	.w2(32'h39f254e7),
	.w3(32'h3c2258e1),
	.w4(32'hbb387328),
	.w5(32'hbb310480),
	.w6(32'h3c42936f),
	.w7(32'hba2791e0),
	.w8(32'hb9fa6848),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6ce9b),
	.w1(32'h39d26d74),
	.w2(32'hb98fb1fb),
	.w3(32'h39a15747),
	.w4(32'h39a67744),
	.w5(32'h373bc78e),
	.w6(32'h390a58a4),
	.w7(32'hb91ee879),
	.w8(32'hb8b78d8e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae1eab),
	.w1(32'hb92de245),
	.w2(32'hb9429e97),
	.w3(32'hb997a5f1),
	.w4(32'hb90fe00e),
	.w5(32'hb909d5aa),
	.w6(32'hb9a33e76),
	.w7(32'hb94212d1),
	.w8(32'hb95676c9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e6ed0),
	.w1(32'hba41d189),
	.w2(32'h3abec5d7),
	.w3(32'h390dce61),
	.w4(32'hbb0fa58e),
	.w5(32'hbb8a5c22),
	.w6(32'h3b3caa81),
	.w7(32'h3a829d1d),
	.w8(32'h3acedb50),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a535037),
	.w1(32'hbb1fe3cf),
	.w2(32'hb8e1705b),
	.w3(32'h39feb225),
	.w4(32'hbb563267),
	.w5(32'hba6ebb35),
	.w6(32'h3a855b6b),
	.w7(32'hbb105a1e),
	.w8(32'h3967cefd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccec1e),
	.w1(32'hba63ccba),
	.w2(32'hba222932),
	.w3(32'h3baff46d),
	.w4(32'hbb28f07d),
	.w5(32'hbb54cf79),
	.w6(32'h3bfbdc86),
	.w7(32'hba9225e5),
	.w8(32'hb9057221),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886e1c2),
	.w1(32'hb86471f3),
	.w2(32'hb818d3ef),
	.w3(32'hb8678934),
	.w4(32'hb86bc557),
	.w5(32'hb7e2f5f0),
	.w6(32'hb89f1fd0),
	.w7(32'hb8a4f293),
	.w8(32'hb868e62b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7338fc8),
	.w1(32'h36392def),
	.w2(32'hb88726e3),
	.w3(32'hb85b754d),
	.w4(32'hb882e179),
	.w5(32'hb8ca1b8e),
	.w6(32'hb8a18912),
	.w7(32'hb8431325),
	.w8(32'hb9127451),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c5b70),
	.w1(32'hb94e8ad6),
	.w2(32'hb900e783),
	.w3(32'h3b1fc928),
	.w4(32'hba68312b),
	.w5(32'hba8a11e0),
	.w6(32'h3b4ad93f),
	.w7(32'hb98630d3),
	.w8(32'h38a5bcaa),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67bc3a),
	.w1(32'h399d2d17),
	.w2(32'h392b526c),
	.w3(32'h3b525d69),
	.w4(32'hba33f8b7),
	.w5(32'hba7b6d3a),
	.w6(32'h3b458f10),
	.w7(32'hb9c1c018),
	.w8(32'hb9ea7fa8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e3533),
	.w1(32'h38bbafcc),
	.w2(32'h392a3181),
	.w3(32'hb86f5e4d),
	.w4(32'h381a7655),
	.w5(32'hb92c2097),
	.w6(32'h391829bc),
	.w7(32'h39116888),
	.w8(32'h3a034020),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a368b70),
	.w1(32'h3a8c07d9),
	.w2(32'h3abfd724),
	.w3(32'h3aa846e0),
	.w4(32'h3accf464),
	.w5(32'h3b11d177),
	.w6(32'h389db78a),
	.w7(32'h3902bd16),
	.w8(32'h38288039),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd27e96),
	.w1(32'hba0c18d1),
	.w2(32'hbb0bb7a9),
	.w3(32'h3b67eb48),
	.w4(32'hbb0d7048),
	.w5(32'hbb26d57d),
	.w6(32'h3a86fc56),
	.w7(32'hba9147a3),
	.w8(32'hbadf8e05),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63224f),
	.w1(32'hbb6e529a),
	.w2(32'hba026b3d),
	.w3(32'h3c49a615),
	.w4(32'hbbfa489a),
	.w5(32'hbb83edcf),
	.w6(32'h3c66b48a),
	.w7(32'hbb368409),
	.w8(32'h3986e115),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd4e5a),
	.w1(32'hbbc282d3),
	.w2(32'hb93d1d7e),
	.w3(32'h3bdccdd9),
	.w4(32'hbc0edc86),
	.w5(32'hbba5db65),
	.w6(32'h3c3b2586),
	.w7(32'hbb86adad),
	.w8(32'h3ae9a707),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f311c),
	.w1(32'h3a474643),
	.w2(32'h39fb638d),
	.w3(32'h3b0791d5),
	.w4(32'hb9c12257),
	.w5(32'hba677bf2),
	.w6(32'h3b1e1e44),
	.w7(32'h3a38130b),
	.w8(32'h3880921d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb800bf13),
	.w1(32'h39241d5d),
	.w2(32'h38e5ba42),
	.w3(32'hb85fa30d),
	.w4(32'h3903ad8a),
	.w5(32'h387466cc),
	.w6(32'hb8f44ea9),
	.w7(32'h37a212d2),
	.w8(32'hb81e5f09),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c8b87),
	.w1(32'hb906907c),
	.w2(32'hb950ad92),
	.w3(32'hb9828767),
	.w4(32'hb86ac369),
	.w5(32'hb8c19838),
	.w6(32'hb99495e3),
	.w7(32'hb91ad2a8),
	.w8(32'hb96733b3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c9aa9),
	.w1(32'hbab89b26),
	.w2(32'hba58398a),
	.w3(32'h3a2788d2),
	.w4(32'hb9be5171),
	.w5(32'h3a67ba66),
	.w6(32'hba1b9616),
	.w7(32'hb9082e47),
	.w8(32'h3ad29419),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e9571),
	.w1(32'h3a411d06),
	.w2(32'h3b4fb0dd),
	.w3(32'h3c200758),
	.w4(32'h3ad1d941),
	.w5(32'h3a8c9b31),
	.w6(32'h3c31a670),
	.w7(32'h3b903773),
	.w8(32'h3b80c937),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fc328),
	.w1(32'hb95b2c45),
	.w2(32'hb78e1d07),
	.w3(32'h3bf74628),
	.w4(32'hbb2e4590),
	.w5(32'hbb1fdc2a),
	.w6(32'h3c1741d5),
	.w7(32'hbaa8647c),
	.w8(32'hba1950ee),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ace16),
	.w1(32'hb914aa24),
	.w2(32'hba2d7261),
	.w3(32'h3c0c6fc7),
	.w4(32'hbb28b94b),
	.w5(32'hbb8820d5),
	.w6(32'h3c27f01f),
	.w7(32'hbab599f4),
	.w8(32'hbac1663b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c146e24),
	.w1(32'h39b28663),
	.w2(32'h3896ce05),
	.w3(32'h3c05d07b),
	.w4(32'h385da40b),
	.w5(32'hbac28af9),
	.w6(32'h3bfd5ca6),
	.w7(32'h379ff9bc),
	.w8(32'h3a06e801),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac51c95),
	.w1(32'h3b7457b5),
	.w2(32'h3bc8ea66),
	.w3(32'h3b272117),
	.w4(32'h3ba6c57e),
	.w5(32'h3bd408e8),
	.w6(32'h3a3a234c),
	.w7(32'h3b328899),
	.w8(32'h3b3808ca),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e54c9b),
	.w1(32'h38f4e079),
	.w2(32'h394d8f64),
	.w3(32'hb8669ee9),
	.w4(32'h38e1d995),
	.w5(32'h38b49780),
	.w6(32'hb858ae8b),
	.w7(32'h38bbd657),
	.w8(32'h398f68c5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c737fc),
	.w1(32'h39a419cc),
	.w2(32'h39d5fb2b),
	.w3(32'h394b4bc3),
	.w4(32'h39c7f32a),
	.w5(32'h3a0cb80c),
	.w6(32'h39894d3d),
	.w7(32'h3a0ac16d),
	.w8(32'h3a6e0012),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07157f),
	.w1(32'hb8cfba1e),
	.w2(32'hb92d9a19),
	.w3(32'hba216666),
	.w4(32'hb90b5dbc),
	.w5(32'hb86b5551),
	.w6(32'hb9eeeed9),
	.w7(32'h386ff34e),
	.w8(32'h398186e8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd64212),
	.w1(32'h3a8d4cd3),
	.w2(32'h3a500efe),
	.w3(32'h3baf9457),
	.w4(32'h39e65c6c),
	.w5(32'h361336d4),
	.w6(32'h3b981714),
	.w7(32'h39ee422a),
	.w8(32'hb697d60c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af92360),
	.w1(32'h3a4c870a),
	.w2(32'h3a145bb5),
	.w3(32'h3ae15cea),
	.w4(32'h3a57fe08),
	.w5(32'h3a534fb5),
	.w6(32'h3aadffdc),
	.w7(32'h39ce5db5),
	.w8(32'h3997d5b4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1c881),
	.w1(32'h3a85cbc0),
	.w2(32'h3b80ed78),
	.w3(32'h3bc0f5d1),
	.w4(32'h3ab34bf5),
	.w5(32'h3ac83f74),
	.w6(32'h3b9c077d),
	.w7(32'hb7c0f0fb),
	.w8(32'h3aa2b580),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac503fa),
	.w1(32'h397b31df),
	.w2(32'h39f572d6),
	.w3(32'h3ae12812),
	.w4(32'h3a205943),
	.w5(32'h3a8c6929),
	.w6(32'h3af0ad91),
	.w7(32'h39ad018d),
	.w8(32'h39dd4234),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947c11f),
	.w1(32'h393d1c3d),
	.w2(32'h369fc3e8),
	.w3(32'h3877314b),
	.w4(32'h370363bf),
	.w5(32'hb8b4f941),
	.w6(32'h390d4e2e),
	.w7(32'h389bb7fa),
	.w8(32'hb7f241ee),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ef1508),
	.w1(32'h37808047),
	.w2(32'h37a36568),
	.w3(32'hb7b14896),
	.w4(32'hb75d20f6),
	.w5(32'h37a0537d),
	.w6(32'hb822b8df),
	.w7(32'hb77d566e),
	.w8(32'h3774de51),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e865b),
	.w1(32'h38680f86),
	.w2(32'h39cfda99),
	.w3(32'h38d286d0),
	.w4(32'h38cbb5fd),
	.w5(32'h3988a944),
	.w6(32'h39dc7b5a),
	.w7(32'h3996b16c),
	.w8(32'h39ad9f19),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb804a2ec),
	.w1(32'hba697a27),
	.w2(32'hb93c7bc4),
	.w3(32'hb9a16d54),
	.w4(32'hbacdc023),
	.w5(32'hba59c15c),
	.w6(32'h39dd750b),
	.w7(32'hba40ca83),
	.w8(32'hb96009e0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f8a7f),
	.w1(32'h364a96a0),
	.w2(32'hb8c470a4),
	.w3(32'hb8c60ef4),
	.w4(32'hb9a499ea),
	.w5(32'hb994160a),
	.w6(32'h39ae9268),
	.w7(32'h38d8bde8),
	.w8(32'h39c0f1ff),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc01ba8),
	.w1(32'h3b0145f3),
	.w2(32'h3b10a64b),
	.w3(32'h3bb2e55e),
	.w4(32'h3b0636ea),
	.w5(32'h3ad6c20b),
	.w6(32'h3b9ad1ab),
	.w7(32'h3af6c4d1),
	.w8(32'h3a845c40),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf4913),
	.w1(32'h3ad8d9d8),
	.w2(32'h3a59760f),
	.w3(32'h3b9f74a5),
	.w4(32'h3b395237),
	.w5(32'h39405473),
	.w6(32'h3b8f324e),
	.w7(32'h3b011bfc),
	.w8(32'h3aa62bd1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a72dc7),
	.w1(32'h37216866),
	.w2(32'hb75886ea),
	.w3(32'hb896fc21),
	.w4(32'h37af581c),
	.w5(32'hb73396ee),
	.w6(32'hb8c1baa7),
	.w7(32'hb787fd58),
	.w8(32'hb8217c8d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abdb9d),
	.w1(32'hb6b303f4),
	.w2(32'hb7fe0c36),
	.w3(32'hb8a16cfb),
	.w4(32'h35e2df48),
	.w5(32'hb79e679b),
	.w6(32'hb8d9eac4),
	.w7(32'hb81c16c4),
	.w8(32'hb85ed389),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a2b76),
	.w1(32'hb8932d89),
	.w2(32'hb6ee7335),
	.w3(32'hb9569a9d),
	.w4(32'hb9062830),
	.w5(32'hb8faea58),
	.w6(32'hb96b0b8f),
	.w7(32'hb93e42ff),
	.w8(32'hb9377b99),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a1d83),
	.w1(32'hb87c82a0),
	.w2(32'hb89278ce),
	.w3(32'hb93ff014),
	.w4(32'hb865fdc0),
	.w5(32'hb874ac57),
	.w6(32'hb95359b6),
	.w7(32'hb8a899e1),
	.w8(32'hb8b5b1c7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b913c6f),
	.w1(32'h3b217a13),
	.w2(32'h3b668b94),
	.w3(32'h3bb55d65),
	.w4(32'h3b9b85c3),
	.w5(32'hb9003a15),
	.w6(32'h3b983a9c),
	.w7(32'h3b72b6df),
	.w8(32'h3b699cba),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c399125),
	.w1(32'h3b24ff72),
	.w2(32'h3b207b80),
	.w3(32'h3c1452de),
	.w4(32'h39c5defb),
	.w5(32'h3a6a56ee),
	.w6(32'h3c32f7c4),
	.w7(32'hb8c20019),
	.w8(32'h39f5ed08),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bcc51),
	.w1(32'h3a6148ac),
	.w2(32'h3b35c9fa),
	.w3(32'h3c42b4da),
	.w4(32'h3ab1923a),
	.w5(32'h3b223ee6),
	.w6(32'h3c4b53df),
	.w7(32'h3b195849),
	.w8(32'h3b5aac27),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bfa43),
	.w1(32'hbb4b00f9),
	.w2(32'h3a39aaed),
	.w3(32'h3c3c6470),
	.w4(32'hbbbc047f),
	.w5(32'hbb2624c1),
	.w6(32'h3c8ad3e5),
	.w7(32'hba5a4ded),
	.w8(32'h3b07944f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9315e00),
	.w1(32'h3738488a),
	.w2(32'hb82ddf07),
	.w3(32'hb92bd023),
	.w4(32'h37b4cd27),
	.w5(32'hb5ba7e40),
	.w6(32'hb94f2cae),
	.w7(32'hb804193c),
	.w8(32'hb8992cb5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993cf0a),
	.w1(32'hb7fcae20),
	.w2(32'hb8d464be),
	.w3(32'hb98c3ac7),
	.w4(32'hb7189c34),
	.w5(32'hb8bbfd23),
	.w6(32'hb9ae63c9),
	.w7(32'hb8d0b3ef),
	.w8(32'hb92eccca),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97901d4),
	.w1(32'h387bf50f),
	.w2(32'hb7d91c1c),
	.w3(32'hb970e508),
	.w4(32'h38c809d5),
	.w5(32'h36a832af),
	.w6(32'hb9a46c4b),
	.w7(32'h37059acf),
	.w8(32'hb8acbe47),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0ded5),
	.w1(32'h38c79036),
	.w2(32'h397a28c9),
	.w3(32'h3ad9f851),
	.w4(32'h3a0fcbdc),
	.w5(32'h3a2deb89),
	.w6(32'h3ad791e3),
	.w7(32'h3a14b4c9),
	.w8(32'h3a0bfc8e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9631d67),
	.w1(32'hb82551d6),
	.w2(32'hb859392b),
	.w3(32'hb9569914),
	.w4(32'h37b36417),
	.w5(32'hb6db27c2),
	.w6(32'hb986eadd),
	.w7(32'hb83e80d2),
	.w8(32'hb88eb64f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a821a53),
	.w1(32'h3a1f5595),
	.w2(32'h3947db27),
	.w3(32'h3b20279e),
	.w4(32'h3b353f8d),
	.w5(32'h3a5a0e68),
	.w6(32'h3a245344),
	.w7(32'h3ade2954),
	.w8(32'h3a5b1446),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1e6d0),
	.w1(32'h3b36b2de),
	.w2(32'h3af53ef8),
	.w3(32'h3bcea719),
	.w4(32'h3b57f2c4),
	.w5(32'h3b8e7b8c),
	.w6(32'h3ba399a0),
	.w7(32'h3b9dd9e4),
	.w8(32'h3b0d0c4f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba209ff),
	.w1(32'h3a1d27ce),
	.w2(32'h39ce772a),
	.w3(32'h3b83184b),
	.w4(32'hbab4be3e),
	.w5(32'hbafab192),
	.w6(32'h3b6cb4ae),
	.w7(32'hba9614aa),
	.w8(32'hba84d5a5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85b00d),
	.w1(32'h3941c17d),
	.w2(32'h3a30fc06),
	.w3(32'h3b866df6),
	.w4(32'h39b9ecbc),
	.w5(32'h39d54d00),
	.w6(32'h3ba0e417),
	.w7(32'h3a5a8f75),
	.w8(32'h39c33c38),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8154398),
	.w1(32'hb91f8c95),
	.w2(32'h3a500bb5),
	.w3(32'h3a835b98),
	.w4(32'h3a7685a3),
	.w5(32'h3a14499b),
	.w6(32'h3a029de0),
	.w7(32'h39f4b17a),
	.w8(32'h3ae83279),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967cc2),
	.w1(32'hb7f76dc6),
	.w2(32'hb9d0b0b9),
	.w3(32'h3b7b98b0),
	.w4(32'hba3f8045),
	.w5(32'hbac2c8a0),
	.w6(32'h3b87ee87),
	.w7(32'hb9b655a5),
	.w8(32'hb9e0833a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae071bc),
	.w1(32'h3a9f2ad6),
	.w2(32'h3ab51280),
	.w3(32'h3b0ed087),
	.w4(32'h3b076a85),
	.w5(32'h3b0e527d),
	.w6(32'h3a8e614f),
	.w7(32'h3a713b34),
	.w8(32'h3a3a088a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d7e596),
	.w1(32'hb73f2795),
	.w2(32'hb772de08),
	.w3(32'hb7a95ed4),
	.w4(32'hb6cfc9df),
	.w5(32'hb752ba09),
	.w6(32'hb7f546c7),
	.w7(32'hb771246d),
	.w8(32'hb7b41a95),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h330e11a5),
	.w1(32'h37c10920),
	.w2(32'h37182c5a),
	.w3(32'hb7a3c95b),
	.w4(32'h34f80827),
	.w5(32'hb7ceeaca),
	.w6(32'hb7d9c253),
	.w7(32'h36af026f),
	.w8(32'hb7209b54),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b97850),
	.w1(32'hb9302f65),
	.w2(32'hb9656c28),
	.w3(32'h38deb593),
	.w4(32'hb88cbd88),
	.w5(32'hb91820a2),
	.w6(32'hb882547e),
	.w7(32'hb9605ac7),
	.w8(32'hb88bb876),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78b1464),
	.w1(32'h39613d48),
	.w2(32'h385c0d05),
	.w3(32'hb8629d3a),
	.w4(32'hb6e3df43),
	.w5(32'hb9970107),
	.w6(32'h399e0397),
	.w7(32'h39922f39),
	.w8(32'h390ad349),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef4ac7),
	.w1(32'hba43339a),
	.w2(32'hbadaae36),
	.w3(32'h3bd1f5b6),
	.w4(32'hbb02d1b0),
	.w5(32'hbb610447),
	.w6(32'h3bce7870),
	.w7(32'hbad10462),
	.w8(32'hbaf508dc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9560911),
	.w1(32'hb970bbf5),
	.w2(32'h39933227),
	.w3(32'hb9bbb243),
	.w4(32'hba5ee853),
	.w5(32'hba8f464b),
	.w6(32'h396abdc9),
	.w7(32'h39a7cbba),
	.w8(32'h39286972),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e8467),
	.w1(32'h3a847710),
	.w2(32'h3a29dfb4),
	.w3(32'h3b0e5784),
	.w4(32'hba4aa6d8),
	.w5(32'hbaf0ac18),
	.w6(32'h3b438556),
	.w7(32'hb9f05862),
	.w8(32'hba7b482c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3278e),
	.w1(32'h3a4950af),
	.w2(32'h3ac5d2ae),
	.w3(32'h3bec5dba),
	.w4(32'h3b639aab),
	.w5(32'h3b318a33),
	.w6(32'h3be206d3),
	.w7(32'h3b54f38f),
	.w8(32'h3b0872c5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada51ee),
	.w1(32'hbb3acc5d),
	.w2(32'h37e96c43),
	.w3(32'h3b0186ee),
	.w4(32'hbb861751),
	.w5(32'hbb30f581),
	.w6(32'h3b4b32fa),
	.w7(32'hbaf0b635),
	.w8(32'h3784870f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b773e58),
	.w1(32'h3aed1610),
	.w2(32'h3a9bc660),
	.w3(32'h3b7c060e),
	.w4(32'h3acab759),
	.w5(32'hbaa49be6),
	.w6(32'h3b7525fd),
	.w7(32'h3b4dfc5e),
	.w8(32'h3b6a3e08),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f53ce),
	.w1(32'h3943a4af),
	.w2(32'h3a24f0ce),
	.w3(32'h3b230d4f),
	.w4(32'hba96a828),
	.w5(32'hbb143cbf),
	.w6(32'h3ba27922),
	.w7(32'h3a32f428),
	.w8(32'hb9834061),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24ba8d),
	.w1(32'h3a98fe8d),
	.w2(32'h3aab5ba2),
	.w3(32'h3bfd666d),
	.w4(32'h371be946),
	.w5(32'hba84eb32),
	.w6(32'h3c0b81bc),
	.w7(32'h3a6e7e67),
	.w8(32'hb8a254f7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83b5f9),
	.w1(32'h3a4ddb82),
	.w2(32'h383d370c),
	.w3(32'h3b5bb28b),
	.w4(32'hb924ac68),
	.w5(32'hbb318ddc),
	.w6(32'h3b32117b),
	.w7(32'hb9689d11),
	.w8(32'hba947ea8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdee5b5),
	.w1(32'h3939fd8d),
	.w2(32'h3a852ade),
	.w3(32'h3b86b2ed),
	.w4(32'hbb33fe87),
	.w5(32'hbb23819c),
	.w6(32'h3bc78b9e),
	.w7(32'hba3d9391),
	.w8(32'hb9fbd319),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f04d8),
	.w1(32'hb88fa4c7),
	.w2(32'hb988373b),
	.w3(32'hb9c09cce),
	.w4(32'h36a587e3),
	.w5(32'hb72ea9b3),
	.w6(32'hb7ee2c16),
	.w7(32'h390f35e0),
	.w8(32'hb8bcaff4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb9c55),
	.w1(32'h3a95c1c0),
	.w2(32'h3b1f0e2a),
	.w3(32'h3bd1225f),
	.w4(32'hb94f3e3c),
	.w5(32'h3a03cb60),
	.w6(32'h3c035d9a),
	.w7(32'h3ad548f3),
	.w8(32'h3b24cb0f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b086a75),
	.w1(32'hbb3f3c5e),
	.w2(32'hb9ade57f),
	.w3(32'h3b579629),
	.w4(32'hbad380e4),
	.w5(32'hb9683d38),
	.w6(32'h3b2e6f87),
	.w7(32'h3a25ed28),
	.w8(32'h3b6d69bf),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09fe2f),
	.w1(32'h3b31bc8f),
	.w2(32'h3b3e38d9),
	.w3(32'h3b9aee5f),
	.w4(32'h3a395eed),
	.w5(32'hbabca24e),
	.w6(32'h3b3409ec),
	.w7(32'h3a07b389),
	.w8(32'hbaa0393d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30face),
	.w1(32'h39447ec2),
	.w2(32'hbac3ed9a),
	.w3(32'h3bf0364e),
	.w4(32'hbba78155),
	.w5(32'hbba3321a),
	.w6(32'h3bed7cee),
	.w7(32'hb9f3e3d8),
	.w8(32'hba314d9a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf50786),
	.w1(32'h3a1a2cac),
	.w2(32'h3a0ca5cd),
	.w3(32'h3bcbf0ce),
	.w4(32'hbaa638b9),
	.w5(32'hba2c1dd4),
	.w6(32'h3c0be0df),
	.w7(32'h3954a788),
	.w8(32'h39ea9687),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b476576),
	.w1(32'h3b1980e2),
	.w2(32'h3a842c8e),
	.w3(32'h3b473afd),
	.w4(32'h3b123dc7),
	.w5(32'h39c83d64),
	.w6(32'hb9e6f487),
	.w7(32'h3a10d15b),
	.w8(32'h3a5f7233),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26063e),
	.w1(32'hb929dc89),
	.w2(32'hba84085c),
	.w3(32'h389e33b7),
	.w4(32'hb8d7f052),
	.w5(32'hb9b35219),
	.w6(32'h37c6c72e),
	.w7(32'hb96c93b6),
	.w8(32'hb90f4b34),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05158e),
	.w1(32'h3b31a9f8),
	.w2(32'hba0d4812),
	.w3(32'h3b9117f0),
	.w4(32'h3b335fce),
	.w5(32'hbb18c1a4),
	.w6(32'hbaab6244),
	.w7(32'hbab9edcb),
	.w8(32'hbb69fa6d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967e227),
	.w1(32'hbac7999c),
	.w2(32'h39c5dcf9),
	.w3(32'h3a6670e9),
	.w4(32'hba72deec),
	.w5(32'h3ac3033b),
	.w6(32'h3a3d29b6),
	.w7(32'h3a0689db),
	.w8(32'h3b10eb7a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b2e79),
	.w1(32'hb89afe3f),
	.w2(32'h37ce18e4),
	.w3(32'hb89cedcf),
	.w4(32'hb9429e44),
	.w5(32'hb8860b11),
	.w6(32'hb8ef8fa0),
	.w7(32'hb989c2b2),
	.w8(32'hb7e91d98),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af11831),
	.w1(32'h39849d93),
	.w2(32'h3a3e1555),
	.w3(32'h3ab09542),
	.w4(32'h3903dd81),
	.w5(32'hb9c726cc),
	.w6(32'h3abddd68),
	.w7(32'h39626e22),
	.w8(32'hb965b977),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34ac13),
	.w1(32'h39f44309),
	.w2(32'h3aa7233d),
	.w3(32'h3b3c4494),
	.w4(32'h3a6aff8c),
	.w5(32'h3ac40172),
	.w6(32'h3b4a0a42),
	.w7(32'h3ae50ccd),
	.w8(32'h3aee2ef3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9acaa5),
	.w1(32'hb9ed540b),
	.w2(32'h396f8778),
	.w3(32'h3ba7b179),
	.w4(32'hba23cae1),
	.w5(32'hba26a6d5),
	.w6(32'h3bc3a798),
	.w7(32'hba1dadc1),
	.w8(32'h38b295d4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af607b3),
	.w1(32'h3993a854),
	.w2(32'hb9cbf242),
	.w3(32'h3ac19118),
	.w4(32'hbaf04cc4),
	.w5(32'hbb176cb3),
	.w6(32'h3b0c4fd2),
	.w7(32'hbabf93d4),
	.w8(32'hba20da90),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b822427),
	.w1(32'hb92f0499),
	.w2(32'hba53556c),
	.w3(32'h3b27ed82),
	.w4(32'hbaca7157),
	.w5(32'hba9be678),
	.w6(32'h3b1e2043),
	.w7(32'hba827ba0),
	.w8(32'hb98b188d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c63af),
	.w1(32'hba7f809e),
	.w2(32'h3a22bdae),
	.w3(32'h3b8c0b87),
	.w4(32'hba48def2),
	.w5(32'h3ab4aa56),
	.w6(32'h3b981b61),
	.w7(32'hba8b8785),
	.w8(32'h38f14bef),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcdbd9),
	.w1(32'h3ad7a3ef),
	.w2(32'h3b2e63e6),
	.w3(32'h3b89baeb),
	.w4(32'h3a58194d),
	.w5(32'hbaa08708),
	.w6(32'h3b7e957c),
	.w7(32'h3a8fb88e),
	.w8(32'h3a4d9bd5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75f484),
	.w1(32'hba4ba293),
	.w2(32'hbacb05ad),
	.w3(32'h3b60cb13),
	.w4(32'hba93fc22),
	.w5(32'hbacb5979),
	.w6(32'h3b85a74f),
	.w7(32'hba75bc29),
	.w8(32'hba615ed8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce2925),
	.w1(32'h38b9a238),
	.w2(32'h382605cc),
	.w3(32'h38b43df6),
	.w4(32'h38aa02b7),
	.w5(32'h37a9b00e),
	.w6(32'h3830b471),
	.w7(32'h383f3f14),
	.w8(32'hb64da0fe),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ae66f),
	.w1(32'h39d0f8c6),
	.w2(32'h38f0c5de),
	.w3(32'h39c4fb82),
	.w4(32'h38ffb208),
	.w5(32'hb85f1c63),
	.w6(32'h39ad27ce),
	.w7(32'hb7dcbabc),
	.w8(32'hb8ad7ad2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bbe3b6),
	.w1(32'hb89d74c2),
	.w2(32'h37ede724),
	.w3(32'h38c681f0),
	.w4(32'hb8d0b480),
	.w5(32'hb8ab3160),
	.w6(32'h38e2a239),
	.w7(32'hb88ec29a),
	.w8(32'hb83db612),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929ae93),
	.w1(32'hb8043573),
	.w2(32'hb90fbfed),
	.w3(32'hb929bb25),
	.w4(32'hb8867105),
	.w5(32'h375d4b4a),
	.w6(32'hb96de711),
	.w7(32'hb92005c8),
	.w8(32'hb8d9a6e8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc32ac4),
	.w1(32'hba467481),
	.w2(32'hba9f6c28),
	.w3(32'h3b96d3b8),
	.w4(32'hbad972f7),
	.w5(32'hbae39318),
	.w6(32'h3bb7dca5),
	.w7(32'hba878992),
	.w8(32'hba4f2525),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a153d4a),
	.w1(32'hb982a3ed),
	.w2(32'hb9556118),
	.w3(32'h398a9614),
	.w4(32'hb91a8041),
	.w5(32'hb8b6a128),
	.w6(32'h39c6dde5),
	.w7(32'hb93cdaf9),
	.w8(32'h37f67a7c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9770fdb),
	.w1(32'h39dff56a),
	.w2(32'h3ab41eeb),
	.w3(32'h3a2817b8),
	.w4(32'h3aa35173),
	.w5(32'h3abcb619),
	.w6(32'hb9fb60dc),
	.w7(32'h3a2d9aa7),
	.w8(32'h3a8686e7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8a7e9),
	.w1(32'h39cc548b),
	.w2(32'h3a837365),
	.w3(32'h3baacb31),
	.w4(32'hbb269c8b),
	.w5(32'hba8f7939),
	.w6(32'h3bb341de),
	.w7(32'hbab57c1c),
	.w8(32'h394e79fd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2e026),
	.w1(32'hb8b96adc),
	.w2(32'hb8adb514),
	.w3(32'hb924d07d),
	.w4(32'hb8c77bde),
	.w5(32'hb8caf4d5),
	.w6(32'hb94e6d1e),
	.w7(32'hb90b500d),
	.w8(32'hb883b89f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8faef16),
	.w1(32'h38019558),
	.w2(32'h39a60264),
	.w3(32'hb9e64c1a),
	.w4(32'hb86573d7),
	.w5(32'h37b1174e),
	.w6(32'hb800b21e),
	.w7(32'h39651574),
	.w8(32'h39d4e544),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd30b5),
	.w1(32'hb8717513),
	.w2(32'hb7cfc702),
	.w3(32'hb89f24b9),
	.w4(32'hb86264c8),
	.w5(32'hb7cdda26),
	.w6(32'hb89c499a),
	.w7(32'hb8863ffe),
	.w8(32'hb85123a0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911d126),
	.w1(32'hb8e7f908),
	.w2(32'hb794c215),
	.w3(32'hb967e18c),
	.w4(32'hba0ee6fd),
	.w5(32'hb9e6da0b),
	.w6(32'h37a8beb8),
	.w7(32'hb88f4d44),
	.w8(32'h38de58d0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b867ac2),
	.w1(32'h3b8df859),
	.w2(32'h3b6745fe),
	.w3(32'h3b3a8c3b),
	.w4(32'h3b65defc),
	.w5(32'h3b7a1f8c),
	.w6(32'h3b00a8f8),
	.w7(32'h3a238f48),
	.w8(32'h39dd2405),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babfc8c),
	.w1(32'h382abc82),
	.w2(32'h3ad00651),
	.w3(32'h3b8be0e1),
	.w4(32'h39480907),
	.w5(32'hb9bb3449),
	.w6(32'h3b935068),
	.w7(32'h39a654d8),
	.w8(32'h3adc3d4b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d6125),
	.w1(32'h3a1363b9),
	.w2(32'h39ac5a6c),
	.w3(32'h39610e5b),
	.w4(32'h39fe23a3),
	.w5(32'h354e1ca1),
	.w6(32'hb88d2a26),
	.w7(32'h39a090d8),
	.w8(32'h39ccc68b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8fd24),
	.w1(32'h3a8f1925),
	.w2(32'h3ac523ca),
	.w3(32'h3aff9928),
	.w4(32'h3a287be9),
	.w5(32'h3ade27e0),
	.w6(32'h3b2aba39),
	.w7(32'h3a179730),
	.w8(32'h3aa37d40),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb632e),
	.w1(32'hb89cd045),
	.w2(32'hb7a4e890),
	.w3(32'h3aa85b7a),
	.w4(32'hba202461),
	.w5(32'hba1df12a),
	.w6(32'h3a7ee581),
	.w7(32'hba2400c9),
	.w8(32'hba01fff5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b584a7a),
	.w1(32'h3a257637),
	.w2(32'h39ebdc5e),
	.w3(32'h3b3297f0),
	.w4(32'h3a1183ec),
	.w5(32'hb7da5029),
	.w6(32'h3b5d0394),
	.w7(32'h39e5047b),
	.w8(32'hb92982fb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc16142),
	.w1(32'h3a55b94d),
	.w2(32'h3a32dfe4),
	.w3(32'h3b6cefac),
	.w4(32'hbadf479a),
	.w5(32'hbb4037ca),
	.w6(32'h3b6b2f01),
	.w7(32'hba36243b),
	.w8(32'hba87d251),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8abbd9),
	.w1(32'h3aed3f69),
	.w2(32'h3b650544),
	.w3(32'h3b8fab02),
	.w4(32'h3aedaa0b),
	.w5(32'h3afdf11b),
	.w6(32'h3b699be8),
	.w7(32'h3b0a8b9a),
	.w8(32'h3b58e97b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f87e3),
	.w1(32'hb9101e8f),
	.w2(32'hba15e581),
	.w3(32'h3b738bc2),
	.w4(32'hba845813),
	.w5(32'hbab4c7b7),
	.w6(32'h3b829250),
	.w7(32'hba49ae58),
	.w8(32'hba60d416),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81f7e8),
	.w1(32'h3a9aa287),
	.w2(32'h3a85f24c),
	.w3(32'h3b2f0532),
	.w4(32'hba1a31fd),
	.w5(32'hb9eb46ea),
	.w6(32'h3b0a2313),
	.w7(32'h3a9452b5),
	.w8(32'h3a96c0ad),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7df7b8),
	.w1(32'hb97f94a5),
	.w2(32'h3a56f235),
	.w3(32'h3ba06ca2),
	.w4(32'h3a3ba753),
	.w5(32'h3a9c8bd9),
	.w6(32'h3b4bfa73),
	.w7(32'h357b5d48),
	.w8(32'h395a76b0),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba81684),
	.w1(32'h3a0fe4ce),
	.w2(32'hba46665a),
	.w3(32'h3b5e4f80),
	.w4(32'hba677e4c),
	.w5(32'hbb2919e9),
	.w6(32'h3b91c87c),
	.w7(32'hb9a0efdb),
	.w8(32'hbae2aa0b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bda5a),
	.w1(32'h3aa9df36),
	.w2(32'h3ad1b15c),
	.w3(32'h3b3e1585),
	.w4(32'h3a1b49a6),
	.w5(32'h3a2d1a6e),
	.w6(32'h3b2f8f48),
	.w7(32'h3aaf716e),
	.w8(32'h3b1e48aa),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae969f7),
	.w1(32'h3907347d),
	.w2(32'hb8839717),
	.w3(32'h3aa80af1),
	.w4(32'hb9e65982),
	.w5(32'hba2aa314),
	.w6(32'h3ae4228d),
	.w7(32'hb78bb53d),
	.w8(32'hb91e1ac4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8903f),
	.w1(32'hbb63fc77),
	.w2(32'hbafb0ca7),
	.w3(32'h3b90e124),
	.w4(32'hbbac0ad2),
	.w5(32'hbb36b615),
	.w6(32'h3bc59a15),
	.w7(32'hbb72c9cf),
	.w8(32'hb8ced3ba),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c8381),
	.w1(32'h3a3254c2),
	.w2(32'hba6337ae),
	.w3(32'h3b4476f0),
	.w4(32'h390e7216),
	.w5(32'hbac69492),
	.w6(32'h3b528557),
	.w7(32'hb92be17c),
	.w8(32'hba772596),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3806889d),
	.w1(32'h3848d20c),
	.w2(32'h38861132),
	.w3(32'h3778bc02),
	.w4(32'h38318333),
	.w5(32'h388b00b8),
	.w6(32'h37733e28),
	.w7(32'h37fc21f2),
	.w8(32'h37d40174),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb866e2d2),
	.w1(32'hb7fae1ea),
	.w2(32'h383da2c0),
	.w3(32'hb6f04159),
	.w4(32'h37923b17),
	.w5(32'h38b2ef56),
	.w6(32'hb883fb35),
	.w7(32'hb8b2c893),
	.w8(32'hb7a1cab6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb114a),
	.w1(32'hba3df50b),
	.w2(32'hba56a4c5),
	.w3(32'h3a681d81),
	.w4(32'hba067442),
	.w5(32'hba5d6a79),
	.w6(32'h39fb8aef),
	.w7(32'hba381eaf),
	.w8(32'hb9f636c0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba044bd),
	.w1(32'hb6a5b287),
	.w2(32'hba0e7742),
	.w3(32'h3b480fda),
	.w4(32'hbafb8549),
	.w5(32'hbad88feb),
	.w6(32'h3b724bc6),
	.w7(32'hb966d1c9),
	.w8(32'hba32344b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc51aaa),
	.w1(32'hb7e6e2fc),
	.w2(32'h3a89523a),
	.w3(32'h3bc2b1db),
	.w4(32'h3a1d6756),
	.w5(32'h39c9288e),
	.w6(32'h3bc56fd3),
	.w7(32'hb923ed9f),
	.w8(32'h379842ae),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb817bf5a),
	.w1(32'h3819a73e),
	.w2(32'h37f168d7),
	.w3(32'hb79ce0df),
	.w4(32'h37a99063),
	.w5(32'h37a3242d),
	.w6(32'h37b1f970),
	.w7(32'h38085235),
	.w8(32'h35f2e9eb),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb689c),
	.w1(32'h397acd1d),
	.w2(32'h3a04a9d5),
	.w3(32'h3ba66812),
	.w4(32'h398fee16),
	.w5(32'hb887b6a8),
	.w6(32'h3bbe3908),
	.w7(32'h3a660f37),
	.w8(32'h3a91c596),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b649503),
	.w1(32'h3a74fa74),
	.w2(32'h39123ce1),
	.w3(32'h3b2b1d78),
	.w4(32'h39a55ee4),
	.w5(32'hba9cdd71),
	.w6(32'h3b51dac2),
	.w7(32'h394ef42f),
	.w8(32'hb9a16575),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc5b0a),
	.w1(32'h3b649feb),
	.w2(32'h3b62ab57),
	.w3(32'h3b3773e9),
	.w4(32'h3b27b1b8),
	.w5(32'h3b0ad06b),
	.w6(32'hba0a0095),
	.w7(32'h3aa073c6),
	.w8(32'h3b1ba2e1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c3889),
	.w1(32'hbab969fe),
	.w2(32'hba06d520),
	.w3(32'h3b5b84f1),
	.w4(32'hbb45ffda),
	.w5(32'hbb0fa69f),
	.w6(32'h3bcf11c6),
	.w7(32'hbaab0c7e),
	.w8(32'h3a9daf69),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae76f71),
	.w1(32'h389563dc),
	.w2(32'hb933d69a),
	.w3(32'h3a8ecdc1),
	.w4(32'hb9ad08e0),
	.w5(32'hba46673a),
	.w6(32'h3a931920),
	.w7(32'hba8374e9),
	.w8(32'hb9875e95),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b2291),
	.w1(32'hba5eeb0e),
	.w2(32'hba58c017),
	.w3(32'hba036e23),
	.w4(32'hb9da5c30),
	.w5(32'hb9e91403),
	.w6(32'hba150adf),
	.w7(32'hba04828e),
	.w8(32'h38428eee),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aca32),
	.w1(32'hb9fd8154),
	.w2(32'hb9fd3690),
	.w3(32'h3b687080),
	.w4(32'hba8ec4e4),
	.w5(32'hba90b222),
	.w6(32'h3b9fb5ff),
	.w7(32'hba0c7bf4),
	.w8(32'h39c6a5c9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb5eae),
	.w1(32'hbb4230f0),
	.w2(32'hbb0a186a),
	.w3(32'h3b5ee434),
	.w4(32'hbb908c30),
	.w5(32'hbb1b84f3),
	.w6(32'h3b596818),
	.w7(32'hbb587f84),
	.w8(32'hba4cbf53),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f75ab),
	.w1(32'hbae532b2),
	.w2(32'h39ab42f6),
	.w3(32'h3b16f6f4),
	.w4(32'hbb2e1f74),
	.w5(32'hba0e87ed),
	.w6(32'h3b452c40),
	.w7(32'hbac5c5b4),
	.w8(32'h3a2d84c5),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994e476),
	.w1(32'h3832c670),
	.w2(32'h393f56d3),
	.w3(32'h3a16b7e7),
	.w4(32'h39c9f1ac),
	.w5(32'h39cee3f7),
	.w6(32'h3980692a),
	.w7(32'h3a0a1c42),
	.w8(32'h39e908a0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3802dafe),
	.w1(32'hb904d703),
	.w2(32'hb80955c9),
	.w3(32'hb82040ec),
	.w4(32'hb991eafd),
	.w5(32'hb9858d6b),
	.w6(32'hb8ff3ea9),
	.w7(32'hb9321f39),
	.w8(32'h3708cc93),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fab30),
	.w1(32'h3ab83b49),
	.w2(32'h3aebffb0),
	.w3(32'h3b242a13),
	.w4(32'hb8deb2fb),
	.w5(32'h3989f578),
	.w6(32'h3b2b8f60),
	.w7(32'h3a147a89),
	.w8(32'h3a941c14),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcc758),
	.w1(32'h38966246),
	.w2(32'h39ed3e73),
	.w3(32'hb93c4306),
	.w4(32'h38873031),
	.w5(32'h39bf8b66),
	.w6(32'hb9e7cd47),
	.w7(32'hb60f3932),
	.w8(32'h39975197),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f80f9),
	.w1(32'h39304cea),
	.w2(32'hb7acc625),
	.w3(32'h3b36aa16),
	.w4(32'hb8a03b10),
	.w5(32'hba5fa059),
	.w6(32'h3b6c4c97),
	.w7(32'hb976c6cf),
	.w8(32'hb90c1e0e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a648c),
	.w1(32'hb96379ee),
	.w2(32'h37d5b5d0),
	.w3(32'h38bbca7d),
	.w4(32'hb90c810e),
	.w5(32'h393ca53a),
	.w6(32'h37e113fb),
	.w7(32'hb8d4773a),
	.w8(32'h38a3a605),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99d3fb),
	.w1(32'hba5332cd),
	.w2(32'h3a9bbdba),
	.w3(32'h3a72f7e8),
	.w4(32'hba910611),
	.w5(32'h3a87b9f8),
	.w6(32'h3b2b8666),
	.w7(32'hb79e0c97),
	.w8(32'h3b03e558),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db75d8),
	.w1(32'hb8fc0404),
	.w2(32'hb8a81466),
	.w3(32'hb95062ec),
	.w4(32'hb922241b),
	.w5(32'hb8804f75),
	.w6(32'hb963b8e4),
	.w7(32'hb92fce7f),
	.w8(32'hb856ced1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa50ef),
	.w1(32'hb97294ee),
	.w2(32'hb8c616db),
	.w3(32'hb954e945),
	.w4(32'hb93f7d1a),
	.w5(32'hb8c23cbe),
	.w6(32'hb915a0cd),
	.w7(32'hb91c0c0d),
	.w8(32'h38da036d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40f12d),
	.w1(32'hb9525f51),
	.w2(32'hba595637),
	.w3(32'h3ae9651a),
	.w4(32'hbaecb313),
	.w5(32'hbae65eb6),
	.w6(32'h3b18e40c),
	.w7(32'hbaa50206),
	.w8(32'hba8ec2f4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c268ab6),
	.w1(32'h3b0651cc),
	.w2(32'h3a1851ef),
	.w3(32'h3c1702dc),
	.w4(32'h3b137262),
	.w5(32'h3ac8fdff),
	.w6(32'h3c113b84),
	.w7(32'h3a8a8d3d),
	.w8(32'h3a8170cd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86b943),
	.w1(32'hbaf1e211),
	.w2(32'h3884c9e9),
	.w3(32'h3a3bbbd6),
	.w4(32'hbb3ab5a5),
	.w5(32'hba598ddd),
	.w6(32'h3ac14789),
	.w7(32'hbaed1f09),
	.w8(32'h3908299f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f8a66),
	.w1(32'hb9ff64e7),
	.w2(32'hba0595da),
	.w3(32'h3b6f37ed),
	.w4(32'hbadf1c5a),
	.w5(32'hbab8663f),
	.w6(32'h3b83d863),
	.w7(32'hbadd6e30),
	.w8(32'hba00cfbd),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c907ef),
	.w1(32'hba03172d),
	.w2(32'h38b50c14),
	.w3(32'h3a0249c5),
	.w4(32'hb9acc463),
	.w5(32'hba34c634),
	.w6(32'h39d14ccb),
	.w7(32'hba36e6c9),
	.w8(32'hba57ca10),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a2aac),
	.w1(32'h3a4b9d18),
	.w2(32'h3bb4df24),
	.w3(32'h3c0721d5),
	.w4(32'h3a840f05),
	.w5(32'h3b420cfe),
	.w6(32'h3c30b216),
	.w7(32'h3bb0e21c),
	.w8(32'h3bbab31a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf116b),
	.w1(32'h3a68d19c),
	.w2(32'h3ace3d49),
	.w3(32'h3ba54ad2),
	.w4(32'hba56b3a7),
	.w5(32'hb98f77ea),
	.w6(32'h3bb20293),
	.w7(32'h399090cb),
	.w8(32'h3a50c3cb),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc94e95),
	.w1(32'h3a22ce00),
	.w2(32'h3ac1657b),
	.w3(32'h3b9d6627),
	.w4(32'h3a1fb4c2),
	.w5(32'h396be369),
	.w6(32'h3bab00e3),
	.w7(32'h39735113),
	.w8(32'h3a437600),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944e719),
	.w1(32'hb91e14f4),
	.w2(32'hb90d3641),
	.w3(32'hb94cf36c),
	.w4(32'hb972b887),
	.w5(32'hb982e2bb),
	.w6(32'hb955a865),
	.w7(32'hb995b47a),
	.w8(32'hb9cd944d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854477),
	.w1(32'h39f5d554),
	.w2(32'h398bda13),
	.w3(32'h3b3c853b),
	.w4(32'hba3af8e2),
	.w5(32'hbade9bdd),
	.w6(32'h3b26d4e6),
	.w7(32'hba560e2f),
	.w8(32'hba7daaac),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f167b),
	.w1(32'hb7b11226),
	.w2(32'hb7d7898c),
	.w3(32'hb91390fe),
	.w4(32'hb6dc8c4c),
	.w5(32'hb7d0ba64),
	.w6(32'hb91bab39),
	.w7(32'hb7ffd81b),
	.w8(32'hb8832916),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17cd35),
	.w1(32'hba36e2b9),
	.w2(32'hb7b2167b),
	.w3(32'h3a0666cd),
	.w4(32'hba4d1b15),
	.w5(32'hb9f65252),
	.w6(32'h3a8ec47f),
	.w7(32'h38f855ff),
	.w8(32'h3981ed69),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fcd24),
	.w1(32'h3a033604),
	.w2(32'h399d3972),
	.w3(32'h39e493d0),
	.w4(32'hb8f14f85),
	.w5(32'h3831d696),
	.w6(32'h3a17fa21),
	.w7(32'hb98b6eae),
	.w8(32'h39653440),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ab28),
	.w1(32'hb9cc1b57),
	.w2(32'h3afa5780),
	.w3(32'h3b6f1916),
	.w4(32'hb839a140),
	.w5(32'h3a246882),
	.w6(32'h3b686041),
	.w7(32'h3a09c050),
	.w8(32'h3af526d3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb841d664),
	.w1(32'hb6e7656f),
	.w2(32'hb7d10c4f),
	.w3(32'hb83d3384),
	.w4(32'hb6132caa),
	.w5(32'hb7892652),
	.w6(32'hb858a762),
	.w7(32'hb7a66841),
	.w8(32'hb80c2242),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a10265),
	.w1(32'h34c7a66f),
	.w2(32'h385e4c87),
	.w3(32'hb7667d0d),
	.w4(32'h3889f400),
	.w5(32'h38c65212),
	.w6(32'hb8871eb6),
	.w7(32'hb72942df),
	.w8(32'h382b33b2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08cebc),
	.w1(32'hb8e823c0),
	.w2(32'h38fce63e),
	.w3(32'h3af6a9f8),
	.w4(32'hba087116),
	.w5(32'hba8ee53b),
	.w6(32'h3ac38647),
	.w7(32'hba8559aa),
	.w8(32'hba43e9bd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58f726),
	.w1(32'hba79a1d5),
	.w2(32'hb7c32026),
	.w3(32'h3b82e397),
	.w4(32'hbaa29fc8),
	.w5(32'hbabfa184),
	.w6(32'h3b66491f),
	.w7(32'hb9fb0dfe),
	.w8(32'hb9d433ea),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8f397),
	.w1(32'hba13867c),
	.w2(32'hba9d525a),
	.w3(32'h3ae88632),
	.w4(32'h39b67dc0),
	.w5(32'h393ccd44),
	.w6(32'hb98776df),
	.w7(32'hb98d1706),
	.w8(32'hb97b1414),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6b35e),
	.w1(32'hb9005f11),
	.w2(32'h391691aa),
	.w3(32'h39fdf520),
	.w4(32'h39d050b9),
	.w5(32'h39fc06c9),
	.w6(32'h3a5021a0),
	.w7(32'h39c96956),
	.w8(32'h3a8607ef),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39e1d4),
	.w1(32'h3b7a56b3),
	.w2(32'h3c0bfe19),
	.w3(32'h3c41d8f9),
	.w4(32'h3b942162),
	.w5(32'h3be09a94),
	.w6(32'h3c18eb38),
	.w7(32'h3b574073),
	.w8(32'h3bc0f8e3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fbb5b),
	.w1(32'hbb4cd2a1),
	.w2(32'hba0a2449),
	.w3(32'h3c27ad4e),
	.w4(32'hbbaf5f78),
	.w5(32'hbbac2377),
	.w6(32'h3c1ffa19),
	.w7(32'hbb941c69),
	.w8(32'hbb352049),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a4536),
	.w1(32'h394d184e),
	.w2(32'h397fcf91),
	.w3(32'hb7c8807c),
	.w4(32'h3a1ab494),
	.w5(32'h3a8899e1),
	.w6(32'hb97529fa),
	.w7(32'h3a52db69),
	.w8(32'h3aaf57f8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b0e8b9),
	.w1(32'h380c2129),
	.w2(32'h38103fdd),
	.w3(32'hb7b24a36),
	.w4(32'h381be723),
	.w5(32'h3840f6b7),
	.w6(32'hb84088dc),
	.w7(32'h3744619b),
	.w8(32'h37e107c6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70ead3d),
	.w1(32'h38fc712f),
	.w2(32'h3987eaa5),
	.w3(32'h38986cc3),
	.w4(32'h3956723a),
	.w5(32'h39ab9469),
	.w6(32'h38307f5d),
	.w7(32'h38f50709),
	.w8(32'h399a6cc5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90296ec),
	.w1(32'hb7f64ac7),
	.w2(32'hb800d935),
	.w3(32'hb8c42c66),
	.w4(32'h35edcbda),
	.w5(32'hb61b1497),
	.w6(32'hb8f5425e),
	.w7(32'hb7d31a47),
	.w8(32'hb7ed0f17),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d6ece),
	.w1(32'h3a64b167),
	.w2(32'h3ab872fa),
	.w3(32'h3a60fb7a),
	.w4(32'h3ae5b6ea),
	.w5(32'h3ada7aee),
	.w6(32'hb9a010b8),
	.w7(32'h3aa94333),
	.w8(32'h3abed9fe),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840508),
	.w1(32'h3a254f39),
	.w2(32'hbacde9b9),
	.w3(32'h3b698439),
	.w4(32'hb8f2a194),
	.w5(32'hbb02eeb0),
	.w6(32'h3b93da58),
	.w7(32'h3a2be3c9),
	.w8(32'hb84eddde),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0652a2),
	.w1(32'h3acaccc8),
	.w2(32'h3ac451e2),
	.w3(32'h3bd2932d),
	.w4(32'hbb02698e),
	.w5(32'hbb0124d6),
	.w6(32'h3be4ee6f),
	.w7(32'hba306a74),
	.w8(32'hbacea989),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a850c65),
	.w1(32'hba2ad836),
	.w2(32'hb8932b3a),
	.w3(32'h3a0936ca),
	.w4(32'hbaab2f06),
	.w5(32'hba862a43),
	.w6(32'h3aa81b9c),
	.w7(32'hba3482a3),
	.w8(32'hb977fc44),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74d60b),
	.w1(32'h3bc7195f),
	.w2(32'h3bb160b6),
	.w3(32'h3b3304e2),
	.w4(32'h3bfd3204),
	.w5(32'h3afad5a5),
	.w6(32'h3b871625),
	.w7(32'h3c14c1f3),
	.w8(32'h3a71ee67),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb731d),
	.w1(32'hbc1d04fe),
	.w2(32'h3b2f2169),
	.w3(32'hba5a1f8c),
	.w4(32'hbbd985ee),
	.w5(32'h3c48ea90),
	.w6(32'h3af66716),
	.w7(32'h3b9b9c66),
	.w8(32'h3c01f2d5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83af30),
	.w1(32'hbc163f91),
	.w2(32'h3aedfddd),
	.w3(32'h3b840928),
	.w4(32'hbc26d61a),
	.w5(32'hbb67ecef),
	.w6(32'h3a9b35cf),
	.w7(32'hbc1debd1),
	.w8(32'h3a95796a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae862e),
	.w1(32'h3b915735),
	.w2(32'h3bd6eee0),
	.w3(32'hba2bb355),
	.w4(32'h3bb8b463),
	.w5(32'h3c976083),
	.w6(32'h3b215214),
	.w7(32'h3a878c15),
	.w8(32'h3c09c893),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f998a),
	.w1(32'h3ada798f),
	.w2(32'hbb20cbde),
	.w3(32'hbb868af1),
	.w4(32'h3b4ff5e0),
	.w5(32'h3b3ca5ba),
	.w6(32'hba008eff),
	.w7(32'h3b38caab),
	.w8(32'h396953f0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b705936),
	.w1(32'hbbc76a61),
	.w2(32'hbaf0ee02),
	.w3(32'h3a4ec1a5),
	.w4(32'h3b51fee9),
	.w5(32'h3c12bce1),
	.w6(32'h3b3bf3dc),
	.w7(32'hb8f9747a),
	.w8(32'hbb8899ab),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f94f5),
	.w1(32'hbb7b0a31),
	.w2(32'hbb685ecc),
	.w3(32'hbb41a776),
	.w4(32'hbc49a292),
	.w5(32'hbb763165),
	.w6(32'h3a00b55b),
	.w7(32'hbbf3f6c6),
	.w8(32'h3b699947),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd3f74),
	.w1(32'hba569748),
	.w2(32'h39cba397),
	.w3(32'h3b88bc8d),
	.w4(32'hbb06300a),
	.w5(32'hbbd50710),
	.w6(32'h3c5079cd),
	.w7(32'h3b1c220a),
	.w8(32'h3abc3aa0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb259562),
	.w1(32'h3cc14386),
	.w2(32'h3c683945),
	.w3(32'hbac71dce),
	.w4(32'h3cd57d15),
	.w5(32'h3c618ee8),
	.w6(32'hbaf94e1b),
	.w7(32'h3bb50a27),
	.w8(32'h3c7523af),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1cc62),
	.w1(32'h3a621867),
	.w2(32'h3a96abe5),
	.w3(32'h3c9b36cf),
	.w4(32'hbbbc0d90),
	.w5(32'h3a2021cd),
	.w6(32'h3c6931d3),
	.w7(32'hbb0e66c1),
	.w8(32'h3a04c94c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69b107),
	.w1(32'h3a1f1ff1),
	.w2(32'hbb1304e2),
	.w3(32'h3b4ea2e4),
	.w4(32'hbb4d68b4),
	.w5(32'hbbbef319),
	.w6(32'hba32d270),
	.w7(32'h3badd829),
	.w8(32'hbb75cd72),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902fa98),
	.w1(32'h3bcd297e),
	.w2(32'hbb76c7b4),
	.w3(32'h391bae35),
	.w4(32'h3bd87440),
	.w5(32'hbc2c589e),
	.w6(32'h393f1389),
	.w7(32'h3c1ff960),
	.w8(32'h3b271177),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d85e),
	.w1(32'hbb68ea3e),
	.w2(32'h3bd3113f),
	.w3(32'h3b8f1937),
	.w4(32'hbaef3e18),
	.w5(32'h3c35f357),
	.w6(32'h3b92b6f3),
	.w7(32'hbaa9072c),
	.w8(32'h3bed4e11),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab20b06),
	.w1(32'h3a8e911f),
	.w2(32'h3c250da6),
	.w3(32'h3b238b4c),
	.w4(32'h3a442ae5),
	.w5(32'hb9c21032),
	.w6(32'h3b6adff2),
	.w7(32'h3c001d07),
	.w8(32'h37f5df3f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ed2bb),
	.w1(32'hbbb56064),
	.w2(32'hbadf420e),
	.w3(32'h3c62638a),
	.w4(32'hbb02bf5d),
	.w5(32'h3c3ebb27),
	.w6(32'h3c55c2d1),
	.w7(32'h3c19ed7e),
	.w8(32'hba909127),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79c6e0),
	.w1(32'hb9ce37db),
	.w2(32'hba1ed174),
	.w3(32'h3c31be6b),
	.w4(32'hbb99e6af),
	.w5(32'h3c6b4544),
	.w6(32'h3b0d26e6),
	.w7(32'hbbf545d6),
	.w8(32'hba318f23),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20e2a1),
	.w1(32'hb9a68993),
	.w2(32'h3c283acc),
	.w3(32'hbac6e0e0),
	.w4(32'h3b815b24),
	.w5(32'h3c66e834),
	.w6(32'h3c123e56),
	.w7(32'h3b779169),
	.w8(32'h3af3fce9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8a3ea),
	.w1(32'hbc4d3c2a),
	.w2(32'h3aee8592),
	.w3(32'h3ad685ee),
	.w4(32'hbc598398),
	.w5(32'hbb8f750a),
	.w6(32'hbb08bf84),
	.w7(32'hbc3819de),
	.w8(32'hba5dd081),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b19a0),
	.w1(32'hbb6ce002),
	.w2(32'hbb99daa5),
	.w3(32'hbb41b699),
	.w4(32'hbc353d80),
	.w5(32'hbbd24866),
	.w6(32'hbc501768),
	.w7(32'hbc176bba),
	.w8(32'hba2b4121),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb549063),
	.w1(32'hbbb2d073),
	.w2(32'hbb99fa21),
	.w3(32'h3abb28a4),
	.w4(32'hbbe4268f),
	.w5(32'hbb07912c),
	.w6(32'h3a2ceacc),
	.w7(32'h3bbdbe14),
	.w8(32'h3b22db94),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1898aa),
	.w1(32'h3bcf94a0),
	.w2(32'h3aecf145),
	.w3(32'h3bd4ea26),
	.w4(32'h3c725d8e),
	.w5(32'hbb885506),
	.w6(32'hbb0e1ffb),
	.w7(32'h3be97643),
	.w8(32'h3ba25ebe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc130d7),
	.w1(32'h3b449a51),
	.w2(32'h3bffd69f),
	.w3(32'hbb27d69c),
	.w4(32'h3bbba273),
	.w5(32'h3be458c6),
	.w6(32'h3b84a1a8),
	.w7(32'h3a70c161),
	.w8(32'h3c2c3503),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13a928),
	.w1(32'h3a09d30a),
	.w2(32'hbb908f7a),
	.w3(32'h3b9ed9f4),
	.w4(32'h3c3248cb),
	.w5(32'hbade7602),
	.w6(32'hb9a0b782),
	.w7(32'hbba90552),
	.w8(32'hbbc53b37),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b12b9),
	.w1(32'hbb8ded88),
	.w2(32'hbb9471f9),
	.w3(32'h3b50e8c5),
	.w4(32'h3a2ccea6),
	.w5(32'h3b4f4570),
	.w6(32'h3b7fa4a1),
	.w7(32'h3b33efc9),
	.w8(32'h3a9c645b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96e431),
	.w1(32'h3b766be1),
	.w2(32'hbae43a3c),
	.w3(32'h3c0dcbc6),
	.w4(32'h3b5e5552),
	.w5(32'hbc09f8d0),
	.w6(32'h3b241cfd),
	.w7(32'h3b8f2713),
	.w8(32'h3b01a582),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc92de),
	.w1(32'hbb90e990),
	.w2(32'hbc3b08b8),
	.w3(32'h3abde6f6),
	.w4(32'hbc3e5250),
	.w5(32'hbc4516fe),
	.w6(32'h3b320516),
	.w7(32'hbc15a621),
	.w8(32'hbc5f3f5e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9163f7),
	.w1(32'h3c9a2b85),
	.w2(32'hbcd169e2),
	.w3(32'hba1bfae4),
	.w4(32'h3cb270a7),
	.w5(32'hbcdaa96e),
	.w6(32'hbc0c3224),
	.w7(32'h3c5c96f3),
	.w8(32'hbc69f531),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe7b1c),
	.w1(32'hbbc47d6e),
	.w2(32'hbbce86dc),
	.w3(32'hb9236311),
	.w4(32'hbc91c3ec),
	.w5(32'h3c7715c0),
	.w6(32'h3c186fb4),
	.w7(32'hbc85e533),
	.w8(32'hbb60733d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51c953),
	.w1(32'h3c18c720),
	.w2(32'h3c6eab2d),
	.w3(32'h3a402d90),
	.w4(32'h3bb5672d),
	.w5(32'h3c817307),
	.w6(32'h3b021b14),
	.w7(32'h3b44546e),
	.w8(32'h3c3a8035),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12173e),
	.w1(32'hbc216ae7),
	.w2(32'hba054784),
	.w3(32'hbb80f138),
	.w4(32'hbb2ab047),
	.w5(32'hbae1d763),
	.w6(32'hba360fa1),
	.w7(32'hbbbfaf0d),
	.w8(32'hb95dfa19),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa1f09),
	.w1(32'hbb2207d6),
	.w2(32'hbc4bdbb8),
	.w3(32'h3ba6bb16),
	.w4(32'h3be3a30d),
	.w5(32'hbbf1c6df),
	.w6(32'h3c078114),
	.w7(32'hbc1192db),
	.w8(32'hbb428adc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bf45a),
	.w1(32'hbbdb3ae2),
	.w2(32'hbbd335de),
	.w3(32'h3966cd03),
	.w4(32'hbc022341),
	.w5(32'hbc0d0365),
	.w6(32'h3bd5cd22),
	.w7(32'hbbf5f2b7),
	.w8(32'hbb8cb17a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3571c),
	.w1(32'hbc1a0211),
	.w2(32'hbc141881),
	.w3(32'hbbbe51d7),
	.w4(32'hbc0405c0),
	.w5(32'h3b418214),
	.w6(32'hbc057df6),
	.w7(32'h392de22d),
	.w8(32'h3aef7960),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57b4f0),
	.w1(32'h3a96cc06),
	.w2(32'hbc06d947),
	.w3(32'hbb6f92a7),
	.w4(32'h3b88e24a),
	.w5(32'hbbae5ddd),
	.w6(32'h3b966364),
	.w7(32'hbb0f8e6b),
	.w8(32'hbba3c4a4),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e33d13),
	.w1(32'h3b276146),
	.w2(32'h3c167aef),
	.w3(32'h3a1ac381),
	.w4(32'h3a42c9eb),
	.w5(32'h3cb546bd),
	.w6(32'h39ba774e),
	.w7(32'hbb24f0c5),
	.w8(32'h3bf8bff7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc051958),
	.w1(32'hb9fa66cd),
	.w2(32'h3be245a8),
	.w3(32'hbc097ba7),
	.w4(32'h3bafba3b),
	.w5(32'h3cded5dd),
	.w6(32'hbc18b2e0),
	.w7(32'h3ca54934),
	.w8(32'h3c6b4c62),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba02b99),
	.w1(32'hbb23c4ca),
	.w2(32'h3b98e42b),
	.w3(32'h3c826144),
	.w4(32'hbb06ae9e),
	.w5(32'hb9fdcef9),
	.w6(32'h3baea893),
	.w7(32'hbb329010),
	.w8(32'h3bbdd70e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98ed81),
	.w1(32'h3c5019a6),
	.w2(32'h3c8870f6),
	.w3(32'h3b2e9c90),
	.w4(32'h3c903914),
	.w5(32'h3b8f50f8),
	.w6(32'h3ba48b09),
	.w7(32'h3c7407ce),
	.w8(32'h3be09390),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b2725),
	.w1(32'hb9225267),
	.w2(32'hbc49a33c),
	.w3(32'h3c52de53),
	.w4(32'h3a9ecc3d),
	.w5(32'hbb393240),
	.w6(32'h3c1cef88),
	.w7(32'h3a4116e8),
	.w8(32'hbb5b0733),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd57c1b),
	.w1(32'hba7e85b5),
	.w2(32'h3c138da9),
	.w3(32'hbc09b7bf),
	.w4(32'hbb2cfbf9),
	.w5(32'h3c859b96),
	.w6(32'hbbd4836f),
	.w7(32'hbb56688c),
	.w8(32'h3b8ebbc2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9380dc),
	.w1(32'h3bafe532),
	.w2(32'hbad6cb78),
	.w3(32'h3bf3b523),
	.w4(32'h3ca7eebe),
	.w5(32'h3b097d6f),
	.w6(32'h3c2ac288),
	.w7(32'h3cdfbd04),
	.w8(32'hbb17c5c5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c469304),
	.w1(32'h3c4a3add),
	.w2(32'h3c124628),
	.w3(32'h3b873350),
	.w4(32'h3cc8861b),
	.w5(32'hbc0151ff),
	.w6(32'h39216b5d),
	.w7(32'h39b14e7d),
	.w8(32'h38d790ff),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40c352),
	.w1(32'h3aecdca6),
	.w2(32'h3abaf5a8),
	.w3(32'h3bfadaba),
	.w4(32'h3b9a7d82),
	.w5(32'h3ba23511),
	.w6(32'h3b84baf4),
	.w7(32'h3c40daeb),
	.w8(32'hb9c93a4d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e651e),
	.w1(32'h3a712fe9),
	.w2(32'hbb8f6f38),
	.w3(32'h3ba0831d),
	.w4(32'hbb410a17),
	.w5(32'h3c406797),
	.w6(32'h3c0be620),
	.w7(32'h3b9f96e4),
	.w8(32'h3bacfa7b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64ae44),
	.w1(32'h3b04616f),
	.w2(32'h3bbc3a73),
	.w3(32'hbbe52481),
	.w4(32'hbab1234b),
	.w5(32'h3b85658e),
	.w6(32'h3a114f70),
	.w7(32'h3bca2f4f),
	.w8(32'h3bab5e5a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f21f5),
	.w1(32'h3a2c7441),
	.w2(32'hbb9a327c),
	.w3(32'hbb81ef8a),
	.w4(32'hbabc860f),
	.w5(32'hbbbf7d82),
	.w6(32'hbb8a1dcd),
	.w7(32'hbb20d8ef),
	.w8(32'hbb7613fa),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc29e66),
	.w1(32'hba33d3b4),
	.w2(32'h3c33879e),
	.w3(32'hba8b610c),
	.w4(32'hbaf4a624),
	.w5(32'h3c47c142),
	.w6(32'hbbb23846),
	.w7(32'hb82354df),
	.w8(32'h3bef1a4f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e5c0),
	.w1(32'h3b40cd53),
	.w2(32'h391386d8),
	.w3(32'h3b8c04cd),
	.w4(32'h3b5a4b66),
	.w5(32'hba202d95),
	.w6(32'h3c0e8a67),
	.w7(32'h3bdf2797),
	.w8(32'hbb8fb34e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c1d32),
	.w1(32'h3b6fd55c),
	.w2(32'h39f76585),
	.w3(32'h3c2c3689),
	.w4(32'hbafe26d5),
	.w5(32'hbc1c133e),
	.w6(32'h3bda313a),
	.w7(32'h3c18b315),
	.w8(32'h3c067c6c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39083b),
	.w1(32'h3c785fb5),
	.w2(32'h3ae74236),
	.w3(32'h3c1b7b25),
	.w4(32'h3c740ae8),
	.w5(32'h3bfe4021),
	.w6(32'h3c0a4a13),
	.w7(32'hbb9544a3),
	.w8(32'h3b39f9b3),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a7e53),
	.w1(32'hbbc543c4),
	.w2(32'h3b42bb44),
	.w3(32'h3af5be1c),
	.w4(32'h3aa3d77e),
	.w5(32'h3a9aed44),
	.w6(32'h3b240896),
	.w7(32'hbb5920de),
	.w8(32'hbc11f56b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a1eb6),
	.w1(32'hbbe2eb07),
	.w2(32'h389c5047),
	.w3(32'hbb32f8a8),
	.w4(32'hbc0840ae),
	.w5(32'h3abb9907),
	.w6(32'hbbceb78b),
	.w7(32'h3b1d28ff),
	.w8(32'h3bb8b9c0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b753215),
	.w1(32'hbbdfab67),
	.w2(32'hbbeb9621),
	.w3(32'h3b042e65),
	.w4(32'hbb5aef7c),
	.w5(32'hbb69f996),
	.w6(32'h3b05682b),
	.w7(32'hbb171aad),
	.w8(32'hbc5434db),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe19c05),
	.w1(32'hbbf4cb38),
	.w2(32'hbbbd38af),
	.w3(32'hbc1b6164),
	.w4(32'hbc8f08fa),
	.w5(32'h3c15113b),
	.w6(32'hbb721502),
	.w7(32'hbbe83bfd),
	.w8(32'hbbb30b6f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57fadd),
	.w1(32'hba91aa32),
	.w2(32'hbc1f14f1),
	.w3(32'hbbadf743),
	.w4(32'hbbee947d),
	.w5(32'h3c5d7755),
	.w6(32'hbb931d28),
	.w7(32'hbb1ab308),
	.w8(32'hbae0f197),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cb654),
	.w1(32'hbc240739),
	.w2(32'hbba632dc),
	.w3(32'hbc595bab),
	.w4(32'hbc95171a),
	.w5(32'hbc4e59bf),
	.w6(32'hbbfacb16),
	.w7(32'hbb9ab2ac),
	.w8(32'hbbce1719),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b883fd1),
	.w1(32'hb8d490ee),
	.w2(32'h3c843b38),
	.w3(32'hbb064b38),
	.w4(32'h3b9949b1),
	.w5(32'h3c73ded3),
	.w6(32'hb8d4e664),
	.w7(32'h3c0e968e),
	.w8(32'h3c32e534),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c242f84),
	.w1(32'h3b8add9c),
	.w2(32'hba2101c7),
	.w3(32'h3acd8c0a),
	.w4(32'hba3a3cc4),
	.w5(32'h3b3a032d),
	.w6(32'hbaf1505b),
	.w7(32'h3a12f3fb),
	.w8(32'h3afd8ff7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5da70),
	.w1(32'hbb968244),
	.w2(32'h3bb7bebc),
	.w3(32'h3c1ff538),
	.w4(32'h3c3c1d39),
	.w5(32'h3c7506c3),
	.w6(32'h3c11d49d),
	.w7(32'h3ba7ef16),
	.w8(32'hbbd20aa2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule