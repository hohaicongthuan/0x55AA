module layer_10_featuremap_53(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc362ba0),
	.w1(32'h3bd680bc),
	.w2(32'hbbd7a915),
	.w3(32'hba927508),
	.w4(32'hbba0a949),
	.w5(32'hbb50c322),
	.w6(32'h3b46d641),
	.w7(32'hbbc97aea),
	.w8(32'h3b54698d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58ece3),
	.w1(32'hbc1def0e),
	.w2(32'h3b5edeba),
	.w3(32'h3b084312),
	.w4(32'hbc382b88),
	.w5(32'hbc076283),
	.w6(32'h3beeeef1),
	.w7(32'hbb6adc27),
	.w8(32'hbc15220c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c8b0c),
	.w1(32'h3a3add22),
	.w2(32'hbad67918),
	.w3(32'hbc174f39),
	.w4(32'hbc697410),
	.w5(32'hbb4472b7),
	.w6(32'hbc80c54a),
	.w7(32'hbc244d1b),
	.w8(32'hbc410f9c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa53128),
	.w1(32'h3b569e61),
	.w2(32'h3ad1c6b3),
	.w3(32'hba1962a1),
	.w4(32'hba656e1d),
	.w5(32'h3b0ba2cc),
	.w6(32'h3a9c2406),
	.w7(32'h3b0ca2ec),
	.w8(32'hba515cd4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affd351),
	.w1(32'hbb8845ad),
	.w2(32'h3a0b00de),
	.w3(32'h3c1fce6a),
	.w4(32'h3bcf3d78),
	.w5(32'h3c200fb5),
	.w6(32'h3bb713ea),
	.w7(32'h3c0d87f6),
	.w8(32'h3be93eb3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f167e),
	.w1(32'hbbb6a450),
	.w2(32'h3c1bcdfc),
	.w3(32'h3adfa81c),
	.w4(32'hbb811262),
	.w5(32'hbb8b443c),
	.w6(32'h3c0fb009),
	.w7(32'hbb3a7360),
	.w8(32'h3aa5bcce),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a9e47),
	.w1(32'h3c093802),
	.w2(32'h3b612e0a),
	.w3(32'hbcd54ffa),
	.w4(32'hbc3c3991),
	.w5(32'h3c2c0224),
	.w6(32'hbc8addd9),
	.w7(32'hbb26d82d),
	.w8(32'h3b800dac),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3646ff),
	.w1(32'h3b2062dd),
	.w2(32'h3bc35150),
	.w3(32'h3c4ea146),
	.w4(32'h3c60b9e2),
	.w5(32'h3c1b9f47),
	.w6(32'h3c14ba52),
	.w7(32'h3c85a503),
	.w8(32'h3c3a1ae5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdec4e7),
	.w1(32'h3afe5bf3),
	.w2(32'h3bf9b057),
	.w3(32'h3c8c752d),
	.w4(32'h3bf62358),
	.w5(32'h3a68d7b5),
	.w6(32'h3b31c584),
	.w7(32'hb73e6bf4),
	.w8(32'hbb768c2a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13d242),
	.w1(32'h3c0cb42a),
	.w2(32'hbc9fb984),
	.w3(32'h3b071c66),
	.w4(32'hba5d8097),
	.w5(32'hbc8a4dd6),
	.w6(32'h3b0582fe),
	.w7(32'hbbaab61c),
	.w8(32'hbcbc6784),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f27f6),
	.w1(32'hbc7d7b0f),
	.w2(32'h38030b81),
	.w3(32'hbb1376f8),
	.w4(32'hbc14ac41),
	.w5(32'h3b371ced),
	.w6(32'hbc67c0ce),
	.w7(32'hbc851629),
	.w8(32'h39500620),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a6d5e),
	.w1(32'hbbcced0f),
	.w2(32'hbba2a84c),
	.w3(32'hbba261f6),
	.w4(32'hbbb1b0cc),
	.w5(32'hbb8ce63c),
	.w6(32'hbbe1929e),
	.w7(32'hbb8dd410),
	.w8(32'h3b65e4ac),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ee76),
	.w1(32'hbbaebe82),
	.w2(32'hbafdcbbf),
	.w3(32'hbbf614d0),
	.w4(32'hbbfc2c5c),
	.w5(32'hba7eeac5),
	.w6(32'hbad9d2d2),
	.w7(32'h39932759),
	.w8(32'hbb029b8d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0db258),
	.w1(32'hbc291012),
	.w2(32'h3ba2fa38),
	.w3(32'hbc71bcf0),
	.w4(32'hbc57a91d),
	.w5(32'h3b313e12),
	.w6(32'hbc413124),
	.w7(32'hbbd25460),
	.w8(32'hbaceb259),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ebc76),
	.w1(32'h3c3a01f5),
	.w2(32'h3a9bad7d),
	.w3(32'h3c1a367f),
	.w4(32'hbac1409d),
	.w5(32'h3b67cea8),
	.w6(32'hbb1cc9e6),
	.w7(32'hbb8b25b2),
	.w8(32'h3c0dc89a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87c310),
	.w1(32'hbbde2a3a),
	.w2(32'hbb6aee8b),
	.w3(32'h3bbec6b0),
	.w4(32'hbbcd7338),
	.w5(32'hbb72deda),
	.w6(32'h3c8f88fb),
	.w7(32'h3bb8cfee),
	.w8(32'hbb7f3ea3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a6bde),
	.w1(32'h3b5f634d),
	.w2(32'hbbbcd2d1),
	.w3(32'h3bd367d7),
	.w4(32'h3bbf2db0),
	.w5(32'hbbd840d1),
	.w6(32'h3afddc3c),
	.w7(32'h3b8a6018),
	.w8(32'hbac9224f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa605f9),
	.w1(32'h3c2dd946),
	.w2(32'hbb017de5),
	.w3(32'h3b6413b8),
	.w4(32'h3c9dcf5a),
	.w5(32'hb9938dbd),
	.w6(32'h3c48ecd5),
	.w7(32'h3cb649b4),
	.w8(32'h3b56ecce),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba39774),
	.w1(32'hb8b790cc),
	.w2(32'hbb9b738b),
	.w3(32'hb92f4041),
	.w4(32'hbb714503),
	.w5(32'h3a471daf),
	.w6(32'h3b4ce8a3),
	.w7(32'hbb4dbca3),
	.w8(32'h3b07e090),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba69ce2),
	.w1(32'h3bd995d5),
	.w2(32'hbb8cd44c),
	.w3(32'hbc1a164c),
	.w4(32'hbb69f81a),
	.w5(32'hbbad07a3),
	.w6(32'hbbf4d75f),
	.w7(32'hbb6f2086),
	.w8(32'hbb972055),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f7f7b),
	.w1(32'hbbd2ebaa),
	.w2(32'h3ace4e4d),
	.w3(32'h3aa52954),
	.w4(32'hbbe18ea0),
	.w5(32'hbb32e1fe),
	.w6(32'h3a8b48a6),
	.w7(32'hbbade0ab),
	.w8(32'hbc32ebe1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ea2c5),
	.w1(32'hbc290878),
	.w2(32'h3aa4b276),
	.w3(32'hbb5b5d8b),
	.w4(32'hbc076e44),
	.w5(32'hba862c93),
	.w6(32'hbc1e2e02),
	.w7(32'hbc1872bc),
	.w8(32'h3b8e94d9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd66e16),
	.w1(32'h3c8bab8e),
	.w2(32'h3b669d0d),
	.w3(32'h3b5549e9),
	.w4(32'h3c3f9748),
	.w5(32'h3c5a2d84),
	.w6(32'h3c5ad931),
	.w7(32'h3c728e0b),
	.w8(32'h3c3307f7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf2613),
	.w1(32'hbb0d00ee),
	.w2(32'hbba1bf21),
	.w3(32'h3ce0effe),
	.w4(32'h3c4c73ba),
	.w5(32'hbbdc485c),
	.w6(32'h3c84da1e),
	.w7(32'h3b4c1ef8),
	.w8(32'hbc07e66c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6c169),
	.w1(32'hba81debf),
	.w2(32'hbc01a26e),
	.w3(32'hbb84e8d6),
	.w4(32'hbc634a55),
	.w5(32'h3bc127ad),
	.w6(32'hbc4a7878),
	.w7(32'hbc4eb42b),
	.w8(32'hb80739df),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb20fbb),
	.w1(32'h3b02cf24),
	.w2(32'hbb0b6b2c),
	.w3(32'h3c43d06f),
	.w4(32'h3bb3fa11),
	.w5(32'h3bc0e53b),
	.w6(32'h3bedf7e0),
	.w7(32'h3b813022),
	.w8(32'hbb5b12dd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabbbd6),
	.w1(32'hbb1925e4),
	.w2(32'h3a3a5be0),
	.w3(32'h3bb52a22),
	.w4(32'h3b9b3327),
	.w5(32'h39a7da50),
	.w6(32'h3b6ef80f),
	.w7(32'h39283808),
	.w8(32'h3a068702),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9fcf6),
	.w1(32'h3a9c8a82),
	.w2(32'h3a99c5db),
	.w3(32'hbb3a05f5),
	.w4(32'hbb0e4772),
	.w5(32'hb9013bb3),
	.w6(32'hbbdd8516),
	.w7(32'hbb319554),
	.w8(32'h3b23906f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35f66a),
	.w1(32'h3b292db5),
	.w2(32'h3a463a92),
	.w3(32'hba92e4a8),
	.w4(32'h3b0f6286),
	.w5(32'h3a0cdf92),
	.w6(32'h3aa3e840),
	.w7(32'h3a9c3c1e),
	.w8(32'hb9f32ee6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9858c56),
	.w1(32'h3b0c53cd),
	.w2(32'hbaa7b4e0),
	.w3(32'h3a7e9aa9),
	.w4(32'hbbb7ebcb),
	.w5(32'hba6dcc5e),
	.w6(32'h3b5115eb),
	.w7(32'hbc1bf6c5),
	.w8(32'hbb434258),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20480c),
	.w1(32'hbae3df33),
	.w2(32'hbb24d127),
	.w3(32'hba178111),
	.w4(32'hbb9208c6),
	.w5(32'hbb8b0716),
	.w6(32'hbb345168),
	.w7(32'hbbcbd612),
	.w8(32'hbb7358e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907cbae),
	.w1(32'h3b7cb0bf),
	.w2(32'hbb32d039),
	.w3(32'h3b3d0fde),
	.w4(32'h39c6c039),
	.w5(32'hba0747c9),
	.w6(32'h3ac7e2c9),
	.w7(32'h3ba2f742),
	.w8(32'h3abda0b3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23a0ca),
	.w1(32'h39777f8c),
	.w2(32'h3b38b533),
	.w3(32'h3a9b4be5),
	.w4(32'hba0492fe),
	.w5(32'h3b000006),
	.w6(32'h3af5a97d),
	.w7(32'hbbc67754),
	.w8(32'h3ac7e3c4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e1c44),
	.w1(32'h3ad69267),
	.w2(32'h3babbf9f),
	.w3(32'h3b680375),
	.w4(32'h3a64c1f0),
	.w5(32'h3b705eb6),
	.w6(32'h3b5dffd0),
	.w7(32'h3a3d0f46),
	.w8(32'h3b48e8c5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b972139),
	.w1(32'hbae6a662),
	.w2(32'hba9e5dd4),
	.w3(32'hb88243db),
	.w4(32'hbc15b976),
	.w5(32'hbaec2a6c),
	.w6(32'hbbdbffa9),
	.w7(32'hbc354632),
	.w8(32'hbaa62881),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab27fb5),
	.w1(32'hba399520),
	.w2(32'hbaaff17b),
	.w3(32'hbaf1ff04),
	.w4(32'h3a95e11a),
	.w5(32'hbbb12aae),
	.w6(32'hba2ec945),
	.w7(32'h3b2e554e),
	.w8(32'hbaa10ab9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fcf45),
	.w1(32'h3aa1e9bd),
	.w2(32'hbb8b199a),
	.w3(32'hbc086afa),
	.w4(32'hbb928161),
	.w5(32'hbb2a9532),
	.w6(32'h38f2522f),
	.w7(32'h3803d6f7),
	.w8(32'h3b1d67af),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c61a8),
	.w1(32'hbb3727ab),
	.w2(32'hbb4c8b39),
	.w3(32'hbb397308),
	.w4(32'hbc792212),
	.w5(32'hbc185ad5),
	.w6(32'hbc041cc8),
	.w7(32'hbc47f746),
	.w8(32'hbbffd27c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0856f),
	.w1(32'hbbda05ac),
	.w2(32'hbc0e8a35),
	.w3(32'hbbf4ab77),
	.w4(32'hbc132a44),
	.w5(32'hbbb495f0),
	.w6(32'hbc77d9dc),
	.w7(32'hbc107219),
	.w8(32'hbab9ebf2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf0c2b),
	.w1(32'hba141940),
	.w2(32'hba8f928f),
	.w3(32'hbb9f8e64),
	.w4(32'h3bac2146),
	.w5(32'hbb198db7),
	.w6(32'h3a63bdcd),
	.w7(32'h3c287e49),
	.w8(32'hbb1b1032),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b482a),
	.w1(32'hb96e7f0d),
	.w2(32'h3b033bb8),
	.w3(32'h3b2964d2),
	.w4(32'h3ad5e63e),
	.w5(32'hbb135dc7),
	.w6(32'h3ae8d2ab),
	.w7(32'hbab4f944),
	.w8(32'hbac37bc3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5be70),
	.w1(32'hb9d48457),
	.w2(32'h3b317206),
	.w3(32'hba843d0d),
	.w4(32'h3aad78b6),
	.w5(32'h3c271a1b),
	.w6(32'hba0dea6f),
	.w7(32'h39d844c5),
	.w8(32'h3bce9861),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afcba2),
	.w1(32'h3a781d03),
	.w2(32'hbb1b501c),
	.w3(32'h3ab00cb2),
	.w4(32'hbb84c182),
	.w5(32'hbb189662),
	.w6(32'h3b73f37a),
	.w7(32'hbb9cc620),
	.w8(32'hbafef772),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5be2d),
	.w1(32'h3b8f32aa),
	.w2(32'hbaf6a3da),
	.w3(32'h3bced899),
	.w4(32'hb92c3c37),
	.w5(32'hbb2967d9),
	.w6(32'h3b049e22),
	.w7(32'hbb4b4319),
	.w8(32'h3b786ab0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf7160),
	.w1(32'h3bf13ba8),
	.w2(32'h3baf7446),
	.w3(32'h3bc66f35),
	.w4(32'h3bd90273),
	.w5(32'h3ba79fa9),
	.w6(32'h3c0e332d),
	.w7(32'h3b41c46a),
	.w8(32'h3a1ed5a2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0dafb),
	.w1(32'h3c35dd56),
	.w2(32'hbba70966),
	.w3(32'h3c76aaf7),
	.w4(32'h3c520f24),
	.w5(32'hbb411926),
	.w6(32'h3c01b88b),
	.w7(32'h3abbdccf),
	.w8(32'hbb7d18ba),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b990f46),
	.w1(32'hbac6482e),
	.w2(32'h3ba1f730),
	.w3(32'hbb2af509),
	.w4(32'hbb4266a1),
	.w5(32'h3bdd2494),
	.w6(32'hb9427669),
	.w7(32'hbadc8554),
	.w8(32'h3bcf513d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9795c3),
	.w1(32'hba01a42f),
	.w2(32'h3c297ae8),
	.w3(32'h3b03d4a2),
	.w4(32'h3b146f62),
	.w5(32'h3b994671),
	.w6(32'h3bb20630),
	.w7(32'h3c09d733),
	.w8(32'h3bb65f1f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3ae1f),
	.w1(32'hb87fa787),
	.w2(32'hbafda152),
	.w3(32'h39651386),
	.w4(32'hba35da24),
	.w5(32'hbafc2504),
	.w6(32'hba85d310),
	.w7(32'hba869525),
	.w8(32'h370e00f2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab54a8b),
	.w1(32'hbaa6eafa),
	.w2(32'hba02e4a6),
	.w3(32'hbb1251bc),
	.w4(32'h3b963f22),
	.w5(32'h3bb736ae),
	.w6(32'h3809ab21),
	.w7(32'h3bdbbb63),
	.w8(32'h3bd81a6a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac205f0),
	.w1(32'hbbda59cb),
	.w2(32'hb9b3d6ef),
	.w3(32'hbbaf0761),
	.w4(32'hbb5cfda4),
	.w5(32'h3ac398ff),
	.w6(32'hba20c9b6),
	.w7(32'h3baeacfb),
	.w8(32'h3a967b85),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94b403),
	.w1(32'h3c0ea8a3),
	.w2(32'h3ac3603b),
	.w3(32'h3c0759dd),
	.w4(32'h3c525458),
	.w5(32'hba8d12c3),
	.w6(32'h3c1de7b9),
	.w7(32'h3bdd7488),
	.w8(32'h3ba752ac),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ae8c),
	.w1(32'hbaa2ffe2),
	.w2(32'h3b3963af),
	.w3(32'hbba1cf74),
	.w4(32'hbb4b832c),
	.w5(32'h39ca6d39),
	.w6(32'h3b397f15),
	.w7(32'h3c4c666f),
	.w8(32'h3b74ea3e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb80227),
	.w1(32'h3bd10158),
	.w2(32'h3b888a18),
	.w3(32'h3be73623),
	.w4(32'h3bc0a42c),
	.w5(32'hbad5fdc2),
	.w6(32'h3c25637d),
	.w7(32'h3c07face),
	.w8(32'hb9d82f77),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe11103),
	.w1(32'h3b130d8d),
	.w2(32'hb8a36b4e),
	.w3(32'hba81b835),
	.w4(32'h3becd440),
	.w5(32'hbaf88eca),
	.w6(32'h3aed3ee4),
	.w7(32'h3bff585a),
	.w8(32'hba82b12a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933cfce),
	.w1(32'h3b7ecc45),
	.w2(32'hba06775d),
	.w3(32'hbb77e432),
	.w4(32'h3a9ce239),
	.w5(32'hbb6b8b23),
	.w6(32'h3b635bd0),
	.w7(32'h3b8507b6),
	.w8(32'hbaffdb6f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae337d),
	.w1(32'hbaf6a116),
	.w2(32'hb9cc3384),
	.w3(32'h391f56e6),
	.w4(32'h39ef8dd1),
	.w5(32'h3a1b05b7),
	.w6(32'h3a60d333),
	.w7(32'h3b5cdccb),
	.w8(32'h3a95d5d6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388cd1ed),
	.w1(32'hba09db52),
	.w2(32'hba9b2dce),
	.w3(32'h3b91a74c),
	.w4(32'h3b1d0265),
	.w5(32'hbaba7e72),
	.w6(32'h3b6a650b),
	.w7(32'hb9826b3f),
	.w8(32'h3b6c8e88),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c92c5),
	.w1(32'hba56dab5),
	.w2(32'hb8e50c0f),
	.w3(32'hbb60954b),
	.w4(32'h3a0bf9f6),
	.w5(32'h38dc8dae),
	.w6(32'h3a9ab144),
	.w7(32'h3bb736de),
	.w8(32'hbb02de5e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fb83f),
	.w1(32'h3ae144b2),
	.w2(32'hbaec4be2),
	.w3(32'h3ae848ea),
	.w4(32'h3b532a4b),
	.w5(32'hba0d1dc0),
	.w6(32'h3a7ff0e8),
	.w7(32'hba60d4aa),
	.w8(32'h3b08cf73),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1cdd4),
	.w1(32'h3a2d22ba),
	.w2(32'h3be5a504),
	.w3(32'hb98563c0),
	.w4(32'h3bbf1178),
	.w5(32'h3bb464ee),
	.w6(32'h3b523970),
	.w7(32'h3c05da99),
	.w8(32'h3bc43ccc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986d8c),
	.w1(32'h3afc42c4),
	.w2(32'h3beb5a79),
	.w3(32'h3c1c0ce4),
	.w4(32'h386dcc48),
	.w5(32'h3bb0d8ee),
	.w6(32'h3b3b5cbb),
	.w7(32'h38a28b52),
	.w8(32'hba8a162e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15a6f9),
	.w1(32'h38f4c34d),
	.w2(32'hb9d1ba4c),
	.w3(32'hbbfc938a),
	.w4(32'hbc2cb1eb),
	.w5(32'hbb042f6c),
	.w6(32'hbc41890e),
	.w7(32'hbc394f51),
	.w8(32'hbb4a4c45),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50db49),
	.w1(32'h3aa7e11a),
	.w2(32'hbb39de48),
	.w3(32'hbb613347),
	.w4(32'hb88d3c59),
	.w5(32'hbc0888f4),
	.w6(32'hbb7e3cf4),
	.w7(32'hbb1bb61d),
	.w8(32'hbc19ba8e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb555dbf),
	.w1(32'hbacd64e1),
	.w2(32'hba81bd00),
	.w3(32'hb98afd79),
	.w4(32'h3a252989),
	.w5(32'hbabd7a4f),
	.w6(32'hbb7f5fec),
	.w7(32'h3b4c7fed),
	.w8(32'hbac87cf7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9831184),
	.w1(32'h3a6f7c17),
	.w2(32'h3aa62760),
	.w3(32'hb9a79a62),
	.w4(32'h3afd80c6),
	.w5(32'h3a43a9a6),
	.w6(32'h394bee0a),
	.w7(32'h3b2c9e34),
	.w8(32'h3a8e5299),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7c69f),
	.w1(32'hb9a1723a),
	.w2(32'hbc036089),
	.w3(32'h3a3658b3),
	.w4(32'hbb29bab9),
	.w5(32'hbc0359e6),
	.w6(32'h3a0ba880),
	.w7(32'h39f604ad),
	.w8(32'hbb3d8547),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb752c06),
	.w1(32'hbc04316a),
	.w2(32'hbc0d0a28),
	.w3(32'hbbd88ea4),
	.w4(32'h3b316c9f),
	.w5(32'hba8e1650),
	.w6(32'h39bb412e),
	.w7(32'h3bc9c5db),
	.w8(32'h3ada6ebe),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb250730),
	.w1(32'h3ab2fb20),
	.w2(32'h3af64ea3),
	.w3(32'hbad350a1),
	.w4(32'h3b6c78df),
	.w5(32'h3a9f7d85),
	.w6(32'h3bdfad7c),
	.w7(32'h3c42f54f),
	.w8(32'h3b4d865d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b315797),
	.w1(32'h3adb3305),
	.w2(32'h3a0e3588),
	.w3(32'hbad6b767),
	.w4(32'hbbcb69bd),
	.w5(32'h399c1d44),
	.w6(32'hbb74220c),
	.w7(32'hbbccc22d),
	.w8(32'hbb163ae2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33934a),
	.w1(32'hbac4b317),
	.w2(32'h3a7e3f42),
	.w3(32'hbb853c8d),
	.w4(32'hbab9b616),
	.w5(32'h3add6256),
	.w6(32'hbb7dd174),
	.w7(32'hbaf8f3c4),
	.w8(32'hb981ef4b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03dea0),
	.w1(32'hbb9ae68d),
	.w2(32'hbb508e40),
	.w3(32'h3af79738),
	.w4(32'hbab89293),
	.w5(32'hbba24369),
	.w6(32'h3b06dd4b),
	.w7(32'h3b009ab6),
	.w8(32'hbb903769),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab196d),
	.w1(32'hbb89dfa1),
	.w2(32'h3b2a4329),
	.w3(32'hbafe4517),
	.w4(32'h3b2dd67c),
	.w5(32'h3c054b3f),
	.w6(32'hbb68180b),
	.w7(32'h3aff277b),
	.w8(32'h3c027d3c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e9a44),
	.w1(32'hbb543ba9),
	.w2(32'h3a9c3e7f),
	.w3(32'h3c15097a),
	.w4(32'hbbc88f4d),
	.w5(32'h3aa471ac),
	.w6(32'h3a298af0),
	.w7(32'hbc3c8f57),
	.w8(32'h3b38e55a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a327d),
	.w1(32'h3a173341),
	.w2(32'h3ae56cec),
	.w3(32'h396e107b),
	.w4(32'hba014f8a),
	.w5(32'h3a0df639),
	.w6(32'hba501500),
	.w7(32'hba1ff6f3),
	.w8(32'hb9802171),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12791f),
	.w1(32'h3b45cbe5),
	.w2(32'h39e1d4a1),
	.w3(32'h3ae24043),
	.w4(32'h3acf3dfb),
	.w5(32'hbbfc6983),
	.w6(32'h3ac80392),
	.w7(32'h3b747194),
	.w8(32'h389e3c5c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb04ae6),
	.w1(32'h3aec3f75),
	.w2(32'hba528013),
	.w3(32'hbc1ae557),
	.w4(32'h3bbc09a9),
	.w5(32'hbb9c7cef),
	.w6(32'hbb90aadd),
	.w7(32'h3c4e1130),
	.w8(32'hbb417a38),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb928b8a),
	.w1(32'hbb47bc74),
	.w2(32'hbbb2fd93),
	.w3(32'hbbd32269),
	.w4(32'hbb3e94ea),
	.w5(32'hbb2607fb),
	.w6(32'hbc0a8127),
	.w7(32'hba12aa25),
	.w8(32'h39301129),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ceb41),
	.w1(32'hbaca4e11),
	.w2(32'h3b79dd30),
	.w3(32'h3b059312),
	.w4(32'hba805d04),
	.w5(32'h3b0da310),
	.w6(32'h3b8e879b),
	.w7(32'h3b5c7e71),
	.w8(32'h3b43d807),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc2691),
	.w1(32'h3a754844),
	.w2(32'hba32adbc),
	.w3(32'h39a8e17e),
	.w4(32'hb790017a),
	.w5(32'h392ef5b3),
	.w6(32'hba494ab7),
	.w7(32'h3a84abcc),
	.w8(32'h3ae03972),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5eed5e),
	.w1(32'h3aa8e84b),
	.w2(32'h3b4310fe),
	.w3(32'h3b11def3),
	.w4(32'hb9856bcd),
	.w5(32'h3aab80c1),
	.w6(32'h3b8728b9),
	.w7(32'h3b22770b),
	.w8(32'h3aa1ac48),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba066da9),
	.w1(32'h3a389ce3),
	.w2(32'h3bc0c174),
	.w3(32'hb9f2149a),
	.w4(32'hba1e2d22),
	.w5(32'h3ae1a005),
	.w6(32'h37a149d2),
	.w7(32'hba9cf2ad),
	.w8(32'hba304222),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab27088),
	.w1(32'hb88b65b1),
	.w2(32'hbb76e81a),
	.w3(32'hbb9c10b9),
	.w4(32'h3b1868b3),
	.w5(32'h3a92d71b),
	.w6(32'hbabfa54c),
	.w7(32'hba9101de),
	.w8(32'hbb9077cd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92b9dd),
	.w1(32'hbb809209),
	.w2(32'h3b472940),
	.w3(32'h3b057127),
	.w4(32'hbb9a8804),
	.w5(32'hbb65daf8),
	.w6(32'hbb92b1de),
	.w7(32'h3b199dd0),
	.w8(32'hbbae6bae),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e5938),
	.w1(32'h3b6bf0ae),
	.w2(32'hbaba86b1),
	.w3(32'hbb6cb416),
	.w4(32'h3a8cc05a),
	.w5(32'h3b3e38f9),
	.w6(32'hbb49408f),
	.w7(32'hba66cda5),
	.w8(32'h3bc57170),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b6b8a),
	.w1(32'h3b0a93c7),
	.w2(32'h39f72345),
	.w3(32'h3be6e0fc),
	.w4(32'h3c08a8bd),
	.w5(32'hb871fc01),
	.w6(32'h3c34c6b2),
	.w7(32'h3bd0af26),
	.w8(32'h3806e063),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5d884),
	.w1(32'h3b0471ae),
	.w2(32'h3a2d5175),
	.w3(32'hb7a5e6e2),
	.w4(32'h3afff848),
	.w5(32'hbae16de2),
	.w6(32'h3a656914),
	.w7(32'h3b9e8cbf),
	.w8(32'hb9a7be2f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e59882),
	.w1(32'hba503a7f),
	.w2(32'hbb87b460),
	.w3(32'h3a6782ab),
	.w4(32'hba81557b),
	.w5(32'h3af8e0a5),
	.w6(32'h3a0b4d67),
	.w7(32'hbaf97c49),
	.w8(32'h3ba2a730),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9086fe),
	.w1(32'hba6e6ee3),
	.w2(32'h3b8e06a2),
	.w3(32'hbb242ce1),
	.w4(32'h3a002f40),
	.w5(32'hba2c1f00),
	.w6(32'h3b953fd1),
	.w7(32'h3b0bc9d6),
	.w8(32'hbb869714),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca5ba7),
	.w1(32'h3bd45b91),
	.w2(32'h3bffba1e),
	.w3(32'hb8d28a8a),
	.w4(32'h3ae90c7c),
	.w5(32'h3b82fa5b),
	.w6(32'h3ba0eb2d),
	.w7(32'h3b8db371),
	.w8(32'h3bdb8c7c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfc7b1),
	.w1(32'h3b890dc3),
	.w2(32'hbae7c296),
	.w3(32'hbb72fa4e),
	.w4(32'hba584561),
	.w5(32'hbb094ba6),
	.w6(32'hbb473fa0),
	.w7(32'h3b208899),
	.w8(32'h3a6dc5c1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae38211),
	.w1(32'h3ace6c99),
	.w2(32'h3b8de5bc),
	.w3(32'hbbdfe59c),
	.w4(32'h3b3c0cc9),
	.w5(32'h3a6a8c9b),
	.w6(32'hbb11e1df),
	.w7(32'h3c19ea98),
	.w8(32'h39d2b0a3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac805ae),
	.w1(32'h39cc54cd),
	.w2(32'hb9dbd593),
	.w3(32'hb731eff3),
	.w4(32'hba90243a),
	.w5(32'h38fd4cac),
	.w6(32'hba8430c6),
	.w7(32'hbb3d516f),
	.w8(32'hb9bc2ad2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0af55d),
	.w1(32'h3c137f8d),
	.w2(32'h3b93ca6a),
	.w3(32'h3bf97061),
	.w4(32'h3bad403b),
	.w5(32'hbaff6edd),
	.w6(32'h3bd7a8f5),
	.w7(32'h3bc39a58),
	.w8(32'h3b40b1d1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7a6b5),
	.w1(32'hbb55ff0e),
	.w2(32'hbadc7864),
	.w3(32'hbbce5f32),
	.w4(32'hbb945f51),
	.w5(32'h3a939094),
	.w6(32'hb9dcb372),
	.w7(32'h3b9d4484),
	.w8(32'h3b1f8f7c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabdcde),
	.w1(32'hb9d1787c),
	.w2(32'hbb85e197),
	.w3(32'h3b8b143f),
	.w4(32'h3c18c9d9),
	.w5(32'hbb2ca60a),
	.w6(32'h3b010911),
	.w7(32'hb92ab96c),
	.w8(32'hbb7d32ca),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920957),
	.w1(32'hbaab1c2d),
	.w2(32'h3c225985),
	.w3(32'hbadb07fb),
	.w4(32'hb8804900),
	.w5(32'h3c1e7a9a),
	.w6(32'hbbda0440),
	.w7(32'h3ab2ea16),
	.w8(32'h3b8b390c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9e854),
	.w1(32'h3b10abfa),
	.w2(32'hba3c18f4),
	.w3(32'hbb6eeb37),
	.w4(32'hba18f491),
	.w5(32'h3b971490),
	.w6(32'hbb74a1f8),
	.w7(32'hbbc6ccec),
	.w8(32'h3bc2cf93),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58b380),
	.w1(32'hbb2a4b17),
	.w2(32'hbbd139bb),
	.w3(32'hbbbf2261),
	.w4(32'hbbdd1baa),
	.w5(32'h39c27602),
	.w6(32'hbb2b415f),
	.w7(32'h3b261707),
	.w8(32'h3c29a1b6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6082b2),
	.w1(32'h3c0b530d),
	.w2(32'h3953e497),
	.w3(32'hb9c30af8),
	.w4(32'h3c3fa609),
	.w5(32'h3938b365),
	.w6(32'h3bcd988b),
	.w7(32'h3c7dd38f),
	.w8(32'h3bd787e6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93318c),
	.w1(32'h3bbb33c8),
	.w2(32'hbb073b68),
	.w3(32'h3c388271),
	.w4(32'hbba3d080),
	.w5(32'hbc6cdff3),
	.w6(32'h3ae101bf),
	.w7(32'hbc50f597),
	.w8(32'hbc2a5bcb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1f174),
	.w1(32'hbae41ef7),
	.w2(32'h3b2979f8),
	.w3(32'hb98caf39),
	.w4(32'h3ad5bedd),
	.w5(32'h3baa5c20),
	.w6(32'h3bf40dfc),
	.w7(32'h3b9f240d),
	.w8(32'h3aa119c8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b20dd),
	.w1(32'h3a7e0195),
	.w2(32'h3ac99189),
	.w3(32'hbb000e8b),
	.w4(32'hbb2a7957),
	.w5(32'h39fc9156),
	.w6(32'hbb4a0823),
	.w7(32'hbb0c6376),
	.w8(32'h3ad032ac),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4cde4),
	.w1(32'hbbd01f7f),
	.w2(32'hbbce4577),
	.w3(32'hbba36a19),
	.w4(32'hbb8b0659),
	.w5(32'hbc0a9a81),
	.w6(32'hbb8fcf3c),
	.w7(32'hbbef1207),
	.w8(32'hbabebe75),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba190dc),
	.w1(32'h3c18d2df),
	.w2(32'h3c594c8b),
	.w3(32'h3bbefa20),
	.w4(32'h3c4966c9),
	.w5(32'h3bebb04e),
	.w6(32'h3c06535d),
	.w7(32'h3ca5f619),
	.w8(32'h3c3910c5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f24aa),
	.w1(32'hbb4882f8),
	.w2(32'h3a452fbb),
	.w3(32'hbb39c30d),
	.w4(32'hba8f60a5),
	.w5(32'h3ae5e8c7),
	.w6(32'hbb331e33),
	.w7(32'hbbb06a31),
	.w8(32'h393497e9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb755bee),
	.w1(32'hbb3db1b2),
	.w2(32'hbaf3e44a),
	.w3(32'hbb5ff0d3),
	.w4(32'h3a079aae),
	.w5(32'hb8539733),
	.w6(32'hbb0f724c),
	.w7(32'h3906cae3),
	.w8(32'hbb0d01a2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe275c),
	.w1(32'hbb5dfb7d),
	.w2(32'h3b6fd0da),
	.w3(32'h3aa73852),
	.w4(32'hbb5415cf),
	.w5(32'hbb51630d),
	.w6(32'h3aab623a),
	.w7(32'h3a6daad4),
	.w8(32'hbb73551d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dd2bb),
	.w1(32'hbb41d345),
	.w2(32'hbbfffa5d),
	.w3(32'hbba412e2),
	.w4(32'hbb8d8eee),
	.w5(32'hbb28fb08),
	.w6(32'hbbbb1ef3),
	.w7(32'hbc158fd0),
	.w8(32'hba802f42),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adda2d7),
	.w1(32'hbb42add3),
	.w2(32'h3c142aee),
	.w3(32'h3b6e595e),
	.w4(32'hbb2263ab),
	.w5(32'h3c74d8ca),
	.w6(32'h3b165271),
	.w7(32'hbb7824eb),
	.w8(32'h3bcfef3a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49312a),
	.w1(32'h3bd3b718),
	.w2(32'h3b52d9ab),
	.w3(32'h3bb48920),
	.w4(32'hbb4483f2),
	.w5(32'h3bc0f4c4),
	.w6(32'hbc210c62),
	.w7(32'hbc0c9def),
	.w8(32'h3b9e17fa),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b984c4b),
	.w1(32'hbbba943a),
	.w2(32'h3b519eb4),
	.w3(32'h3b63e471),
	.w4(32'hbb265628),
	.w5(32'h3bd00541),
	.w6(32'h3a65e8e3),
	.w7(32'hbb49851e),
	.w8(32'h3b5a9d65),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b449b46),
	.w1(32'hbb564123),
	.w2(32'hbb02a43d),
	.w3(32'h3b66a088),
	.w4(32'hbbca1227),
	.w5(32'h39767103),
	.w6(32'hbae3c448),
	.w7(32'hbc2e0ff6),
	.w8(32'h3af0dd31),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a939983),
	.w1(32'hb9ebb0df),
	.w2(32'h3a620629),
	.w3(32'h3c213f96),
	.w4(32'h38a41737),
	.w5(32'hba90e907),
	.w6(32'h3c262e37),
	.w7(32'h3b96bb60),
	.w8(32'h3a1616c5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9240e44),
	.w1(32'h3b0ed4d9),
	.w2(32'h3a5c2c3a),
	.w3(32'hbb473944),
	.w4(32'hbb6f4b36),
	.w5(32'hba728921),
	.w6(32'hbac40cb0),
	.w7(32'hbb7acb2d),
	.w8(32'h399e9ab0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa59416),
	.w1(32'h3ab509ad),
	.w2(32'h3b2f3b79),
	.w3(32'h39f84fb6),
	.w4(32'h3ab725e6),
	.w5(32'hba9a9900),
	.w6(32'h3b06a3cf),
	.w7(32'h3b345d58),
	.w8(32'hba8c49e2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85b4e2),
	.w1(32'hbac7e779),
	.w2(32'h3b32b504),
	.w3(32'hba421bbd),
	.w4(32'hbafc1194),
	.w5(32'h3aa4185c),
	.w6(32'h3a99bbfc),
	.w7(32'h3b7e1811),
	.w8(32'h3bde0ead),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c4f25),
	.w1(32'h3b387114),
	.w2(32'hbb101965),
	.w3(32'h3a5427d4),
	.w4(32'h3a87c0e7),
	.w5(32'hbbe9265e),
	.w6(32'h3bea66dc),
	.w7(32'h3b93aab6),
	.w8(32'hbb15088f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb725211),
	.w1(32'h3aad3c5c),
	.w2(32'hbb8a70ad),
	.w3(32'hbb4f8790),
	.w4(32'hba67442e),
	.w5(32'hbbac80f0),
	.w6(32'hbb8e18b4),
	.w7(32'h39e5b432),
	.w8(32'h3ae0c8cc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbe5da),
	.w1(32'h3a0e3e6c),
	.w2(32'h3b01eed3),
	.w3(32'hbaed5c23),
	.w4(32'hbb3f2047),
	.w5(32'h3b962664),
	.w6(32'h3b9f1102),
	.w7(32'hbb3af736),
	.w8(32'hb90e91e2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8ff57),
	.w1(32'h3b99a91f),
	.w2(32'h3ab424ea),
	.w3(32'hbb515725),
	.w4(32'hbba85824),
	.w5(32'h3998783c),
	.w6(32'hbbe6d14b),
	.w7(32'hbc2e7032),
	.w8(32'hba96741a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e6679),
	.w1(32'h3a035c54),
	.w2(32'h3a3569a9),
	.w3(32'h3a6b02cc),
	.w4(32'h38fac9fc),
	.w5(32'hba046ce7),
	.w6(32'h3a09c1df),
	.w7(32'hb9fe3e6e),
	.w8(32'h3a028a5c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a345059),
	.w1(32'hbac8a03d),
	.w2(32'h3b06333e),
	.w3(32'h3a05d3a1),
	.w4(32'hbb88aed0),
	.w5(32'hba3507d4),
	.w6(32'hbb157fb6),
	.w7(32'hbbb3337d),
	.w8(32'h3ad860a8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3638c6),
	.w1(32'hbc1beba0),
	.w2(32'h3adb1e3a),
	.w3(32'hbb31a966),
	.w4(32'hbc19516a),
	.w5(32'h38e67056),
	.w6(32'hbbbeb119),
	.w7(32'hbc1a5065),
	.w8(32'hba468f78),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92e193),
	.w1(32'hb9a6849b),
	.w2(32'h38844df9),
	.w3(32'hbaae1c48),
	.w4(32'hbb364efa),
	.w5(32'h3afc5ce7),
	.w6(32'hbb0d5324),
	.w7(32'hbb8d24c1),
	.w8(32'h3b921d3d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba30f6c),
	.w1(32'hbb1d7c18),
	.w2(32'hbbc496ee),
	.w3(32'hb91ed2c8),
	.w4(32'hbb6f5a47),
	.w5(32'hbb8bed2c),
	.w6(32'h3b1a994e),
	.w7(32'h3a0f8d95),
	.w8(32'hb927eec3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d3621),
	.w1(32'hbb359fcf),
	.w2(32'hbb2ebd08),
	.w3(32'hbb774b8d),
	.w4(32'hbb726009),
	.w5(32'hbbc77c38),
	.w6(32'h3b083452),
	.w7(32'h3b0c4edb),
	.w8(32'hba3ba6b9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0558da),
	.w1(32'hbbc0750e),
	.w2(32'hba495308),
	.w3(32'hbc0bbd43),
	.w4(32'h3b903b67),
	.w5(32'hba469414),
	.w6(32'h3b970481),
	.w7(32'h3ba5a692),
	.w8(32'h398c7608),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886db9),
	.w1(32'h3b945b51),
	.w2(32'h3be45af5),
	.w3(32'h3b1a49b9),
	.w4(32'h3c09e57c),
	.w5(32'h3a98f744),
	.w6(32'h3b49f0f1),
	.w7(32'h3c36265a),
	.w8(32'hbb2dc850),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dae6e),
	.w1(32'hbb3b0248),
	.w2(32'h3b36bfd4),
	.w3(32'hbb92e533),
	.w4(32'hbad4026f),
	.w5(32'h3b4376fa),
	.w6(32'hbb08758b),
	.w7(32'h3b205de3),
	.w8(32'h3ba9f0fd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b898fd9),
	.w1(32'h3b3fc71d),
	.w2(32'h3a37e787),
	.w3(32'h3c09a4d4),
	.w4(32'hbb9184b2),
	.w5(32'h3c03e020),
	.w6(32'hbb58534f),
	.w7(32'hbc1b9039),
	.w8(32'h3b97d734),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0e825),
	.w1(32'h3a3b5a29),
	.w2(32'hbb25643d),
	.w3(32'h3b4bdcef),
	.w4(32'hbba989d9),
	.w5(32'h3a4019a4),
	.w6(32'h3858e033),
	.w7(32'hbc0f47c6),
	.w8(32'hbb96ae2d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b204afb),
	.w1(32'h3bcbd8d9),
	.w2(32'hba0d8fa4),
	.w3(32'h3b1b71d9),
	.w4(32'h3c047ce9),
	.w5(32'hbae798e1),
	.w6(32'hba4ad073),
	.w7(32'h3b725c61),
	.w8(32'h3ace932e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba048b08),
	.w1(32'hb98dd3e3),
	.w2(32'h3b43d01b),
	.w3(32'h3a893eae),
	.w4(32'h3b2a616c),
	.w5(32'hba553184),
	.w6(32'h3c2bc432),
	.w7(32'h3b4c1e0d),
	.w8(32'h3a73de5b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9bfec),
	.w1(32'h3b933b23),
	.w2(32'h3b85222f),
	.w3(32'h3b179ada),
	.w4(32'h3b867121),
	.w5(32'h3918cb39),
	.w6(32'h3b986e13),
	.w7(32'h3baff722),
	.w8(32'h3b1ba3c7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961cc6e),
	.w1(32'h3a693347),
	.w2(32'h3a8e0194),
	.w3(32'hba0b52c8),
	.w4(32'hbab34786),
	.w5(32'h398f7ef7),
	.w6(32'h3b1f998a),
	.w7(32'hbb26dadf),
	.w8(32'hbb244792),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b834f84),
	.w1(32'hbaf4c2fa),
	.w2(32'h3b7ae248),
	.w3(32'h3b01921e),
	.w4(32'hb8afd8bc),
	.w5(32'h3ab44507),
	.w6(32'h3abfa60d),
	.w7(32'h3b749966),
	.w8(32'h3b8006b3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf14660),
	.w1(32'h3b9c8fef),
	.w2(32'h3b607cd7),
	.w3(32'hbaf66c3e),
	.w4(32'h3c2eec7b),
	.w5(32'h3a0c6a17),
	.w6(32'h3c13f152),
	.w7(32'h3c8cd218),
	.w8(32'h3b1da480),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903839e),
	.w1(32'hb8b3ca4c),
	.w2(32'hbb10a59c),
	.w3(32'hba340055),
	.w4(32'hbacb1b79),
	.w5(32'h3b55de0c),
	.w6(32'hb95f0316),
	.w7(32'hbb184992),
	.w8(32'h3bf2ae47),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73dd9c),
	.w1(32'h3af842f2),
	.w2(32'h39d6b446),
	.w3(32'h3b8dce5d),
	.w4(32'hbae7d6fa),
	.w5(32'hb94dcfc2),
	.w6(32'h3bffb56b),
	.w7(32'hba937293),
	.w8(32'h3925175f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c1497),
	.w1(32'h3ac561b2),
	.w2(32'h3bff022a),
	.w3(32'h3ad7e719),
	.w4(32'h3a8a1ec5),
	.w5(32'h3b7f4d7a),
	.w6(32'h3a822a65),
	.w7(32'h394e5290),
	.w8(32'h3bd779a9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba098b8),
	.w1(32'h3bd12d3f),
	.w2(32'hbb6b5938),
	.w3(32'h3bba3950),
	.w4(32'h3adb6ea8),
	.w5(32'hba90d2a7),
	.w6(32'h3b4b47f9),
	.w7(32'h38e6e8d3),
	.w8(32'hbb96cd9f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2dd06),
	.w1(32'h3b0686aa),
	.w2(32'h3ae452e1),
	.w3(32'h3b3085b6),
	.w4(32'h3c2ed872),
	.w5(32'h3aab638e),
	.w6(32'h3a1bc6ed),
	.w7(32'h3b89fb90),
	.w8(32'h3b879f46),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3262a2),
	.w1(32'h3a74227e),
	.w2(32'h3a8b238f),
	.w3(32'h3af83eda),
	.w4(32'h3a511aa0),
	.w5(32'h3a4f463b),
	.w6(32'h3bb0c9de),
	.w7(32'h3b816a7c),
	.w8(32'h3a8a70e9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13d293),
	.w1(32'h39e6ab0d),
	.w2(32'h3b98b08d),
	.w3(32'h395226d6),
	.w4(32'h366a978c),
	.w5(32'h3a7bfbd1),
	.w6(32'h39b6e05f),
	.w7(32'hba3aeb54),
	.w8(32'h3a1c3ccb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a698dc7),
	.w1(32'h3a6aa76b),
	.w2(32'h3b97f129),
	.w3(32'hbb1af8fb),
	.w4(32'hbb59a7a0),
	.w5(32'h3c1a5930),
	.w6(32'hbb9e8ec8),
	.w7(32'hbb908c20),
	.w8(32'h3b686afb),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdce1df),
	.w1(32'h3ba7501f),
	.w2(32'h3aea25c2),
	.w3(32'h3c116b97),
	.w4(32'h3af88842),
	.w5(32'h3b508880),
	.w6(32'h3b13af1e),
	.w7(32'hb95e15e8),
	.w8(32'h3ae64b4a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e4123),
	.w1(32'h394e2ec7),
	.w2(32'h3b3dcc38),
	.w3(32'h3a4524bc),
	.w4(32'hba076d8d),
	.w5(32'h3b47326e),
	.w6(32'hbb12f49d),
	.w7(32'hbb907ca6),
	.w8(32'h3b3bf0c1),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad13b2e),
	.w1(32'h3aa3c0b7),
	.w2(32'h3bef1595),
	.w3(32'hb91115e5),
	.w4(32'hb9c67d34),
	.w5(32'h3bebea91),
	.w6(32'h3b1d137f),
	.w7(32'h3971731a),
	.w8(32'hbab84e41),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e71c5),
	.w1(32'h3bb2fe88),
	.w2(32'h3b816b93),
	.w3(32'h3ba3f877),
	.w4(32'hbb185b45),
	.w5(32'h3b6d5411),
	.w6(32'hbbaa452f),
	.w7(32'hbbcc40fc),
	.w8(32'h3a2903fc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7a27c),
	.w1(32'hba8de991),
	.w2(32'h39665d1c),
	.w3(32'h3a54549b),
	.w4(32'hba75dc14),
	.w5(32'h3b61d651),
	.w6(32'hbaa89e5c),
	.w7(32'hbbe7ee77),
	.w8(32'h3bc013be),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394da480),
	.w1(32'h3a70f03f),
	.w2(32'h3be47f44),
	.w3(32'h399f6e41),
	.w4(32'h3a5e5290),
	.w5(32'h3bfeee7e),
	.w6(32'h3b2342c1),
	.w7(32'h3b965fbe),
	.w8(32'h3be722d3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55f3b6),
	.w1(32'h3b45b299),
	.w2(32'h3be379d9),
	.w3(32'h3bcabca7),
	.w4(32'hb9d164f0),
	.w5(32'h3b9edb49),
	.w6(32'h3baaa22f),
	.w7(32'h3b88552b),
	.w8(32'h3a159d43),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1318ff),
	.w1(32'hbbc9dc99),
	.w2(32'hbacedcba),
	.w3(32'hbb1ed9d4),
	.w4(32'hbbc1e531),
	.w5(32'hbb809ace),
	.w6(32'hbbe9a159),
	.w7(32'hbc1af3b9),
	.w8(32'hbb8a2ad7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e0c72),
	.w1(32'hbacb9496),
	.w2(32'hbb7ddd5d),
	.w3(32'hbbfdd7ee),
	.w4(32'hbb8244e2),
	.w5(32'hbbd28299),
	.w6(32'hbc108dd0),
	.w7(32'h3b183d21),
	.w8(32'hbb50779d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f16da),
	.w1(32'h3a972fff),
	.w2(32'h3a540c94),
	.w3(32'hb88a6e34),
	.w4(32'hba9b83c2),
	.w5(32'h3a1ed60e),
	.w6(32'h390ab27e),
	.w7(32'hbb1ef8a4),
	.w8(32'h3a27fe17),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eb120),
	.w1(32'h3b06883c),
	.w2(32'h39e071fd),
	.w3(32'h3b57c514),
	.w4(32'h3b571ef5),
	.w5(32'hbbe30112),
	.w6(32'hbaaee765),
	.w7(32'h3ab68c12),
	.w8(32'hbb23c7ff),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae06469),
	.w1(32'hbaaa5069),
	.w2(32'hba084ad8),
	.w3(32'hbb9c435d),
	.w4(32'hbb48f716),
	.w5(32'hbaa99a72),
	.w6(32'hbbb7b6fb),
	.w7(32'hbaf2f297),
	.w8(32'hba02f76a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9f857),
	.w1(32'h3b896de6),
	.w2(32'h3af6c060),
	.w3(32'hba690778),
	.w4(32'h3b236ad7),
	.w5(32'h3b116c74),
	.w6(32'h39b07e7a),
	.w7(32'h3b5139f4),
	.w8(32'hb9a567fc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25f507),
	.w1(32'hb9175941),
	.w2(32'h3ade2312),
	.w3(32'h3b40c9b5),
	.w4(32'h3b88dd09),
	.w5(32'hbadedcb7),
	.w6(32'hba8f643b),
	.w7(32'h3abb3cc4),
	.w8(32'h3a1e311f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a3e270),
	.w1(32'h3aeb1aa9),
	.w2(32'hbba9b2ec),
	.w3(32'h3b49f2be),
	.w4(32'h3a9b45b5),
	.w5(32'hbbe27aa9),
	.w6(32'h3b56f00f),
	.w7(32'h3a232580),
	.w8(32'hbba3a54a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1d0ab),
	.w1(32'hbb3172a1),
	.w2(32'h3b1d58ad),
	.w3(32'hbbd51d37),
	.w4(32'hbb805498),
	.w5(32'hba7869ff),
	.w6(32'hbbd635b8),
	.w7(32'hbb7ae4c3),
	.w8(32'hbb3987ff),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08531f),
	.w1(32'hbaa8c5b1),
	.w2(32'h39be3086),
	.w3(32'h3a2e3466),
	.w4(32'hbb6c95e6),
	.w5(32'h3a789172),
	.w6(32'h3a05535f),
	.w7(32'hbbb297b7),
	.w8(32'hba5ee364),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6977aa),
	.w1(32'hba557c72),
	.w2(32'h3adfea71),
	.w3(32'h3b062082),
	.w4(32'h398c4f59),
	.w5(32'h3aa9808f),
	.w6(32'h3ab077ee),
	.w7(32'h3a8b04aa),
	.w8(32'h3aa5d97d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22b0bf),
	.w1(32'hbc1ac325),
	.w2(32'hbb21fad0),
	.w3(32'hbc0db308),
	.w4(32'hbc163e4f),
	.w5(32'hbb09087c),
	.w6(32'hbbf3e5ed),
	.w7(32'hbbb44f2f),
	.w8(32'h3aa808e5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ea22),
	.w1(32'hba9fbb95),
	.w2(32'h394f80b9),
	.w3(32'hbba83f65),
	.w4(32'hbb38eae6),
	.w5(32'hb9232c6b),
	.w6(32'hbba0ba97),
	.w7(32'hbb37a71c),
	.w8(32'hba771ff9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d26d1),
	.w1(32'h3b81a2ff),
	.w2(32'hbbd6f9d9),
	.w3(32'hbb034417),
	.w4(32'h3a952d08),
	.w5(32'hbbd82ba5),
	.w6(32'hbb17dbf6),
	.w7(32'hb9213b67),
	.w8(32'hbb84ba34),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b598116),
	.w1(32'h3bc70c03),
	.w2(32'hba9ff2f0),
	.w3(32'h39e8fe43),
	.w4(32'hbb0a9e8b),
	.w5(32'hbb690289),
	.w6(32'h3acf22bb),
	.w7(32'hbb3805c1),
	.w8(32'hbb8e7a41),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac37f41),
	.w1(32'h3a712d95),
	.w2(32'hba1d24b4),
	.w3(32'h3b17b061),
	.w4(32'h3b76f76f),
	.w5(32'hbb6f3430),
	.w6(32'h3bd31f60),
	.w7(32'h3b9ff73c),
	.w8(32'h3b922691),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c1604),
	.w1(32'hbabaf8a9),
	.w2(32'hba8d4859),
	.w3(32'hbb9582ac),
	.w4(32'hbb33ebc8),
	.w5(32'hbab63647),
	.w6(32'hbb27493e),
	.w7(32'hbaaf187c),
	.w8(32'hba3ceaea),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b0b26),
	.w1(32'h3b9a229e),
	.w2(32'h3b664733),
	.w3(32'h3a94416f),
	.w4(32'hbad1e84c),
	.w5(32'h3b53272d),
	.w6(32'h3aa7a357),
	.w7(32'hbb295578),
	.w8(32'h3aa44cfa),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa18c7),
	.w1(32'h39b058a4),
	.w2(32'h3b526fca),
	.w3(32'h3b4a514d),
	.w4(32'h3ae0933c),
	.w5(32'h3a96e0b2),
	.w6(32'h3aa51102),
	.w7(32'h3aae2946),
	.w8(32'hba291429),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c036181),
	.w1(32'h3c5f1a37),
	.w2(32'hbb53a868),
	.w3(32'h3b47e942),
	.w4(32'h3c20c90f),
	.w5(32'hbc207528),
	.w6(32'h3b5dbf76),
	.w7(32'h3c4e1c89),
	.w8(32'hbbb3dce0),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea8e78),
	.w1(32'h3b8f0397),
	.w2(32'h3b84cbaa),
	.w3(32'hbb8b8991),
	.w4(32'h3ab9f3f3),
	.w5(32'hb7d0d328),
	.w6(32'hba74f33e),
	.w7(32'h3b5c6e6d),
	.w8(32'h3a431555),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b609ed1),
	.w1(32'h3b4c5751),
	.w2(32'h3b44fb48),
	.w3(32'hb95d7d90),
	.w4(32'hbb18df97),
	.w5(32'h3b06b988),
	.w6(32'h3b2b6930),
	.w7(32'hbb194269),
	.w8(32'h3b9660d2),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37a8be),
	.w1(32'h3b481b85),
	.w2(32'h3ad43383),
	.w3(32'h39c7fd9b),
	.w4(32'h3a3d2d1f),
	.w5(32'h3a1947f3),
	.w6(32'h3b153fa9),
	.w7(32'h3b8dfb40),
	.w8(32'hba2fbd67),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75ec62),
	.w1(32'h3ab6c406),
	.w2(32'hbb52d04d),
	.w3(32'h3bcea53a),
	.w4(32'h3b274b4d),
	.w5(32'hbb23fb12),
	.w6(32'h3bf1a5d8),
	.w7(32'h3b541c0b),
	.w8(32'h3a10d8e8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45edcf),
	.w1(32'hbab438cd),
	.w2(32'h3af54b94),
	.w3(32'hbb988a8f),
	.w4(32'h39a8cd73),
	.w5(32'h3a9ae7c8),
	.w6(32'hba85aa72),
	.w7(32'h3a57c2fa),
	.w8(32'h3ab1bbbd),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba378b44),
	.w1(32'hba6b9b60),
	.w2(32'hba61e262),
	.w3(32'hbb1269fc),
	.w4(32'hba2b318c),
	.w5(32'hbb626150),
	.w6(32'hbb1c433b),
	.w7(32'hba97e035),
	.w8(32'hbb6bc1b1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab78a74),
	.w1(32'h3b1084f1),
	.w2(32'hbab57e3f),
	.w3(32'hbb28306c),
	.w4(32'h3b983ea6),
	.w5(32'h3b4894de),
	.w6(32'h3a9a3683),
	.w7(32'h3c1f4284),
	.w8(32'hbb2a6fec),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbaf6b),
	.w1(32'hbb4cafa0),
	.w2(32'h3aa663f0),
	.w3(32'h3a5f6706),
	.w4(32'hbb81ce28),
	.w5(32'h3accbceb),
	.w6(32'hbab97e2f),
	.w7(32'hbb559103),
	.w8(32'h3a4b7b67),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa92652),
	.w1(32'hba82f14e),
	.w2(32'h3acdfd69),
	.w3(32'h3b0a4a89),
	.w4(32'h3a93d2e5),
	.w5(32'h399bd677),
	.w6(32'h3a85d12e),
	.w7(32'h3b0cd0dc),
	.w8(32'hbab124c2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9770b3a),
	.w1(32'hba7da6b3),
	.w2(32'hba7c798c),
	.w3(32'hba5c18c8),
	.w4(32'h3acaf914),
	.w5(32'hbb74fd76),
	.w6(32'hbaebd7f4),
	.w7(32'hbad268fb),
	.w8(32'h392ce803),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39644b0d),
	.w1(32'hba83a468),
	.w2(32'hbb5b8cb4),
	.w3(32'hbad32577),
	.w4(32'hbb5a3845),
	.w5(32'hbbdb7567),
	.w6(32'h3a709686),
	.w7(32'hba11fa8d),
	.w8(32'hbb3e4943),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb146a86),
	.w1(32'hba1cd685),
	.w2(32'h3b972ee9),
	.w3(32'hbbee0d24),
	.w4(32'hbb5d26cd),
	.w5(32'h3b90be3c),
	.w6(32'hbc03de66),
	.w7(32'h3af57aed),
	.w8(32'h3bc7ed0b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a6e24),
	.w1(32'hb5b4ae80),
	.w2(32'hbabbe639),
	.w3(32'h3b0fbd52),
	.w4(32'hbb0d197d),
	.w5(32'hbaebf673),
	.w6(32'h3b641e79),
	.w7(32'hba886190),
	.w8(32'hbaaf2279),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba850bad),
	.w1(32'h3c3aadb1),
	.w2(32'h3bc641e7),
	.w3(32'hba425cab),
	.w4(32'h3c1fc031),
	.w5(32'h3b975a65),
	.w6(32'hbac9efda),
	.w7(32'h3c01117d),
	.w8(32'h3bc4451a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc30c3),
	.w1(32'h3c1c6dff),
	.w2(32'h3bf83c6f),
	.w3(32'h3b3af1c2),
	.w4(32'h3bc2698b),
	.w5(32'h3c151a7e),
	.w6(32'h3c053988),
	.w7(32'h3c0377fb),
	.w8(32'h3c2a5b79),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1b5de),
	.w1(32'h3b0be0d3),
	.w2(32'h3ac99209),
	.w3(32'hba2305ea),
	.w4(32'hbc41f424),
	.w5(32'hbb4cb0f8),
	.w6(32'hbacdd4c8),
	.w7(32'hbc0a3cc1),
	.w8(32'h39666794),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb319),
	.w1(32'hba25fef7),
	.w2(32'hbb986b5f),
	.w3(32'hbb1b148f),
	.w4(32'hbb1398fd),
	.w5(32'h3a000ef0),
	.w6(32'h38f58a1e),
	.w7(32'h3ad8e5a3),
	.w8(32'hba8f4e38),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dd192),
	.w1(32'hbb3ab410),
	.w2(32'hba26084d),
	.w3(32'hb9df4497),
	.w4(32'hbad5d99a),
	.w5(32'hbade5cb0),
	.w6(32'hbaef5e6d),
	.w7(32'hbb31e378),
	.w8(32'hbaa886f0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7f7ef),
	.w1(32'h3af741fb),
	.w2(32'hba199f96),
	.w3(32'hb8bff868),
	.w4(32'h3890e215),
	.w5(32'hbb4ef6a3),
	.w6(32'hba40072c),
	.w7(32'hba8513c4),
	.w8(32'hb9c5862f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1525d3),
	.w1(32'hbb3e2f67),
	.w2(32'h38d75759),
	.w3(32'hbaa84fff),
	.w4(32'hba9fe0a2),
	.w5(32'hb9b140f6),
	.w6(32'hbb242033),
	.w7(32'hbadba21e),
	.w8(32'h3812fcd2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a8f4a),
	.w1(32'hbb12e221),
	.w2(32'hb98979cd),
	.w3(32'hbb10fb41),
	.w4(32'hbab51669),
	.w5(32'h3944c01e),
	.w6(32'hbabab5f1),
	.w7(32'hba7f9ff4),
	.w8(32'h3aca578a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0024ee),
	.w1(32'h3b2bd607),
	.w2(32'hbb1666d3),
	.w3(32'h3a5e0e2f),
	.w4(32'h3b73d2b4),
	.w5(32'h390f32c6),
	.w6(32'hb802d865),
	.w7(32'h3b82d145),
	.w8(32'h3a93ce69),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ca253),
	.w1(32'hbae22cb0),
	.w2(32'hba59335d),
	.w3(32'hbb82e575),
	.w4(32'hbb490e2a),
	.w5(32'hbb8b8845),
	.w6(32'hbbd80e63),
	.w7(32'hbbec435e),
	.w8(32'hbb61e16d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d6d71),
	.w1(32'hb9e324a8),
	.w2(32'h3b1e0868),
	.w3(32'hbab58588),
	.w4(32'hbaeb9ef3),
	.w5(32'h3b4c3556),
	.w6(32'hba0807b9),
	.w7(32'hb997cf03),
	.w8(32'h3b4c953c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b187d81),
	.w1(32'h3b9df576),
	.w2(32'h3bd617e2),
	.w3(32'h3b333614),
	.w4(32'h3b5cc744),
	.w5(32'h3be2ce36),
	.w6(32'h3b8a425f),
	.w7(32'h3b8978f1),
	.w8(32'h3bd05065),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae8a61),
	.w1(32'h3c3cfd06),
	.w2(32'h3b26e14c),
	.w3(32'h3b366841),
	.w4(32'h3c1162d0),
	.w5(32'h39e7897a),
	.w6(32'h3b647150),
	.w7(32'h3c1a16f1),
	.w8(32'h3a86111b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebd3dc),
	.w1(32'h3b05b7fd),
	.w2(32'hbb9bb604),
	.w3(32'h3a6df629),
	.w4(32'h3aec99e6),
	.w5(32'hbaa7cb8e),
	.w6(32'h3aa34cab),
	.w7(32'h3a0db765),
	.w8(32'hbae74c37),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75194f),
	.w1(32'h3b250795),
	.w2(32'h3ae1989f),
	.w3(32'hbb3fbe70),
	.w4(32'h3a917b40),
	.w5(32'h3ab64de0),
	.w6(32'hbb1135b0),
	.w7(32'h3a874143),
	.w8(32'hba579cd4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c4375),
	.w1(32'hbb2ff26a),
	.w2(32'h3ba8c0b5),
	.w3(32'hbab80815),
	.w4(32'hbb3efa14),
	.w5(32'h3bab966b),
	.w6(32'hbb1d8be8),
	.w7(32'hbb18f246),
	.w8(32'h3b71ee2a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf33b2a),
	.w1(32'h3bfa36e5),
	.w2(32'h3a84333c),
	.w3(32'h3c1ffaa2),
	.w4(32'h3c086b49),
	.w5(32'h3aaed08f),
	.w6(32'h3c0ef27c),
	.w7(32'h3c02409f),
	.w8(32'h3a4174e8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafad948),
	.w1(32'hbb6611bc),
	.w2(32'h3b6a9a45),
	.w3(32'hbbac0413),
	.w4(32'hbbbf7e26),
	.w5(32'h3b0aca11),
	.w6(32'hbb8d1b0b),
	.w7(32'hbb79cf8b),
	.w8(32'hb931ca7f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d974b),
	.w1(32'h3a2a3446),
	.w2(32'h3a91df8c),
	.w3(32'h3861555c),
	.w4(32'hb9df8c3a),
	.w5(32'h3b15de84),
	.w6(32'hbac96192),
	.w7(32'hbb8ea1aa),
	.w8(32'h3a4e4d7a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4192bd),
	.w1(32'h3a7e9b5e),
	.w2(32'hbb0b2c26),
	.w3(32'hba5884f4),
	.w4(32'h3b48547a),
	.w5(32'hbafe1b59),
	.w6(32'hb9f493ad),
	.w7(32'hba984334),
	.w8(32'hba955705),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21aa70),
	.w1(32'hba158312),
	.w2(32'hbafa5fa9),
	.w3(32'hbbaa4fdb),
	.w4(32'hbab6fb87),
	.w5(32'hbb0babbf),
	.w6(32'hbb5cb4e9),
	.w7(32'hbba549fd),
	.w8(32'hbb399d3c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a687d),
	.w1(32'h3b79b578),
	.w2(32'h3b739036),
	.w3(32'h3a63c5ec),
	.w4(32'h3b0a58b2),
	.w5(32'h3b620247),
	.w6(32'h3aad15ad),
	.w7(32'h3ae93bba),
	.w8(32'h3b6b39e3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f4459),
	.w1(32'h3b537c63),
	.w2(32'hbaeba3a4),
	.w3(32'h3b114d5f),
	.w4(32'h3b1bbc34),
	.w5(32'hbac71d16),
	.w6(32'h3a74280f),
	.w7(32'h3afb8555),
	.w8(32'hbaac6a26),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b5202),
	.w1(32'h3b2799f1),
	.w2(32'hbb6d0e7a),
	.w3(32'hbabc902e),
	.w4(32'h3b0936bc),
	.w5(32'hbb354677),
	.w6(32'hbb082e8f),
	.w7(32'h3aa5794e),
	.w8(32'hbadc6def),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba721a1f),
	.w1(32'hbb44cf16),
	.w2(32'h3aa0f57f),
	.w3(32'hb9247aa4),
	.w4(32'hbb1d880b),
	.w5(32'h3b0ff9d5),
	.w6(32'hbb091d06),
	.w7(32'hbb0e04b4),
	.w8(32'h3ac54a78),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb267de2),
	.w1(32'h39e9367e),
	.w2(32'hbae0304a),
	.w3(32'hbbe10511),
	.w4(32'h3b114428),
	.w5(32'h38f178d4),
	.w6(32'hbaeff4ad),
	.w7(32'h3a4a5081),
	.w8(32'h3b157543),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb86d90),
	.w1(32'h3bc72f0a),
	.w2(32'hbb0cc229),
	.w3(32'h393453cc),
	.w4(32'h3b675c8a),
	.w5(32'hbaeafa84),
	.w6(32'h3c0b9ac4),
	.w7(32'h3bb21301),
	.w8(32'h3b66a299),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf3b83),
	.w1(32'hbb302deb),
	.w2(32'hbb169caf),
	.w3(32'hbb1c06c4),
	.w4(32'hbb9542f1),
	.w5(32'hbadb1b00),
	.w6(32'hbadfceb5),
	.w7(32'hbb912fe5),
	.w8(32'hbb2024f6),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9697b4),
	.w1(32'hbbd67a5e),
	.w2(32'hb901d8c0),
	.w3(32'hbb8d6e8c),
	.w4(32'hbbcf832c),
	.w5(32'hb9552ad1),
	.w6(32'hbbd09b2d),
	.w7(32'hbb9b5377),
	.w8(32'h3b22df0f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a56c8),
	.w1(32'h3a59e196),
	.w2(32'hb9d7f300),
	.w3(32'h3b299350),
	.w4(32'h3b0ad984),
	.w5(32'h3b0092c0),
	.w6(32'h3b33cde9),
	.w7(32'h3a8417d1),
	.w8(32'h3ab2f8a0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c96d29),
	.w1(32'hbaa7b261),
	.w2(32'hba859113),
	.w3(32'hba0d8606),
	.w4(32'hbb20e04e),
	.w5(32'hba9e4283),
	.w6(32'h3a8bd7f9),
	.w7(32'h3b04afcc),
	.w8(32'hba944496),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9366e7),
	.w1(32'hbbaf4b27),
	.w2(32'hba04b317),
	.w3(32'hbbf48c3f),
	.w4(32'hbb3fdfbf),
	.w5(32'h3b126b6b),
	.w6(32'hbb7da7dc),
	.w7(32'hbb577525),
	.w8(32'h3b941d01),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d478b),
	.w1(32'h3c141149),
	.w2(32'h3bdd6b71),
	.w3(32'h3bbb4319),
	.w4(32'h3c09cf44),
	.w5(32'h3b4c5957),
	.w6(32'h3bd109f3),
	.w7(32'h3c5d6a9f),
	.w8(32'h3b938c47),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a085dda),
	.w1(32'h3a3885d6),
	.w2(32'h3b82da1c),
	.w3(32'hbb1a3f09),
	.w4(32'h3b0c0096),
	.w5(32'h3b76350e),
	.w6(32'h3a412a0d),
	.w7(32'h3b824219),
	.w8(32'h3ba929ce),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e05a),
	.w1(32'h3b6b768a),
	.w2(32'h3bae1f58),
	.w3(32'h3b0017b9),
	.w4(32'h3a933161),
	.w5(32'h3b8417ad),
	.w6(32'h39671c46),
	.w7(32'hb8eb7364),
	.w8(32'h3b4fdec5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20d4fb),
	.w1(32'h3bee7d71),
	.w2(32'hbaa5ca82),
	.w3(32'h3be91119),
	.w4(32'h3b59344c),
	.w5(32'hb887946e),
	.w6(32'h3bb1e527),
	.w7(32'h3b62080a),
	.w8(32'h39b8af49),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a331414),
	.w1(32'hbb14b874),
	.w2(32'hba6c70c8),
	.w3(32'h3a941573),
	.w4(32'hba7602bb),
	.w5(32'hbb22e5a6),
	.w6(32'hbb26930e),
	.w7(32'hbb247e06),
	.w8(32'hbb11ed0a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980340c),
	.w1(32'hb9f0ad49),
	.w2(32'hbb5b0221),
	.w3(32'h391b42ee),
	.w4(32'hba247b7c),
	.w5(32'hbb302c78),
	.w6(32'h38744204),
	.w7(32'h3ac28580),
	.w8(32'hbab61e4f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb121e),
	.w1(32'hbb8e7aa5),
	.w2(32'h3b26acdf),
	.w3(32'hbbde8be1),
	.w4(32'hbb43a254),
	.w5(32'hba1dcaae),
	.w6(32'hbb97b36c),
	.w7(32'h3a40e591),
	.w8(32'h3afccba1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1e1ad),
	.w1(32'hbaa18996),
	.w2(32'h3b24ccbe),
	.w3(32'h3ab439e5),
	.w4(32'hbaa2a117),
	.w5(32'h3ad0ec74),
	.w6(32'h3ae980fa),
	.w7(32'hbb39e8b2),
	.w8(32'hb97f4b7c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0c5c9),
	.w1(32'hbae605cb),
	.w2(32'h3be1574e),
	.w3(32'hb9c166d1),
	.w4(32'h3a867d1b),
	.w5(32'h3c032d50),
	.w6(32'hbbaf13c1),
	.w7(32'h3b4da658),
	.w8(32'h3bd691af),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb98e5),
	.w1(32'h3bd1ada5),
	.w2(32'hbaece9b8),
	.w3(32'h3b9d7544),
	.w4(32'h3bc9897e),
	.w5(32'h3a8520b7),
	.w6(32'h3c050b8d),
	.w7(32'h3bd0a48a),
	.w8(32'hb943daa7),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaab521),
	.w1(32'hbbbd633c),
	.w2(32'hbacd0f5a),
	.w3(32'h3a34e5c5),
	.w4(32'h3a98b676),
	.w5(32'hba369aaf),
	.w6(32'hbb147643),
	.w7(32'hbb62ef6d),
	.w8(32'hbb7776a0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf99d90),
	.w1(32'h396786d4),
	.w2(32'hba2329cc),
	.w3(32'hbb109f2a),
	.w4(32'hbabfda02),
	.w5(32'h39abd5e3),
	.w6(32'hbb376da0),
	.w7(32'h39be9b71),
	.w8(32'hbac68505),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20796a),
	.w1(32'hba72538e),
	.w2(32'hb9ac7d21),
	.w3(32'hba194b63),
	.w4(32'h3b296d01),
	.w5(32'h3a7aae55),
	.w6(32'h3a9a3149),
	.w7(32'h3ba1f969),
	.w8(32'h3b87ed4b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac929e5),
	.w1(32'h3a2d7dc2),
	.w2(32'h3a274cfc),
	.w3(32'h3ac1d133),
	.w4(32'h3aba2fa2),
	.w5(32'hbaf6bade),
	.w6(32'h3ae72668),
	.w7(32'h3b69ea9d),
	.w8(32'h39f3d8c9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb728ce8),
	.w1(32'hbb846f11),
	.w2(32'h3a835762),
	.w3(32'hbbcbd5b1),
	.w4(32'hbb48b650),
	.w5(32'h3ac820ef),
	.w6(32'hbb9c21f7),
	.w7(32'h39ae7eb1),
	.w8(32'h3a550673),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab66ee7),
	.w1(32'h3b00cd70),
	.w2(32'h3a8f64e2),
	.w3(32'h3ac8bd14),
	.w4(32'h3a4207ef),
	.w5(32'hb9912dca),
	.w6(32'h3a855bcd),
	.w7(32'h3a8018cc),
	.w8(32'h39e160a6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe67aa),
	.w1(32'h3a1dc3c4),
	.w2(32'hbb27708e),
	.w3(32'hbb2a2f8b),
	.w4(32'h3b08b85e),
	.w5(32'hbb662c2f),
	.w6(32'hbb5abf0e),
	.w7(32'h3a57d9fe),
	.w8(32'hba341d41),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb27fd2),
	.w1(32'hbbafcc8b),
	.w2(32'hbb84bcc4),
	.w3(32'hbb7e93c4),
	.w4(32'hbb0f9348),
	.w5(32'hbb0ca7fa),
	.w6(32'hbacf7d9f),
	.w7(32'hb8000a34),
	.w8(32'h39af5842),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b2a48),
	.w1(32'hbaa6220c),
	.w2(32'hba3001c8),
	.w3(32'hba2533cb),
	.w4(32'h3b20c238),
	.w5(32'hbaa5026a),
	.w6(32'hbb7553f5),
	.w7(32'h3a1405db),
	.w8(32'h3b13c6e1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb4c3e),
	.w1(32'hbaac168f),
	.w2(32'h3a74afb4),
	.w3(32'hb8b092bb),
	.w4(32'hba4c91b7),
	.w5(32'h3a345609),
	.w6(32'h3b0aedac),
	.w7(32'h3abc0596),
	.w8(32'h3a9fb1e7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bf223),
	.w1(32'hbb43bb40),
	.w2(32'hba37211c),
	.w3(32'h3b034496),
	.w4(32'h3a3022d4),
	.w5(32'h3a86647d),
	.w6(32'h3b44ceef),
	.w7(32'h3ab603f5),
	.w8(32'h3aa621ae),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994d669),
	.w1(32'h3b75e0b9),
	.w2(32'hb9b8ea26),
	.w3(32'hba3d61b4),
	.w4(32'hbad7eb6a),
	.w5(32'hbaac0d85),
	.w6(32'h3b81b307),
	.w7(32'h3b750cc3),
	.w8(32'h3a162866),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6eeb0),
	.w1(32'h3b1fdb56),
	.w2(32'h3ae114e4),
	.w3(32'hba438792),
	.w4(32'hba2f1af8),
	.w5(32'h3a81c782),
	.w6(32'hbaee3217),
	.w7(32'hbb391261),
	.w8(32'h3a32a7dd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7d72b),
	.w1(32'h3b1584f1),
	.w2(32'hbabcfeb1),
	.w3(32'h3b3958fd),
	.w4(32'h3b3ec94e),
	.w5(32'hbb0d7423),
	.w6(32'h3b9b5b1d),
	.w7(32'h3b7ea266),
	.w8(32'hbad04579),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4becf3),
	.w1(32'h3b0bdebc),
	.w2(32'h39f02b3f),
	.w3(32'hba1d574c),
	.w4(32'h3ac12e1b),
	.w5(32'h3a3d44e4),
	.w6(32'h3b2d5532),
	.w7(32'h3b8d8985),
	.w8(32'h3a349c35),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c9b1c),
	.w1(32'h3abc5afe),
	.w2(32'h3b59c18e),
	.w3(32'h3a3f5191),
	.w4(32'h3b0bd014),
	.w5(32'h3a9183b8),
	.w6(32'h3afc4478),
	.w7(32'h3b2d3840),
	.w8(32'hba68b33c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b441564),
	.w1(32'h3b65226c),
	.w2(32'hbaa38f83),
	.w3(32'h3ab52dcc),
	.w4(32'h3b0ec158),
	.w5(32'hba5c2bb6),
	.w6(32'hba6e3542),
	.w7(32'h3aa9c00d),
	.w8(32'hba8180aa),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a366d),
	.w1(32'hbb37540d),
	.w2(32'hb808327f),
	.w3(32'hba894b45),
	.w4(32'hbb06b8dd),
	.w5(32'hba8ac196),
	.w6(32'hba0dfc5f),
	.w7(32'hbb2f3c19),
	.w8(32'hbb41f803),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e75b6),
	.w1(32'h3931a698),
	.w2(32'h3a3bdcaf),
	.w3(32'h3ac62ccd),
	.w4(32'hbaaeefd4),
	.w5(32'h3aac4543),
	.w6(32'h3b68beb8),
	.w7(32'h3afff84a),
	.w8(32'hbac2d77c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390212b3),
	.w1(32'hba8b0289),
	.w2(32'h3a700317),
	.w3(32'hb9cf133e),
	.w4(32'h3a144272),
	.w5(32'hbaf3da39),
	.w6(32'h3a1cf874),
	.w7(32'hb8ba0f99),
	.w8(32'h39cc082b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4e12),
	.w1(32'hbb3414ce),
	.w2(32'hb97628ab),
	.w3(32'hbb60ea9d),
	.w4(32'hbb2ae9be),
	.w5(32'hba946a21),
	.w6(32'hbb115b49),
	.w7(32'hbb85ca53),
	.w8(32'h3932aea7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afd6f5),
	.w1(32'h3a8134ff),
	.w2(32'h3b446b61),
	.w3(32'hb9fdbe83),
	.w4(32'hb9aa92b6),
	.w5(32'h3b167721),
	.w6(32'h390ddb30),
	.w7(32'hba411d23),
	.w8(32'h3af52eda),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaedbbb),
	.w1(32'h3afa7b3b),
	.w2(32'h3b08abe6),
	.w3(32'hb9112c39),
	.w4(32'h3a9a72f0),
	.w5(32'h3b1d1c5a),
	.w6(32'h39ae1c54),
	.w7(32'h3abbfbda),
	.w8(32'h3aabbc52),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ae467),
	.w1(32'h3a6e450a),
	.w2(32'hb961c9fc),
	.w3(32'hba87796e),
	.w4(32'h3ad20b44),
	.w5(32'h395f737f),
	.w6(32'hbb1def76),
	.w7(32'h3a38d274),
	.w8(32'hb91c296f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fd4d15),
	.w1(32'hbb0ecb7a),
	.w2(32'h385c7936),
	.w3(32'hba196718),
	.w4(32'hbb42b3cb),
	.w5(32'hba361fa3),
	.w6(32'hbafef259),
	.w7(32'hbb793644),
	.w8(32'hbb73f004),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b411d),
	.w1(32'hbb07b2e3),
	.w2(32'h3ba67d1e),
	.w3(32'hba425f88),
	.w4(32'hbb7ff5a7),
	.w5(32'hb95c26f7),
	.w6(32'h3b9dc82c),
	.w7(32'h3a945a80),
	.w8(32'hb904da6e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf596f4),
	.w1(32'hba2b0fca),
	.w2(32'hbb2f76f7),
	.w3(32'hbbe6445f),
	.w4(32'hbb2d1d00),
	.w5(32'hbb5a9d34),
	.w6(32'hbb7ac40e),
	.w7(32'h3b84897f),
	.w8(32'hbb2eef0f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23eaf7),
	.w1(32'h3b95522c),
	.w2(32'hbace4ffd),
	.w3(32'h3a8eafb4),
	.w4(32'h3afe322d),
	.w5(32'hbb4e632f),
	.w6(32'h3b0f1ec7),
	.w7(32'h3b41b17b),
	.w8(32'hba82fd8f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule